H   �V�\V�/@                        �V�\V�/@                        �V�\V�/@H      H   H   H            j����������΢��+�j��5���	���ȿ%8����7�D�꾂S���7�3但L��-�)��ƼE�\���ݻ�+�Gwɸ��:>w;��0;��?;}�F;+I;��I;�I;�I;G�I;�gI;NI;�;I;�/I;�(I;�&I;�(I;�/I;�;I;NI;�gI;G�I;�I;�I;��I;+I;}�F;��?;��0;>w;��:Gwɸ�+���ݻE�\��Ƽ-�)��L��3��7��S��D�꾧�7�%8����ȿ��	��5�+�j�΢����������      ��������B��Z�����c�321�#X��ÿhڇ�q�3��s��7��74�i�Gى���&�-Nür�X�?�ػ��%���J�΁�:�a;z�0;��?;8�F;�1I;�I;b�I;	�I;l�I;xgI;�MI;R;I;�/I;~(I;�&I;~(I;�/I;R;I;�MI;xgI;l�I;	�I;b�I;�I;�1I;8�F;��?;z�0;�a;΁�:��J���%�?�ػr�X�-Nü��&�Gى�i�74��7���s�q�3�hڇ��ÿ#X�321���c�Z����B�����      �����B����C��s�P���#�I�������x|��'�YD־�X��s�)�&Խ�Ă�\<�^_���-M�j ˻_����8ϑ�:�;J2;/u@;��F;�EI;��I;+�I;F�I;%�I;�eI;YLI;c:I;�.I;�'I;�%I;�'I;�.I;c:I;YLI;�eI;%�I;F�I;+�I;��I;�EI;��F;/u@;J2;�;ϑ�:��8_��j ˻�-M�^_��\<��Ă�&Խs�)��X��YD־�'��x|����I�����#�s�P�C�����B��      ΢��Z���C���/]��5�L���,ݿ)8��nm_��K��t��Y�s�'>����J�o��3��۩��:��T�������9�d�:�;;�^4;%gA;:7G;�cI;%�I;P�I;v�I;��I;JcI;7JI;�8I;l-I;�&I;�$I;�&I;l-I;�8I;7JI;JcI;��I;v�I;P�I;%�I;�cI;:7G;%gA;�^4;�;;�d�:��9����T���:��۩��3�J�o����'>�Y�s��t���K�nm_�)8���,ݿL���5��/]�C��Z���      +�j���c�s�P��5���o��E���gڇ�Dv<�&���q���_S��������+T��� �P$��+H#�W���r3���:Ư�:Q�;67;��B;��G;ֆI;6�I;��I;�I;��I;�_I;eGI;�6I;�+I;*%I;#I;*%I;�+I;�6I;eGI;�_I;��I;�I;��I;6�I;ֆI;��G;��B;67;Q�;Ư�:�:r3��W���+H#�P$���� �+T���������_S�q��&���Dv<�gڇ�E���o�����5�s�P���c�      �5�321���#�L��o���ÿ�ҕ�Z������̾�X����0�3�8W����5��zܼ������m�s��Y\�[�n:���:��%;��9;��C;.H;1�I;1�I;$�I;��I;�zI;-[I;�CI;�3I;L)I;8#I;8!I;8#I;L)I;�3I;�CI;-[I;�zI;��I;$�I;1�I;1�I;.H;��C;��9;��%;���:[�n:�Y\�m�s��������zܼ��5�8W��3佃�0��X����̾���Z��ҕ��ÿo��L����#�321�      ��	�#X�I����,ݿE����ҕ� �d��'�?��#���{�W����t���C�o��G��*���Q�(�ػ�0�>�~���:��;M,;p=;VAE;��H;��I;��I;h�I;�I;�sI;�UI;�?I;�0I;�&I;� I;�I;� I;�&I;�0I;�?I;�UI;�sI;�I;h�I;��I;��I;��H;VAE;p=;M,;��;��:>�~��0�(�ػ�Q��*���G�C�o�t������{�W�#���?�꾊'� �d��ҕ�E����,ݿI���#X�      ��ȿ�ÿ���)8��gڇ�Z��'�����l8��Y�s�0�&�`�9{??�W�A琼�G#��7���Vܺ��9U�:��;8K2;b@;��F;I;��I;��I;o�I;d�I;�kI;�OI;u;I;-I;�#I;CI;dI;CI;�#I;-I;u;I;�OI;�kI;d�I;o�I;��I;��I;I;��F;b@;8K2;��;U�:��9�Vܺ�7���G#�A琼W�{??�9`�0�&�Y�s�l8�������'�Z�gڇ�)8������ÿ      %8��hڇ��x|�nm_�Dv<����?��l8��'6~�r74��l������Inc�G��_��3�\�A:�VZ�� >���n:Z��:
#;�8;ܿB;��G;�wI;��I;��I;��I;��I;ZcI;�II;�6I;5)I;W I;lI;�I;lI;W I;5)I;�6I;�II;ZcI;��I;��I;��I;��I;�wI;��G;ܿB;�8;
#;Z��:��n:� >�VZ�A:�3�\�_��G��Inc������l��r74�'6~�l8��?�꾎��Dv<�nm_��x|�hڇ�      ��7�q�3��'��K�&�����̾#���Y�s�r74����*N���|��)�_zܼZ��� � ��R����C9釹:-�;-;$=;�E; �H;n�I;M�I;��I;ǤI;<zI;�ZI;�BI;q1I;2%I;�I;II;�I;II;�I;2%I;q1I;�BI;�ZI;<zI;ǤI;��I;M�I;n�I; �H;�E;$=;-;-�;釹:�C9R��� ��� �Z��_zܼ�)��|�*N�����r74�Y�s�#�����̾&����K��'�q�3�      D���s�YD־�t��q���X��{�W�0�&��l��*N���Ă�|�5�׃���Q��#�A���ػ��G�$&/�6f:`�:Õ;x�5;�8A;\�F;�)I;��I;��I;+�I;}�I;QnI;�QI;�;I;4,I;� I;aI;I;�I;I;aI;� I;4,I;�;I;�QI;QnI;}�I;+�I;��I;��I;�)I;\�F;�8A;x�5;Õ;`�:6f:$&/���G���ػ#�A��Q��׃��|�5��Ă�*N���l��0�&�{�W��X��q���t��YD־�s�      �S���7���X��Y�s��_S���0����`ང����|�|�5����۩���X�fc �����5����9!��:��;�,;�K<;vnD;&-H;�I;��I;��I;t�I;q�I;YbI;{HI;�4I;�&I;eI;�I;�I;�I;�I;�I;eI;�&I;�4I;{HI;YbI;q�I;t�I;��I;��I;�I;&-H;vnD;�K<;�,;��;!��:��9�5�����fc ���X�۩����|�5��|�����`ས����0��_S�Y�s��X���7��      �7�74�s�)�'>����3�t���9Inc��)�׃��۩��a�2R�ݒ��&O���ȸ$��:��;�#;��6;gA;��F;�I;Y�I;��I;0�I;��I;�tI;�VI;�?I;%.I;|!I;2I;I;�I;wI;�I;I;2I;|!I;%.I;�?I;�VI;�tI;��I;0�I;��I;Y�I;�I;��F;gA;��6;�#;��;$��:��ȸ&O�ݒ��2R��a�۩�׃���)�Inc�9t���3����'>�s�)�74�      3�i�&Խ�������8W��C�o�{??�G��_zܼ�Q����X�2R�07������Ϲ��n:�k�:!=;��0;�>;KE;qRH;c�I;��I;�I;[�I;x�I;�eI;DKI;�6I;'I;$I;I;{I;8I;Y
I;8I;{I;I;$I;'I;�6I;DKI;�eI;x�I;[�I;�I;��I;c�I;qRH;KE;�>;��0;!=;�k�:��n:�Ϲ���07��2R���X��Q��_zܼG��{??�C�o�8W���������&Խi�      �L��Gى��Ă�J�o�+T���5��G�W�_��Z��#�A�fc �ݒ��������6�J:sj�:�d;2,;��:;"4C;+kG;DI;�I;��I;��I;��I;�uI;�WI;a@I;�.I;+!I;�I;�I;�
I;I;eI;I;�
I;�I;�I;+!I;�.I;a@I;�WI;�uI;��I;��I;��I;�I;DI;+kG;"4C;��:;2,;�d;sj�:6�J:������ݒ��fc �#�A�Z��_��W��G���5�+T�J�o��Ă�Gى�      -�)���&�\<��3��� ��zܼ�*��A琼3�\�� ���ػ���&O��Ϲ6�J:xh�:u�;��(;�d8;��A;*�F;��H;=�I;��I;!�I;�I;|�I;zdI;�JI;36I;�&I;I;&I;�I;{I;�I;@I;�I;{I;�I;&I;I;�&I;36I;�JI;zdI;|�I;�I;!�I;��I;=�I;��H;*�F;��A;�d8;��(;u�;xh�:6�J:�Ϲ&O������ػ� �3�\�A琼�*���zܼ�� ��3�\<���&�      �Ƽ-Nü^_���۩�P$������Q��G#�A:� ����G��5����ȸ��n:sj�:u�;*�';�7;�u@;;�E;-uH;�I;��I;��I;]�I;��I;�pI;�TI;I>I;�,I;�I;,I;�I;�I;YI;I;7I;I;YI;�I;�I;,I;�I;�,I;I>I;�TI;�pI;��I;]�I;��I;��I;�I;-uH;;�E;�u@;�7;*�';u�;sj�:��n:��ȸ�5����G� ��A:�G#��Q����P$���۩�^_��-Nü      E�\�r�X��-M��:�+H#����(�ػ�7��VZ�R���$&/���9$��:�k�:�d;��(;�7;�@;:\E;�,H;OvI;��I;��I;��I;ܡI;�{I;�]I;�EI;3I;b$I;�I;�I;[	I;UI;7I;@�H;��H;@�H;7I;UI;[	I;�I;�I;b$I;3I;�EI;�]I;�{I;ܡI;��I;��I;��I;OvI;�,H;:\E;�@;�7;��(;�d;�k�:$��:��9$&/�R���VZ��7��(�ػ���+H#��:��-M�r�X�      ��ݻ?�ػj ˻�T��W���m�s��0��Vܺ� >��C96f:!��:��;!=;2,;�d8;�u@;:\E;HH;aI;*�I;��I;X�I;��I;y�I;fI;MI;�8I;)I;~I;�I;I;II;I;Y�H;��H;��H;��H;Y�H;I;II;I;�I;~I;)I;�8I;MI;fI;y�I;��I;X�I;��I;*�I;aI;HH;:\E;�u@;�d8;2,;!=;��;!��:6f:�C9� >��Vܺ�0�m�s�W����T��j ˻?�ػ      �+���%�_�����r3���Y\�>�~���9��n:釹:`�:��;�#;��0;��:;��A;;�E;�,H;aI;��I;��I;��I;!�I;͌I;�lI;SI; >I;I-I;�I;kI;I;tI;�I;�H;��H;�H;��H;�H;��H;�H;�I;tI;I;kI;�I;I-I; >I;SI;�lI;͌I;!�I;��I;��I;��I;aI;�,H;;�E;��A;��:;��0;�#;��;`�:釹:��n:��9>�~��Y\�r3�����_����%�      Gwɸ��J���8��9�:[�n:��:U�:Z��:-�;Õ;�,;��6;�>;"4C;*�F;-uH;OvI;*�I;��I;O�I;ݷI;n�I;�qI;�WI;JBI;1I;<#I;�I;�I;�I;XI;Q�H;?�H;��H;��H;��H;��H;��H;?�H;Q�H;XI;�I;�I;�I;<#I;1I;JBI;�WI;�qI;n�I;ݷI;O�I;��I;*�I;OvI;-uH;*�F;"4C;�>;��6;�,;Õ;-�;Z��:U�:��:[�n:�:��9��8��J�      ��:΁�:ϑ�:�d�:Ư�:���:��;��;
#;-;x�5;�K<;gA;KE;+kG;��H;�I;��I;��I;��I;ݷI;	�I;tI;�ZI;gEI;�3I;�%I;FI;�I;b	I;}I;��H;�H;��H;��H;��H;x�H;��H;��H;��H;�H;��H;}I;b	I;�I;FI;�%I;�3I;gEI;�ZI;tI;	�I;ݷI;��I;��I;��I;�I;��H;+kG;KE;gA;�K<;x�5;-;
#;��;��;���:Ư�:�d�:ϑ�:΁�:      >w;�a;�;�;;Q�;��%;M,;8K2;�8;$=;�8A;vnD;��F;qRH;DI;=�I;��I;��I;X�I;!�I;n�I;tI;u[I;�FI;�5I;�'I;�I;TI;�
I;]I;V�H;��H;]�H;�H;��H;��H;��H;��H;��H;�H;]�H;��H;V�H;]I;�
I;TI;�I;�'I;�5I;�FI;u[I;tI;n�I;!�I;X�I;��I;��I;=�I;DI;qRH;��F;vnD;�8A;$=;�8;8K2;M,;��%;Q�;�;;�;�a;      ��0;z�0;J2;�^4;67;��9;p=;b@;ܿB;�E;\�F;&-H;�I;c�I;�I;��I;��I;��I;��I;͌I;�qI;�ZI;�FI;36I;�(I;I;hI;�I;@I;��H;��H;��H;
�H; �H;��H;�H;��H;�H;��H; �H;
�H;��H;��H;��H;@I;�I;hI;I;�(I;36I;�FI;�ZI;�qI;͌I;��I;��I;��I;��I;�I;c�I;�I;&-H;\�F;�E;ܿB;b@;p=;��9;67;�^4;J2;z�0;      ��?;��?;/u@;%gA;��B;��C;VAE;��F;��G; �H;�)I;�I;Y�I;��I;��I;!�I;]�I;ܡI;y�I;�lI;�WI;gEI;�5I;�(I;qI;�I;HI;�I;� I;D�H;��H;��H;��H;7�H;�H;u�H;=�H;u�H;�H;7�H;��H;��H;��H;D�H;� I;�I;HI;�I;qI;�(I;�5I;gEI;�WI;�lI;y�I;ܡI;]�I;!�I;��I;��I;Y�I;�I;�)I; �H;��G;��F;VAE;��C;��B;%gA;/u@;��?;      }�F;8�F;��F;:7G;��G;.H;��H;I;�wI;n�I;��I;��I;��I;�I;��I;�I;��I;�{I;fI;SI;JBI;�3I;�'I;I;�I;�I;CI;� I;{�H;��H;�H;��H;��H;��H;��H; �H;��H; �H;��H;��H;��H;��H;�H;��H;{�H;� I;CI;�I;�I;I;�'I;�3I;JBI;SI;fI;�{I;��I;�I;��I;�I;��I;��I;��I;n�I;�wI;I;��H;.H;��G;:7G;��F;8�F;      +I;�1I;�EI;�cI;ֆI;1�I;��I;��I;��I;M�I;��I;��I;0�I;[�I;��I;|�I;�pI;�]I;MI; >I;1I;�%I;�I;hI;HI;CI;� I;��H;�H;	�H;��H;��H;D�H;(�H;3�H;��H;��H;��H;3�H;(�H;D�H;��H;��H;	�H;�H;��H;� I;CI;HI;hI;�I;�%I;1I; >I;MI;�]I;�pI;|�I;��I;[�I;0�I;��I;��I;M�I;��I;��I;��I;1�I;ֆI;�cI;�EI;�1I;      ��I;�I;��I;%�I;6�I;1�I;��I;��I;��I;��I;+�I;t�I;��I;x�I;�uI;zdI;�TI;�EI;�8I;I-I;<#I;FI;TI;�I;�I;� I;��H;?�H;'�H;��H;��H;�H;��H;��H;(�H;��H;��H;��H;(�H;��H;��H;�H;��H;��H;'�H;?�H;��H;� I;�I;�I;TI;FI;<#I;I-I;�8I;�EI;�TI;zdI;�uI;x�I;��I;t�I;+�I;��I;��I;��I;��I;1�I;6�I;%�I;��I;�I;      �I;b�I;+�I;P�I;��I;$�I;h�I;o�I;��I;ǤI;}�I;q�I;�tI;�eI;�WI;�JI;I>I;3I;)I;�I;�I;�I;�
I;@I;� I;{�H;�H;'�H;��H;��H;��H;��H;[�H;��H;A�H;��H;��H;��H;A�H;��H;[�H;��H;��H;��H;��H;'�H;�H;{�H;� I;@I;�
I;�I;�I;�I;)I;3I;I>I;�JI;�WI;�eI;�tI;q�I;}�I;ǤI;��I;o�I;h�I;$�I;��I;P�I;+�I;b�I;      �I;	�I;F�I;v�I;�I;��I;�I;d�I;��I;<zI;QnI;YbI;�VI;DKI;a@I;36I;�,I;b$I;~I;kI;�I;b	I;]I;��H;D�H;��H;	�H;��H;��H;��H;��H;O�H;e�H;��H;'�H;��H;��H;��H;'�H;��H;e�H;O�H;��H;��H;��H;��H;	�H;��H;D�H;��H;]I;b	I;�I;kI;~I;b$I;�,I;36I;a@I;DKI;�VI;YbI;QnI;<zI;��I;d�I;�I;��I;�I;v�I;F�I;	�I;      G�I;l�I;%�I;��I;��I;�zI;�sI;�kI;ZcI;�ZI;�QI;{HI;�?I;�6I;�.I;�&I;�I;�I;�I;I;�I;}I;V�H;��H;��H;�H;��H;��H;��H;��H;C�H;>�H;��H;��H;p�H;N�H;4�H;N�H;p�H;��H;��H;>�H;C�H;��H;��H;��H;��H;�H;��H;��H;V�H;}I;�I;I;�I;�I;�I;�&I;�.I;�6I;�?I;{HI;�QI;�ZI;ZcI;�kI;�sI;�zI;��I;��I;%�I;l�I;      �gI;xgI;�eI;JcI;�_I;-[I;�UI;�OI;�II;�BI;�;I;�4I;%.I;'I;+!I;I;,I;�I;I;tI;XI;��H;��H;��H;��H;��H;��H;�H;��H;O�H;>�H;��H;��H;7�H;��H;��H;��H;��H;��H;7�H;��H;��H;>�H;O�H;��H;�H;��H;��H;��H;��H;��H;��H;XI;tI;I;�I;,I;I;+!I;'I;%.I;�4I;�;I;�BI;�II;�OI;�UI;-[I;�_I;JcI;�eI;xgI;      NI;�MI;YLI;7JI;eGI;�CI;�?I;u;I;�6I;q1I;4,I;�&I;|!I;$I;�I;&I;�I;[	I;II;�I;Q�H;�H;]�H;
�H;��H;��H;D�H;��H;[�H;e�H;��H;��H;�H;��H;{�H;;�H;2�H;;�H;{�H;��H;�H;��H;��H;e�H;[�H;��H;D�H;��H;��H;
�H;]�H;�H;Q�H;�I;II;[	I;�I;&I;�I;$I;|!I;�&I;4,I;q1I;�6I;u;I;�?I;�CI;eGI;7JI;YLI;�MI;      �;I;R;I;c:I;�8I;�6I;�3I;�0I;-I;5)I;2%I;� I;eI;2I;I;�I;�I;�I;UI;I;�H;?�H;��H;�H; �H;7�H;��H;(�H;��H;��H;��H;��H;7�H;��H;W�H;�H;��H;��H;��H;�H;W�H;��H;7�H;��H;��H;��H;��H;(�H;��H;7�H; �H;�H;��H;?�H;�H;I;UI;�I;�I;�I;I;2I;eI;� I;2%I;5)I;-I;�0I;�3I;�6I;�8I;c:I;R;I;      �/I;�/I;�.I;l-I;�+I;L)I;�&I;�#I;W I;�I;aI;�I;I;{I;�
I;{I;YI;7I;Y�H;��H;��H;��H;��H;��H;�H;��H;3�H;(�H;A�H;'�H;p�H;��H;{�H;�H;��H;��H;��H;��H;��H;�H;{�H;��H;p�H;'�H;A�H;(�H;3�H;��H;�H;��H;��H;��H;��H;��H;Y�H;7I;YI;{I;�
I;{I;I;�I;aI;�I;W I;�#I;�&I;L)I;�+I;l-I;�.I;�/I;      �(I;~(I;�'I;�&I;*%I;8#I;� I;CI;lI;II;I;�I;�I;8I;I;�I;I;@�H;��H;�H;��H;��H;��H;�H;u�H; �H;��H;��H;��H;��H;N�H;��H;;�H;��H;��H;o�H;i�H;o�H;��H;��H;;�H;��H;N�H;��H;��H;��H;��H; �H;u�H;�H;��H;��H;��H;�H;��H;@�H;I;�I;I;8I;�I;�I;I;II;lI;CI;� I;8#I;*%I;�&I;�'I;~(I;      �&I;�&I;�%I;�$I;#I;8!I;�I;dI;�I;�I;�I;�I;wI;Y
I;eI;@I;7I;��H;��H;��H;��H;x�H;��H;��H;=�H;��H;��H;��H;��H;��H;4�H;��H;2�H;��H;��H;i�H;L�H;i�H;��H;��H;2�H;��H;4�H;��H;��H;��H;��H;��H;=�H;��H;��H;x�H;��H;��H;��H;��H;7I;@I;eI;Y
I;wI;�I;�I;�I;�I;dI;�I;8!I;#I;�$I;�%I;�&I;      �(I;~(I;�'I;�&I;*%I;8#I;� I;CI;lI;II;I;�I;�I;8I;I;�I;I;@�H;��H;�H;��H;��H;��H;�H;u�H; �H;��H;��H;��H;��H;N�H;��H;;�H;��H;��H;o�H;i�H;o�H;��H;��H;;�H;��H;N�H;��H;��H;��H;��H; �H;u�H;�H;��H;��H;��H;�H;��H;@�H;I;�I;I;8I;�I;�I;I;II;lI;CI;� I;8#I;*%I;�&I;�'I;~(I;      �/I;�/I;�.I;l-I;�+I;L)I;�&I;�#I;W I;�I;aI;�I;I;{I;�
I;{I;YI;7I;Y�H;��H;��H;��H;��H;��H;�H;��H;3�H;(�H;A�H;'�H;p�H;��H;{�H;�H;��H;��H;��H;��H;��H;�H;{�H;��H;p�H;'�H;A�H;(�H;3�H;��H;�H;��H;��H;��H;��H;��H;Y�H;7I;YI;{I;�
I;{I;I;�I;aI;�I;W I;�#I;�&I;L)I;�+I;l-I;�.I;�/I;      �;I;R;I;c:I;�8I;�6I;�3I;�0I;-I;5)I;2%I;� I;eI;2I;I;�I;�I;�I;UI;I;�H;?�H;��H;�H; �H;7�H;��H;(�H;��H;��H;��H;��H;7�H;��H;W�H;�H;��H;��H;��H;�H;W�H;��H;7�H;��H;��H;��H;��H;(�H;��H;7�H; �H;�H;��H;?�H;�H;I;UI;�I;�I;�I;I;2I;eI;� I;2%I;5)I;-I;�0I;�3I;�6I;�8I;c:I;R;I;      NI;�MI;YLI;7JI;eGI;�CI;�?I;u;I;�6I;q1I;4,I;�&I;|!I;$I;�I;&I;�I;[	I;II;�I;Q�H;�H;]�H;
�H;��H;��H;D�H;��H;[�H;e�H;��H;��H;�H;��H;{�H;;�H;2�H;;�H;{�H;��H;�H;��H;��H;e�H;[�H;��H;D�H;��H;��H;
�H;]�H;�H;Q�H;�I;II;[	I;�I;&I;�I;$I;|!I;�&I;4,I;q1I;�6I;u;I;�?I;�CI;eGI;7JI;YLI;�MI;      �gI;xgI;�eI;JcI;�_I;-[I;�UI;�OI;�II;�BI;�;I;�4I;%.I;'I;+!I;I;,I;�I;I;tI;XI;��H;��H;��H;��H;��H;��H;�H;��H;O�H;>�H;��H;��H;7�H;��H;��H;��H;��H;��H;7�H;��H;��H;>�H;O�H;��H;�H;��H;��H;��H;��H;��H;��H;XI;tI;I;�I;,I;I;+!I;'I;%.I;�4I;�;I;�BI;�II;�OI;�UI;-[I;�_I;JcI;�eI;xgI;      G�I;l�I;%�I;��I;��I;�zI;�sI;�kI;ZcI;�ZI;�QI;{HI;�?I;�6I;�.I;�&I;�I;�I;�I;I;�I;}I;V�H;��H;��H;�H;��H;��H;��H;��H;C�H;>�H;��H;��H;p�H;N�H;4�H;N�H;p�H;��H;��H;>�H;C�H;��H;��H;��H;��H;�H;��H;��H;V�H;}I;�I;I;�I;�I;�I;�&I;�.I;�6I;�?I;{HI;�QI;�ZI;ZcI;�kI;�sI;�zI;��I;��I;%�I;l�I;      �I;	�I;F�I;v�I;�I;��I;�I;d�I;��I;<zI;QnI;YbI;�VI;DKI;a@I;36I;�,I;b$I;~I;kI;�I;b	I;]I;��H;D�H;��H;	�H;��H;��H;��H;��H;O�H;e�H;��H;'�H;��H;��H;��H;'�H;��H;e�H;O�H;��H;��H;��H;��H;	�H;��H;D�H;��H;]I;b	I;�I;kI;~I;b$I;�,I;36I;a@I;DKI;�VI;YbI;QnI;<zI;��I;d�I;�I;��I;�I;v�I;F�I;	�I;      �I;b�I;+�I;P�I;��I;$�I;h�I;o�I;��I;ǤI;}�I;q�I;�tI;�eI;�WI;�JI;I>I;3I;)I;�I;�I;�I;�
I;@I;� I;{�H;�H;'�H;��H;��H;��H;��H;[�H;��H;A�H;��H;��H;��H;A�H;��H;[�H;��H;��H;��H;��H;'�H;�H;{�H;� I;@I;�
I;�I;�I;�I;)I;3I;I>I;�JI;�WI;�eI;�tI;q�I;}�I;ǤI;��I;o�I;h�I;$�I;��I;P�I;+�I;b�I;      ��I;�I;��I;%�I;6�I;1�I;��I;��I;��I;��I;+�I;t�I;��I;x�I;�uI;zdI;�TI;�EI;�8I;I-I;<#I;FI;TI;�I;�I;� I;��H;?�H;'�H;��H;��H;�H;��H;��H;(�H;��H;��H;��H;(�H;��H;��H;�H;��H;��H;'�H;?�H;��H;� I;�I;�I;TI;FI;<#I;I-I;�8I;�EI;�TI;zdI;�uI;x�I;��I;t�I;+�I;��I;��I;��I;��I;1�I;6�I;%�I;��I;�I;      +I;�1I;�EI;�cI;ֆI;1�I;��I;��I;��I;M�I;��I;��I;0�I;[�I;��I;|�I;�pI;�]I;MI; >I;1I;�%I;�I;hI;HI;CI;� I;��H;�H;	�H;��H;��H;D�H;(�H;3�H;��H;��H;��H;3�H;(�H;D�H;��H;��H;	�H;�H;��H;� I;CI;HI;hI;�I;�%I;1I; >I;MI;�]I;�pI;|�I;��I;[�I;0�I;��I;��I;M�I;��I;��I;��I;1�I;ֆI;�cI;�EI;�1I;      }�F;8�F;��F;:7G;��G;.H;��H;I;�wI;n�I;��I;��I;��I;�I;��I;�I;��I;�{I;fI;SI;JBI;�3I;�'I;I;�I;�I;CI;� I;{�H;��H;�H;��H;��H;��H;��H; �H;��H; �H;��H;��H;��H;��H;�H;��H;{�H;� I;CI;�I;�I;I;�'I;�3I;JBI;SI;fI;�{I;��I;�I;��I;�I;��I;��I;��I;n�I;�wI;I;��H;.H;��G;:7G;��F;8�F;      ��?;��?;/u@;%gA;��B;��C;VAE;��F;��G; �H;�)I;�I;Y�I;��I;��I;!�I;]�I;ܡI;y�I;�lI;�WI;gEI;�5I;�(I;qI;�I;HI;�I;� I;D�H;��H;��H;��H;7�H;�H;u�H;=�H;u�H;�H;7�H;��H;��H;��H;D�H;� I;�I;HI;�I;qI;�(I;�5I;gEI;�WI;�lI;y�I;ܡI;]�I;!�I;��I;��I;Y�I;�I;�)I; �H;��G;��F;VAE;��C;��B;%gA;/u@;��?;      ��0;z�0;J2;�^4;67;��9;p=;b@;ܿB;�E;\�F;&-H;�I;c�I;�I;��I;��I;��I;��I;͌I;�qI;�ZI;�FI;36I;�(I;I;hI;�I;@I;��H;��H;��H;
�H; �H;��H;�H;��H;�H;��H; �H;
�H;��H;��H;��H;@I;�I;hI;I;�(I;36I;�FI;�ZI;�qI;͌I;��I;��I;��I;��I;�I;c�I;�I;&-H;\�F;�E;ܿB;b@;p=;��9;67;�^4;J2;z�0;      >w;�a;�;�;;Q�;��%;M,;8K2;�8;$=;�8A;vnD;��F;qRH;DI;=�I;��I;��I;X�I;!�I;n�I;tI;u[I;�FI;�5I;�'I;�I;TI;�
I;]I;V�H;��H;]�H;�H;��H;��H;��H;��H;��H;�H;]�H;��H;V�H;]I;�
I;TI;�I;�'I;�5I;�FI;u[I;tI;n�I;!�I;X�I;��I;��I;=�I;DI;qRH;��F;vnD;�8A;$=;�8;8K2;M,;��%;Q�;�;;�;�a;      ��:΁�:ϑ�:�d�:Ư�:���:��;��;
#;-;x�5;�K<;gA;KE;+kG;��H;�I;��I;��I;��I;ݷI;	�I;tI;�ZI;gEI;�3I;�%I;FI;�I;b	I;}I;��H;�H;��H;��H;��H;x�H;��H;��H;��H;�H;��H;}I;b	I;�I;FI;�%I;�3I;gEI;�ZI;tI;	�I;ݷI;��I;��I;��I;�I;��H;+kG;KE;gA;�K<;x�5;-;
#;��;��;���:Ư�:�d�:ϑ�:΁�:      Gwɸ��J���8��9�:[�n:��:U�:Z��:-�;Õ;�,;��6;�>;"4C;*�F;-uH;OvI;*�I;��I;O�I;ݷI;n�I;�qI;�WI;JBI;1I;<#I;�I;�I;�I;XI;Q�H;?�H;��H;��H;��H;��H;��H;?�H;Q�H;XI;�I;�I;�I;<#I;1I;JBI;�WI;�qI;n�I;ݷI;O�I;��I;*�I;OvI;-uH;*�F;"4C;�>;��6;�,;Õ;-�;Z��:U�:��:[�n:�:��9��8��J�      �+���%�_�����r3���Y\�>�~���9��n:釹:`�:��;�#;��0;��:;��A;;�E;�,H;aI;��I;��I;��I;!�I;͌I;�lI;SI; >I;I-I;�I;kI;I;tI;�I;�H;��H;�H;��H;�H;��H;�H;�I;tI;I;kI;�I;I-I; >I;SI;�lI;͌I;!�I;��I;��I;��I;aI;�,H;;�E;��A;��:;��0;�#;��;`�:釹:��n:��9>�~��Y\�r3�����_����%�      ��ݻ?�ػj ˻�T��W���m�s��0��Vܺ� >��C96f:!��:��;!=;2,;�d8;�u@;:\E;HH;aI;*�I;��I;X�I;��I;y�I;fI;MI;�8I;)I;~I;�I;I;II;I;Y�H;��H;��H;��H;Y�H;I;II;I;�I;~I;)I;�8I;MI;fI;y�I;��I;X�I;��I;*�I;aI;HH;:\E;�u@;�d8;2,;!=;��;!��:6f:�C9� >��Vܺ�0�m�s�W����T��j ˻?�ػ      E�\�r�X��-M��:�+H#����(�ػ�7��VZ�R���$&/���9$��:�k�:�d;��(;�7;�@;:\E;�,H;OvI;��I;��I;��I;ܡI;�{I;�]I;�EI;3I;b$I;�I;�I;[	I;UI;7I;@�H;��H;@�H;7I;UI;[	I;�I;�I;b$I;3I;�EI;�]I;�{I;ܡI;��I;��I;��I;OvI;�,H;:\E;�@;�7;��(;�d;�k�:$��:��9$&/�R���VZ��7��(�ػ���+H#��:��-M�r�X�      �Ƽ-Nü^_���۩�P$������Q��G#�A:� ����G��5����ȸ��n:sj�:u�;*�';�7;�u@;;�E;-uH;�I;��I;��I;]�I;��I;�pI;�TI;I>I;�,I;�I;,I;�I;�I;YI;I;7I;I;YI;�I;�I;,I;�I;�,I;I>I;�TI;�pI;��I;]�I;��I;��I;�I;-uH;;�E;�u@;�7;*�';u�;sj�:��n:��ȸ�5����G� ��A:�G#��Q����P$���۩�^_��-Nü      -�)���&�\<��3��� ��zܼ�*��A琼3�\�� ���ػ���&O��Ϲ6�J:xh�:u�;��(;�d8;��A;*�F;��H;=�I;��I;!�I;�I;|�I;zdI;�JI;36I;�&I;I;&I;�I;{I;�I;@I;�I;{I;�I;&I;I;�&I;36I;�JI;zdI;|�I;�I;!�I;��I;=�I;��H;*�F;��A;�d8;��(;u�;xh�:6�J:�Ϲ&O������ػ� �3�\�A琼�*���zܼ�� ��3�\<���&�      �L��Gى��Ă�J�o�+T���5��G�W�_��Z��#�A�fc �ݒ��������6�J:sj�:�d;2,;��:;"4C;+kG;DI;�I;��I;��I;��I;�uI;�WI;a@I;�.I;+!I;�I;�I;�
I;I;eI;I;�
I;�I;�I;+!I;�.I;a@I;�WI;�uI;��I;��I;��I;�I;DI;+kG;"4C;��:;2,;�d;sj�:6�J:������ݒ��fc �#�A�Z��_��W��G���5�+T�J�o��Ă�Gى�      3�i�&Խ�������8W��C�o�{??�G��_zܼ�Q����X�2R�07������Ϲ��n:�k�:!=;��0;�>;KE;qRH;c�I;��I;�I;[�I;x�I;�eI;DKI;�6I;'I;$I;I;{I;8I;Y
I;8I;{I;I;$I;'I;�6I;DKI;�eI;x�I;[�I;�I;��I;c�I;qRH;KE;�>;��0;!=;�k�:��n:�Ϲ���07��2R���X��Q��_zܼG��{??�C�o�8W���������&Խi�      �7�74�s�)�'>����3�t���9Inc��)�׃��۩��a�2R�ݒ��&O���ȸ$��:��;�#;��6;gA;��F;�I;Y�I;��I;0�I;��I;�tI;�VI;�?I;%.I;|!I;2I;I;�I;wI;�I;I;2I;|!I;%.I;�?I;�VI;�tI;��I;0�I;��I;Y�I;�I;��F;gA;��6;�#;��;$��:��ȸ&O�ݒ��2R��a�۩�׃���)�Inc�9t���3����'>�s�)�74�      �S���7���X��Y�s��_S���0����`ང����|�|�5����۩���X�fc �����5����9!��:��;�,;�K<;vnD;&-H;�I;��I;��I;t�I;q�I;YbI;{HI;�4I;�&I;eI;�I;�I;�I;�I;�I;eI;�&I;�4I;{HI;YbI;q�I;t�I;��I;��I;�I;&-H;vnD;�K<;�,;��;!��:��9�5�����fc ���X�۩����|�5��|�����`ས����0��_S�Y�s��X���7��      D���s�YD־�t��q���X��{�W�0�&��l��*N���Ă�|�5�׃���Q��#�A���ػ��G�$&/�6f:`�:Õ;x�5;�8A;\�F;�)I;��I;��I;+�I;}�I;QnI;�QI;�;I;4,I;� I;aI;I;�I;I;aI;� I;4,I;�;I;�QI;QnI;}�I;+�I;��I;��I;�)I;\�F;�8A;x�5;Õ;`�:6f:$&/���G���ػ#�A��Q��׃��|�5��Ă�*N���l��0�&�{�W��X��q���t��YD־�s�      ��7�q�3��'��K�&�����̾#���Y�s�r74����*N���|��)�_zܼZ��� � ��R����C9釹:-�;-;$=;�E; �H;n�I;M�I;��I;ǤI;<zI;�ZI;�BI;q1I;2%I;�I;II;�I;II;�I;2%I;q1I;�BI;�ZI;<zI;ǤI;��I;M�I;n�I; �H;�E;$=;-;-�;釹:�C9R��� ��� �Z��_zܼ�)��|�*N�����r74�Y�s�#�����̾&����K��'�q�3�      %8��hڇ��x|�nm_�Dv<����?��l8��'6~�r74��l������Inc�G��_��3�\�A:�VZ�� >���n:Z��:
#;�8;ܿB;��G;�wI;��I;��I;��I;��I;ZcI;�II;�6I;5)I;W I;lI;�I;lI;W I;5)I;�6I;�II;ZcI;��I;��I;��I;��I;�wI;��G;ܿB;�8;
#;Z��:��n:� >�VZ�A:�3�\�_��G��Inc������l��r74�'6~�l8��?�꾎��Dv<�nm_��x|�hڇ�      ��ȿ�ÿ���)8��gڇ�Z��'�����l8��Y�s�0�&�`�9{??�W�A琼�G#��7���Vܺ��9U�:��;8K2;b@;��F;I;��I;��I;o�I;d�I;�kI;�OI;u;I;-I;�#I;CI;dI;CI;�#I;-I;u;I;�OI;�kI;d�I;o�I;��I;��I;I;��F;b@;8K2;��;U�:��9�Vܺ�7���G#�A琼W�{??�9`�0�&�Y�s�l8�������'�Z�gڇ�)8������ÿ      ��	�#X�I����,ݿE����ҕ� �d��'�?��#���{�W����t���C�o��G��*���Q�(�ػ�0�>�~���:��;M,;p=;VAE;��H;��I;��I;h�I;�I;�sI;�UI;�?I;�0I;�&I;� I;�I;� I;�&I;�0I;�?I;�UI;�sI;�I;h�I;��I;��I;��H;VAE;p=;M,;��;��:>�~��0�(�ػ�Q��*���G�C�o�t������{�W�#���?�꾊'� �d��ҕ�E����,ݿI���#X�      �5�321���#�L��o���ÿ�ҕ�Z������̾�X����0�3�8W����5��zܼ������m�s��Y\�[�n:���:��%;��9;��C;.H;1�I;1�I;$�I;��I;�zI;-[I;�CI;�3I;L)I;8#I;8!I;8#I;L)I;�3I;�CI;-[I;�zI;��I;$�I;1�I;1�I;.H;��C;��9;��%;���:[�n:�Y\�m�s��������zܼ��5�8W��3佃�0��X����̾���Z��ҕ��ÿo��L����#�321�      +�j���c�s�P��5���o��E���gڇ�Dv<�&���q���_S��������+T��� �P$��+H#�W���r3���:Ư�:Q�;67;��B;��G;ֆI;6�I;��I;�I;��I;�_I;eGI;�6I;�+I;*%I;#I;*%I;�+I;�6I;eGI;�_I;��I;�I;��I;6�I;ֆI;��G;��B;67;Q�;Ư�:�:r3��W���+H#�P$���� �+T���������_S�q��&���Dv<�gڇ�E���o�����5�s�P���c�      ΢��Z���C���/]��5�L���,ݿ)8��nm_��K��t��Y�s�'>����J�o��3��۩��:��T�������9�d�:�;;�^4;%gA;:7G;�cI;%�I;P�I;v�I;��I;JcI;7JI;�8I;l-I;�&I;�$I;�&I;l-I;�8I;7JI;JcI;��I;v�I;P�I;%�I;�cI;:7G;%gA;�^4;�;;�d�:��9����T���:��۩��3�J�o����'>�Y�s��t���K�nm_�)8���,ݿL���5��/]�C��Z���      �����B����C��s�P���#�I�������x|��'�YD־�X��s�)�&Խ�Ă�\<�^_���-M�j ˻_����8ϑ�:�;J2;/u@;��F;�EI;��I;+�I;F�I;%�I;�eI;YLI;c:I;�.I;�'I;�%I;�'I;�.I;c:I;YLI;�eI;%�I;F�I;+�I;��I;�EI;��F;/u@;J2;�;ϑ�:��8_��j ˻�-M�^_��\<��Ă�&Խs�)��X��YD־�'��x|����I�����#�s�P�C�����B��      ��������B��Z�����c�321�#X��ÿhڇ�q�3��s��7��74�i�Gى���&�-Nür�X�?�ػ��%���J�΁�:�a;z�0;��?;8�F;�1I;�I;b�I;	�I;l�I;xgI;�MI;R;I;�/I;~(I;�&I;~(I;�/I;R;I;�MI;xgI;l�I;	�I;b�I;�I;�1I;8�F;��?;z�0;�a;΁�:��J���%�?�ػr�X�-Nü��&�Gى�i�74��7���s�q�3�hڇ��ÿ#X�321���c�Z����B�����      A(��o'���o��L�d��X1�|x�Ŀ����3�v���x����4�s��b+���'�"�ü�yY�mlٻq&���p�W��:^;��0;��?;�F;tI;�I;��I;H�I;��I;ucI;�JI;�8I;�-I;�&I;�$I;�&I;�-I;�8I;�JI;ucI;��I;H�I;��I;�I;tI;�F;��?;��0;^;W��:��p�q&�mlٻ�yY�"�ü�'�b+��s����4��x��v���3����Ŀ|x��X1�d�L��o��o'��      o'���X��c^�������]]���,�N9�3g��S�����/����o��j1��hܽ���-$��l��,}U��Ի!���-���:;�41;��?;l�F;N&I;��I;6�I;Y�I;ąI;�bI;\JI;�8I;E-I;�&I;�$I;�&I;E-I;�8I;\JI;�bI;ąI;Y�I;6�I;��I;N&I;l�F;��?;�41;;��:��-�!��Ի,}U��l���-$����hܽj1��o���྘�/�S���3g��N9���,��]]�����c^���X��      �o��c^���ē��4z�1K�e��M��$ﱿQ�v��X#���Ѿń�	�&�x�нk̀�r��������I� ǻ�5��9�
�:W�; �2;��@;�F;:I;�I;�I;��I;��I;qaI;II;�7I;~,I;�%I;�#I;�%I;~,I;�7I;II;qaI;��I;��I;�I;�I;:I;�F;��@; �2;W�;�
�:�9�5� ǻ��I�����r��k̀�x�н	�&�ń���Ѿ�X#�Q�v�$ﱿM��e��1K��4z��ē�c^��      L������4z���V��X1��<�pؿ����RZ��	�(���KUo����fy��?l�l�S����7������𺞽�9��:��;\�4;�sA;�1G;�WI;��I;r�I;)�I;�I;�^I;GI;A6I;+I;�$I;�"I;�$I;+I;A6I;GI;�^I;�I;)�I;r�I;��I;�WI;�1G;�sA;\�4;��;��:���9�𺙼����7�S��l�?l�fy�����KUo�(����	��RZ����pؿ�<��X1���V��4z�����      d��]]�1K��X1�Xf���kQ��S���Z58��A���נ���O���h什�Q�,���cߓ��� �W��~谺�":��:# ;�/7;�B;_�G;{I;�I;��I;ԦI;\{I;Y[I;hDI;;4I;X)I;Q#I;G!I;Q#I;X)I;;4I;hDI;Y[I;\{I;ԦI;��I;�I;{I;_�G;�B;�/7;# ;��:�":~谺W���� �cߓ�,����Q�h什����O��נ��A��Z58�S���kQ����Xf��X1�1K��]]�      �X1���,�e���<���2g��c_���U�˂�ՌȾ	ń�-�-�q��Y ��8�2�/?ټ��{�G"��n��O���u:�O ;�&;5":;[�C;!%H;0�I;C�I;��I;�I;�uI;�VI;AI;�1I;3'I;c!I;|I;c!I;3'I;�1I;AI;�VI;�uI;�I;��I;C�I;0�I;!%H;[�C;5":;�&;�O ;��u:�O��n�G"���{�/?ټ8�2�Y ��q��-�-�	ń�ՌȾ˂��U�c_��2g���<�e����,�      |x�N9�M��pؿkQ��c_��4�_��X#�p���f��<�S�{�����-l�T�-w��f�M�#�Ի�+��LT���:�d;�[,;/=;�AE;|�H;��I;��I;��I;֕I;�nI;�QI;/=I;{.I;�$I;I;bI;I;�$I;{.I;/=I;�QI;�nI;֕I;��I;��I;��I;|�H;�AE;/=;�[,;�d;��:�LT��+�#�Իf�M�-w��T�-l�����{�<�S��f��p���X#�4�_�c_��kQ��pؿM��N9�      Ŀ3g��$ﱿ���S����U��X#�s��d���JUo�
�#��hܽ����n<����`���Ӊ �<❻K�Ժ�l�9p��:�U;�2;�@;s�F;�I;�I;b�I;J�I;��I;$gI;.LI;�8I;+I;�!I;�I;�I;�I;�!I;+I;�8I;.LI;$gI;��I;J�I;b�I;�I;�I;s�F;�@;�2;�U;p��:�l�9K�Ժ<❻Ӊ �`�������n<�����hܽ
�#�JUo�d���s���X#��U�S������$ﱿ3g��      ���S���Q�v��RZ�Z58�˂�p��d���hoy�`1�gO��d什�`�`��7����yY���컟�T��1���u:��:[~#;-88;�B;��G;lI;,�I;!�I;L�I;��I;�^I;!FI;4I;C'I;�I;�I;)I;�I;�I;C'I;4I;!FI;�^I;��I;L�I;!�I;,�I;lI;��G;�B;-88;[~#;��:��u:�1���T���컷yY�7���`���`�d什gO��`1�hoy�d���p��˂�Z58��RZ�Q�v�S���      �3���/��X#��	��A��ՌȾ�f��JUo�`1�Ӱ���n���x��'��>ټ�@��.l�T���'���39�!�::Q; d-;�.=;�E;~wH;��I;,�I;��I;�I;5uI;�VI;�?I;/I;B#I;_I;�I;SI;�I;_I;B#I;/I;�?I;�VI;5uI;�I;��I;,�I;��I;~wH;�E;�.=; d-;:Q;�!�:�39'��T���.l��@���>ټ�'��x��n��Ӱ��`1�JUo��f��ՌȾ�A���	��X#���/�      v���ྃ�Ѿ(����נ�	ń�<�S�
�#�gO���n��R̀��2�-������>���Ի��B��#�Wm:�E�:n ;��5;�EA;��F;�I;r�I;o�I;ĽI;��I;�iI;�MI;.9I;�)I;I;�I;�I;iI;�I;�I;I;�)I;.9I;�MI;�iI;��I;ĽI;o�I;r�I;�I;��F;�EA;��5;n ;�E�:Wm:�#���B���Ի��>���-���2�R̀��n��gO��
�#�<�S�	ń��נ�(�����Ѿ��      �x���o��ń�KUo���O�-�-�{��hܽd什�x��2��b��yR���|U��2�����%찺�m�9��:C;��,;�g<;�qD;g$H;�I;��I;��I;&�I;%I;�]I;(EI;r2I;�$I;�I;}I;�I;PI;�I;}I;�I;�$I;r2I;(EI;�]I;%I;&�I;��I;��I;�I;g$H;�qD;�g<;��,;C;��:�m�9%찺����2���|U�yR���b���2��x�d什�hܽ{�-�-���O�KUo�ń��o��      ��4�j1�	�&������q�ཌྷ�������`��'�-��yR����]�����V��
[����o����:z�;<~#;/�6;msA;r�F;�I;��I;��I;��I;6�I;�oI;�RI;�<I;�+I;�I;�I;�I;`I;VI;`I;�I;�I;�I;�+I;�<I;�RI;�oI;6�I;��I;��I;��I;�I;r�F;msA;/�6;<~#;z�;���:��o�
[���V�������]�yR��-��'��`��������q�������	�&�j1�      s�ཾhܽx�нfy��h什Y ��-l��n<�`���>ټ�𛼞|U����H᝻�2�������u:hj�:�;|61;j(>;rE;+IH;p�I;��I;��I;�I;��I;zaI;�GI;G4I;~%I;�I;�I;WI;<
I;6	I;<
I;WI;�I;�I;~%I;G4I;�GI;zaI;��I;�I;��I;��I;p�I;+IH;rE;j(>;|61;�;hj�:��u:�����2�H᝻����|U����>ټ`���n<�-l�Y ��h什fy��x�н�hܽ      b+����k̀�?l��Q�8�2�T����7����@����>��2���V���2���� R:���:�;�[,;O;;;C;�dG;w8I;��I;U�I;��I;^�I;�pI;�SI;=I;W,I;KI;�I;�I;�	I;*I;'I;*I;�	I;�I;�I;KI;W,I;=I;�SI;�pI;^�I;��I;U�I;��I;w8I;�dG;;C;O;;�[,;�;���: R:���2��V���2����>��@��7������T�8�2��Q�?l�k̀���      �'��-$�r��l�,���/?ټ-w��`����yY�.l���Ի���
[������ R:���:�Q;�);�8;��A;�F;R�H;I�I;��I;��I;ȨI;$�I;�_I;GI;�3I;�$I;cI;�I;�
I;�I;*I;]I;*I;�I;�
I;�I;cI;�$I;�3I;GI;�_I;$�I;ȨI;��I;��I;I�I;R�H;�F;��A;�8;�);�Q;���: R:����
[�������Ի.l��yY�`���-w��/?ټ,���l�r���-$�      "�ü�l������S��cߓ���{�f�M�Ӊ ����T�����B�%찺��o���u:���:�Q;D�';)07;Մ@;�E;�kH;M�I;��I;��I;+�I;��I;�kI;�PI;C;I;�*I;�I;�I;|I;�I;ZI;CI;� I;CI;ZI;�I;|I;�I;�I;�*I;C;I;�PI;�kI;��I;+�I;��I;��I;M�I;�kH;�E;Մ@;)07;D�';�Q;���:��u:��o�%찺��B�T������Ӊ �f�M���{�cߓ�S�������l��      �yY�,}U���I���7��� �G"�#�Ի<❻��T�'���#��m�9���:hj�:�;�);)07;C@;U\E;�#H;�jI;'�I;r�I;�I;L�I;�vI;�YI;�BI;�0I;g"I;CI;�I;DI;�I;N I;�H;�H;�H;N I;�I;DI;�I;CI;g"I;�0I;�BI;�YI;�vI;L�I;�I;r�I;'�I;�jI;�#H;U\E;C@;)07;�);�;hj�:���:�m�9�#�'���T�<❻#�ԻG"��� ���7���I�,}U�      mlٻ�Ի ǻ����W���n��+�K�Ժ�1��39Wm:��:z�;�;�[,;�8;Մ@;U\E;�	H;iUI;��I;	�I;�I;}�I;#�I;�aI;}II;>6I;�&I;�I;GI;�	I;NI;O I;{�H;��H;��H;��H;{�H;O I;NI;�	I;GI;�I;�&I;>6I;}II;�aI;#�I;}�I;�I;	�I;��I;iUI;�	H;U\E;Մ@;�8;�[,;�;z�;��:Wm:�39�1�K�Ժ�+��n�W������ ǻ�Ի      q&�!��5���~谺�O��LT��l�9��u:�!�:�E�:C;<~#;|61;O;;��A;�E;�#H;iUI;,�I;��I;0�I;��I;�I;-hI;BOI;6;I;+I;3I;�I;�I;�I;� I;F�H;��H;��H;�H;��H;��H;F�H;� I;�I;�I;�I;3I;+I;6;I;BOI;-hI;�I;��I;0�I;��I;,�I;iUI;�#H;�E;��A;O;;|61;<~#;C;�E�:�!�:��u:�l�9�LT��O�~谺���5�!�      ��p���-��9���9�":��u:��:p��:��::Q;n ;��,;/�6;j(>;;C;�F;�kH;�jI;��I;��I;��I;3�I;��I;�lI;�SI;>?I;�.I;8!I;nI;�I;�I;�I;��H;��H;��H;c�H;��H;c�H;��H;��H;��H;�I;�I;�I;nI;8!I;�.I;>?I;�SI;�lI;��I;3�I;��I;��I;��I;�jI;�kH;�F;;C;j(>;/�6;��,;n ;:Q;��:p��:��:��u:�":���9�9��-�      W��:��:�
�:��:��:�O ;�d;�U;[~#; d-;��5;�g<;msA;rE;�dG;R�H;M�I;'�I;	�I;0�I;3�I;�I;!oI;aVI;BI;X1I;�#I;�I;�I;VI;�I;�H;��H;�H;f�H;>�H;��H;>�H;f�H;�H;��H;�H;�I;VI;�I;�I;�#I;X1I;BI;aVI;!oI;�I;3�I;0�I;	�I;'�I;M�I;R�H;�dG;rE;msA;�g<;��5; d-;[~#;�U;�d;�O ;��:��:�
�:��:      ^;;W�;��;# ;�&;�[,;�2;-88;�.=;�EA;�qD;r�F;+IH;w8I;I�I;��I;r�I;�I;��I;��I;!oI;bWI;�CI;3I;r%I;7I;�I;�	I;�I;��H;��H;��H;��H;G�H;V�H;�H;V�H;G�H;��H;��H;��H;��H;�I;�	I;�I;7I;r%I;3I;�CI;bWI;!oI;��I;��I;�I;r�I;��I;I�I;w8I;+IH;r�F;�qD;�EA;�.=;-88;�2;�[,;�&;# ;��;W�;;      ��0;�41; �2;\�4;�/7;5":;/=;�@;�B;�E;��F;g$H;�I;p�I;��I;��I;��I;�I;}�I;�I;�lI;aVI;�CI;�3I;Y&I;DI;I;�
I;II;>�H;A�H;��H;��H;��H;o�H;��H;w�H;��H;o�H;��H;��H;��H;A�H;>�H;II;�
I;I;DI;Y&I;�3I;�CI;aVI;�lI;�I;}�I;�I;��I;��I;��I;p�I;�I;g$H;��F;�E;�B;�@;/=;5":;�/7;\�4; �2;�41;      ��?;��?;��@;�sA;�B;[�C;�AE;s�F;��G;~wH;�I;�I;��I;��I;U�I;��I;+�I;L�I;#�I;-hI;�SI;BI;3I;Y&I;�I;�I;(I;�I;��H;��H;%�H;z�H;p�H;��H;��H;5�H;�H;5�H;��H;��H;p�H;z�H;%�H;��H;��H;�I;(I;�I;�I;Y&I;3I;BI;�SI;-hI;#�I;L�I;+�I;��I;U�I;��I;��I;�I;�I;~wH;��G;s�F;�AE;[�C;�B;�sA;��@;��?;      �F;l�F;�F;�1G;_�G;!%H;|�H;�I;lI;��I;r�I;��I;��I;��I;��I;ȨI;��I;�vI;�aI;BOI;>?I;X1I;r%I;DI;�I;OI;1I; I;��H;T�H;��H;c�H;��H;4�H;e�H;��H;��H;��H;e�H;4�H;��H;c�H;��H;T�H;��H; I;1I;OI;�I;DI;r%I;X1I;>?I;BOI;�aI;�vI;��I;ȨI;��I;��I;��I;��I;r�I;��I;lI;�I;|�H;!%H;_�G;�1G;�F;l�F;      tI;N&I;:I;�WI;{I;0�I;��I;�I;,�I;,�I;o�I;��I;��I;�I;^�I;$�I;�kI;�YI;}II;6;I;�.I;�#I;7I;I;(I;1I; I;��H;}�H;��H;\�H;`�H;��H;��H;�H;��H;w�H;��H;�H;��H;��H;`�H;\�H;��H;}�H;��H; I;1I;(I;I;7I;�#I;�.I;6;I;}II;�YI;�kI;$�I;^�I;�I;��I;��I;o�I;,�I;,�I;�I;��I;0�I;{I;�WI;:I;N&I;      �I;��I;�I;��I;�I;C�I;��I;b�I;!�I;��I;ĽI;&�I;6�I;��I;�pI;�_I;�PI;�BI;>6I;+I;8!I;�I;�I;�
I;�I; I;��H;y�H;��H;b�H;a�H;��H;��H;��H;��H;��H;y�H;��H;��H;��H;��H;��H;a�H;b�H;��H;y�H;��H; I;�I;�
I;�I;�I;8!I;+I;>6I;�BI;�PI;�_I;�pI;��I;6�I;&�I;ĽI;��I;!�I;b�I;��I;C�I;�I;��I;�I;��I;      ��I;6�I;�I;r�I;��I;��I;��I;J�I;L�I;�I;��I;%I;�oI;zaI;�SI;GI;C;I;�0I;�&I;3I;nI;�I;�	I;II;��H;��H;}�H;��H;X�H;[�H;��H;Z�H;K�H;��H;��H;��H;��H;��H;��H;��H;K�H;Z�H;��H;[�H;X�H;��H;}�H;��H;��H;II;�	I;�I;nI;3I;�&I;�0I;C;I;GI;�SI;zaI;�oI;%I;��I;�I;L�I;J�I;��I;��I;��I;r�I;�I;6�I;      H�I;Y�I;��I;)�I;ԦI;�I;֕I;��I;��I;5uI;�iI;�]I;�RI;�GI;=I;�3I;�*I;g"I;�I;�I;�I;VI;�I;>�H;��H;T�H;��H;b�H;[�H;��H;5�H;�H;A�H;��H;�H;��H;��H;��H;�H;��H;A�H;�H;5�H;��H;[�H;b�H;��H;T�H;��H;>�H;�I;VI;�I;�I;�I;g"I;�*I;�3I;=I;�GI;�RI;�]I;�iI;5uI;��I;��I;֕I;�I;ԦI;)�I;��I;Y�I;      ��I;ąI;��I;�I;\{I;�uI;�nI;$gI;�^I;�VI;�MI;(EI;�<I;G4I;W,I;�$I;�I;CI;GI;�I;�I;�I;��H;A�H;%�H;��H;\�H;a�H;��H;5�H;�H;�H;\�H;��H;z�H;7�H;��H;7�H;z�H;��H;\�H;�H;�H;5�H;��H;a�H;\�H;��H;%�H;A�H;��H;�I;�I;�I;GI;CI;�I;�$I;W,I;G4I;�<I;(EI;�MI;�VI;�^I;$gI;�nI;�uI;\{I;�I;��I;ąI;      ucI;�bI;qaI;�^I;Y[I;�VI;�QI;.LI;!FI;�?I;.9I;r2I;�+I;~%I;KI;cI;�I;�I;�	I;�I;�I;�H;��H;��H;z�H;c�H;`�H;��H;Z�H;�H;�H;U�H;��H;,�H;��H;��H;��H;��H;��H;,�H;��H;U�H;�H;�H;Z�H;��H;`�H;c�H;z�H;��H;��H;�H;�I;�I;�	I;�I;�I;cI;KI;~%I;�+I;r2I;.9I;�?I;!FI;.LI;�QI;�VI;Y[I;�^I;qaI;�bI;      �JI;\JI;II;GI;hDI;AI;/=I;�8I;4I;/I;�)I;�$I;�I;�I;�I;�I;|I;DI;NI;� I;��H;��H;��H;��H;p�H;��H;��H;��H;K�H;A�H;\�H;��H;�H;��H;M�H;!�H;3�H;!�H;M�H;��H;�H;��H;\�H;A�H;K�H;��H;��H;��H;p�H;��H;��H;��H;��H;� I;NI;DI;|I;�I;�I;�I;�I;�$I;�)I;/I;4I;�8I;/=I;AI;hDI;GI;II;\JI;      �8I;�8I;�7I;A6I;;4I;�1I;{.I;+I;C'I;B#I;I;�I;�I;�I;�I;�
I;�I;�I;O I;F�H;��H;�H;��H;��H;��H;4�H;��H;��H;��H;��H;��H;,�H;��H;<�H;��H;��H;��H;��H;��H;<�H;��H;,�H;��H;��H;��H;��H;��H;4�H;��H;��H;��H;�H;��H;F�H;O I;�I;�I;�
I;�I;�I;�I;�I;I;B#I;C'I;+I;{.I;�1I;;4I;A6I;�7I;�8I;      �-I;E-I;~,I;+I;X)I;3'I;�$I;�!I;�I;_I;�I;}I;�I;WI;�	I;�I;ZI;N I;{�H;��H;��H;f�H;G�H;o�H;��H;e�H;�H;��H;��H;�H;z�H;��H;M�H;��H;��H;��H;�H;��H;��H;��H;M�H;��H;z�H;�H;��H;��H;�H;e�H;��H;o�H;G�H;f�H;��H;��H;{�H;N I;ZI;�I;�	I;WI;�I;}I;�I;_I;�I;�!I;�$I;3'I;X)I;+I;~,I;E-I;      �&I;�&I;�%I;�$I;Q#I;c!I;I;�I;�I;�I;�I;�I;`I;<
I;*I;*I;CI;�H;��H;��H;c�H;>�H;V�H;��H;5�H;��H;��H;��H;��H;��H;7�H;��H;!�H;��H;��H;k�H;q�H;k�H;��H;��H;!�H;��H;7�H;��H;��H;��H;��H;��H;5�H;��H;V�H;>�H;c�H;��H;��H;�H;CI;*I;*I;<
I;`I;�I;�I;�I;�I;�I;I;c!I;Q#I;�$I;�%I;�&I;      �$I;�$I;�#I;�"I;G!I;|I;bI;�I;)I;SI;iI;PI;VI;6	I;'I;]I;� I;�H;��H;�H;��H;��H;�H;w�H;�H;��H;w�H;y�H;��H;��H;��H;��H;3�H;��H;�H;q�H;w�H;q�H;�H;��H;3�H;��H;��H;��H;��H;y�H;w�H;��H;�H;w�H;�H;��H;��H;�H;��H;�H;� I;]I;'I;6	I;VI;PI;iI;SI;)I;�I;bI;|I;G!I;�"I;�#I;�$I;      �&I;�&I;�%I;�$I;Q#I;c!I;I;�I;�I;�I;�I;�I;`I;<
I;*I;*I;CI;�H;��H;��H;c�H;>�H;V�H;��H;5�H;��H;��H;��H;��H;��H;7�H;��H;!�H;��H;��H;k�H;q�H;k�H;��H;��H;!�H;��H;7�H;��H;��H;��H;��H;��H;5�H;��H;V�H;>�H;c�H;��H;��H;�H;CI;*I;*I;<
I;`I;�I;�I;�I;�I;�I;I;c!I;Q#I;�$I;�%I;�&I;      �-I;E-I;~,I;+I;X)I;3'I;�$I;�!I;�I;_I;�I;}I;�I;WI;�	I;�I;ZI;N I;{�H;��H;��H;f�H;G�H;o�H;��H;e�H;�H;��H;��H;�H;z�H;��H;M�H;��H;��H;��H;�H;��H;��H;��H;M�H;��H;z�H;�H;��H;��H;�H;e�H;��H;o�H;G�H;f�H;��H;��H;{�H;N I;ZI;�I;�	I;WI;�I;}I;�I;_I;�I;�!I;�$I;3'I;X)I;+I;~,I;E-I;      �8I;�8I;�7I;A6I;;4I;�1I;{.I;+I;C'I;B#I;I;�I;�I;�I;�I;�
I;�I;�I;O I;F�H;��H;�H;��H;��H;��H;4�H;��H;��H;��H;��H;��H;,�H;��H;<�H;��H;��H;��H;��H;��H;<�H;��H;,�H;��H;��H;��H;��H;��H;4�H;��H;��H;��H;�H;��H;F�H;O I;�I;�I;�
I;�I;�I;�I;�I;I;B#I;C'I;+I;{.I;�1I;;4I;A6I;�7I;�8I;      �JI;\JI;II;GI;hDI;AI;/=I;�8I;4I;/I;�)I;�$I;�I;�I;�I;�I;|I;DI;NI;� I;��H;��H;��H;��H;p�H;��H;��H;��H;K�H;A�H;\�H;��H;�H;��H;M�H;!�H;3�H;!�H;M�H;��H;�H;��H;\�H;A�H;K�H;��H;��H;��H;p�H;��H;��H;��H;��H;� I;NI;DI;|I;�I;�I;�I;�I;�$I;�)I;/I;4I;�8I;/=I;AI;hDI;GI;II;\JI;      ucI;�bI;qaI;�^I;Y[I;�VI;�QI;.LI;!FI;�?I;.9I;r2I;�+I;~%I;KI;cI;�I;�I;�	I;�I;�I;�H;��H;��H;z�H;c�H;`�H;��H;Z�H;�H;�H;U�H;��H;,�H;��H;��H;��H;��H;��H;,�H;��H;U�H;�H;�H;Z�H;��H;`�H;c�H;z�H;��H;��H;�H;�I;�I;�	I;�I;�I;cI;KI;~%I;�+I;r2I;.9I;�?I;!FI;.LI;�QI;�VI;Y[I;�^I;qaI;�bI;      ��I;ąI;��I;�I;\{I;�uI;�nI;$gI;�^I;�VI;�MI;(EI;�<I;G4I;W,I;�$I;�I;CI;GI;�I;�I;�I;��H;A�H;%�H;��H;\�H;a�H;��H;5�H;�H;�H;\�H;��H;z�H;7�H;��H;7�H;z�H;��H;\�H;�H;�H;5�H;��H;a�H;\�H;��H;%�H;A�H;��H;�I;�I;�I;GI;CI;�I;�$I;W,I;G4I;�<I;(EI;�MI;�VI;�^I;$gI;�nI;�uI;\{I;�I;��I;ąI;      H�I;Y�I;��I;)�I;ԦI;�I;֕I;��I;��I;5uI;�iI;�]I;�RI;�GI;=I;�3I;�*I;g"I;�I;�I;�I;VI;�I;>�H;��H;T�H;��H;b�H;[�H;��H;5�H;�H;A�H;��H;�H;��H;��H;��H;�H;��H;A�H;�H;5�H;��H;[�H;b�H;��H;T�H;��H;>�H;�I;VI;�I;�I;�I;g"I;�*I;�3I;=I;�GI;�RI;�]I;�iI;5uI;��I;��I;֕I;�I;ԦI;)�I;��I;Y�I;      ��I;6�I;�I;r�I;��I;��I;��I;J�I;L�I;�I;��I;%I;�oI;zaI;�SI;GI;C;I;�0I;�&I;3I;nI;�I;�	I;II;��H;��H;}�H;��H;X�H;[�H;��H;Z�H;K�H;��H;��H;��H;��H;��H;��H;��H;K�H;Z�H;��H;[�H;X�H;��H;}�H;��H;��H;II;�	I;�I;nI;3I;�&I;�0I;C;I;GI;�SI;zaI;�oI;%I;��I;�I;L�I;J�I;��I;��I;��I;r�I;�I;6�I;      �I;��I;�I;��I;�I;C�I;��I;b�I;!�I;��I;ĽI;&�I;6�I;��I;�pI;�_I;�PI;�BI;>6I;+I;8!I;�I;�I;�
I;�I; I;��H;y�H;��H;b�H;a�H;��H;��H;��H;��H;��H;y�H;��H;��H;��H;��H;��H;a�H;b�H;��H;y�H;��H; I;�I;�
I;�I;�I;8!I;+I;>6I;�BI;�PI;�_I;�pI;��I;6�I;&�I;ĽI;��I;!�I;b�I;��I;C�I;�I;��I;�I;��I;      tI;N&I;:I;�WI;{I;0�I;��I;�I;,�I;,�I;o�I;��I;��I;�I;^�I;$�I;�kI;�YI;}II;6;I;�.I;�#I;7I;I;(I;1I; I;��H;}�H;��H;\�H;`�H;��H;��H;�H;��H;w�H;��H;�H;��H;��H;`�H;\�H;��H;}�H;��H; I;1I;(I;I;7I;�#I;�.I;6;I;}II;�YI;�kI;$�I;^�I;�I;��I;��I;o�I;,�I;,�I;�I;��I;0�I;{I;�WI;:I;N&I;      �F;l�F;�F;�1G;_�G;!%H;|�H;�I;lI;��I;r�I;��I;��I;��I;��I;ȨI;��I;�vI;�aI;BOI;>?I;X1I;r%I;DI;�I;OI;1I; I;��H;T�H;��H;c�H;��H;4�H;e�H;��H;��H;��H;e�H;4�H;��H;c�H;��H;T�H;��H; I;1I;OI;�I;DI;r%I;X1I;>?I;BOI;�aI;�vI;��I;ȨI;��I;��I;��I;��I;r�I;��I;lI;�I;|�H;!%H;_�G;�1G;�F;l�F;      ��?;��?;��@;�sA;�B;[�C;�AE;s�F;��G;~wH;�I;�I;��I;��I;U�I;��I;+�I;L�I;#�I;-hI;�SI;BI;3I;Y&I;�I;�I;(I;�I;��H;��H;%�H;z�H;p�H;��H;��H;5�H;�H;5�H;��H;��H;p�H;z�H;%�H;��H;��H;�I;(I;�I;�I;Y&I;3I;BI;�SI;-hI;#�I;L�I;+�I;��I;U�I;��I;��I;�I;�I;~wH;��G;s�F;�AE;[�C;�B;�sA;��@;��?;      ��0;�41; �2;\�4;�/7;5":;/=;�@;�B;�E;��F;g$H;�I;p�I;��I;��I;��I;�I;}�I;�I;�lI;aVI;�CI;�3I;Y&I;DI;I;�
I;II;>�H;A�H;��H;��H;��H;o�H;��H;w�H;��H;o�H;��H;��H;��H;A�H;>�H;II;�
I;I;DI;Y&I;�3I;�CI;aVI;�lI;�I;}�I;�I;��I;��I;��I;p�I;�I;g$H;��F;�E;�B;�@;/=;5":;�/7;\�4; �2;�41;      ^;;W�;��;# ;�&;�[,;�2;-88;�.=;�EA;�qD;r�F;+IH;w8I;I�I;��I;r�I;�I;��I;��I;!oI;bWI;�CI;3I;r%I;7I;�I;�	I;�I;��H;��H;��H;��H;G�H;V�H;�H;V�H;G�H;��H;��H;��H;��H;�I;�	I;�I;7I;r%I;3I;�CI;bWI;!oI;��I;��I;�I;r�I;��I;I�I;w8I;+IH;r�F;�qD;�EA;�.=;-88;�2;�[,;�&;# ;��;W�;;      W��:��:�
�:��:��:�O ;�d;�U;[~#; d-;��5;�g<;msA;rE;�dG;R�H;M�I;'�I;	�I;0�I;3�I;�I;!oI;aVI;BI;X1I;�#I;�I;�I;VI;�I;�H;��H;�H;f�H;>�H;��H;>�H;f�H;�H;��H;�H;�I;VI;�I;�I;�#I;X1I;BI;aVI;!oI;�I;3�I;0�I;	�I;'�I;M�I;R�H;�dG;rE;msA;�g<;��5; d-;[~#;�U;�d;�O ;��:��:�
�:��:      ��p���-��9���9�":��u:��:p��:��::Q;n ;��,;/�6;j(>;;C;�F;�kH;�jI;��I;��I;��I;3�I;��I;�lI;�SI;>?I;�.I;8!I;nI;�I;�I;�I;��H;��H;��H;c�H;��H;c�H;��H;��H;��H;�I;�I;�I;nI;8!I;�.I;>?I;�SI;�lI;��I;3�I;��I;��I;��I;�jI;�kH;�F;;C;j(>;/�6;��,;n ;:Q;��:p��:��:��u:�":���9�9��-�      q&�!��5���~谺�O��LT��l�9��u:�!�:�E�:C;<~#;|61;O;;��A;�E;�#H;iUI;,�I;��I;0�I;��I;�I;-hI;BOI;6;I;+I;3I;�I;�I;�I;� I;F�H;��H;��H;�H;��H;��H;F�H;� I;�I;�I;�I;3I;+I;6;I;BOI;-hI;�I;��I;0�I;��I;,�I;iUI;�#H;�E;��A;O;;|61;<~#;C;�E�:�!�:��u:�l�9�LT��O�~谺���5�!�      mlٻ�Ի ǻ����W���n��+�K�Ժ�1��39Wm:��:z�;�;�[,;�8;Մ@;U\E;�	H;iUI;��I;	�I;�I;}�I;#�I;�aI;}II;>6I;�&I;�I;GI;�	I;NI;O I;{�H;��H;��H;��H;{�H;O I;NI;�	I;GI;�I;�&I;>6I;}II;�aI;#�I;}�I;�I;	�I;��I;iUI;�	H;U\E;Մ@;�8;�[,;�;z�;��:Wm:�39�1�K�Ժ�+��n�W������ ǻ�Ի      �yY�,}U���I���7��� �G"�#�Ի<❻��T�'���#��m�9���:hj�:�;�);)07;C@;U\E;�#H;�jI;'�I;r�I;�I;L�I;�vI;�YI;�BI;�0I;g"I;CI;�I;DI;�I;N I;�H;�H;�H;N I;�I;DI;�I;CI;g"I;�0I;�BI;�YI;�vI;L�I;�I;r�I;'�I;�jI;�#H;U\E;C@;)07;�);�;hj�:���:�m�9�#�'���T�<❻#�ԻG"��� ���7���I�,}U�      "�ü�l������S��cߓ���{�f�M�Ӊ ����T�����B�%찺��o���u:���:�Q;D�';)07;Մ@;�E;�kH;M�I;��I;��I;+�I;��I;�kI;�PI;C;I;�*I;�I;�I;|I;�I;ZI;CI;� I;CI;ZI;�I;|I;�I;�I;�*I;C;I;�PI;�kI;��I;+�I;��I;��I;M�I;�kH;�E;Մ@;)07;D�';�Q;���:��u:��o�%찺��B�T������Ӊ �f�M���{�cߓ�S�������l��      �'��-$�r��l�,���/?ټ-w��`����yY�.l���Ի���
[������ R:���:�Q;�);�8;��A;�F;R�H;I�I;��I;��I;ȨI;$�I;�_I;GI;�3I;�$I;cI;�I;�
I;�I;*I;]I;*I;�I;�
I;�I;cI;�$I;�3I;GI;�_I;$�I;ȨI;��I;��I;I�I;R�H;�F;��A;�8;�);�Q;���: R:����
[�������Ի.l��yY�`���-w��/?ټ,���l�r���-$�      b+����k̀�?l��Q�8�2�T����7����@����>��2���V���2���� R:���:�;�[,;O;;;C;�dG;w8I;��I;U�I;��I;^�I;�pI;�SI;=I;W,I;KI;�I;�I;�	I;*I;'I;*I;�	I;�I;�I;KI;W,I;=I;�SI;�pI;^�I;��I;U�I;��I;w8I;�dG;;C;O;;�[,;�;���: R:���2��V���2����>��@��7������T�8�2��Q�?l�k̀���      s�ཾhܽx�нfy��h什Y ��-l��n<�`���>ټ�𛼞|U����H᝻�2�������u:hj�:�;|61;j(>;rE;+IH;p�I;��I;��I;�I;��I;zaI;�GI;G4I;~%I;�I;�I;WI;<
I;6	I;<
I;WI;�I;�I;~%I;G4I;�GI;zaI;��I;�I;��I;��I;p�I;+IH;rE;j(>;|61;�;hj�:��u:�����2�H᝻����|U����>ټ`���n<�-l�Y ��h什fy��x�н�hܽ      ��4�j1�	�&������q�ཌྷ�������`��'�-��yR����]�����V��
[����o����:z�;<~#;/�6;msA;r�F;�I;��I;��I;��I;6�I;�oI;�RI;�<I;�+I;�I;�I;�I;`I;VI;`I;�I;�I;�I;�+I;�<I;�RI;�oI;6�I;��I;��I;��I;�I;r�F;msA;/�6;<~#;z�;���:��o�
[���V�������]�yR��-��'��`��������q�������	�&�j1�      �x���o��ń�KUo���O�-�-�{��hܽd什�x��2��b��yR���|U��2�����%찺�m�9��:C;��,;�g<;�qD;g$H;�I;��I;��I;&�I;%I;�]I;(EI;r2I;�$I;�I;}I;�I;PI;�I;}I;�I;�$I;r2I;(EI;�]I;%I;&�I;��I;��I;�I;g$H;�qD;�g<;��,;C;��:�m�9%찺����2���|U�yR���b���2��x�d什�hܽ{�-�-���O�KUo�ń��o��      v���ྃ�Ѿ(����נ�	ń�<�S�
�#�gO���n��R̀��2�-������>���Ի��B��#�Wm:�E�:n ;��5;�EA;��F;�I;r�I;o�I;ĽI;��I;�iI;�MI;.9I;�)I;I;�I;�I;iI;�I;�I;I;�)I;.9I;�MI;�iI;��I;ĽI;o�I;r�I;�I;��F;�EA;��5;n ;�E�:Wm:�#���B���Ի��>���-���2�R̀��n��gO��
�#�<�S�	ń��נ�(�����Ѿ��      �3���/��X#��	��A��ՌȾ�f��JUo�`1�Ӱ���n���x��'��>ټ�@��.l�T���'���39�!�::Q; d-;�.=;�E;~wH;��I;,�I;��I;�I;5uI;�VI;�?I;/I;B#I;_I;�I;SI;�I;_I;B#I;/I;�?I;�VI;5uI;�I;��I;,�I;��I;~wH;�E;�.=; d-;:Q;�!�:�39'��T���.l��@���>ټ�'��x��n��Ӱ��`1�JUo��f��ՌȾ�A���	��X#���/�      ���S���Q�v��RZ�Z58�˂�p��d���hoy�`1�gO��d什�`�`��7����yY���컟�T��1���u:��:[~#;-88;�B;��G;lI;,�I;!�I;L�I;��I;�^I;!FI;4I;C'I;�I;�I;)I;�I;�I;C'I;4I;!FI;�^I;��I;L�I;!�I;,�I;lI;��G;�B;-88;[~#;��:��u:�1���T���컷yY�7���`���`�d什gO��`1�hoy�d���p��˂�Z58��RZ�Q�v�S���      Ŀ3g��$ﱿ���S����U��X#�s��d���JUo�
�#��hܽ����n<����`���Ӊ �<❻K�Ժ�l�9p��:�U;�2;�@;s�F;�I;�I;b�I;J�I;��I;$gI;.LI;�8I;+I;�!I;�I;�I;�I;�!I;+I;�8I;.LI;$gI;��I;J�I;b�I;�I;�I;s�F;�@;�2;�U;p��:�l�9K�Ժ<❻Ӊ �`�������n<�����hܽ
�#�JUo�d���s���X#��U�S������$ﱿ3g��      |x�N9�M��pؿkQ��c_��4�_��X#�p���f��<�S�{�����-l�T�-w��f�M�#�Ի�+��LT���:�d;�[,;/=;�AE;|�H;��I;��I;��I;֕I;�nI;�QI;/=I;{.I;�$I;I;bI;I;�$I;{.I;/=I;�QI;�nI;֕I;��I;��I;��I;|�H;�AE;/=;�[,;�d;��:�LT��+�#�Իf�M�-w��T�-l�����{�<�S��f��p���X#�4�_�c_��kQ��pؿM��N9�      �X1���,�e���<���2g��c_���U�˂�ՌȾ	ń�-�-�q��Y ��8�2�/?ټ��{�G"��n��O���u:�O ;�&;5":;[�C;!%H;0�I;C�I;��I;�I;�uI;�VI;AI;�1I;3'I;c!I;|I;c!I;3'I;�1I;AI;�VI;�uI;�I;��I;C�I;0�I;!%H;[�C;5":;�&;�O ;��u:�O��n�G"���{�/?ټ8�2�Y ��q��-�-�	ń�ՌȾ˂��U�c_��2g���<�e����,�      d��]]�1K��X1�Xf���kQ��S���Z58��A���נ���O���h什�Q�,���cߓ��� �W��~谺�":��:# ;�/7;�B;_�G;{I;�I;��I;ԦI;\{I;Y[I;hDI;;4I;X)I;Q#I;G!I;Q#I;X)I;;4I;hDI;Y[I;\{I;ԦI;��I;�I;{I;_�G;�B;�/7;# ;��:�":~谺W���� �cߓ�,����Q�h什����O��נ��A��Z58�S���kQ����Xf��X1�1K��]]�      L������4z���V��X1��<�pؿ����RZ��	�(���KUo����fy��?l�l�S����7������𺞽�9��:��;\�4;�sA;�1G;�WI;��I;r�I;)�I;�I;�^I;GI;A6I;+I;�$I;�"I;�$I;+I;A6I;GI;�^I;�I;)�I;r�I;��I;�WI;�1G;�sA;\�4;��;��:���9�𺙼����7�S��l�?l�fy�����KUo�(����	��RZ����pؿ�<��X1���V��4z�����      �o��c^���ē��4z�1K�e��M��$ﱿQ�v��X#���Ѿń�	�&�x�нk̀�r��������I� ǻ�5��9�
�:W�; �2;��@;�F;:I;�I;�I;��I;��I;qaI;II;�7I;~,I;�%I;�#I;�%I;~,I;�7I;II;qaI;��I;��I;�I;�I;:I;�F;��@; �2;W�;�
�:�9�5� ǻ��I�����r��k̀�x�н	�&�ń���Ѿ�X#�Q�v�$ﱿM��e��1K��4z��ē�c^��      o'���X��c^�������]]���,�N9�3g��S�����/����o��j1��hܽ���-$��l��,}U��Ի!���-���:;�41;��?;l�F;N&I;��I;6�I;Y�I;ąI;�bI;\JI;�8I;E-I;�&I;�$I;�&I;E-I;�8I;\JI;�bI;ąI;Y�I;6�I;��I;N&I;l�F;��?;�41;;��:��-�!��Ի,}U��l���-$����hܽj1��o���྘�/�S���3g��N9���,��]]�����c^���X��      ����,������Q���F�Q�Ù$�.���~�7�}�E(�>�׾�T���L+���սr����@L��jO�9�ͻ�����l8�m�:��;T�1;��?;uF;r�H;��I;��I;��I;�uI;�VI;�@I;1I;�&I;� I;I;� I;�&I;1I;�@I;�VI;�uI;��I;��I;��I;r�H;uF;��?;T�1;��;�m�:��l8���9�ͻjO�@L����r����ս�L+��T��>�׾E(�7�}�~�.���Ù$�F�Q�Q��������,��      �,��^�� P���{��K��x �����n�����w��$���Ҿf��� (���ѽٷ��7����%�K��ɻ��ۀ�8���:��;��1;@;��F;.I;�I;3�I;ĝI;�tI;NVI;�@I;�0I;�&I;� I;�I;� I;�&I;�0I;�@I;NVI;�tI;ĝI;3�I;�I;.I;��F;@;��1;��;���:ۀ�8���ɻ%�K����7�ٷ����ѽ (�f�����Ҿ�$���w�n��������x ��K��{� P��^��      ���� P�������d���;� ����㿰���#f�b��ž��z���C�ƽ40v�e5�R����o@�	���pj��Pu9]I�:=\;�63;?�@;�F;WI;��I;{�I;o�I;�rI;�TI;^?I;0I;&I;, I;LI;, I;&I;0I;^?I;�TI;�rI;o�I;{�I;��I;WI;�F;?�@;�63;=\;]I�:�Pu9pj�	����o@�R���e5�40v�C�ƽ����z�žb��#f�������� ����;���d���� P��      Q����{���d��F�Ù$�7����ɿ,蒿��K�O���j�� Zb�H�8�����a����`���&�.�!e��X�غ¨�9�W�:UW;�15;?�A;� G;Z6I;��I;k�I;m�I;�oI;�RI;�=I;�.I;�$I;AI;NI;AI;�$I;�.I;�=I;�RI;�oI;m�I;k�I;��I;Z6I;� G;?�A;�15;UW;�W�:¨�9X�غ!e��&�.�`��������a�8���H� Zb��j��O����K�,蒿��ɿ7��Ù$��F���d��{�      F�Q��K���;�Ù$��;
��޿�����w�o,���澝���(�D������I��3�G�����N��Ǩ�2��;�����9:���:�m!;��7;ڸB;}�G;	YI;K�I;��I;ؑI;�kI;�OI;4;I;�,I;3#I;�I;�I;�I;3#I;�,I;4;I;�OI;�kI;ؑI;��I;K�I;	YI;}�G;ڸB;��7;�m!;���:��9:;���2��Ǩ��N�����3�G��I������(�D��������o,���w�����޿�;
�Ù$���;��K�      Ù$��x � ��7���޿m���ǅ����F�{�
��~����z��$���ս$���P2+���ϼXPp����K�]��*�!��:,�;�7';��:;�C;+H;�|I;?�I;��I;��I;�fI;�KI;98I;V*I;D!I;I;GI;I;D!I;V*I;98I;�KI;�fI;��I;��I;?�I;�|I;+H;�C;��:;�7';,�;!��:�*�K�]����XPp���ϼP2+�$�����ս�$���z��~��{�
���F�ǅ��m����޿7�� ���x �      .���������㿆�ɿ���ǅ����P�b��:�׾�`��U�H����@��a�a�"���"D�Hɻ�!������U�:�~;�H-;G{=;ABE;ȄH;)�I;��I;��I;ւI;�`I;BGI;�4I;�'I;�I; I;oI; I;�I;�'I;�4I;BGI;�`I;ւI;��I;��I;)�I;ȄH;ABE;G{=;�H-;�~;�U�:�����!�Hɻ"D��"��a�a��@����U�H��`��:�׾b����P�ǅ�������ɿ��㿯���      ~�n�������,蒿��w���F�b��Ȱ�����Yb�+����ѽ�%��'D4����@X��ʨ��H���轺G��9ap�:�; 93;:P@;�uF;8�H;%�I;��I;��I;�yI;�YI;2BI;�0I;�$I;dI;�I;@I;�I;dI;�$I;�0I;2BI;�YI;�yI;��I;��I;%�I;8�H;�uF;:P@; 93;�;ap�:G��9�轺�H��ʨ�@X�����'D4��%����ѽ+���Yb����Ȱ�b����F���w�,蒿����n���      7�}���w�#f���K�o,�{�
�:�׾�����k���'�lz꽥I���;V�LM�*����iO��G�opE����a�:S� ;��$;˳8;q�B;�G;UJI;1�I;9�I;a�I;*pI;�RI;�<I;�,I;%!I;�I;9I;�I;9I;�I;%!I;�,I;�<I;�RI;*pI;a�I;9�I;1�I;UJI;�G;q�B;˳8;��$;S� ;a�:���opE��G��iO�*���LM��;V��I��lz���'���k����:�׾{�
�o,���K�#f���w�      E(��$�b��O������~���`���Yb���'��U�N$��S�m�5����ϼ0�����`�����غ�0�9b��: F;�F.;2{=;aE;�[H;A�I;��I;��I;�I;$fI;%KI;7I;%(I;�I;�I;�I;DI;�I;�I;�I;%(I;7I;%KI;$fI;�I;��I;��I;A�I;�[H;aE;2{=;�F.; F;b��:�0�9��غ`������0����ϼ5��S�m�N$���U���'��Yb��`���~�����O��b���$�      >�׾��Ҿž�j��������z�U�H�+��lz�N$��0v�!2+����9�� �5�-ɻ54�0�����:���:Mn!;*O6;(kA;��F;��H;��I;��I;�I;j|I;�[I;~CI;%1I;�#I;�I;jI;�I;�I;�I;jI;�I;�#I;%1I;~CI;�[I;j|I;�I;��I;��I;��H;��F;(kA;*O6;Mn!;���:���:0��54�-ɻ �5�9�����!2+�0v�N$��lz�+��U�H���z������j��ž��Ҿ      �T��f�����z� Zb�(�D��$�����ѽ�I��S�m�!2+��������K��ﻚ�p�=������9KR�:�.;��-;��<;iyD;uH;�lI;�I;��I;��I;�nI;�QI;�;I;!+I;�I;*I;NI;�I;�I;�I;NI;*I;�I;!+I;�;I;�QI;�nI;��I;��I;�I;�lI;uH;iyD;��<;��-;�.;KR�:���9=�����p��ﻍ�K������!2+�S�m��I����ѽ���$�(�D� Zb���z�f���      �L+� (���H�������ս�@���%���;V�5���������MS�������{F�ܺn8o�:�;��$;^7;J�A;��F;�H;��I;��I;��I;��I;uaI;�GI;-4I;A%I;HI;ZI;
I;�	I;	I;�	I;
I;ZI;HI;A%I;-4I;�GI;uaI;��I;��I;��I;��I;�H;��F;J�A;^7;��$;�;o�:ܺn8{F⺧������MS�������5���;V��%���@����ս����H��� (�      ��ս��ѽC�ƽ8����I��$���a�a�'D4�LM���ϼ9����K�����G��^g�x�o���:�@�:�X;��1;jk>;�
E;
/H;;pI;"�I;�I;��I; rI;�TI;>I;�,I;}I;�I;�I;�	I;.I;MI;.I;�	I;�I;�I;}I;�,I;>I;�TI; rI;��I;�I;"�I;;pI;
/H;�
E;jk>;��1;�X;�@�:��:x�o�^g��G�������K�9����ϼLM�'D4�a�a�$����I��8���C�ƽ��ѽ      r��ٷ��40v���a�3�G�P2+�"�����*���0�� �5��ﻧ��^g��ହ�g:]�:�;0H-;2f;;NC;)RG;�I;�I;@�I;�I;$�I;+bI;�HI;�4I;�%I;�I;PI;�
I;�I;eI;sI;eI;�I;�
I;PI;�I;�%I;�4I;�HI;+bI;$�I;�I;@�I;�I;�I;)RG;NC;2f;;0H-;�;]�:�g:�ହ^g������ �5�0��*������"��P2+�3�G���a�40v�ٷ��      ��7�e5���������ϼ�@X���iO����-ɻ��p�{F�x�o��g:^�:YF;�*;�9;��A;�tF;;�H;�I;��I;ȺI;d�I;�oI;SSI;n=I;9,I;�I;�I;I;pI;�I;�I;� I;�I;�I;pI;I;�I;�I;9,I;n=I;SSI;�oI;d�I;ȺI;��I;�I;;�H;�tF;��A;�9;�*;YF;^�:�g:x�o�{F⺚�p�-ɻ����iO�@X�����ϼ������e5�7�      @L�����R���`����N��XPp�"D�ʨ��G�`���54�=���ܺn8��:]�:YF;�(;��7;u�@;��E;mPH;5lI;��I;�I;��I;B|I;�]I;�EI;�2I;�#I;zI;�I;		I;(I;� I; �H;g�H; �H;� I;(I;		I;�I;zI;�#I;�2I;�EI;�]I;B|I;��I;�I;��I;5lI;mPH;��E;u�@;��7;�(;YF;]�:��:ܺn8=���54�`����G�ʨ�"D�XPp��N��`���R������      jO�%�K��o@�&�.�Ǩ����Hɻ�H��opE���غ0�����9o�:�@�:�;�*;��7;�O@;�[E;H;�HI;��I;��I;)�I;|�I;YgI;�MI;z9I;W)I;�I;�I;�
I;,I;'I;G�H;r�H;��H;r�H;G�H;'I;,I;�
I;�I;�I;W)I;z9I;�MI;YgI;|�I;)�I;��I;��I;�HI;H;�[E;�O@;��7;�*;�;�@�:o�:���90����غopE��H��Hɻ���Ǩ�&�.��o@�%�K�      9�ͻ�ɻ	���!e��2��K�]��!��轺����0�9���:KR�:�;�X;0H-;�9;u�@;�[E;��G;P4I;ճI;d�I;��I;l�I;�oI;�TI;q?I;M.I;� I;�I;YI;�I;�I;6�H;��H;,�H;��H;,�H;��H;6�H;�I;�I;YI;�I;� I;M.I;q?I;�TI;�oI;l�I;��I;d�I;ճI;P4I;��G;�[E;u�@;�9;0H-;�X;�;KR�:���:�0�9����轺�!�K�]�2��!e��	����ɻ      �����pj�X�غ;����*�����G��9a�:b��:���:�.;��$;��1;2f;;��A;��E;H;P4I;W�I;��I;m�I;��I;�uI;sZI;xDI;�2I;K$I;�I;�I;hI;�I;��H;s�H;7�H;��H;��H;��H;7�H;s�H;��H;�I;hI;�I;�I;K$I;�2I;xDI;sZI;�uI;��I;m�I;��I;W�I;P4I;H;��E;��A;2f;;��1;��$;�.;���:b��:a�:G��9�����*�;���X�غpj���      ��l8ۀ�8�Pu9¨�9��9:!��:�U�:ap�:S� ; F;Mn!;��-;^7;jk>;NC;�tF;mPH;�HI;ճI;��I;ϺI;әI;�yI;�^I;aHI;d6I;|'I;uI;�I;0
I;�I;>�H;��H;��H;�H;��H;��H;��H;�H;��H;��H;>�H;�I;0
I;�I;uI;|'I;d6I;aHI;�^I;�yI;әI;ϺI;��I;ճI;�HI;mPH;�tF;NC;jk>;^7;��-;Mn!; F;S� ;ap�:�U�:!��:��9:¨�9�Pu9ۀ�8      �m�:���:]I�:�W�:���:,�;�~;�;��$;�F.;*O6;��<;J�A;�
E;)RG;;�H;5lI;��I;d�I;m�I;әI;�zI;�`I;�JI;�8I;�)I;�I;�I;�I;9I; I;�H;��H;{�H; �H;�H;��H;�H; �H;{�H;��H;�H; I;9I;�I;�I;�I;�)I;�8I;�JI;�`I;�zI;әI;m�I;d�I;��I;5lI;;�H;)RG;�
E;J�A;��<;*O6;�F.;��$;�;�~;,�;���:�W�:]I�:���:      ��;��;=\;UW;�m!;�7';�H-; 93;˳8;2{=;(kA;iyD;��F;
/H;�I;�I;��I;��I;��I;��I;�yI;�`I;�KI;4:I;+I;EI;8I;I;MI;� I;��H;�H;w�H;~�H;�H;a�H;2�H;a�H;�H;~�H;w�H;�H;��H;� I;MI;I;8I;EI;+I;4:I;�KI;�`I;�yI;��I;��I;��I;��I;�I;�I;
/H;��F;iyD;(kA;2{=;˳8; 93;�H-;�7';�m!;UW;=\;��;      T�1;��1;�63;�15;��7;��:;G{=;:P@;q�B;aE;��F;uH;�H;;pI;�I;��I;�I;)�I;l�I;�uI;�^I;�JI;4:I;�+I; I;+I;�I;*I;�I;�H;��H;~�H;4�H;��H;z�H;��H;��H;��H;z�H;��H;4�H;~�H;��H;�H;�I;*I;�I;+I; I;�+I;4:I;�JI;�^I;�uI;l�I;)�I;�I;��I;�I;;pI;�H;uH;��F;aE;q�B;:P@;G{=;��:;��7;�15;�63;��1;      ��?;@;?�@;?�A;ڸB;�C;ABE;�uF;�G;�[H;��H;�lI;��I;"�I;@�I;ȺI;��I;|�I;�oI;sZI;aHI;�8I;+I; I;�I;sI;�I;I;s�H;��H;��H;;�H;d�H;��H;��H;f�H;=�H;f�H;��H;��H;d�H;;�H;��H;��H;s�H;I;�I;sI;�I; I;+I;�8I;aHI;sZI;�oI;|�I;��I;ȺI;@�I;"�I;��I;�lI;��H;�[H;�G;�uF;ABE;�C;ڸB;?�A;?�@;@;      uF;��F;�F;� G;}�G;+H;ȄH;8�H;UJI;A�I;��I;�I;��I;�I;�I;d�I;B|I;YgI;�TI;xDI;d6I;�)I;EI;+I;sI;�I;ZI;��H;��H;��H;6�H;I�H;��H;j�H;��H;$�H;��H;$�H;��H;j�H;��H;I�H;6�H;��H;��H;��H;ZI;�I;sI;+I;EI;�)I;d6I;xDI;�TI;YgI;B|I;d�I;�I;�I;��I;�I;��I;A�I;UJI;8�H;ȄH;+H;}�G;� G;�F;��F;      r�H;.I;WI;Z6I;	YI;�|I;)�I;%�I;1�I;��I;��I;��I;��I;��I;$�I;�oI;�]I;�MI;q?I;�2I;|'I;�I;8I;�I;�I;ZI;��H;2�H;��H;@�H;1�H;s�H;%�H;#�H;��H;�H;��H;�H;��H;#�H;%�H;s�H;1�H;@�H;��H;2�H;��H;ZI;�I;�I;8I;�I;|'I;�2I;q?I;�MI;�]I;�oI;$�I;��I;��I;��I;��I;��I;1�I;%�I;)�I;�|I;	YI;Z6I;WI;.I;      ��I;�I;��I;��I;K�I;?�I;��I;��I;9�I;��I;�I;��I;��I; rI;+bI;SSI;�EI;z9I;M.I;K$I;uI;�I;I;*I;I;��H;2�H;�H;L�H;-�H;d�H;��H;��H;
�H;b�H;�H;��H;�H;b�H;
�H;��H;��H;d�H;-�H;L�H;�H;2�H;��H;I;*I;I;�I;uI;K$I;M.I;z9I;�EI;SSI;+bI; rI;��I;��I;�I;��I;9�I;��I;��I;?�I;K�I;��I;��I;�I;      ��I;3�I;{�I;k�I;��I;��I;��I;��I;a�I;�I;j|I;�nI;uaI;�TI;�HI;n=I;�2I;W)I;� I;�I;�I;�I;MI;�I;s�H;��H;��H;L�H;8�H;a�H;��H;��H;��H;�H;��H;<�H;4�H;<�H;��H;�H;��H;��H;��H;a�H;8�H;L�H;��H;��H;s�H;�I;MI;�I;�I;�I;� I;W)I;�2I;n=I;�HI;�TI;uaI;�nI;j|I;�I;a�I;��I;��I;��I;��I;k�I;{�I;3�I;      ��I;ĝI;o�I;m�I;ؑI;��I;ւI;�yI;*pI;$fI;�[I;�QI;�GI;>I;�4I;9,I;�#I;�I;�I;�I;0
I;9I;� I;�H;��H;��H;@�H;-�H;a�H;��H;��H;��H;��H;!�H;��H;��H;c�H;��H;��H;!�H;��H;��H;��H;��H;a�H;-�H;@�H;��H;��H;�H;� I;9I;0
I;�I;�I;�I;�#I;9,I;�4I;>I;�GI;�QI;�[I;$fI;*pI;�yI;ւI;��I;ؑI;m�I;o�I;ĝI;      �uI;�tI;�rI;�oI;�kI;�fI;�`I;�YI;�RI;%KI;~CI;�;I;-4I;�,I;�%I;�I;zI;�I;YI;hI;�I; I;��H;��H;��H;6�H;1�H;d�H;��H;��H;��H;��H;��H;c�H;�H;��H;��H;��H;�H;c�H;��H;��H;��H;��H;��H;d�H;1�H;6�H;��H;��H;��H; I;�I;hI;YI;�I;zI;�I;�%I;�,I;-4I;�;I;~CI;%KI;�RI;�YI;�`I;�fI;�kI;�oI;�rI;�tI;      �VI;NVI;�TI;�RI;�OI;�KI;BGI;2BI;�<I;7I;%1I;!+I;A%I;}I;�I;�I;�I;�
I;�I;�I;>�H;�H;�H;~�H;;�H;I�H;s�H;��H;��H;��H;��H;��H;J�H;��H;��H;J�H;P�H;J�H;��H;��H;J�H;��H;��H;��H;��H;��H;s�H;I�H;;�H;~�H;�H;�H;>�H;�I;�I;�
I;�I;�I;�I;}I;A%I;!+I;%1I;7I;�<I;2BI;BGI;�KI;�OI;�RI;�TI;NVI;      �@I;�@I;^?I;�=I;4;I;98I;�4I;�0I;�,I;%(I;�#I;�I;HI;�I;PI;I;		I;,I;�I;��H;��H;��H;w�H;4�H;d�H;��H;%�H;��H;��H;��H;��H;J�H;��H;d�H;�H;��H;��H;��H;�H;d�H;��H;J�H;��H;��H;��H;��H;%�H;��H;d�H;4�H;w�H;��H;��H;��H;�I;,I;		I;I;PI;�I;HI;�I;�#I;%(I;�,I;�0I;�4I;98I;4;I;�=I;^?I;�@I;      1I;�0I;0I;�.I;�,I;V*I;�'I;�$I;%!I;�I;�I;*I;ZI;�I;�
I;pI;(I;'I;6�H;s�H;��H;{�H;~�H;��H;��H;j�H;#�H;
�H;�H;!�H;c�H;��H;d�H;��H;��H;��H;��H;��H;��H;��H;d�H;��H;c�H;!�H;�H;
�H;#�H;j�H;��H;��H;~�H;{�H;��H;s�H;6�H;'I;(I;pI;�
I;�I;ZI;*I;�I;�I;%!I;�$I;�'I;V*I;�,I;�.I;0I;�0I;      �&I;�&I;&I;�$I;3#I;D!I;�I;dI;�I;�I;jI;NI;
I;�	I;�I;�I;� I;G�H;��H;7�H;�H; �H;�H;z�H;��H;��H;��H;b�H;��H;��H;�H;��H;�H;��H;��H;d�H;[�H;d�H;��H;��H;�H;��H;�H;��H;��H;b�H;��H;��H;��H;z�H;�H; �H;�H;7�H;��H;G�H;� I;�I;�I;�	I;
I;NI;jI;�I;�I;dI;�I;D!I;3#I;�$I;&I;�&I;      � I;� I;, I;AI;�I;I; I;�I;9I;�I;�I;�I;�	I;.I;eI;�I; �H;r�H;,�H;��H;��H;�H;a�H;��H;f�H;$�H;�H;�H;<�H;��H;��H;J�H;��H;��H;d�H;2�H;/�H;2�H;d�H;��H;��H;J�H;��H;��H;<�H;�H;�H;$�H;f�H;��H;a�H;�H;��H;��H;,�H;r�H; �H;�I;eI;.I;�	I;�I;�I;�I;9I;�I; I;I;�I;AI;, I;� I;      I;�I;LI;NI;�I;GI;oI;@I;�I;DI;�I;�I;	I;MI;sI;� I;g�H;��H;��H;��H;��H;��H;2�H;��H;=�H;��H;��H;��H;4�H;c�H;��H;P�H;��H;��H;[�H;/�H;�H;/�H;[�H;��H;��H;P�H;��H;c�H;4�H;��H;��H;��H;=�H;��H;2�H;��H;��H;��H;��H;��H;g�H;� I;sI;MI;	I;�I;�I;DI;�I;@I;oI;GI;�I;NI;LI;�I;      � I;� I;, I;AI;�I;I; I;�I;9I;�I;�I;�I;�	I;.I;eI;�I; �H;r�H;,�H;��H;��H;�H;a�H;��H;f�H;$�H;�H;�H;<�H;��H;��H;J�H;��H;��H;d�H;2�H;/�H;2�H;d�H;��H;��H;J�H;��H;��H;<�H;�H;�H;$�H;f�H;��H;a�H;�H;��H;��H;,�H;r�H; �H;�I;eI;.I;�	I;�I;�I;�I;9I;�I; I;I;�I;AI;, I;� I;      �&I;�&I;&I;�$I;3#I;D!I;�I;dI;�I;�I;jI;NI;
I;�	I;�I;�I;� I;G�H;��H;7�H;�H; �H;�H;z�H;��H;��H;��H;b�H;��H;��H;�H;��H;�H;��H;��H;d�H;[�H;d�H;��H;��H;�H;��H;�H;��H;��H;b�H;��H;��H;��H;z�H;�H; �H;�H;7�H;��H;G�H;� I;�I;�I;�	I;
I;NI;jI;�I;�I;dI;�I;D!I;3#I;�$I;&I;�&I;      1I;�0I;0I;�.I;�,I;V*I;�'I;�$I;%!I;�I;�I;*I;ZI;�I;�
I;pI;(I;'I;6�H;s�H;��H;{�H;~�H;��H;��H;j�H;#�H;
�H;�H;!�H;c�H;��H;d�H;��H;��H;��H;��H;��H;��H;��H;d�H;��H;c�H;!�H;�H;
�H;#�H;j�H;��H;��H;~�H;{�H;��H;s�H;6�H;'I;(I;pI;�
I;�I;ZI;*I;�I;�I;%!I;�$I;�'I;V*I;�,I;�.I;0I;�0I;      �@I;�@I;^?I;�=I;4;I;98I;�4I;�0I;�,I;%(I;�#I;�I;HI;�I;PI;I;		I;,I;�I;��H;��H;��H;w�H;4�H;d�H;��H;%�H;��H;��H;��H;��H;J�H;��H;d�H;�H;��H;��H;��H;�H;d�H;��H;J�H;��H;��H;��H;��H;%�H;��H;d�H;4�H;w�H;��H;��H;��H;�I;,I;		I;I;PI;�I;HI;�I;�#I;%(I;�,I;�0I;�4I;98I;4;I;�=I;^?I;�@I;      �VI;NVI;�TI;�RI;�OI;�KI;BGI;2BI;�<I;7I;%1I;!+I;A%I;}I;�I;�I;�I;�
I;�I;�I;>�H;�H;�H;~�H;;�H;I�H;s�H;��H;��H;��H;��H;��H;J�H;��H;��H;J�H;P�H;J�H;��H;��H;J�H;��H;��H;��H;��H;��H;s�H;I�H;;�H;~�H;�H;�H;>�H;�I;�I;�
I;�I;�I;�I;}I;A%I;!+I;%1I;7I;�<I;2BI;BGI;�KI;�OI;�RI;�TI;NVI;      �uI;�tI;�rI;�oI;�kI;�fI;�`I;�YI;�RI;%KI;~CI;�;I;-4I;�,I;�%I;�I;zI;�I;YI;hI;�I; I;��H;��H;��H;6�H;1�H;d�H;��H;��H;��H;��H;��H;c�H;�H;��H;��H;��H;�H;c�H;��H;��H;��H;��H;��H;d�H;1�H;6�H;��H;��H;��H; I;�I;hI;YI;�I;zI;�I;�%I;�,I;-4I;�;I;~CI;%KI;�RI;�YI;�`I;�fI;�kI;�oI;�rI;�tI;      ��I;ĝI;o�I;m�I;ؑI;��I;ւI;�yI;*pI;$fI;�[I;�QI;�GI;>I;�4I;9,I;�#I;�I;�I;�I;0
I;9I;� I;�H;��H;��H;@�H;-�H;a�H;��H;��H;��H;��H;!�H;��H;��H;c�H;��H;��H;!�H;��H;��H;��H;��H;a�H;-�H;@�H;��H;��H;�H;� I;9I;0
I;�I;�I;�I;�#I;9,I;�4I;>I;�GI;�QI;�[I;$fI;*pI;�yI;ւI;��I;ؑI;m�I;o�I;ĝI;      ��I;3�I;{�I;k�I;��I;��I;��I;��I;a�I;�I;j|I;�nI;uaI;�TI;�HI;n=I;�2I;W)I;� I;�I;�I;�I;MI;�I;s�H;��H;��H;L�H;8�H;a�H;��H;��H;��H;�H;��H;<�H;4�H;<�H;��H;�H;��H;��H;��H;a�H;8�H;L�H;��H;��H;s�H;�I;MI;�I;�I;�I;� I;W)I;�2I;n=I;�HI;�TI;uaI;�nI;j|I;�I;a�I;��I;��I;��I;��I;k�I;{�I;3�I;      ��I;�I;��I;��I;K�I;?�I;��I;��I;9�I;��I;�I;��I;��I; rI;+bI;SSI;�EI;z9I;M.I;K$I;uI;�I;I;*I;I;��H;2�H;�H;L�H;-�H;d�H;��H;��H;
�H;b�H;�H;��H;�H;b�H;
�H;��H;��H;d�H;-�H;L�H;�H;2�H;��H;I;*I;I;�I;uI;K$I;M.I;z9I;�EI;SSI;+bI; rI;��I;��I;�I;��I;9�I;��I;��I;?�I;K�I;��I;��I;�I;      r�H;.I;WI;Z6I;	YI;�|I;)�I;%�I;1�I;��I;��I;��I;��I;��I;$�I;�oI;�]I;�MI;q?I;�2I;|'I;�I;8I;�I;�I;ZI;��H;2�H;��H;@�H;1�H;s�H;%�H;#�H;��H;�H;��H;�H;��H;#�H;%�H;s�H;1�H;@�H;��H;2�H;��H;ZI;�I;�I;8I;�I;|'I;�2I;q?I;�MI;�]I;�oI;$�I;��I;��I;��I;��I;��I;1�I;%�I;)�I;�|I;	YI;Z6I;WI;.I;      uF;��F;�F;� G;}�G;+H;ȄH;8�H;UJI;A�I;��I;�I;��I;�I;�I;d�I;B|I;YgI;�TI;xDI;d6I;�)I;EI;+I;sI;�I;ZI;��H;��H;��H;6�H;I�H;��H;j�H;��H;$�H;��H;$�H;��H;j�H;��H;I�H;6�H;��H;��H;��H;ZI;�I;sI;+I;EI;�)I;d6I;xDI;�TI;YgI;B|I;d�I;�I;�I;��I;�I;��I;A�I;UJI;8�H;ȄH;+H;}�G;� G;�F;��F;      ��?;@;?�@;?�A;ڸB;�C;ABE;�uF;�G;�[H;��H;�lI;��I;"�I;@�I;ȺI;��I;|�I;�oI;sZI;aHI;�8I;+I; I;�I;sI;�I;I;s�H;��H;��H;;�H;d�H;��H;��H;f�H;=�H;f�H;��H;��H;d�H;;�H;��H;��H;s�H;I;�I;sI;�I; I;+I;�8I;aHI;sZI;�oI;|�I;��I;ȺI;@�I;"�I;��I;�lI;��H;�[H;�G;�uF;ABE;�C;ڸB;?�A;?�@;@;      T�1;��1;�63;�15;��7;��:;G{=;:P@;q�B;aE;��F;uH;�H;;pI;�I;��I;�I;)�I;l�I;�uI;�^I;�JI;4:I;�+I; I;+I;�I;*I;�I;�H;��H;~�H;4�H;��H;z�H;��H;��H;��H;z�H;��H;4�H;~�H;��H;�H;�I;*I;�I;+I; I;�+I;4:I;�JI;�^I;�uI;l�I;)�I;�I;��I;�I;;pI;�H;uH;��F;aE;q�B;:P@;G{=;��:;��7;�15;�63;��1;      ��;��;=\;UW;�m!;�7';�H-; 93;˳8;2{=;(kA;iyD;��F;
/H;�I;�I;��I;��I;��I;��I;�yI;�`I;�KI;4:I;+I;EI;8I;I;MI;� I;��H;�H;w�H;~�H;�H;a�H;2�H;a�H;�H;~�H;w�H;�H;��H;� I;MI;I;8I;EI;+I;4:I;�KI;�`I;�yI;��I;��I;��I;��I;�I;�I;
/H;��F;iyD;(kA;2{=;˳8; 93;�H-;�7';�m!;UW;=\;��;      �m�:���:]I�:�W�:���:,�;�~;�;��$;�F.;*O6;��<;J�A;�
E;)RG;;�H;5lI;��I;d�I;m�I;әI;�zI;�`I;�JI;�8I;�)I;�I;�I;�I;9I; I;�H;��H;{�H; �H;�H;��H;�H; �H;{�H;��H;�H; I;9I;�I;�I;�I;�)I;�8I;�JI;�`I;�zI;әI;m�I;d�I;��I;5lI;;�H;)RG;�
E;J�A;��<;*O6;�F.;��$;�;�~;,�;���:�W�:]I�:���:      ��l8ۀ�8�Pu9¨�9��9:!��:�U�:ap�:S� ; F;Mn!;��-;^7;jk>;NC;�tF;mPH;�HI;ճI;��I;ϺI;әI;�yI;�^I;aHI;d6I;|'I;uI;�I;0
I;�I;>�H;��H;��H;�H;��H;��H;��H;�H;��H;��H;>�H;�I;0
I;�I;uI;|'I;d6I;aHI;�^I;�yI;әI;ϺI;��I;ճI;�HI;mPH;�tF;NC;jk>;^7;��-;Mn!; F;S� ;ap�:�U�:!��:��9:¨�9�Pu9ۀ�8      �����pj�X�غ;����*�����G��9a�:b��:���:�.;��$;��1;2f;;��A;��E;H;P4I;W�I;��I;m�I;��I;�uI;sZI;xDI;�2I;K$I;�I;�I;hI;�I;��H;s�H;7�H;��H;��H;��H;7�H;s�H;��H;�I;hI;�I;�I;K$I;�2I;xDI;sZI;�uI;��I;m�I;��I;W�I;P4I;H;��E;��A;2f;;��1;��$;�.;���:b��:a�:G��9�����*�;���X�غpj���      9�ͻ�ɻ	���!e��2��K�]��!��轺����0�9���:KR�:�;�X;0H-;�9;u�@;�[E;��G;P4I;ճI;d�I;��I;l�I;�oI;�TI;q?I;M.I;� I;�I;YI;�I;�I;6�H;��H;,�H;��H;,�H;��H;6�H;�I;�I;YI;�I;� I;M.I;q?I;�TI;�oI;l�I;��I;d�I;ճI;P4I;��G;�[E;u�@;�9;0H-;�X;�;KR�:���:�0�9����轺�!�K�]�2��!e��	����ɻ      jO�%�K��o@�&�.�Ǩ����Hɻ�H��opE���غ0�����9o�:�@�:�;�*;��7;�O@;�[E;H;�HI;��I;��I;)�I;|�I;YgI;�MI;z9I;W)I;�I;�I;�
I;,I;'I;G�H;r�H;��H;r�H;G�H;'I;,I;�
I;�I;�I;W)I;z9I;�MI;YgI;|�I;)�I;��I;��I;�HI;H;�[E;�O@;��7;�*;�;�@�:o�:���90����غopE��H��Hɻ���Ǩ�&�.��o@�%�K�      @L�����R���`����N��XPp�"D�ʨ��G�`���54�=���ܺn8��:]�:YF;�(;��7;u�@;��E;mPH;5lI;��I;�I;��I;B|I;�]I;�EI;�2I;�#I;zI;�I;		I;(I;� I; �H;g�H; �H;� I;(I;		I;�I;zI;�#I;�2I;�EI;�]I;B|I;��I;�I;��I;5lI;mPH;��E;u�@;��7;�(;YF;]�:��:ܺn8=���54�`����G�ʨ�"D�XPp��N��`���R������      ��7�e5���������ϼ�@X���iO����-ɻ��p�{F�x�o��g:^�:YF;�*;�9;��A;�tF;;�H;�I;��I;ȺI;d�I;�oI;SSI;n=I;9,I;�I;�I;I;pI;�I;�I;� I;�I;�I;pI;I;�I;�I;9,I;n=I;SSI;�oI;d�I;ȺI;��I;�I;;�H;�tF;��A;�9;�*;YF;^�:�g:x�o�{F⺚�p�-ɻ����iO�@X�����ϼ������e5�7�      r��ٷ��40v���a�3�G�P2+�"�����*���0�� �5��ﻧ��^g��ହ�g:]�:�;0H-;2f;;NC;)RG;�I;�I;@�I;�I;$�I;+bI;�HI;�4I;�%I;�I;PI;�
I;�I;eI;sI;eI;�I;�
I;PI;�I;�%I;�4I;�HI;+bI;$�I;�I;@�I;�I;�I;)RG;NC;2f;;0H-;�;]�:�g:�ହ^g������ �5�0��*������"��P2+�3�G���a�40v�ٷ��      ��ս��ѽC�ƽ8����I��$���a�a�'D4�LM���ϼ9����K�����G��^g�x�o���:�@�:�X;��1;jk>;�
E;
/H;;pI;"�I;�I;��I; rI;�TI;>I;�,I;}I;�I;�I;�	I;.I;MI;.I;�	I;�I;�I;}I;�,I;>I;�TI; rI;��I;�I;"�I;;pI;
/H;�
E;jk>;��1;�X;�@�:��:x�o�^g��G�������K�9����ϼLM�'D4�a�a�$����I��8���C�ƽ��ѽ      �L+� (���H�������ս�@���%���;V�5���������MS�������{F�ܺn8o�:�;��$;^7;J�A;��F;�H;��I;��I;��I;��I;uaI;�GI;-4I;A%I;HI;ZI;
I;�	I;	I;�	I;
I;ZI;HI;A%I;-4I;�GI;uaI;��I;��I;��I;��I;�H;��F;J�A;^7;��$;�;o�:ܺn8{F⺧������MS�������5���;V��%���@����ս����H��� (�      �T��f�����z� Zb�(�D��$�����ѽ�I��S�m�!2+��������K��ﻚ�p�=������9KR�:�.;��-;��<;iyD;uH;�lI;�I;��I;��I;�nI;�QI;�;I;!+I;�I;*I;NI;�I;�I;�I;NI;*I;�I;!+I;�;I;�QI;�nI;��I;��I;�I;�lI;uH;iyD;��<;��-;�.;KR�:���9=�����p��ﻍ�K������!2+�S�m��I����ѽ���$�(�D� Zb���z�f���      >�׾��Ҿž�j��������z�U�H�+��lz�N$��0v�!2+����9�� �5�-ɻ54�0�����:���:Mn!;*O6;(kA;��F;��H;��I;��I;�I;j|I;�[I;~CI;%1I;�#I;�I;jI;�I;�I;�I;jI;�I;�#I;%1I;~CI;�[I;j|I;�I;��I;��I;��H;��F;(kA;*O6;Mn!;���:���:0��54�-ɻ �5�9�����!2+�0v�N$��lz�+��U�H���z������j��ž��Ҿ      E(��$�b��O������~���`���Yb���'��U�N$��S�m�5����ϼ0�����`�����غ�0�9b��: F;�F.;2{=;aE;�[H;A�I;��I;��I;�I;$fI;%KI;7I;%(I;�I;�I;�I;DI;�I;�I;�I;%(I;7I;%KI;$fI;�I;��I;��I;A�I;�[H;aE;2{=;�F.; F;b��:�0�9��غ`������0����ϼ5��S�m�N$���U���'��Yb��`���~�����O��b���$�      7�}���w�#f���K�o,�{�
�:�׾�����k���'�lz꽥I���;V�LM�*����iO��G�opE����a�:S� ;��$;˳8;q�B;�G;UJI;1�I;9�I;a�I;*pI;�RI;�<I;�,I;%!I;�I;9I;�I;9I;�I;%!I;�,I;�<I;�RI;*pI;a�I;9�I;1�I;UJI;�G;q�B;˳8;��$;S� ;a�:���opE��G��iO�*���LM��;V��I��lz���'���k����:�׾{�
�o,���K�#f���w�      ~�n�������,蒿��w���F�b��Ȱ�����Yb�+����ѽ�%��'D4����@X��ʨ��H���轺G��9ap�:�; 93;:P@;�uF;8�H;%�I;��I;��I;�yI;�YI;2BI;�0I;�$I;dI;�I;@I;�I;dI;�$I;�0I;2BI;�YI;�yI;��I;��I;%�I;8�H;�uF;:P@; 93;�;ap�:G��9�轺�H��ʨ�@X�����'D4��%����ѽ+���Yb����Ȱ�b����F���w�,蒿����n���      .���������㿆�ɿ���ǅ����P�b��:�׾�`��U�H����@��a�a�"���"D�Hɻ�!������U�:�~;�H-;G{=;ABE;ȄH;)�I;��I;��I;ւI;�`I;BGI;�4I;�'I;�I; I;oI; I;�I;�'I;�4I;BGI;�`I;ւI;��I;��I;)�I;ȄH;ABE;G{=;�H-;�~;�U�:�����!�Hɻ"D��"��a�a��@����U�H��`��:�׾b����P�ǅ�������ɿ��㿯���      Ù$��x � ��7���޿m���ǅ����F�{�
��~����z��$���ս$���P2+���ϼXPp����K�]��*�!��:,�;�7';��:;�C;+H;�|I;?�I;��I;��I;�fI;�KI;98I;V*I;D!I;I;GI;I;D!I;V*I;98I;�KI;�fI;��I;��I;?�I;�|I;+H;�C;��:;�7';,�;!��:�*�K�]����XPp���ϼP2+�$�����ս�$���z��~��{�
���F�ǅ��m����޿7�� ���x �      F�Q��K���;�Ù$��;
��޿�����w�o,���澝���(�D������I��3�G�����N��Ǩ�2��;�����9:���:�m!;��7;ڸB;}�G;	YI;K�I;��I;ؑI;�kI;�OI;4;I;�,I;3#I;�I;�I;�I;3#I;�,I;4;I;�OI;�kI;ؑI;��I;K�I;	YI;}�G;ڸB;��7;�m!;���:��9:;���2��Ǩ��N�����3�G��I������(�D��������o,���w�����޿�;
�Ù$���;��K�      Q����{���d��F�Ù$�7����ɿ,蒿��K�O���j�� Zb�H�8�����a����`���&�.�!e��X�غ¨�9�W�:UW;�15;?�A;� G;Z6I;��I;k�I;m�I;�oI;�RI;�=I;�.I;�$I;AI;NI;AI;�$I;�.I;�=I;�RI;�oI;m�I;k�I;��I;Z6I;� G;?�A;�15;UW;�W�:¨�9X�غ!e��&�.�`��������a�8���H� Zb��j��O����K�,蒿��ɿ7��Ù$��F���d��{�      ���� P�������d���;� ����㿰���#f�b��ž��z���C�ƽ40v�e5�R����o@�	���pj��Pu9]I�:=\;�63;?�@;�F;WI;��I;{�I;o�I;�rI;�TI;^?I;0I;&I;, I;LI;, I;&I;0I;^?I;�TI;�rI;o�I;{�I;��I;WI;�F;?�@;�63;=\;]I�:�Pu9pj�	����o@�R���e5�40v�C�ƽ����z�žb��#f�������� ����;���d���� P��      �,��^�� P���{��K��x �����n�����w��$���Ҿf��� (���ѽٷ��7����%�K��ɻ��ۀ�8���:��;��1;@;��F;.I;�I;3�I;ĝI;�tI;NVI;�@I;�0I;�&I;� I;�I;� I;�&I;�0I;�@I;NVI;�tI;ĝI;3�I;�I;.I;��F;@;��1;��;���:ۀ�8���ɻ%�K����7�ٷ����ѽ (�f�����Ҿ�$���w�n��������x ��K��{� P��^��      ݶ��O���ά��(�_���7�w�}߿���~,b��V�*l¾Fx�c.���Ž��t�6�����*�?��N�����sx9���:��;��2;T?@;�eF;C�H;��I;��I;8{I;�ZI;�BI;"1I;�$I;�I;�I;NI;�I;�I;�$I;"1I;�BI;�ZI;8{I;��I;��I;C�H;�eF;T?@;��2;��;���:�sx9���N��*�?����6����t���Žc.�Fx�*l¾�V�~,b����}߿w���7�(�_�ά��O���      O���A���}��+Y��3�����$ڿ"����\����(���s��3�9�����p�p�p���<<����f������9{��:�;V$3;ho@;yF;��H;�I;�I;�zI;rZI;yBI;�0I;s$I;EI;tI; I;tI;EI;s$I;�0I;yBI;rZI;�zI;�I;�I;��H;yF;ho@;V$3;�;{��:���9f�������<<�p��p���p�9����3��s�(�������\�"���$ڿ����3��+Y�}�A���      ά��}�8tf��lG�Ң%��p�*�ʿV����>M����S����d�ɤ�̷�9�d��
��I��@�1����� ��ݤ�9���:M;�T4;��@;�F;@�H; �I;ۙI;�xI;�XI;aAI;�/I;�#I;�I;�I;�I;�I;�I;�#I;�/I;aAI;�XI;�xI;ۙI; �I;@�H;�F;��@;�T4;M;���:ݤ�9 ������@�1��I���
�9�d�̷�ɤ��d�S�������>M�V���*�ʿ�p�Ң%��lG�8tf�}�      (�_��+Y��lG�f.�w���꿭���J䂿��5���󾋰��M�N�W��V��-�Q�*�������;i!��g��-󳺍:��:�;e06;��A;tG;I;Z�I;��I;�uI;pVI;�?I;�.I;�"I;�I;'I;�I;'I;�I;�"I;�.I;�?I;pVI;�uI;��I;Z�I;I;tG;��A;e06;�;��:�:-��g��;i!�����*���-�Q�V��W��M�N���������5�J䂿�������w�f.��lG��+Y�      ��7��3�Ң%�w��<����ſ�����\�9����Ͼ����`�3����z����9�z�ἷ���z��8}�ht�F�^:�)�:΢#;��8;��B;ArG;�$I;јI;�I;#qI;6SI;=I;�,I;0!I;nI;I;�I;I;nI;0!I;�,I;=I;6SI;#qI;�I;јI;�$I;ArG;��B;��8;΢#;�)�:F�^:ht��8}��z����z�Ἁ�9��z����`�3�������Ͼ9����\������ſ�<��w�Ң%��3�      w�����p������ſ!��{Ps���1�-r���d���d�}I�҈Ž��}�l*�gC��W�^�RC�g�D�,N๩��:��;�);-6;;JD;e�G;kGI;ΜI;ǎI;�kI;OI;�9I;3*I;8I;�I;�I;KI;�I;�I;8I;3*I;�9I;OI;�kI;ǎI;ΜI;kGI;e�G;JD;-6;;�);��;���:,N�g�D�RC�W�^�gC��l*���}�҈Ž}I��d��d��-r����1�{Ps�!����ſ��꿀p����      }߿�$ڿ*�ʿ�������{Ps�MX:����#l¾�ǆ���7����<5��$�Q�����t��85���������8�Ǽ:��;��.;��=;�DE;�XH;�gI;G�I;ڇI;FeI;@JI;D6I;a'I;�I;I;�I;�I;�I;I;�I;a'I;D6I;@JI;FeI;ڇI;G�I;�gI;�XH;�DE;��=;��.;��;�Ǽ:��8������85��t�����$�Q�<5�������7��ǆ�#l¾���MX:�{Ps��������*�ʿ�$ڿ      ���"��V���J䂿��\���1�����J˾睒�C�N�y��L������c�'���Ҽ �|��z�lo�� z��%�&:�N�:˧;�V4;�@;GfF;��H;.�I;A�I;UI;<^I;�DI;%2I;<$I;bI;�I;I;�I;I;�I;bI;<$I;%2I;�DI;<^I;UI;A�I;.�I;��H;GfF;�@;�V4;˧;�N�:%�&: z��lo���z� �|���Ҽc�'����L���y��C�N�睒��J˾�����1���\�J䂿V���"��      ~,b���\��>M���5�9��-r��#l¾睒�"&W��3�<Sؽ�z��fG�����I���?��̻{�-����J��:��;ο&;B{9;�C;�cG;sI;\�I;r�I;quI;�VI;O?I;�-I;� I;�I;yI;�I;�I;�I;yI;�I;� I;�-I;O?I;�VI;quI;r�I;\�I;sI;�cG;�C;B{9;ο&;��;J��:���{�-��̻�?��I�����fG��z��<Sؽ�3�"&W�睒�#l¾-r��9����5��>M���\�      �V������������Ͼ�d���ǆ�C�N��3��c�[����\�@��EC��O�o�Ъ	�t숻1�H��9I��:�g;o�/;\�=;aE;2H;�VI;؜I;�I;�jI;�NI;F9I;)I;=I;�I;I;�I;�
I;�I;I;�I;=I;)I;F9I;�NI;�jI;�I;؜I;�VI;2H;aE;\�=;o�/;�g;I��:H��91�t숻Ъ	�O�o�EC��@����\�[���cཱ3�C�N��ǆ��d����Ͼ���������      *l¾(��S������������d���7�y��<Sؽ[�� �d�P*�kּI\����'�����S������
�:�Y;�#;Y<7;M�A;2�F;{�H;��I;�I;րI;	`I;�FI;3I;B$I;�I;�I;vI;h	I;iI;h	I;vI;�I;�I;B$I;3I;�FI;	`I;րI;�I;��I;{�H;2�F;M�A;Y<7;�#;�Y;�
�:�����S������'�I\��kּP*� �d�[��<Sؽy����7��d���������S���(��      Fx��s��d�M�N�`�3�}I����L����z����\�P*�'�ݼe���k<<���ڻ��V��gt�p�&:���:[B;�;/;nC=;��D;��G;8I;�I;ÓI;3sI;IUI;}>I;�,I;�I;�I;xI;�	I;I;.I;I;�	I;xI;�I;�I;�,I;}>I;IUI;3sI;ÓI;�I;8I;��G;��D;nC=;�;/;[B;���:p�&:�gt���V���ڻk<<�e���'�ݼP*���\��z��L������}I�`�3�M�N��d��s�      c.��3�ɤ�W����҈Ž<5�����fG�@��kּe���:yC�?�X7}�񮼺C�x9���:%	;N�&;�:8;��A;��F;ϸH;WxI;��I;�I;PeI;�JI;m6I;�&I;�I;�I;uI;/I;�I;�I;�I;/I;uI;�I;�I;�&I;m6I;�JI;PeI;�I;��I;WxI;ϸH;��F;��A;�:8;N�&;%	;���:C�x9񮼺X7}�?�:yC�e���kּ@��fG����<5��҈Ž��W��ɤ��3�      ��Ž9���̷�V���z����}�$�Q�c�'����EC��I\��k<<�?��n�� ��xU�b��:Y��:,�;�&3;��>;�E;�H;};I;�I;ÔI;�uI;�WI;�@I;�.I;� I;�I;I;oI;I;<I;�I;<I;I;oI;I;�I;� I;�.I;�@I;�WI;�uI;ÔI;�I;};I;�H;�E;��>;�&3;,�;Y��:b��:xU� ���n��?�k<<�I\��EC�����c�'�$�Q���}��z��V��̷�9���      ��t���p�9�d�-�Q���9�l*������Ҽ�I��O�o���'���ڻX7}� ��wH��߄:�k�:��;�.;5<;�nC;^6G;��H;�I;��I;�I;;eI;^KI;7I;�&I;�I;�I;h
I;cI;�I;��H;l�H;��H;�I;cI;h
I;�I;�I;�&I;7I;^KI;;eI;�I;��I;�I;��H;^6G;�nC;5<;�.;��;�k�:�߄:wH� ��X7}���ڻ��'�O�o��I����Ҽ���l*���9�-�Q�9�d���p�      6��p��
�*���z��gC���t�� �|��?�Ъ	������V�񮼺xU��߄:��:�g;6�+;�9;��A;�eF;w�H;�^I;��I;��I; rI;�UI;�?I;�-I; I;uI;'I;�I;�I;i�H;��H;�H;��H;i�H;�I;�I;'I;uI; I;�-I;�?I;�UI; rI;��I;��I;�^I;w�H;�eF;��A;�9;6�+;�g;��:�߄:xU�񮼺��V����Ъ	��?� �|��t��gC��z��*����
�p�      ���p���I���������W�^�85��z��̻t숻�S��gt�C�x9b��:�k�:�g;y�*;�8;�@;��E;W'H;�7I;ߒI;2�I;o}I;�_I;�GI;�4I;y%I;�I;QI;	I;�I;��H;�H;i�H;��H;i�H;�H;��H;�I;	I;QI;�I;y%I;�4I;�GI;�_I;o}I;2�I;ߒI;�7I;W'H;��E;�@;�8;y�*;�g;�k�:b��:C�x9�gt��S�t숻�̻�z�85�W�^���������I��p��      *�?��<<�@�1�;i!��z�RC����lo��{�-�1򳺵���p�&:���:Y��:��;6�+;�8;W�@;]E;��G;eI;	�I;l�I;P�I;�hI;TOI;";I;�*I;�I;�I;nI;EI;� I;��H;��H;d�H;��H;d�H;��H;��H;� I;EI;nI;�I;�I;�*I;";I;TOI;�hI;P�I;l�I;	�I;eI;��G;]E;W�@;�8;6�+;��;Y��:���:p�&:����1�{�-�lo�����RC��z�;i!�@�1��<<�      �N����������g���8}�g�D���� z�����H��9�
�:���:%	;,�;�.;�9;�@;]E;��G;\I;�~I;#�I;g�I;�oI;�UI;�@I;�/I;�!I;�I;I;I;�I;��H;s�H;��H;r�H;��H;r�H;��H;s�H;��H;�I;I;I;�I;�!I;�/I;�@I;�UI;�oI;g�I;#�I;�~I;\I;��G;]E;�@;�9;�.;,�;%	;���:�
�:H��9��� z�����g�D��8}��g���������      ��f��� ��-�ht�,N���8%�&:J��:I��:�Y;[B;N�&;�&3;5<;��A;��E;��G;\I;v{I;ߛI;��I;�tI;�ZI;*EI;�3I;D%I;�I;bI;�I;I;O�H;��H;I�H;��H;��H;0�H;��H;��H;I�H;��H;O�H;I;�I;bI;�I;D%I;�3I;*EI;�ZI;�tI;��I;ߛI;v{I;\I;��G;��E;��A;5<;�&3;N�&;[B;�Y;I��:J��:%�&:��8,N�ht�-� ��f���      �sx9���9ݤ�9�:F�^:���:�Ǽ:�N�:��;�g;�#;�;/;�:8;��>;�nC;�eF;W'H;eI;�~I;ߛI;ːI;wI;�]I;QHI;�6I;(I;"I;�I;�
I;\I;b�H;]�H;h�H;L�H;��H;��H;��H;��H;��H;L�H;h�H;]�H;b�H;\I;�
I;�I;"I;(I;�6I;QHI;�]I;wI;ːI;ߛI;�~I;eI;W'H;�eF;�nC;��>;�:8;�;/;�#;�g;��;�N�:�Ǽ:���:F�^:�:ݤ�9���9      ���:{��:���:��:�)�:��;��;˧;ο&;o�/;Y<7;nC=;��A;�E;^6G;w�H;�7I;	�I;#�I;��I;wI;�^I;�II;�8I;*I;I;LI;QI;�I;L I;�H;��H;*�H;M�H;��H;�H;��H;�H;��H;M�H;*�H;��H;�H;L I;�I;QI;LI;I;*I;�8I;�II;�^I;wI;��I;#�I;	�I;�7I;w�H;^6G;�E;��A;nC=;Y<7;o�/;ο&;˧;��;��;�)�:��:���:{��:      ��;�;M;�;΢#;�);��.;�V4;B{9;\�=;M�A;��D;��F;�H;��H;�^I;ߒI;l�I;g�I;�tI;�]I;�II;=9I;5+I;UI;�I;gI;�I;4I;��H;�H;F�H;�H;z�H;o�H;��H;b�H;��H;o�H;z�H;�H;F�H;�H;��H;4I;�I;gI;�I;UI;5+I;=9I;�II;�]I;�tI;g�I;l�I;ߒI;�^I;��H;�H;��F;��D;M�A;\�=;B{9;�V4;��.;�);΢#;�;M;�;      ��2;V$3;�T4;e06;��8;-6;;��=;�@;�C;aE;2�F;��G;ϸH;};I;�I;��I;2�I;P�I;�oI;�ZI;QHI;�8I;5+I;�I;5I;2I;iI;�I;Y�H;s�H;q�H;:�H;L�H;��H;��H;i�H;�H;i�H;��H;��H;L�H;:�H;q�H;s�H;Y�H;�I;iI;2I;5I;�I;5+I;�8I;QHI;�ZI;�oI;P�I;2�I;��I;�I;};I;ϸH;��G;2�F;aE;�C;�@;��=;-6;;��8;e06;�T4;V$3;      T?@;ho@;��@;��A;��B;JD;�DE;GfF;�cG;2H;{�H;8I;WxI;�I;��I;��I;o}I;�hI;�UI;*EI;�6I;*I;UI;5I;tI;�I;QI;��H;��H;��H;-�H;0�H;��H;}�H;��H;,�H;	�H;,�H;��H;}�H;��H;0�H;-�H;��H;��H;��H;QI;�I;tI;5I;UI;*I;�6I;*EI;�UI;�hI;o}I;��I;��I;�I;WxI;8I;{�H;2H;�cG;GfF;�DE;JD;��B;��A;��@;ho@;      �eF;yF;�F;tG;ArG;e�G;�XH;��H;sI;�VI;��I;�I;��I;ÔI;�I; rI;�_I;TOI;�@I;�3I;(I;I;�I;2I;�I;jI;��H;�H;��H;a�H;?�H;q�H;#�H;9�H;|�H;�H;�H;�H;|�H;9�H;#�H;q�H;?�H;a�H;��H;�H;��H;jI;�I;2I;�I;I;(I;�3I;�@I;TOI;�_I; rI;�I;ÔI;��I;�I;��I;�VI;sI;��H;�XH;e�G;ArG;tG;�F;yF;      C�H;��H;@�H;I;�$I;kGI;�gI;.�I;\�I;؜I;�I;ÓI;�I;�uI;;eI;�UI;�GI;";I;�/I;D%I;"I;LI;gI;iI;QI;��H;�H;��H;r�H;@�H;{�H; �H;��H;�H;q�H;�H;�H;�H;q�H;�H;��H; �H;{�H;@�H;r�H;��H;�H;��H;QI;iI;gI;LI;"I;D%I;�/I;";I;�GI;�UI;;eI;�uI;�I;ÓI;�I;؜I;\�I;.�I;�gI;kGI;�$I;I;@�H;��H;      ��I;�I; �I;Z�I;јI;ΜI;G�I;A�I;r�I;�I;րI;3sI;PeI;�WI;^KI;�?I;�4I;�*I;�!I;�I;�I;QI;�I;�I;��H;�H;��H;k�H;Q�H;j�H;��H;��H;��H;�H;��H;H�H;1�H;H�H;��H;�H;��H;��H;��H;j�H;Q�H;k�H;��H;�H;��H;�I;�I;QI;�I;�I;�!I;�*I;�4I;�?I;^KI;�WI;PeI;3sI;րI;�I;r�I;A�I;G�I;ΜI;јI;Z�I; �I;�I;      ��I;�I;ۙI;��I;�I;ǎI;ڇI;UI;quI;�jI;	`I;IUI;�JI;�@I;7I;�-I;y%I;�I;�I;bI;�
I;�I;4I;Y�H;��H;��H;r�H;Q�H;i�H;��H;��H;��H;��H;,�H;��H;��H;Y�H;��H;��H;,�H;��H;��H;��H;��H;i�H;Q�H;r�H;��H;��H;Y�H;4I;�I;�
I;bI;�I;�I;y%I;�-I;7I;�@I;�JI;IUI;	`I;�jI;quI;UI;ڇI;ǎI;�I;��I;ۙI;�I;      8{I;�zI;�xI;�uI;#qI;�kI;FeI;<^I;�VI;�NI;�FI;}>I;m6I;�.I;�&I; I;�I;�I;I;�I;\I;L I;��H;s�H;��H;a�H;@�H;j�H;��H;��H;��H;��H;�H;��H;�H;��H;��H;��H;�H;��H;�H;��H;��H;��H;��H;j�H;@�H;a�H;��H;s�H;��H;L I;\I;�I;I;�I;�I; I;�&I;�.I;m6I;}>I;�FI;�NI;�VI;<^I;FeI;�kI;#qI;�uI;�xI;�zI;      �ZI;rZI;�XI;pVI;6SI;OI;@JI;�DI;O?I;F9I;3I;�,I;�&I;� I;�I;uI;QI;nI;I;I;b�H;�H;�H;q�H;-�H;?�H;{�H;��H;��H;��H;��H;��H;_�H;��H;|�H;c�H;Z�H;c�H;|�H;��H;_�H;��H;��H;��H;��H;��H;{�H;?�H;-�H;q�H;�H;�H;b�H;I;I;nI;QI;uI;�I;� I;�&I;�,I;3I;F9I;O?I;�DI;@JI;OI;6SI;pVI;�XI;rZI;      �BI;yBI;aAI;�?I;=I;�9I;D6I;%2I;�-I;)I;B$I;�I;�I;�I;�I;'I;	I;EI;�I;O�H;]�H;��H;F�H;:�H;0�H;q�H; �H;��H;��H;��H;��H;I�H;��H;U�H;�H;��H;��H;��H;�H;U�H;��H;I�H;��H;��H;��H;��H; �H;q�H;0�H;:�H;F�H;��H;]�H;O�H;�I;EI;	I;'I;�I;�I;�I;�I;B$I;)I;�-I;%2I;D6I;�9I;=I;�?I;aAI;yBI;      "1I;�0I;�/I;�.I;�,I;3*I;a'I;<$I;� I;=I;�I;�I;�I;I;h
I;�I;�I;� I;��H;��H;h�H;*�H;�H;L�H;��H;#�H;��H;��H;��H;�H;_�H;��H;8�H;��H;��H;��H;t�H;��H;��H;��H;8�H;��H;_�H;�H;��H;��H;��H;#�H;��H;L�H;�H;*�H;h�H;��H;��H;� I;�I;�I;h
I;I;�I;�I;�I;=I;� I;<$I;a'I;3*I;�,I;�.I;�/I;�0I;      �$I;s$I;�#I;�"I;0!I;8I;�I;bI;�I;�I;�I;xI;uI;oI;cI;�I;��H;��H;s�H;I�H;L�H;M�H;z�H;��H;}�H;9�H;�H;�H;,�H;��H;��H;U�H;��H;��H;b�H;@�H;(�H;@�H;b�H;��H;��H;U�H;��H;��H;,�H;�H;�H;9�H;}�H;��H;z�H;M�H;L�H;I�H;s�H;��H;��H;�I;cI;oI;uI;xI;�I;�I;�I;bI;�I;8I;0!I;�"I;�#I;s$I;      �I;EI;�I;�I;nI;�I;I;�I;yI;I;vI;�	I;/I;I;�I;i�H;�H;��H;��H;��H;��H;��H;o�H;��H;��H;|�H;q�H;��H;��H;�H;|�H;�H;��H;b�H;�H;�H;�H;�H;�H;b�H;��H;�H;|�H;�H;��H;��H;q�H;|�H;��H;��H;o�H;��H;��H;��H;��H;��H;�H;i�H;�I;I;/I;�	I;vI;I;yI;�I;I;�I;nI;�I;�I;EI;      �I;tI;�I;'I;I;�I;�I;I;�I;�I;h	I;I;�I;<I;��H;��H;i�H;d�H;r�H;��H;��H;�H;��H;i�H;,�H;�H;�H;H�H;��H;��H;c�H;��H;��H;@�H;�H;��H;��H;��H;�H;@�H;��H;��H;c�H;��H;��H;H�H;�H;�H;,�H;i�H;��H;�H;��H;��H;r�H;d�H;i�H;��H;��H;<I;�I;I;h	I;�I;�I;I;�I;�I;I;'I;�I;tI;      NI; I;�I;�I;�I;KI;�I;�I;�I;�
I;iI;.I;�I;�I;l�H;�H;��H;��H;��H;0�H;��H;��H;b�H;�H;	�H;�H;�H;1�H;Y�H;��H;Z�H;��H;t�H;(�H;�H;��H;��H;��H;�H;(�H;t�H;��H;Z�H;��H;Y�H;1�H;�H;�H;	�H;�H;b�H;��H;��H;0�H;��H;��H;��H;�H;l�H;�I;�I;.I;iI;�
I;�I;�I;�I;KI;�I;�I;�I; I;      �I;tI;�I;'I;I;�I;�I;I;�I;�I;h	I;I;�I;<I;��H;��H;i�H;d�H;r�H;��H;��H;�H;��H;i�H;,�H;�H;�H;H�H;��H;��H;c�H;��H;��H;@�H;�H;��H;��H;��H;�H;@�H;��H;��H;c�H;��H;��H;H�H;�H;�H;,�H;i�H;��H;�H;��H;��H;r�H;d�H;i�H;��H;��H;<I;�I;I;h	I;�I;�I;I;�I;�I;I;'I;�I;tI;      �I;EI;�I;�I;nI;�I;I;�I;yI;I;vI;�	I;/I;I;�I;i�H;�H;��H;��H;��H;��H;��H;o�H;��H;��H;|�H;q�H;��H;��H;�H;|�H;�H;��H;b�H;�H;�H;�H;�H;�H;b�H;��H;�H;|�H;�H;��H;��H;q�H;|�H;��H;��H;o�H;��H;��H;��H;��H;��H;�H;i�H;�I;I;/I;�	I;vI;I;yI;�I;I;�I;nI;�I;�I;EI;      �$I;s$I;�#I;�"I;0!I;8I;�I;bI;�I;�I;�I;xI;uI;oI;cI;�I;��H;��H;s�H;I�H;L�H;M�H;z�H;��H;}�H;9�H;�H;�H;,�H;��H;��H;U�H;��H;��H;b�H;@�H;(�H;@�H;b�H;��H;��H;U�H;��H;��H;,�H;�H;�H;9�H;}�H;��H;z�H;M�H;L�H;I�H;s�H;��H;��H;�I;cI;oI;uI;xI;�I;�I;�I;bI;�I;8I;0!I;�"I;�#I;s$I;      "1I;�0I;�/I;�.I;�,I;3*I;a'I;<$I;� I;=I;�I;�I;�I;I;h
I;�I;�I;� I;��H;��H;h�H;*�H;�H;L�H;��H;#�H;��H;��H;��H;�H;_�H;��H;8�H;��H;��H;��H;t�H;��H;��H;��H;8�H;��H;_�H;�H;��H;��H;��H;#�H;��H;L�H;�H;*�H;h�H;��H;��H;� I;�I;�I;h
I;I;�I;�I;�I;=I;� I;<$I;a'I;3*I;�,I;�.I;�/I;�0I;      �BI;yBI;aAI;�?I;=I;�9I;D6I;%2I;�-I;)I;B$I;�I;�I;�I;�I;'I;	I;EI;�I;O�H;]�H;��H;F�H;:�H;0�H;q�H; �H;��H;��H;��H;��H;I�H;��H;U�H;�H;��H;��H;��H;�H;U�H;��H;I�H;��H;��H;��H;��H; �H;q�H;0�H;:�H;F�H;��H;]�H;O�H;�I;EI;	I;'I;�I;�I;�I;�I;B$I;)I;�-I;%2I;D6I;�9I;=I;�?I;aAI;yBI;      �ZI;rZI;�XI;pVI;6SI;OI;@JI;�DI;O?I;F9I;3I;�,I;�&I;� I;�I;uI;QI;nI;I;I;b�H;�H;�H;q�H;-�H;?�H;{�H;��H;��H;��H;��H;��H;_�H;��H;|�H;c�H;Z�H;c�H;|�H;��H;_�H;��H;��H;��H;��H;��H;{�H;?�H;-�H;q�H;�H;�H;b�H;I;I;nI;QI;uI;�I;� I;�&I;�,I;3I;F9I;O?I;�DI;@JI;OI;6SI;pVI;�XI;rZI;      8{I;�zI;�xI;�uI;#qI;�kI;FeI;<^I;�VI;�NI;�FI;}>I;m6I;�.I;�&I; I;�I;�I;I;�I;\I;L I;��H;s�H;��H;a�H;@�H;j�H;��H;��H;��H;��H;�H;��H;�H;��H;��H;��H;�H;��H;�H;��H;��H;��H;��H;j�H;@�H;a�H;��H;s�H;��H;L I;\I;�I;I;�I;�I; I;�&I;�.I;m6I;}>I;�FI;�NI;�VI;<^I;FeI;�kI;#qI;�uI;�xI;�zI;      ��I;�I;ۙI;��I;�I;ǎI;ڇI;UI;quI;�jI;	`I;IUI;�JI;�@I;7I;�-I;y%I;�I;�I;bI;�
I;�I;4I;Y�H;��H;��H;r�H;Q�H;i�H;��H;��H;��H;��H;,�H;��H;��H;Y�H;��H;��H;,�H;��H;��H;��H;��H;i�H;Q�H;r�H;��H;��H;Y�H;4I;�I;�
I;bI;�I;�I;y%I;�-I;7I;�@I;�JI;IUI;	`I;�jI;quI;UI;ڇI;ǎI;�I;��I;ۙI;�I;      ��I;�I; �I;Z�I;јI;ΜI;G�I;A�I;r�I;�I;րI;3sI;PeI;�WI;^KI;�?I;�4I;�*I;�!I;�I;�I;QI;�I;�I;��H;�H;��H;k�H;Q�H;j�H;��H;��H;��H;�H;��H;H�H;1�H;H�H;��H;�H;��H;��H;��H;j�H;Q�H;k�H;��H;�H;��H;�I;�I;QI;�I;�I;�!I;�*I;�4I;�?I;^KI;�WI;PeI;3sI;րI;�I;r�I;A�I;G�I;ΜI;јI;Z�I; �I;�I;      C�H;��H;@�H;I;�$I;kGI;�gI;.�I;\�I;؜I;�I;ÓI;�I;�uI;;eI;�UI;�GI;";I;�/I;D%I;"I;LI;gI;iI;QI;��H;�H;��H;r�H;@�H;{�H; �H;��H;�H;q�H;�H;�H;�H;q�H;�H;��H; �H;{�H;@�H;r�H;��H;�H;��H;QI;iI;gI;LI;"I;D%I;�/I;";I;�GI;�UI;;eI;�uI;�I;ÓI;�I;؜I;\�I;.�I;�gI;kGI;�$I;I;@�H;��H;      �eF;yF;�F;tG;ArG;e�G;�XH;��H;sI;�VI;��I;�I;��I;ÔI;�I; rI;�_I;TOI;�@I;�3I;(I;I;�I;2I;�I;jI;��H;�H;��H;a�H;?�H;q�H;#�H;9�H;|�H;�H;�H;�H;|�H;9�H;#�H;q�H;?�H;a�H;��H;�H;��H;jI;�I;2I;�I;I;(I;�3I;�@I;TOI;�_I; rI;�I;ÔI;��I;�I;��I;�VI;sI;��H;�XH;e�G;ArG;tG;�F;yF;      T?@;ho@;��@;��A;��B;JD;�DE;GfF;�cG;2H;{�H;8I;WxI;�I;��I;��I;o}I;�hI;�UI;*EI;�6I;*I;UI;5I;tI;�I;QI;��H;��H;��H;-�H;0�H;��H;}�H;��H;,�H;	�H;,�H;��H;}�H;��H;0�H;-�H;��H;��H;��H;QI;�I;tI;5I;UI;*I;�6I;*EI;�UI;�hI;o}I;��I;��I;�I;WxI;8I;{�H;2H;�cG;GfF;�DE;JD;��B;��A;��@;ho@;      ��2;V$3;�T4;e06;��8;-6;;��=;�@;�C;aE;2�F;��G;ϸH;};I;�I;��I;2�I;P�I;�oI;�ZI;QHI;�8I;5+I;�I;5I;2I;iI;�I;Y�H;s�H;q�H;:�H;L�H;��H;��H;i�H;�H;i�H;��H;��H;L�H;:�H;q�H;s�H;Y�H;�I;iI;2I;5I;�I;5+I;�8I;QHI;�ZI;�oI;P�I;2�I;��I;�I;};I;ϸH;��G;2�F;aE;�C;�@;��=;-6;;��8;e06;�T4;V$3;      ��;�;M;�;΢#;�);��.;�V4;B{9;\�=;M�A;��D;��F;�H;��H;�^I;ߒI;l�I;g�I;�tI;�]I;�II;=9I;5+I;UI;�I;gI;�I;4I;��H;�H;F�H;�H;z�H;o�H;��H;b�H;��H;o�H;z�H;�H;F�H;�H;��H;4I;�I;gI;�I;UI;5+I;=9I;�II;�]I;�tI;g�I;l�I;ߒI;�^I;��H;�H;��F;��D;M�A;\�=;B{9;�V4;��.;�);΢#;�;M;�;      ���:{��:���:��:�)�:��;��;˧;ο&;o�/;Y<7;nC=;��A;�E;^6G;w�H;�7I;	�I;#�I;��I;wI;�^I;�II;�8I;*I;I;LI;QI;�I;L I;�H;��H;*�H;M�H;��H;�H;��H;�H;��H;M�H;*�H;��H;�H;L I;�I;QI;LI;I;*I;�8I;�II;�^I;wI;��I;#�I;	�I;�7I;w�H;^6G;�E;��A;nC=;Y<7;o�/;ο&;˧;��;��;�)�:��:���:{��:      �sx9���9ݤ�9�:F�^:���:�Ǽ:�N�:��;�g;�#;�;/;�:8;��>;�nC;�eF;W'H;eI;�~I;ߛI;ːI;wI;�]I;QHI;�6I;(I;"I;�I;�
I;\I;b�H;]�H;h�H;L�H;��H;��H;��H;��H;��H;L�H;h�H;]�H;b�H;\I;�
I;�I;"I;(I;�6I;QHI;�]I;wI;ːI;ߛI;�~I;eI;W'H;�eF;�nC;��>;�:8;�;/;�#;�g;��;�N�:�Ǽ:���:F�^:�:ݤ�9���9      ��f��� ��-�ht�,N���8%�&:J��:I��:�Y;[B;N�&;�&3;5<;��A;��E;��G;\I;v{I;ߛI;��I;�tI;�ZI;*EI;�3I;D%I;�I;bI;�I;I;O�H;��H;I�H;��H;��H;0�H;��H;��H;I�H;��H;O�H;I;�I;bI;�I;D%I;�3I;*EI;�ZI;�tI;��I;ߛI;v{I;\I;��G;��E;��A;5<;�&3;N�&;[B;�Y;I��:J��:%�&:��8,N�ht�-� ��f���      �N����������g���8}�g�D���� z�����H��9�
�:���:%	;,�;�.;�9;�@;]E;��G;\I;�~I;#�I;g�I;�oI;�UI;�@I;�/I;�!I;�I;I;I;�I;��H;s�H;��H;r�H;��H;r�H;��H;s�H;��H;�I;I;I;�I;�!I;�/I;�@I;�UI;�oI;g�I;#�I;�~I;\I;��G;]E;�@;�9;�.;,�;%	;���:�
�:H��9��� z�����g�D��8}��g���������      *�?��<<�@�1�;i!��z�RC����lo��{�-�1򳺵���p�&:���:Y��:��;6�+;�8;W�@;]E;��G;eI;	�I;l�I;P�I;�hI;TOI;";I;�*I;�I;�I;nI;EI;� I;��H;��H;d�H;��H;d�H;��H;��H;� I;EI;nI;�I;�I;�*I;";I;TOI;�hI;P�I;l�I;	�I;eI;��G;]E;W�@;�8;6�+;��;Y��:���:p�&:����1�{�-�lo�����RC��z�;i!�@�1��<<�      ���p���I���������W�^�85��z��̻t숻�S��gt�C�x9b��:�k�:�g;y�*;�8;�@;��E;W'H;�7I;ߒI;2�I;o}I;�_I;�GI;�4I;y%I;�I;QI;	I;�I;��H;�H;i�H;��H;i�H;�H;��H;�I;	I;QI;�I;y%I;�4I;�GI;�_I;o}I;2�I;ߒI;�7I;W'H;��E;�@;�8;y�*;�g;�k�:b��:C�x9�gt��S�t숻�̻�z�85�W�^���������I��p��      6��p��
�*���z��gC���t�� �|��?�Ъ	������V�񮼺xU��߄:��:�g;6�+;�9;��A;�eF;w�H;�^I;��I;��I; rI;�UI;�?I;�-I; I;uI;'I;�I;�I;i�H;��H;�H;��H;i�H;�I;�I;'I;uI; I;�-I;�?I;�UI; rI;��I;��I;�^I;w�H;�eF;��A;�9;6�+;�g;��:�߄:xU�񮼺��V����Ъ	��?� �|��t��gC��z��*����
�p�      ��t���p�9�d�-�Q���9�l*������Ҽ�I��O�o���'���ڻX7}� ��wH��߄:�k�:��;�.;5<;�nC;^6G;��H;�I;��I;�I;;eI;^KI;7I;�&I;�I;�I;h
I;cI;�I;��H;l�H;��H;�I;cI;h
I;�I;�I;�&I;7I;^KI;;eI;�I;��I;�I;��H;^6G;�nC;5<;�.;��;�k�:�߄:wH� ��X7}���ڻ��'�O�o��I����Ҽ���l*���9�-�Q�9�d���p�      ��Ž9���̷�V���z����}�$�Q�c�'����EC��I\��k<<�?��n�� ��xU�b��:Y��:,�;�&3;��>;�E;�H;};I;�I;ÔI;�uI;�WI;�@I;�.I;� I;�I;I;oI;I;<I;�I;<I;I;oI;I;�I;� I;�.I;�@I;�WI;�uI;ÔI;�I;};I;�H;�E;��>;�&3;,�;Y��:b��:xU� ���n��?�k<<�I\��EC�����c�'�$�Q���}��z��V��̷�9���      c.��3�ɤ�W����҈Ž<5�����fG�@��kּe���:yC�?�X7}�񮼺C�x9���:%	;N�&;�:8;��A;��F;ϸH;WxI;��I;�I;PeI;�JI;m6I;�&I;�I;�I;uI;/I;�I;�I;�I;/I;uI;�I;�I;�&I;m6I;�JI;PeI;�I;��I;WxI;ϸH;��F;��A;�:8;N�&;%	;���:C�x9񮼺X7}�?�:yC�e���kּ@��fG����<5��҈Ž��W��ɤ��3�      Fx��s��d�M�N�`�3�}I����L����z����\�P*�'�ݼe���k<<���ڻ��V��gt�p�&:���:[B;�;/;nC=;��D;��G;8I;�I;ÓI;3sI;IUI;}>I;�,I;�I;�I;xI;�	I;I;.I;I;�	I;xI;�I;�I;�,I;}>I;IUI;3sI;ÓI;�I;8I;��G;��D;nC=;�;/;[B;���:p�&:�gt���V���ڻk<<�e���'�ݼP*���\��z��L������}I�`�3�M�N��d��s�      *l¾(��S������������d���7�y��<Sؽ[�� �d�P*�kּI\����'�����S������
�:�Y;�#;Y<7;M�A;2�F;{�H;��I;�I;րI;	`I;�FI;3I;B$I;�I;�I;vI;h	I;iI;h	I;vI;�I;�I;B$I;3I;�FI;	`I;րI;�I;��I;{�H;2�F;M�A;Y<7;�#;�Y;�
�:�����S������'�I\��kּP*� �d�[��<Sؽy����7��d���������S���(��      �V������������Ͼ�d���ǆ�C�N��3��c�[����\�@��EC��O�o�Ъ	�t숻1�H��9I��:�g;o�/;\�=;aE;2H;�VI;؜I;�I;�jI;�NI;F9I;)I;=I;�I;I;�I;�
I;�I;I;�I;=I;)I;F9I;�NI;�jI;�I;؜I;�VI;2H;aE;\�=;o�/;�g;I��:H��91�t숻Ъ	�O�o�EC��@����\�[���cཱ3�C�N��ǆ��d����Ͼ���������      ~,b���\��>M���5�9��-r��#l¾睒�"&W��3�<Sؽ�z��fG�����I���?��̻{�-����J��:��;ο&;B{9;�C;�cG;sI;\�I;r�I;quI;�VI;O?I;�-I;� I;�I;yI;�I;�I;�I;yI;�I;� I;�-I;O?I;�VI;quI;r�I;\�I;sI;�cG;�C;B{9;ο&;��;J��:���{�-��̻�?��I�����fG��z��<Sؽ�3�"&W�睒�#l¾-r��9����5��>M���\�      ���"��V���J䂿��\���1�����J˾睒�C�N�y��L������c�'���Ҽ �|��z�lo�� z��%�&:�N�:˧;�V4;�@;GfF;��H;.�I;A�I;UI;<^I;�DI;%2I;<$I;bI;�I;I;�I;I;�I;bI;<$I;%2I;�DI;<^I;UI;A�I;.�I;��H;GfF;�@;�V4;˧;�N�:%�&: z��lo���z� �|���Ҽc�'����L���y��C�N�睒��J˾�����1���\�J䂿V���"��      }߿�$ڿ*�ʿ�������{Ps�MX:����#l¾�ǆ���7����<5��$�Q�����t��85���������8�Ǽ:��;��.;��=;�DE;�XH;�gI;G�I;ڇI;FeI;@JI;D6I;a'I;�I;I;�I;�I;�I;I;�I;a'I;D6I;@JI;FeI;ڇI;G�I;�gI;�XH;�DE;��=;��.;��;�Ǽ:��8������85��t�����$�Q�<5�������7��ǆ�#l¾���MX:�{Ps��������*�ʿ�$ڿ      w�����p������ſ!��{Ps���1�-r���d���d�}I�҈Ž��}�l*�gC��W�^�RC�g�D�,N๩��:��;�);-6;;JD;e�G;kGI;ΜI;ǎI;�kI;OI;�9I;3*I;8I;�I;�I;KI;�I;�I;8I;3*I;�9I;OI;�kI;ǎI;ΜI;kGI;e�G;JD;-6;;�);��;���:,N�g�D�RC�W�^�gC��l*���}�҈Ž}I��d��d��-r����1�{Ps�!����ſ��꿀p����      ��7��3�Ң%�w��<����ſ�����\�9����Ͼ����`�3����z����9�z�ἷ���z��8}�ht�F�^:�)�:΢#;��8;��B;ArG;�$I;јI;�I;#qI;6SI;=I;�,I;0!I;nI;I;�I;I;nI;0!I;�,I;=I;6SI;#qI;�I;јI;�$I;ArG;��B;��8;΢#;�)�:F�^:ht��8}��z����z�Ἁ�9��z����`�3�������Ͼ9����\������ſ�<��w�Ң%��3�      (�_��+Y��lG�f.�w���꿭���J䂿��5���󾋰��M�N�W��V��-�Q�*�������;i!��g��-󳺍:��:�;e06;��A;tG;I;Z�I;��I;�uI;pVI;�?I;�.I;�"I;�I;'I;�I;'I;�I;�"I;�.I;�?I;pVI;�uI;��I;Z�I;I;tG;��A;e06;�;��:�:-��g��;i!�����*���-�Q�V��W��M�N���������5�J䂿�������w�f.��lG��+Y�      ά��}�8tf��lG�Ң%��p�*�ʿV����>M����S����d�ɤ�̷�9�d��
��I��@�1����� ��ݤ�9���:M;�T4;��@;�F;@�H; �I;ۙI;�xI;�XI;aAI;�/I;�#I;�I;�I;�I;�I;�I;�#I;�/I;aAI;�XI;�xI;ۙI; �I;@�H;�F;��@;�T4;M;���:ݤ�9 ������@�1��I���
�9�d�̷�ɤ��d�S�������>M�V���*�ʿ�p�Ң%��lG�8tf�}�      O���A���}��+Y��3�����$ڿ"����\����(���s��3�9�����p�p�p���<<����f������9{��:�;V$3;ho@;yF;��H;�I;�I;�zI;rZI;yBI;�0I;s$I;EI;tI; I;tI;EI;s$I;�0I;yBI;rZI;�zI;�I;�I;��H;yF;ho@;V$3;�;{��:���9f�������<<�p��p���p�9����3��s�(�������\�"���$ڿ����3��+Y�}�A���      �Aq���i���U�A:�@�����6���q���uA�a5�� ��y^Z�����A���]�����d��|",�6��;�Ѻ���9'��:d�;dX4;p�@;�UF;��H;�FI;�aI;2NI;A9I;�(I;<I;�I;�I;�I;�
I;�I;�I;�I;<I;�(I;A9I;2NI;�aI;�FI;��H;�UF;p�@;dX4;d�;'��:���9;�Ѻ6��|",��d������]��A�����y^Z�� ��a5�uA�q���6�������@�A:���U���i�      ��i���b�T�O�.5�-i������������q<�����e��[
V�FE	�!���IY�s9�Z����(� S����Ⱥ��:���:'�;K�4;h�@;jgF;��H;4HI;�aI;�MI;�8I;�(I;I;~I;�I;{I;x
I;{I;�I;~I;I;�(I;�8I;�MI;�aI;4HI;��H;jgF;h�@;K�4;'�;���:��:��Ⱥ S���(�Z���s9��IY�!��FE	�[
V��e������q<������������-i�.5�T�O���b�      ��U�T�O�B-?�(�'���F�`欿Y�{�aa/���뾙���I����e���ZN�o5��Ǩ��nH�� ������ۧ":��:��;��5;�_A;ٚF;Z�H;;LI;aI;�LI;�7I;(I;aI;I;_I;%I;&
I;%I;_I;I;aI;(I;�7I;�LI;aI;;LI;Z�H;ٚF;�_A;��5;��;��:ۧ":����� ��nH�Ǩ��o5���ZN�e������I�������aa/�Y�{��欿F����(�'�B-?�T�O�      A:�.5�(�'��������dȿ���e$_���Q�Ҿؕ��
�6�����*���`=�P���)��{G��6��B����Q:�:/";�7;�%B;�F;��H;RI;�_I;�JI;C6I;�&I;YI;7I;�I;�
I;�	I;�
I;�I;7I;YI;�&I;C6I;�JI;�_I;RI;��H;�F;�%B;�7;/";�:��Q:B���6��{G��)��P���`=��*�����
�6�ؕ��Q�Ҿ��e$_����dȿ�������(�'�.5�      @�-i�������B�ѿf�������q<��:��a����q����Wн齅���'�ib̼�zl�/���X�{���:��;
�&;٪9;KC;vLG;�H;]XI;�]I;�GI;4I;�$I;I;'I;�I;�	I;�I;�	I;�I;'I;I;�$I;4I;�GI;�]I;]XI;�H;vLG;KC;٪9;
�&;��;�:{���X�/���zl�ib̼��'�齅��Wн����q��a���:��q<����f���B�ѿ������-i�      �������F��dȿf���������O���u]׾w���	�I�����A��C�d�v��֮�<RH�Kkλ �$�z5����:mM;˅+;�<;"3D;�G;�I;�]I;�ZI;DI;H1I;�"I;`I;�I;�I;�I;�I;�I;�I;�I;`I;�"I;H1I;DI;�ZI;�]I;�I;�G;"3D;�<;˅+;mM;���:z5� �$�Kkλ<RH��֮�v�C�d��A�����	�I�w���u]׾����O�����f���dȿF�ῢ��      6��������欿��������O�}x����� ���l���"��ܽ���`=�Ý��l"��R���ۺL��9�=�:�K;��0;͞>;�LE;|"H;�$I;�`I;(VI;�?I;.I;` I;[I;"I;/
I;lI;�I;lI;/
I;"I;[I;` I;.I;�?I;(VI;�`I;�$I;|"H;�LE;͞>;��0;�K;�=�:L��9�ۺ�R��l"����Ý��`=����ܽ��"��l�� �����}x���O��������欿����      q�������Y�{�e$_��q<�������}��w���6�����!��!�h��������� d��.��g_e�VL[���Z:���:�+ ;��5;�A;�UF;˃H;@I;�aI;�PI;;I;e*I;�I;+I;WI;�I;
I;LI;
I;�I;WI;+I;�I;e*I;;I;�PI;�aI;@I;˃H;�UF;�A;��5;�+ ;���:��Z:VL[�g_e��.��� d��������!�h�!�������6�w���}��������q<�e$_�Y�{�����      uA��q<�aa/����:�u]׾� ��w��>�BE	�����ܽ����3�r�꼰���>",�X��4��hAQ�خ�:�L
;�e);݄:;D?C;?G;|�H;fSI;�^I;KJI;6I;t&I;�I;�I;ZI;�I;�I;�I;�I;�I;ZI;�I;�I;t&I;6I;KJI;�^I;fSI;|�H;?G;D?C;݄:;�e);�L
;خ�:hAQ�4��X��>",�����r�꼠�3�ܽ������BE	�>�w��� ��u]׾�:���aa/��q<�      a5�������Q�Ҿ�a��w����l��6�BE	���Ƚk���aG����z֮�C�W����:�k����S`,:���:�;��1;m�>;^E;L�G;BI;G^I;hYI;YCI;�0I;U"I;cI;I;#	I;,I;�I;=I;�I;,I;#	I;I;cI;U"I;�0I;YCI;hYI;G^I;BI;L�G;^E;m�>;��1;�;���:S`,:���:�k����C�W�z֮�����aG�k����ȽBE	��6��l�w����a��Q�Ҿ������      � ���e�����ؕ����q�	�I���"���������k���ZN�c�6¼~�y��$�PR��]� �_�[��:G/;J�&;
w8;��A;��F;��H;?I;aI;�QI;:<I;7+I;�I;I;uI;�I;WI;9I;� I;9I;WI;�I;uI;I;�I;7+I;:<I;�QI;aI;?I;��H;��F;��A;
w8;J�&;G/;�:_�[�]� �PR���$�~�y�6¼c��ZN�k������������"�	�I���q�ؕ������e��      y^Z�[
V��I�
�6�������ܽ!��ܽ���aG�c��ȼ�)����(����H5���,�Z:j�:7R;.&1;��=;ПD;O�G;�H;�WI;9]I;�HI;5I;�%I;�I;�I;�	I;�I;mI;|�H;��H;|�H;mI;�I;�	I;�I;�I;�%I;5I;�HI;9]I;�WI;�H;O�G;ПD;��=;.&1;7R;j�:,�Z:��H5������(��)���ȼc��aG�ܽ��!���ܽ�����
�6��I�[
V�      ���FE	��������Wн�A����!�h���3����6¼�)��ax/�v�һD�X�!%����9���:�=;[e);�_9;�%B;ډF;�|H;�5I;u`I;�TI;�?I;�-I; I;jI;DI;�I;jI;p�H;��H;�H;��H;p�H;jI;�I;DI;jI; I;�-I;�?I;�TI;u`I;�5I;�|H;ډF;�%B;�_9;[e);�=;���:��9!%��D�X�v�һax/��)��6¼�����3�!�h��󑽢A���Wн��콹��FE	�      �A��!��e���*��齅�C�d��`=����r��z֮�~�y���(�v�һk^e�������f9���:X�;m0";A�4;�l?; E;��G;��H;�VI;�]I;(JI;�6I;'I;�I;FI;�	I;=I;7 I;��H;��H;V�H;��H;��H;7 I;=I;�	I;FI;�I;'I;�6I;(JI;�]I;�VI;��H;��G; E;�l?;A�4;m0";X�;���:��f9����k^e�v�һ��(�~�y�z֮�r�꼠���`=�C�d�齅��*��e��!��      �]��IY��ZN��`=���'�v�Ý���������C�W��$����D�X������9�ޚ:���:��;ʷ0;�<;v�C;GG;�H;�>I;P`I;�SI;^?I;1.I;z I;�I;.I;�I;�I;��H;��H;&�H;��H;&�H;��H;��H;�I;�I;.I;�I;z I;1.I;^?I;�SI;P`I;�>I;�H;GG;v�C;�<;ʷ0;��;���:�ޚ:�9����D�X�����$�C�W���������Ý�v���'��`=��ZN��IY�      ���s9�o5��P��ib̼�֮����� d�>",����PR��H5�!%����f9�ޚ:��:5�;��-;��:;KB;_UF;:JH; I;�[I;G[I;�GI;%5I;<&I;6I;�I;8	I;^I;�H;��H;��H;n�H;�H;n�H;��H;��H;�H;^I;8	I;�I;6I;<&I;%5I;�GI;G[I;�[I; I;:JH;_UF;KB;��:;��-;5�;��:�ޚ:��f9!%��H5�PR�����>",�� d�����֮�ib̼P��o5��s9�      �d��Z���Ǩ���)���zl�<RH�l"��.��X��:�k�]� �����9���:���:5�;�-;�9;i`A;ڹE;J�G;��H;#RI;4_I;OI;�;I;�+I;�I;MI;)I;�I;p I;��H;��H;��H;��H;{�H;��H;��H;��H;��H;p I;�I;)I;MI;�I;�+I;�;I;OI;4_I;#RI;��H;J�G;ڹE;i`A;�9;�-;5�;���:���:��9��]� �:�k�X���.��l"�<RH��zl��)��Ǩ��Z���      |",��(�nH�{G�/��Kkλ�R��g_e�4�����_�[�,�Z:���:X�;��;��-;�9;�A;�bE;D�G;��H;tFI;`I;�TI;bAI;�0I;#I;�I;I;�I;I;��H;a�H;��H;!�H;,�H;��H;,�H;!�H;��H;a�H;��H;I;�I;I;�I;#I;�0I;bAI;�TI;`I;tFI;��H;D�G;�bE;�A;�9;��-;��;X�;���:,�Z:_�[����4��g_e��R��Kkλ/��{G�nH��(�      6�� S��� ���6���X� �$��ۺVL[�hAQ�S`,:�:j�:�=;m0";ʷ0;��:;i`A;�bE;�G;��H;�<I;N_I;�XI;FI;5I;�&I;I;�I;
I;�I;��H;�H;5�H;�H;��H;��H;S�H;��H;��H;�H;5�H;�H;��H;�I;
I;�I;I;�&I;5I;FI;�XI;N_I;�<I;��H;�G;�bE;i`A;��:;ʷ0;m0";�=;j�:�:S`,:hAQ�VL[��ۺ �$��X��6��� �� S��      ;�Ѻ��Ⱥ����B��{��z5�L��9��Z:خ�:���:G/;7R;[e);A�4;�<;KB;ڹE;D�G;��H;9I;q^I;�ZI;?II;8I;�)I;�I;I;I;vI;$ I;��H;��H;%�H;C�H;�H;F�H;��H;F�H;�H;C�H;%�H;��H;��H;$ I;vI;I;I;�I;�)I;8I;?II;�ZI;q^I;9I;��H;D�G;ڹE;KB;�<;A�4;[e);7R;G/;���:خ�:��Z:L��9z5�{��B��������Ⱥ      ���9��:ۧ":��Q:�:���:�=�:���:�L
;�;J�&;.&1;�_9;�l?;v�C;_UF;J�G;��H;�<I;q^I;1[I;�JI;1:I;�+I;�I;I;�I;�I;_I;��H;K�H;��H;J�H;��H;��H;��H;��H;��H;��H;��H;J�H;��H;K�H;��H;_I;�I;�I;I;�I;�+I;1:I;�JI;1[I;q^I;�<I;��H;J�G;_UF;v�C;�l?;�_9;.&1;J�&;�;�L
;���:�=�:���:�:��Q:ۧ":��:      '��:���:��:�:��;mM;�K;�+ ;�e);��1;
w8;��=;�%B; E;GG;:JH;��H;tFI;N_I;�ZI;�JI;�:I;-I;H!I;QI;*I;0I;xI;��H;��H;��H;}�H;��H;-�H;Q�H;��H;y�H;��H;Q�H;-�H;��H;}�H;��H;��H;��H;xI;0I;*I;QI;H!I;-I;�:I;�JI;�ZI;N_I;tFI;��H;:JH;GG; E;�%B;��=;
w8;��1;�e);�+ ;�K;mM;��;�:��:���:      d�;'�;��;/";
�&;˅+;��0;��5;݄:;m�>;��A;ПD;ډF;��G;�H; I;#RI;`I;�XI;?II;1:I;-I;�!I;I;�I;	I;BI;]�H;��H;j�H;��H;��H;
�H;��H; �H;��H;p�H;��H; �H;��H;
�H;��H;��H;j�H;��H;]�H;BI;	I;�I;I;�!I;-I;1:I;?II;�XI;`I;#RI; I;�H;��G;ډF;ПD;��A;m�>;݄:;��5;��0;˅+;
�&;/";��;'�;      dX4;K�4;��5;�7;٪9;�<;͞>;�A;D?C;^E;��F;O�G;�|H;��H;�>I;�[I;4_I;�TI;FI;8I;�+I;H!I;I;8I;v	I;�I; �H;��H;��H;��H;��H;�H;��H;��H;��H;��H;u�H;��H;��H;��H;��H;�H;��H;��H;��H;��H; �H;�I;v	I;8I;I;H!I;�+I;8I;FI;�TI;4_I;�[I;�>I;��H;�|H;O�G;��F;^E;D?C;�A;͞>;�<;٪9;�7;��5;K�4;      p�@;h�@;�_A;�%B;KC;"3D;�LE;�UF;?G;L�G;��H;�H;�5I;�VI;P`I;G[I;OI;bAI;5I;�)I;�I;QI;�I;v	I;I;.�H;D�H;��H;0�H;��H;�H;��H;[�H;��H;��H;��H;r�H;��H;��H;��H;[�H;��H;�H;��H;0�H;��H;D�H;.�H;I;v	I;�I;QI;�I;�)I;5I;bAI;OI;G[I;P`I;�VI;�5I;�H;��H;L�G;?G;�UF;�LE;"3D;KC;�%B;�_A;h�@;      �UF;jgF;ٚF;�F;vLG;�G;|"H;˃H;|�H;BI;?I;�WI;u`I;�]I;�SI;�GI;�;I;�0I;�&I;�I;I;*I;	I;�I;.�H;V�H;'�H;i�H;��H;�H;��H;V�H;L�H;��H;�H;��H;��H;��H;�H;��H;L�H;V�H;��H;�H;��H;i�H;'�H;V�H;.�H;�I;	I;*I;I;�I;�&I;�0I;�;I;�GI;�SI;�]I;u`I;�WI;?I;BI;|�H;˃H;|"H;�G;vLG;�F;ٚF;jgF;      ��H;��H;Z�H;��H;�H;�I;�$I;@I;fSI;G^I;aI;9]I;�TI;(JI;^?I;%5I;�+I;#I;I;I;�I;0I;BI; �H;D�H;'�H;\�H;�H;7�H;|�H;6�H;�H;E�H;��H;@�H;��H;��H;��H;@�H;��H;E�H;�H;6�H;|�H;7�H;�H;\�H;'�H;D�H; �H;BI;0I;�I;I;I;#I;�+I;%5I;^?I;(JI;�TI;9]I;aI;G^I;fSI;@I;�$I;�I;�H;��H;Z�H;��H;      �FI;4HI;;LI;RI;]XI;�]I;�`I;�aI;�^I;hYI;�QI;�HI;�?I;�6I;1.I;<&I;�I;�I;�I;I;�I;xI;]�H;��H;��H;i�H;�H;�H;��H;2�H;�H;�H;p�H;��H;|�H;F�H;@�H;F�H;|�H;��H;p�H;�H;�H;2�H;��H;�H;�H;i�H;��H;��H;]�H;xI;�I;I;�I;�I;�I;<&I;1.I;�6I;�?I;�HI;�QI;hYI;�^I;�aI;�`I;�]I;]XI;RI;;LI;4HI;      �aI;�aI;aI;�_I;�]I;�ZI;(VI;�PI;KJI;YCI;:<I;5I;�-I;'I;z I;6I;MI;I;
I;vI;_I;��H;��H;��H;0�H;��H;7�H;��H;)�H;�H; �H;B�H;��H;2�H;��H;��H;��H;��H;��H;2�H;��H;B�H; �H;�H;)�H;��H;7�H;��H;0�H;��H;��H;��H;_I;vI;
I;I;MI;6I;z I;'I;�-I;5I;:<I;YCI;KJI;�PI;(VI;�ZI;�]I;�_I;aI;�aI;      2NI;�MI;�LI;�JI;�GI;DI;�?I;;I;6I;�0I;7+I;�%I; I;�I;�I;�I;)I;�I;�I;$ I;��H;��H;j�H;��H;��H;�H;|�H;2�H;�H;�H;1�H;��H;��H;��H;H�H;(�H;%�H;(�H;H�H;��H;��H;��H;1�H;�H;�H;2�H;|�H;�H;��H;��H;j�H;��H;��H;$ I;�I;�I;)I;�I;�I;�I; I;�%I;7+I;�0I;6I;;I;�?I;DI;�GI;�JI;�LI;�MI;      A9I;�8I;�7I;C6I;4I;H1I;.I;e*I;t&I;U"I;�I;�I;jI;FI;.I;8	I;�I;I;��H;��H;K�H;��H;��H;��H;�H;��H;6�H;�H; �H;1�H;��H;��H;d�H;�H;��H;��H;��H;��H;��H;�H;d�H;��H;��H;1�H; �H;�H;6�H;��H;�H;��H;��H;��H;K�H;��H;��H;I;�I;8	I;.I;FI;jI;�I;�I;U"I;t&I;e*I;.I;H1I;4I;C6I;�7I;�8I;      �(I;�(I;(I;�&I;�$I;�"I;` I;�I;�I;cI;I;�I;DI;�	I;�I;^I;p I;��H;�H;��H;��H;}�H;��H;�H;��H;V�H;�H;�H;B�H;��H;��H;{�H;��H;��H;z�H;T�H;>�H;T�H;z�H;��H;��H;{�H;��H;��H;B�H;�H;�H;V�H;��H;�H;��H;}�H;��H;��H;�H;��H;p I;^I;�I;�	I;DI;�I;I;cI;�I;�I;` I;�"I;�$I;�&I;(I;�(I;      <I;I;aI;YI;I;`I;[I;+I;�I;I;uI;�	I;�I;=I;�I;�H;��H;a�H;5�H;%�H;J�H;��H;
�H;��H;[�H;L�H;E�H;p�H;��H;��H;d�H;��H;��H;[�H;�H;�H;�H;�H;�H;[�H;��H;��H;d�H;��H;��H;p�H;E�H;L�H;[�H;��H;
�H;��H;J�H;%�H;5�H;a�H;��H;�H;�I;=I;�I;�	I;uI;I;�I;+I;[I;`I;I;YI;aI;I;      �I;~I;I;7I;'I;�I;"I;WI;ZI;#	I;�I;�I;jI;7 I;��H;��H;��H;��H;�H;C�H;��H;-�H;��H;��H;��H;��H;��H;��H;2�H;��H;�H;��H;[�H; �H;��H;��H;��H;��H;��H; �H;[�H;��H;�H;��H;2�H;��H;��H;��H;��H;��H;��H;-�H;��H;C�H;�H;��H;��H;��H;��H;7 I;jI;�I;�I;#	I;ZI;WI;"I;�I;'I;7I;I;~I;      �I;�I;_I;�I;�I;�I;/
I;�I;�I;,I;WI;mI;p�H;��H;��H;��H;��H;!�H;��H;�H;��H;Q�H; �H;��H;��H;�H;@�H;|�H;��H;H�H;��H;z�H;�H;��H;��H;��H;��H;��H;��H;��H;�H;z�H;��H;H�H;��H;|�H;@�H;�H;��H;��H; �H;Q�H;��H;�H;��H;!�H;��H;��H;��H;��H;p�H;mI;WI;,I;�I;�I;/
I;�I;�I;�I;_I;�I;      �I;{I;%I;�
I;�	I;�I;lI;
I;�I;�I;9I;|�H;��H;��H;&�H;n�H;��H;,�H;��H;F�H;��H;��H;��H;��H;��H;��H;��H;F�H;��H;(�H;��H;T�H;�H;��H;��H;��H;}�H;��H;��H;��H;�H;T�H;��H;(�H;��H;F�H;��H;��H;��H;��H;��H;��H;��H;F�H;��H;,�H;��H;n�H;&�H;��H;��H;|�H;9I;�I;�I;
I;lI;�I;�	I;�
I;%I;{I;      �
I;x
I;&
I;�	I;�I;�I;�I;LI;�I;=I;� I;��H;�H;V�H;��H;�H;{�H;��H;S�H;��H;��H;y�H;p�H;u�H;r�H;��H;��H;@�H;��H;%�H;��H;>�H;�H;��H;��H;}�H;��H;}�H;��H;��H;�H;>�H;��H;%�H;��H;@�H;��H;��H;r�H;u�H;p�H;y�H;��H;��H;S�H;��H;{�H;�H;��H;V�H;�H;��H;� I;=I;�I;LI;�I;�I;�I;�	I;&
I;x
I;      �I;{I;%I;�
I;�	I;�I;lI;
I;�I;�I;9I;|�H;��H;��H;&�H;n�H;��H;,�H;��H;F�H;��H;��H;��H;��H;��H;��H;��H;F�H;��H;(�H;��H;T�H;�H;��H;��H;��H;}�H;��H;��H;��H;�H;T�H;��H;(�H;��H;F�H;��H;��H;��H;��H;��H;��H;��H;F�H;��H;,�H;��H;n�H;&�H;��H;��H;|�H;9I;�I;�I;
I;lI;�I;�	I;�
I;%I;{I;      �I;�I;_I;�I;�I;�I;/
I;�I;�I;,I;WI;mI;p�H;��H;��H;��H;��H;!�H;��H;�H;��H;Q�H; �H;��H;��H;�H;@�H;|�H;��H;H�H;��H;z�H;�H;��H;��H;��H;��H;��H;��H;��H;�H;z�H;��H;H�H;��H;|�H;@�H;�H;��H;��H; �H;Q�H;��H;�H;��H;!�H;��H;��H;��H;��H;p�H;mI;WI;,I;�I;�I;/
I;�I;�I;�I;_I;�I;      �I;~I;I;7I;'I;�I;"I;WI;ZI;#	I;�I;�I;jI;7 I;��H;��H;��H;��H;�H;C�H;��H;-�H;��H;��H;��H;��H;��H;��H;2�H;��H;�H;��H;[�H; �H;��H;��H;��H;��H;��H; �H;[�H;��H;�H;��H;2�H;��H;��H;��H;��H;��H;��H;-�H;��H;C�H;�H;��H;��H;��H;��H;7 I;jI;�I;�I;#	I;ZI;WI;"I;�I;'I;7I;I;~I;      <I;I;aI;YI;I;`I;[I;+I;�I;I;uI;�	I;�I;=I;�I;�H;��H;a�H;5�H;%�H;J�H;��H;
�H;��H;[�H;L�H;E�H;p�H;��H;��H;d�H;��H;��H;[�H;�H;�H;�H;�H;�H;[�H;��H;��H;d�H;��H;��H;p�H;E�H;L�H;[�H;��H;
�H;��H;J�H;%�H;5�H;a�H;��H;�H;�I;=I;�I;�	I;uI;I;�I;+I;[I;`I;I;YI;aI;I;      �(I;�(I;(I;�&I;�$I;�"I;` I;�I;�I;cI;I;�I;DI;�	I;�I;^I;p I;��H;�H;��H;��H;}�H;��H;�H;��H;V�H;�H;�H;B�H;��H;��H;{�H;��H;��H;z�H;T�H;>�H;T�H;z�H;��H;��H;{�H;��H;��H;B�H;�H;�H;V�H;��H;�H;��H;}�H;��H;��H;�H;��H;p I;^I;�I;�	I;DI;�I;I;cI;�I;�I;` I;�"I;�$I;�&I;(I;�(I;      A9I;�8I;�7I;C6I;4I;H1I;.I;e*I;t&I;U"I;�I;�I;jI;FI;.I;8	I;�I;I;��H;��H;K�H;��H;��H;��H;�H;��H;6�H;�H; �H;1�H;��H;��H;d�H;�H;��H;��H;��H;��H;��H;�H;d�H;��H;��H;1�H; �H;�H;6�H;��H;�H;��H;��H;��H;K�H;��H;��H;I;�I;8	I;.I;FI;jI;�I;�I;U"I;t&I;e*I;.I;H1I;4I;C6I;�7I;�8I;      2NI;�MI;�LI;�JI;�GI;DI;�?I;;I;6I;�0I;7+I;�%I; I;�I;�I;�I;)I;�I;�I;$ I;��H;��H;j�H;��H;��H;�H;|�H;2�H;�H;�H;1�H;��H;��H;��H;H�H;(�H;%�H;(�H;H�H;��H;��H;��H;1�H;�H;�H;2�H;|�H;�H;��H;��H;j�H;��H;��H;$ I;�I;�I;)I;�I;�I;�I; I;�%I;7+I;�0I;6I;;I;�?I;DI;�GI;�JI;�LI;�MI;      �aI;�aI;aI;�_I;�]I;�ZI;(VI;�PI;KJI;YCI;:<I;5I;�-I;'I;z I;6I;MI;I;
I;vI;_I;��H;��H;��H;0�H;��H;7�H;��H;)�H;�H; �H;B�H;��H;2�H;��H;��H;��H;��H;��H;2�H;��H;B�H; �H;�H;)�H;��H;7�H;��H;0�H;��H;��H;��H;_I;vI;
I;I;MI;6I;z I;'I;�-I;5I;:<I;YCI;KJI;�PI;(VI;�ZI;�]I;�_I;aI;�aI;      �FI;4HI;;LI;RI;]XI;�]I;�`I;�aI;�^I;hYI;�QI;�HI;�?I;�6I;1.I;<&I;�I;�I;�I;I;�I;xI;]�H;��H;��H;i�H;�H;�H;��H;2�H;�H;�H;p�H;��H;|�H;F�H;@�H;F�H;|�H;��H;p�H;�H;�H;2�H;��H;�H;�H;i�H;��H;��H;]�H;xI;�I;I;�I;�I;�I;<&I;1.I;�6I;�?I;�HI;�QI;hYI;�^I;�aI;�`I;�]I;]XI;RI;;LI;4HI;      ��H;��H;Z�H;��H;�H;�I;�$I;@I;fSI;G^I;aI;9]I;�TI;(JI;^?I;%5I;�+I;#I;I;I;�I;0I;BI; �H;D�H;'�H;\�H;�H;7�H;|�H;6�H;�H;E�H;��H;@�H;��H;��H;��H;@�H;��H;E�H;�H;6�H;|�H;7�H;�H;\�H;'�H;D�H; �H;BI;0I;�I;I;I;#I;�+I;%5I;^?I;(JI;�TI;9]I;aI;G^I;fSI;@I;�$I;�I;�H;��H;Z�H;��H;      �UF;jgF;ٚF;�F;vLG;�G;|"H;˃H;|�H;BI;?I;�WI;u`I;�]I;�SI;�GI;�;I;�0I;�&I;�I;I;*I;	I;�I;.�H;V�H;'�H;i�H;��H;�H;��H;V�H;L�H;��H;�H;��H;��H;��H;�H;��H;L�H;V�H;��H;�H;��H;i�H;'�H;V�H;.�H;�I;	I;*I;I;�I;�&I;�0I;�;I;�GI;�SI;�]I;u`I;�WI;?I;BI;|�H;˃H;|"H;�G;vLG;�F;ٚF;jgF;      p�@;h�@;�_A;�%B;KC;"3D;�LE;�UF;?G;L�G;��H;�H;�5I;�VI;P`I;G[I;OI;bAI;5I;�)I;�I;QI;�I;v	I;I;.�H;D�H;��H;0�H;��H;�H;��H;[�H;��H;��H;��H;r�H;��H;��H;��H;[�H;��H;�H;��H;0�H;��H;D�H;.�H;I;v	I;�I;QI;�I;�)I;5I;bAI;OI;G[I;P`I;�VI;�5I;�H;��H;L�G;?G;�UF;�LE;"3D;KC;�%B;�_A;h�@;      dX4;K�4;��5;�7;٪9;�<;͞>;�A;D?C;^E;��F;O�G;�|H;��H;�>I;�[I;4_I;�TI;FI;8I;�+I;H!I;I;8I;v	I;�I; �H;��H;��H;��H;��H;�H;��H;��H;��H;��H;u�H;��H;��H;��H;��H;�H;��H;��H;��H;��H; �H;�I;v	I;8I;I;H!I;�+I;8I;FI;�TI;4_I;�[I;�>I;��H;�|H;O�G;��F;^E;D?C;�A;͞>;�<;٪9;�7;��5;K�4;      d�;'�;��;/";
�&;˅+;��0;��5;݄:;m�>;��A;ПD;ډF;��G;�H; I;#RI;`I;�XI;?II;1:I;-I;�!I;I;�I;	I;BI;]�H;��H;j�H;��H;��H;
�H;��H; �H;��H;p�H;��H; �H;��H;
�H;��H;��H;j�H;��H;]�H;BI;	I;�I;I;�!I;-I;1:I;?II;�XI;`I;#RI; I;�H;��G;ډF;ПD;��A;m�>;݄:;��5;��0;˅+;
�&;/";��;'�;      '��:���:��:�:��;mM;�K;�+ ;�e);��1;
w8;��=;�%B; E;GG;:JH;��H;tFI;N_I;�ZI;�JI;�:I;-I;H!I;QI;*I;0I;xI;��H;��H;��H;}�H;��H;-�H;Q�H;��H;y�H;��H;Q�H;-�H;��H;}�H;��H;��H;��H;xI;0I;*I;QI;H!I;-I;�:I;�JI;�ZI;N_I;tFI;��H;:JH;GG; E;�%B;��=;
w8;��1;�e);�+ ;�K;mM;��;�:��:���:      ���9��:ۧ":��Q:�:���:�=�:���:�L
;�;J�&;.&1;�_9;�l?;v�C;_UF;J�G;��H;�<I;q^I;1[I;�JI;1:I;�+I;�I;I;�I;�I;_I;��H;K�H;��H;J�H;��H;��H;��H;��H;��H;��H;��H;J�H;��H;K�H;��H;_I;�I;�I;I;�I;�+I;1:I;�JI;1[I;q^I;�<I;��H;J�G;_UF;v�C;�l?;�_9;.&1;J�&;�;�L
;���:�=�:���:�:��Q:ۧ":��:      ;�Ѻ��Ⱥ����B��{��z5�L��9��Z:خ�:���:G/;7R;[e);A�4;�<;KB;ڹE;D�G;��H;9I;q^I;�ZI;?II;8I;�)I;�I;I;I;vI;$ I;��H;��H;%�H;C�H;�H;F�H;��H;F�H;�H;C�H;%�H;��H;��H;$ I;vI;I;I;�I;�)I;8I;?II;�ZI;q^I;9I;��H;D�G;ڹE;KB;�<;A�4;[e);7R;G/;���:خ�:��Z:L��9z5�{��B��������Ⱥ      6�� S��� ���6���X� �$��ۺVL[�hAQ�S`,:�:j�:�=;m0";ʷ0;��:;i`A;�bE;�G;��H;�<I;N_I;�XI;FI;5I;�&I;I;�I;
I;�I;��H;�H;5�H;�H;��H;��H;S�H;��H;��H;�H;5�H;�H;��H;�I;
I;�I;I;�&I;5I;FI;�XI;N_I;�<I;��H;�G;�bE;i`A;��:;ʷ0;m0";�=;j�:�:S`,:hAQ�VL[��ۺ �$��X��6��� �� S��      |",��(�nH�{G�/��Kkλ�R��g_e�4�����_�[�,�Z:���:X�;��;��-;�9;�A;�bE;D�G;��H;tFI;`I;�TI;bAI;�0I;#I;�I;I;�I;I;��H;a�H;��H;!�H;,�H;��H;,�H;!�H;��H;a�H;��H;I;�I;I;�I;#I;�0I;bAI;�TI;`I;tFI;��H;D�G;�bE;�A;�9;��-;��;X�;���:,�Z:_�[����4��g_e��R��Kkλ/��{G�nH��(�      �d��Z���Ǩ���)���zl�<RH�l"��.��X��:�k�]� �����9���:���:5�;�-;�9;i`A;ڹE;J�G;��H;#RI;4_I;OI;�;I;�+I;�I;MI;)I;�I;p I;��H;��H;��H;��H;{�H;��H;��H;��H;��H;p I;�I;)I;MI;�I;�+I;�;I;OI;4_I;#RI;��H;J�G;ڹE;i`A;�9;�-;5�;���:���:��9��]� �:�k�X���.��l"�<RH��zl��)��Ǩ��Z���      ���s9�o5��P��ib̼�֮����� d�>",����PR��H5�!%����f9�ޚ:��:5�;��-;��:;KB;_UF;:JH; I;�[I;G[I;�GI;%5I;<&I;6I;�I;8	I;^I;�H;��H;��H;n�H;�H;n�H;��H;��H;�H;^I;8	I;�I;6I;<&I;%5I;�GI;G[I;�[I; I;:JH;_UF;KB;��:;��-;5�;��:�ޚ:��f9!%��H5�PR�����>",�� d�����֮�ib̼P��o5��s9�      �]��IY��ZN��`=���'�v�Ý���������C�W��$����D�X������9�ޚ:���:��;ʷ0;�<;v�C;GG;�H;�>I;P`I;�SI;^?I;1.I;z I;�I;.I;�I;�I;��H;��H;&�H;��H;&�H;��H;��H;�I;�I;.I;�I;z I;1.I;^?I;�SI;P`I;�>I;�H;GG;v�C;�<;ʷ0;��;���:�ޚ:�9����D�X�����$�C�W���������Ý�v���'��`=��ZN��IY�      �A��!��e���*��齅�C�d��`=����r��z֮�~�y���(�v�һk^e�������f9���:X�;m0";A�4;�l?; E;��G;��H;�VI;�]I;(JI;�6I;'I;�I;FI;�	I;=I;7 I;��H;��H;V�H;��H;��H;7 I;=I;�	I;FI;�I;'I;�6I;(JI;�]I;�VI;��H;��G; E;�l?;A�4;m0";X�;���:��f9����k^e�v�һ��(�~�y�z֮�r�꼠���`=�C�d�齅��*��e��!��      ���FE	��������Wн�A����!�h���3����6¼�)��ax/�v�һD�X�!%����9���:�=;[e);�_9;�%B;ډF;�|H;�5I;u`I;�TI;�?I;�-I; I;jI;DI;�I;jI;p�H;��H;�H;��H;p�H;jI;�I;DI;jI; I;�-I;�?I;�TI;u`I;�5I;�|H;ډF;�%B;�_9;[e);�=;���:��9!%��D�X�v�һax/��)��6¼�����3�!�h��󑽢A���Wн��콹��FE	�      y^Z�[
V��I�
�6�������ܽ!��ܽ���aG�c��ȼ�)����(����H5���,�Z:j�:7R;.&1;��=;ПD;O�G;�H;�WI;9]I;�HI;5I;�%I;�I;�I;�	I;�I;mI;|�H;��H;|�H;mI;�I;�	I;�I;�I;�%I;5I;�HI;9]I;�WI;�H;O�G;ПD;��=;.&1;7R;j�:,�Z:��H5������(��)���ȼc��aG�ܽ��!���ܽ�����
�6��I�[
V�      � ���e�����ؕ����q�	�I���"���������k���ZN�c�6¼~�y��$�PR��]� �_�[��:G/;J�&;
w8;��A;��F;��H;?I;aI;�QI;:<I;7+I;�I;I;uI;�I;WI;9I;� I;9I;WI;�I;uI;I;�I;7+I;:<I;�QI;aI;?I;��H;��F;��A;
w8;J�&;G/;�:_�[�]� �PR���$�~�y�6¼c��ZN�k������������"�	�I���q�ؕ������e��      a5�������Q�Ҿ�a��w����l��6�BE	���Ƚk���aG����z֮�C�W����:�k����S`,:���:�;��1;m�>;^E;L�G;BI;G^I;hYI;YCI;�0I;U"I;cI;I;#	I;,I;�I;=I;�I;,I;#	I;I;cI;U"I;�0I;YCI;hYI;G^I;BI;L�G;^E;m�>;��1;�;���:S`,:���:�k����C�W�z֮�����aG�k����ȽBE	��6��l�w����a��Q�Ҿ������      uA��q<�aa/����:�u]׾� ��w��>�BE	�����ܽ����3�r�꼰���>",�X��4��hAQ�خ�:�L
;�e);݄:;D?C;?G;|�H;fSI;�^I;KJI;6I;t&I;�I;�I;ZI;�I;�I;�I;�I;�I;ZI;�I;�I;t&I;6I;KJI;�^I;fSI;|�H;?G;D?C;݄:;�e);�L
;خ�:hAQ�4��X��>",�����r�꼠�3�ܽ������BE	�>�w��� ��u]׾�:���aa/��q<�      q�������Y�{�e$_��q<�������}��w���6�����!��!�h��������� d��.��g_e�VL[���Z:���:�+ ;��5;�A;�UF;˃H;@I;�aI;�PI;;I;e*I;�I;+I;WI;�I;
I;LI;
I;�I;WI;+I;�I;e*I;;I;�PI;�aI;@I;˃H;�UF;�A;��5;�+ ;���:��Z:VL[�g_e��.��� d��������!�h�!�������6�w���}��������q<�e$_�Y�{�����      6��������欿��������O�}x����� ���l���"��ܽ���`=�Ý��l"��R���ۺL��9�=�:�K;��0;͞>;�LE;|"H;�$I;�`I;(VI;�?I;.I;` I;[I;"I;/
I;lI;�I;lI;/
I;"I;[I;` I;.I;�?I;(VI;�`I;�$I;|"H;�LE;͞>;��0;�K;�=�:L��9�ۺ�R��l"����Ý��`=����ܽ��"��l�� �����}x���O��������欿����      �������F��dȿf���������O���u]׾w���	�I�����A��C�d�v��֮�<RH�Kkλ �$�z5����:mM;˅+;�<;"3D;�G;�I;�]I;�ZI;DI;H1I;�"I;`I;�I;�I;�I;�I;�I;�I;�I;`I;�"I;H1I;DI;�ZI;�]I;�I;�G;"3D;�<;˅+;mM;���:z5� �$�Kkλ<RH��֮�v�C�d��A�����	�I�w���u]׾����O�����f���dȿF�ῢ��      @�-i�������B�ѿf�������q<��:��a����q����Wн齅���'�ib̼�zl�/���X�{���:��;
�&;٪9;KC;vLG;�H;]XI;�]I;�GI;4I;�$I;I;'I;�I;�	I;�I;�	I;�I;'I;I;�$I;4I;�GI;�]I;]XI;�H;vLG;KC;٪9;
�&;��;�:{���X�/���zl�ib̼��'�齅��Wн����q��a���:��q<����f���B�ѿ������-i�      A:�.5�(�'��������dȿ���e$_���Q�Ҿؕ��
�6�����*���`=�P���)��{G��6��B����Q:�:/";�7;�%B;�F;��H;RI;�_I;�JI;C6I;�&I;YI;7I;�I;�
I;�	I;�
I;�I;7I;YI;�&I;C6I;�JI;�_I;RI;��H;�F;�%B;�7;/";�:��Q:B���6��{G��)��P���`=��*�����
�6�ؕ��Q�Ҿ��e$_����dȿ�������(�'�.5�      ��U�T�O�B-?�(�'���F�`欿Y�{�aa/���뾙���I����e���ZN�o5��Ǩ��nH�� ������ۧ":��:��;��5;�_A;ٚF;Z�H;;LI;aI;�LI;�7I;(I;aI;I;_I;%I;&
I;%I;_I;I;aI;(I;�7I;�LI;aI;;LI;Z�H;ٚF;�_A;��5;��;��:ۧ":����� ��nH�Ǩ��o5���ZN�e������I�������aa/�Y�{��欿F����(�'�B-?�T�O�      ��i���b�T�O�.5�-i������������q<�����e��[
V�FE	�!���IY�s9�Z����(� S����Ⱥ��:���:'�;K�4;h�@;jgF;��H;4HI;�aI;�MI;�8I;�(I;I;~I;�I;{I;x
I;{I;�I;~I;I;�(I;�8I;�MI;�aI;4HI;��H;jgF;h�@;K�4;'�;���:��:��Ⱥ S���(�Z���s9��IY�!��FE	�[
V��e������q<������������-i�.5�T�O���b�      �>���8���*�O������˿�o��<�b�=\�+m־^��K�:��J�&��F�B�F���������/��������>:�r�:do ;�I6;DA;�HF;�MH;�H;!I;�I;I;�I;mI;I;q�H;��H;*�H;��H;q�H;I;mI;�I;I;�I;!I;�H;�MH;�HF;DA;�I6;do ;�r�:��>:�����/���������F��F�B�&���J�K�:�^��+m־=\�<�b��o���˿����O���*���8�      ��8��4��g&�0��2����<ƿ벗��>]����G�Ѿ�p���*7����"W��MR?�	}鼀8����s������6�G:���: !;&�6;'kA;�XF;�SH;s�H;!I;�I;�I;�I;FI;�I;e�H;��H;�H;��H;e�H;�I;FI;�I;�I;�I;!I;s�H;�SH;�XF;'kA;&�6; !;���:6�G:���s������8��	}�MR?�"W�����*7��p��G�Ѿ����>]�벗��<ƿ2���0���g&��4�      ��*��g&��#�o�K[�jL�������M�l5��>ľ
����,��D�撐��5�<�ݼ���q
���x��wk�}�b:�j�:#;ږ7;��A;�F;�cH;�I;\!I;I;oI;AI;�I;�I; �H;x�H;��H;x�H; �H;�I;�I;AI;oI;I;\!I;�I;�cH;�F;��A;ږ7;#;�j�:}�b:�wk���x��q
���<�ݼ�5�撐��Dὤ�,�
���>ľl5���M����jL��K[�o��#��g&�      O�0��o����˿:1��-�y���6��z �����)�l�+��ͽ!�����&���˼_�k�q���l�X��� �ϳ�:o�;(&;�9;��B;�F;�|H;�I;e!I;5I;�I;�
I;qI;EI;��H;"�H;��H;"�H;��H;EI;qI;�
I;�I;5I;e!I;�I;�|H;�F;��B;�9;(&;o�;ϳ�:�� �l�X�q���_�k���˼��&�!����ͽ+�)�l������z ���6�-�y�:1���˿���o�0��      ����2���K[忭˿�T��蟉�s�R�����E۾̗����M�~�	������j��3�"d��ɆO���׻c�/��
�����:��	;$*;k;;�iC;�&G;�H;�I;
!I;�I;�I;�	I;�I;� I;I�H;��H;��H;��H;I�H;� I;�I;�	I;�I;�I;
!I;�I;�H;�&G;�iC;k;;$*;��	;���:�
��c�/���׻ɆO�"d���3���j����~�	���M�̗���E۾���s�R�蟉��T���˿K[�2���      �˿�<ƿjL��:1��蟉��>]���)��$���ճ���{���,�j��$��Q`I��J��-��4/�T,��˻ ��!69	3�:�;o.;0-=;n`D;�G;n�H;�I;? I;`I;SI;�I;�I;��H;��H;�H;d�H;�H;��H;��H;�I;�I;SI;`I;? I;�I;n�H;�G;n`D;0-=;o.;�;	3�:�!69˻ �T,��4/�-���J��Q`I�$��j�齞�,���{��ճ��$����)��>]�蟉�:1��jL���<ƿ      �o��벗����-�y�s�R���)�iv��>ľ�]����I�Tl�~��������&�߮Ҽ
�}�VB�"���������!:=)�:Vy;�3;ki?;�[E;��G;��H;tI;�I;�I;�I;|I;�I;�H;��H;c�H;��H;c�H;��H;�H;�I;|I;�I;�I;�I;tI;��H;��G;�[E;ki?;�3;Vy;=)�:��!:����"���VB�
�}�߮Ҽ��&����~���Tl���I��]���>ľiv���)�s�R�-�y����벗�      <�b��>]���M���6�����$���>ľq��q�Z�+�K9ݽW����L����0F��&�G�\�׻�;�u�Ǌ:�h;5O$;�7;x�A;IF;9BH;��H;�I;mI;wI;I;-I;�I;�H;��H;��H;�H;��H;��H;�H;�I;-I;I;wI;mI;�I;��H;9BH;IF;x�A;�7;5O$;�h;Ǌ:u칹;�\�׻&�G�0F�������L�W��K9ݽ+�q�Z�q���>ľ�$�������6���M��>]�      =\����l5��z ��E۾�ճ��]��q�Z�F?#����A����j�(��Pϼ��������Tnۺi3�9�2�:o�;y�,;��;;B�C;�G;Q�H;�
I;� I;�I;FI;.
I;�I;> I;�H;�H;��H;!�H;��H;�H;�H;> I;�I;.
I;FI;�I;� I;�
I;Q�H;�G;B�C;��;;y�,;o�;�2�:i3�9Tnۺ��������Pϼ(����j��A�����F?#�q�Z��]���ճ��E۾�z �l5����      +m־G�Ѿ�>ľ����̗����{���I�+����V���{�?�/�.���,��c=���һ�@�=� ���k:B�:#a;��3;@i?;v1E;��G;o�H;7I;wI;�I;�I;%I;�I;��H;��H;��H;��H;V�H;��H;��H;��H;��H;�I;%I;�I;�I;wI;7I;o�H;��G;v1E;@i?;��3;#a;B�:��k:=� ��@���һc=��,��.��?�/��{��V�����+���I���{�̗�������>ľG�Ѿ      ^���p��
��)�l���M���,�Tl�K9ݽ�A���{���5��J��;���T[�J?������Q���I�9�:��;9*;4�9;ijB;چF;�MH;��H;I;�I;�I;!I;I;@I;^�H;��H;��H;��H;i�H;��H;��H;��H;^�H;@I;I;!I;�I;�I;I;��H;�MH;چF;ijB;4�9;9*;��;�:�I�9�Q������J?��T[�;���J����5��{��A��K9ݽTl���,���M�)�l�
���p��      K�:��*7���,�+�~�	�j��~���W����j�?�/��J���I��&�k���c.������:Ǌ:�m�:';mq3;1�>;8�D;t�G;R�H;I;. I;�I;�I;�	I;�I;_�H;��H;��H;��H;��H;^�H;��H;��H;��H;��H;_�H;�I;�	I;�I;�I;. I;I;R�H;t�G;8�D;1�>;mq3;';�m�::Ǌ:����c.����&�k��I���J��?�/���j�W��~���j��~�	�+���,��*7�      �J���D��ͽ���$�������L�(��.��;��&�k����I����/��"/�'�>:���:�A;v�,;��:;=�B;�wF;�;H;��H;	I;�I;�I;AI;�I;�I;��H;s�H;4�H;n�H;��H;k�H;��H;n�H;4�H;s�H;��H;�I;�I;AI;�I;�I;	I;��H;�;H;�wF;=�B;��:;v�,;�A;���:'�>:�"/���/��I����&�k�;��.��(����L����$������ͽ�Dὼ��      &��"W��撐�!�����j�Q`I���&����Pϼ�,���T[����I��;��qk�i:g3�:� ; &;�6;� @;C1E;�G;��H;�I;�I;OI;I;�	I;:I;t�H;��H;�H;��H;^�H;��H;D�H;��H;^�H;��H;�H;��H;t�H;:I;�	I;I;OI;�I;�I;��H;�G;C1E;� @;�6; &;� ;g3�:i:�qk�;��I�����T[��,��Pϼ�����&�Q`I���j�!���撐�"W��      F�B�MR?��5���&��3��J��߮Ҽ0F����c=�J?�c.����/��qk����9�ճ:�;J!;l3;��=;��C;*�F;cH;��H;�I;I;�I;#I;�I;�I;C�H;��H;��H;|�H;?�H;|�H;3�H;|�H;?�H;|�H;��H;��H;C�H;�I;�I;#I;�I;I;�I;��H;cH;*�F;��C;��=;l3;J!;�;�ճ:���9�qk���/�c.��J?�c=���0F��߮Ҽ�J���3���&��5�MR?�      F��	}�<�ݼ��˼"d��-��
�}�&�G������һ�������"/�i:�ճ:"�;�a;â0;�<;��B;�HF;uH;,�H;�I;yI;I;8I;Y	I;�I;�H;/�H;T�H;�H;#�H;�H;r�H;5�H;r�H;�H;#�H;�H;T�H;/�H;�H;�I;Y	I;8I;I;yI;�I;,�H;uH;�HF;��B;�<;â0;�a;"�;�ճ:i:�"/���������һ���&�G�
�}�-��"d����˼<�ݼ	}�      �����8����_�k�ɆO�4/�VB�\�׻����@��Q����'�>:g3�:�;�a;��/;=;;J�A;��E;ɾG;��H;�	I;gI;I;�I;�I;�I;� I;��H;;�H;��H;��H;��H;�H;c�H;)�H;c�H;�H;��H;��H;��H;;�H;��H;� I;�I;�I;�I;I;gI;�	I;��H;ɾG;��E;J�A;=;;��/;�a;�;g3�:'�>:���Q���@����\�׻VB�4/�ɆO�_�k����8��      ������q
�q�����׻T,��"����;�Tnۺ=� ��I�9:Ǌ:���:� ;J!;â0;=;;̒A;�oE;|�G;ӍH;��H;�I;9I;ZI; I;�I;oI;��H;=�H;x�H;�H;�H;��H;��H;Z�H;1�H;Z�H;��H;��H;�H;�H;x�H;=�H;��H;oI;�I; I;ZI;9I;�I;��H;ӍH;|�G;�oE;̒A;=;;â0;J!;� ;���::Ǌ:�I�9=� �Tnۺ�;�"���T,����׻q����q
���      �/��s�����x�l�X�c�/�˻ �����u�i3�9��k:�:�m�:�A; &;l3;�<;J�A;�oE;hsG;�{H;-�H;,I;rI;BI;�I;h	I;�I;L�H;I�H;�H;��H;x�H;��H;��H;��H;l�H;\�H;l�H;��H;��H;��H;x�H;��H;�H;I�H;L�H;�I;h	I;�I;BI;rI;,I;-�H;�{H;hsG;�oE;J�A;�<;l3; &;�A;�m�:�:��k:i3�9u칌���˻ �c�/�l�X���x�s���      ��������wk��� ��
���!69��!:Ǌ:�2�:B�:��;';v�,;�6;��=;��B;��E;|�G;�{H;��H;zI;I;�I;WI;�
I;"I;� I;A�H;��H;4�H;��H;�H;��H;��H;��H;}�H;k�H;}�H;��H;��H;��H;�H;��H;4�H;��H;A�H;� I;"I;�
I;WI;�I;I;zI;��H;�{H;|�G;��E;��B;��=;�6;v�,;';��;B�:�2�:Ǌ:��!:�!69�
���� ��wk����      ��>:6�G:}�b:ϳ�:���:	3�:=)�:�h;o�;#a;9*;mq3;��:;� @;��C;�HF;ɾG;ӍH;-�H;zI;I;BI;9I;�I;I;UI;�H;��H;��H;o�H;B�H;��H;��H;��H;	�H;��H;y�H;��H;	�H;��H;��H;��H;B�H;o�H;��H;��H;�H;UI;I;�I;9I;BI;I;zI;-�H;ӍH;ɾG;�HF;��C;� @;��:;mq3;9*;#a;o�;�h;=)�:	3�:���:ϳ�:}�b:6�G:      �r�:���:�j�:o�;��	;�;Vy;5O$;y�,;��3;4�9;1�>;=�B;C1E;*�F;uH;��H;��H;,I;I;BI;�I;6I;�I;�I;��H;�H;F�H;��H;��H;��H;��H;��H;��H;)�H;��H;��H;��H;)�H;��H;��H;��H;��H;��H;��H;F�H;�H;��H;�I;�I;6I;�I;BI;I;,I;��H;��H;uH;*�F;C1E;=�B;1�>;4�9;��3;y�,;5O$;Vy;�;��	;o�;�j�:���:      do ; !;#;(&;$*;o.;�3;�7;��;;@i?;ijB;8�D;�wF;�G;cH;,�H;�	I;�I;rI;�I;9I;6I;�I;QI;4�H;��H;��H; �H;��H;�H;��H;x�H;��H;��H;E�H;�H;��H;�H;E�H;��H;��H;x�H;��H;�H;��H; �H;��H;��H;4�H;QI;�I;6I;9I;�I;rI;�I;�	I;,�H;cH;�G;�wF;8�D;ijB;@i?;��;;�7;�3;o.;$*;(&;#; !;      �I6;&�6;ږ7;�9;k;;0-=;ki?;x�A;B�C;v1E;چF;t�G;�;H;��H;��H;�I;gI;9I;BI;WI;�I;�I;QI;E�H;��H;��H;Y�H;$�H;0�H;��H;~�H;e�H;��H;�H;��H;]�H;:�H;]�H;��H;�H;��H;e�H;~�H;��H;0�H;$�H;Y�H;��H;��H;E�H;QI;�I;�I;WI;BI;9I;gI;�I;��H;��H;�;H;t�G;چF;v1E;B�C;x�A;ki?;0-=;k;;�9;ږ7;&�6;      DA;'kA;��A;��B;�iC;n`D;�[E;IF;�G;��G;�MH;R�H;��H;�I;�I;yI;I;ZI;�I;�
I;I;�I;4�H;��H;��H;w�H;-�H;@�H;��H;��H;`�H;t�H;��H;O�H;��H;��H;��H;��H;��H;O�H;��H;t�H;`�H;��H;��H;@�H;-�H;w�H;��H;��H;4�H;�I;I;�
I;�I;ZI;I;yI;�I;�I;��H;R�H;�MH;��G;�G;IF;�[E;n`D;�iC;��B;��A;'kA;      �HF;�XF;�F;�F;�&G;�G;��G;9BH;Q�H;o�H;��H;I;	I;�I;I;I;�I; I;h	I;"I;UI;��H;��H;��H;w�H;S�H;Z�H;��H;��H;i�H;X�H;��H;&�H;��H;@�H;"�H;�H;"�H;@�H;��H;&�H;��H;X�H;i�H;��H;��H;Z�H;S�H;w�H;��H;��H;��H;UI;"I;h	I; I;�I;I;I;�I;	I;I;��H;o�H;Q�H;9BH;��G;�G;�&G;�F;�F;�XF;      �MH;�SH;�cH;�|H;�H;n�H;��H;��H;�
I;7I;I;. I;�I;OI;�I;8I;�I;�I;�I;� I;�H;�H;��H;Y�H;-�H;Z�H;��H;��H;X�H;Z�H;��H;��H;d�H;��H;��H;��H;��H;��H;��H;��H;d�H;��H;��H;Z�H;X�H;��H;��H;Z�H;-�H;Y�H;��H;�H;�H;� I;�I;�I;�I;8I;�I;OI;�I;. I;I;7I;�
I;��H;��H;n�H;�H;�|H;�cH;�SH;      �H;s�H;�I;�I;�I;�I;tI;�I;� I;wI;�I;�I;�I;I;#I;Y	I;�I;oI;L�H;A�H;��H;F�H; �H;$�H;@�H;��H;��H;k�H;O�H;��H;��H;;�H;��H;{�H;9�H;
�H;�H;
�H;9�H;{�H;��H;;�H;��H;��H;O�H;k�H;��H;��H;@�H;$�H; �H;F�H;��H;A�H;L�H;oI;�I;Y	I;#I;I;�I;�I;�I;wI;� I;�I;tI;�I;�I;�I;�I;s�H;      !I;!I;\!I;e!I;
!I;? I;�I;mI;�I;�I;�I;�I;AI;�	I;�I;�I;� I;��H;I�H;��H;��H;��H;��H;0�H;��H;��H;X�H;O�H;��H;��H;/�H;��H;M�H;��H;��H;��H;��H;��H;��H;��H;M�H;��H;/�H;��H;��H;O�H;X�H;��H;��H;0�H;��H;��H;��H;��H;I�H;��H;� I;�I;�I;�	I;AI;�I;�I;�I;�I;mI;�I;? I;
!I;e!I;\!I;!I;      �I;�I;I;5I;�I;`I;�I;wI;FI;�I;!I;�	I;�I;:I;�I;�H;��H;=�H;�H;4�H;o�H;��H;�H;��H;��H;i�H;Z�H;��H;��H;�H;��H;C�H;��H;��H;f�H;I�H;9�H;I�H;f�H;��H;��H;C�H;��H;�H;��H;��H;Z�H;i�H;��H;��H;�H;��H;o�H;4�H;�H;=�H;��H;�H;�I;:I;�I;�	I;!I;�I;FI;wI;�I;`I;�I;5I;I;�I;      I;�I;oI;�I;�I;SI;�I;I;.
I;%I;I;�I;�I;t�H;C�H;/�H;;�H;x�H;��H;��H;B�H;��H;��H;~�H;`�H;X�H;��H;��H;/�H;��H;'�H;��H;v�H;<�H;	�H;��H;��H;��H;	�H;<�H;v�H;��H;'�H;��H;/�H;��H;��H;X�H;`�H;~�H;��H;��H;B�H;��H;��H;x�H;;�H;/�H;C�H;t�H;�I;�I;I;%I;.
I;I;�I;SI;�I;�I;oI;�I;      �I;�I;AI;�
I;�	I;�I;|I;-I;�I;�I;@I;_�H;��H;��H;��H;T�H;��H;�H;x�H;�H;��H;��H;x�H;e�H;t�H;��H;��H;;�H;��H;C�H;��H;R�H;!�H;��H;��H;��H;��H;��H;��H;��H;!�H;R�H;��H;C�H;��H;;�H;��H;��H;t�H;e�H;x�H;��H;��H;�H;x�H;�H;��H;T�H;��H;��H;��H;_�H;@I;�I;�I;-I;|I;�I;�	I;�
I;AI;�I;      mI;FI;�I;qI;�I;�I;�I;�I;> I;��H;^�H;��H;s�H;�H;��H;�H;��H;�H;��H;��H;��H;��H;��H;��H;��H;&�H;d�H;��H;M�H;��H;v�H;!�H;��H;��H;��H;m�H;f�H;m�H;��H;��H;��H;!�H;v�H;��H;M�H;��H;d�H;&�H;��H;��H;��H;��H;��H;��H;��H;�H;��H;�H;��H;�H;s�H;��H;^�H;��H;> I;�I;�I;�I;�I;qI;�I;FI;      I;�I;�I;EI;� I;��H;�H;�H;�H;��H;��H;��H;4�H;��H;|�H;#�H;��H;��H;��H;��H;��H;��H;��H;�H;O�H;��H;��H;{�H;��H;��H;<�H;��H;��H;n�H;V�H;I�H;9�H;I�H;V�H;n�H;��H;��H;<�H;��H;��H;{�H;��H;��H;O�H;�H;��H;��H;��H;��H;��H;��H;��H;#�H;|�H;��H;4�H;��H;��H;��H;�H;�H;�H;��H;� I;EI;�I;�I;      q�H;e�H; �H;��H;I�H;��H;��H;��H;�H;��H;��H;��H;n�H;^�H;?�H;�H;�H;��H;��H;��H;	�H;)�H;E�H;��H;��H;@�H;��H;9�H;��H;f�H;	�H;��H;��H;V�H;1�H;&�H;(�H;&�H;1�H;V�H;��H;��H;	�H;f�H;��H;9�H;��H;@�H;��H;��H;E�H;)�H;	�H;��H;��H;��H;�H;�H;?�H;^�H;n�H;��H;��H;��H;�H;��H;��H;��H;I�H;��H; �H;e�H;      ��H;��H;x�H;"�H;��H;�H;c�H;��H;��H;��H;��H;��H;��H;��H;|�H;r�H;c�H;Z�H;l�H;}�H;��H;��H;�H;]�H;��H;"�H;��H;
�H;��H;I�H;��H;��H;m�H;I�H;&�H;
�H;�H;
�H;&�H;I�H;m�H;��H;��H;I�H;��H;
�H;��H;"�H;��H;]�H;�H;��H;��H;}�H;l�H;Z�H;c�H;r�H;|�H;��H;��H;��H;��H;��H;��H;��H;c�H;�H;��H;"�H;x�H;��H;      *�H;�H;��H;��H;��H;d�H;��H;�H;!�H;V�H;i�H;^�H;k�H;D�H;3�H;5�H;)�H;1�H;\�H;k�H;y�H;��H;��H;:�H;��H;�H;��H;�H;��H;9�H;��H;��H;f�H;9�H;(�H;�H;�H;�H;(�H;9�H;f�H;��H;��H;9�H;��H;�H;��H;�H;��H;:�H;��H;��H;y�H;k�H;\�H;1�H;)�H;5�H;3�H;D�H;k�H;^�H;i�H;V�H;!�H;�H;��H;d�H;��H;��H;��H;�H;      ��H;��H;x�H;"�H;��H;�H;c�H;��H;��H;��H;��H;��H;��H;��H;|�H;r�H;c�H;Z�H;l�H;}�H;��H;��H;�H;]�H;��H;"�H;��H;
�H;��H;I�H;��H;��H;m�H;I�H;&�H;
�H;�H;
�H;&�H;I�H;m�H;��H;��H;I�H;��H;
�H;��H;"�H;��H;]�H;�H;��H;��H;}�H;l�H;Z�H;c�H;r�H;|�H;��H;��H;��H;��H;��H;��H;��H;c�H;�H;��H;"�H;x�H;��H;      q�H;e�H; �H;��H;I�H;��H;��H;��H;�H;��H;��H;��H;n�H;^�H;?�H;�H;�H;��H;��H;��H;	�H;)�H;E�H;��H;��H;@�H;��H;9�H;��H;f�H;	�H;��H;��H;V�H;1�H;&�H;(�H;&�H;1�H;V�H;��H;��H;	�H;f�H;��H;9�H;��H;@�H;��H;��H;E�H;)�H;	�H;��H;��H;��H;�H;�H;?�H;^�H;n�H;��H;��H;��H;�H;��H;��H;��H;I�H;��H; �H;e�H;      I;�I;�I;EI;� I;��H;�H;�H;�H;��H;��H;��H;4�H;��H;|�H;#�H;��H;��H;��H;��H;��H;��H;��H;�H;O�H;��H;��H;{�H;��H;��H;<�H;��H;��H;n�H;V�H;I�H;9�H;I�H;V�H;n�H;��H;��H;<�H;��H;��H;{�H;��H;��H;O�H;�H;��H;��H;��H;��H;��H;��H;��H;#�H;|�H;��H;4�H;��H;��H;��H;�H;�H;�H;��H;� I;EI;�I;�I;      mI;FI;�I;qI;�I;�I;�I;�I;> I;��H;^�H;��H;s�H;�H;��H;�H;��H;�H;��H;��H;��H;��H;��H;��H;��H;&�H;d�H;��H;M�H;��H;v�H;!�H;��H;��H;��H;m�H;f�H;m�H;��H;��H;��H;!�H;v�H;��H;M�H;��H;d�H;&�H;��H;��H;��H;��H;��H;��H;��H;�H;��H;�H;��H;�H;s�H;��H;^�H;��H;> I;�I;�I;�I;�I;qI;�I;FI;      �I;�I;AI;�
I;�	I;�I;|I;-I;�I;�I;@I;_�H;��H;��H;��H;T�H;��H;�H;x�H;�H;��H;��H;x�H;e�H;t�H;��H;��H;;�H;��H;C�H;��H;R�H;!�H;��H;��H;��H;��H;��H;��H;��H;!�H;R�H;��H;C�H;��H;;�H;��H;��H;t�H;e�H;x�H;��H;��H;�H;x�H;�H;��H;T�H;��H;��H;��H;_�H;@I;�I;�I;-I;|I;�I;�	I;�
I;AI;�I;      I;�I;oI;�I;�I;SI;�I;I;.
I;%I;I;�I;�I;t�H;C�H;/�H;;�H;x�H;��H;��H;B�H;��H;��H;~�H;`�H;X�H;��H;��H;/�H;��H;'�H;��H;v�H;<�H;	�H;��H;��H;��H;	�H;<�H;v�H;��H;'�H;��H;/�H;��H;��H;X�H;`�H;~�H;��H;��H;B�H;��H;��H;x�H;;�H;/�H;C�H;t�H;�I;�I;I;%I;.
I;I;�I;SI;�I;�I;oI;�I;      �I;�I;I;5I;�I;`I;�I;wI;FI;�I;!I;�	I;�I;:I;�I;�H;��H;=�H;�H;4�H;o�H;��H;�H;��H;��H;i�H;Z�H;��H;��H;�H;��H;C�H;��H;��H;f�H;I�H;9�H;I�H;f�H;��H;��H;C�H;��H;�H;��H;��H;Z�H;i�H;��H;��H;�H;��H;o�H;4�H;�H;=�H;��H;�H;�I;:I;�I;�	I;!I;�I;FI;wI;�I;`I;�I;5I;I;�I;      !I;!I;\!I;e!I;
!I;? I;�I;mI;�I;�I;�I;�I;AI;�	I;�I;�I;� I;��H;I�H;��H;��H;��H;��H;0�H;��H;��H;X�H;O�H;��H;��H;/�H;��H;M�H;��H;��H;��H;��H;��H;��H;��H;M�H;��H;/�H;��H;��H;O�H;X�H;��H;��H;0�H;��H;��H;��H;��H;I�H;��H;� I;�I;�I;�	I;AI;�I;�I;�I;�I;mI;�I;? I;
!I;e!I;\!I;!I;      �H;s�H;�I;�I;�I;�I;tI;�I;� I;wI;�I;�I;�I;I;#I;Y	I;�I;oI;L�H;A�H;��H;F�H; �H;$�H;@�H;��H;��H;k�H;O�H;��H;��H;;�H;��H;{�H;9�H;
�H;�H;
�H;9�H;{�H;��H;;�H;��H;��H;O�H;k�H;��H;��H;@�H;$�H; �H;F�H;��H;A�H;L�H;oI;�I;Y	I;#I;I;�I;�I;�I;wI;� I;�I;tI;�I;�I;�I;�I;s�H;      �MH;�SH;�cH;�|H;�H;n�H;��H;��H;�
I;7I;I;. I;�I;OI;�I;8I;�I;�I;�I;� I;�H;�H;��H;Y�H;-�H;Z�H;��H;��H;X�H;Z�H;��H;��H;d�H;��H;��H;��H;��H;��H;��H;��H;d�H;��H;��H;Z�H;X�H;��H;��H;Z�H;-�H;Y�H;��H;�H;�H;� I;�I;�I;�I;8I;�I;OI;�I;. I;I;7I;�
I;��H;��H;n�H;�H;�|H;�cH;�SH;      �HF;�XF;�F;�F;�&G;�G;��G;9BH;Q�H;o�H;��H;I;	I;�I;I;I;�I; I;h	I;"I;UI;��H;��H;��H;w�H;S�H;Z�H;��H;��H;i�H;X�H;��H;&�H;��H;@�H;"�H;�H;"�H;@�H;��H;&�H;��H;X�H;i�H;��H;��H;Z�H;S�H;w�H;��H;��H;��H;UI;"I;h	I; I;�I;I;I;�I;	I;I;��H;o�H;Q�H;9BH;��G;�G;�&G;�F;�F;�XF;      DA;'kA;��A;��B;�iC;n`D;�[E;IF;�G;��G;�MH;R�H;��H;�I;�I;yI;I;ZI;�I;�
I;I;�I;4�H;��H;��H;w�H;-�H;@�H;��H;��H;`�H;t�H;��H;O�H;��H;��H;��H;��H;��H;O�H;��H;t�H;`�H;��H;��H;@�H;-�H;w�H;��H;��H;4�H;�I;I;�
I;�I;ZI;I;yI;�I;�I;��H;R�H;�MH;��G;�G;IF;�[E;n`D;�iC;��B;��A;'kA;      �I6;&�6;ږ7;�9;k;;0-=;ki?;x�A;B�C;v1E;چF;t�G;�;H;��H;��H;�I;gI;9I;BI;WI;�I;�I;QI;E�H;��H;��H;Y�H;$�H;0�H;��H;~�H;e�H;��H;�H;��H;]�H;:�H;]�H;��H;�H;��H;e�H;~�H;��H;0�H;$�H;Y�H;��H;��H;E�H;QI;�I;�I;WI;BI;9I;gI;�I;��H;��H;�;H;t�G;چF;v1E;B�C;x�A;ki?;0-=;k;;�9;ږ7;&�6;      do ; !;#;(&;$*;o.;�3;�7;��;;@i?;ijB;8�D;�wF;�G;cH;,�H;�	I;�I;rI;�I;9I;6I;�I;QI;4�H;��H;��H; �H;��H;�H;��H;x�H;��H;��H;E�H;�H;��H;�H;E�H;��H;��H;x�H;��H;�H;��H; �H;��H;��H;4�H;QI;�I;6I;9I;�I;rI;�I;�	I;,�H;cH;�G;�wF;8�D;ijB;@i?;��;;�7;�3;o.;$*;(&;#; !;      �r�:���:�j�:o�;��	;�;Vy;5O$;y�,;��3;4�9;1�>;=�B;C1E;*�F;uH;��H;��H;,I;I;BI;�I;6I;�I;�I;��H;�H;F�H;��H;��H;��H;��H;��H;��H;)�H;��H;��H;��H;)�H;��H;��H;��H;��H;��H;��H;F�H;�H;��H;�I;�I;6I;�I;BI;I;,I;��H;��H;uH;*�F;C1E;=�B;1�>;4�9;��3;y�,;5O$;Vy;�;��	;o�;�j�:���:      ��>:6�G:}�b:ϳ�:���:	3�:=)�:�h;o�;#a;9*;mq3;��:;� @;��C;�HF;ɾG;ӍH;-�H;zI;I;BI;9I;�I;I;UI;�H;��H;��H;o�H;B�H;��H;��H;��H;	�H;��H;y�H;��H;	�H;��H;��H;��H;B�H;o�H;��H;��H;�H;UI;I;�I;9I;BI;I;zI;-�H;ӍH;ɾG;�HF;��C;� @;��:;mq3;9*;#a;o�;�h;=)�:	3�:���:ϳ�:}�b:6�G:      ��������wk��� ��
���!69��!:Ǌ:�2�:B�:��;';v�,;�6;��=;��B;��E;|�G;�{H;��H;zI;I;�I;WI;�
I;"I;� I;A�H;��H;4�H;��H;�H;��H;��H;��H;}�H;k�H;}�H;��H;��H;��H;�H;��H;4�H;��H;A�H;� I;"I;�
I;WI;�I;I;zI;��H;�{H;|�G;��E;��B;��=;�6;v�,;';��;B�:�2�:Ǌ:��!:�!69�
���� ��wk����      �/��s�����x�l�X�c�/�˻ �����u�i3�9��k:�:�m�:�A; &;l3;�<;J�A;�oE;hsG;�{H;-�H;,I;rI;BI;�I;h	I;�I;L�H;I�H;�H;��H;x�H;��H;��H;��H;l�H;\�H;l�H;��H;��H;��H;x�H;��H;�H;I�H;L�H;�I;h	I;�I;BI;rI;,I;-�H;�{H;hsG;�oE;J�A;�<;l3; &;�A;�m�:�:��k:i3�9u칌���˻ �c�/�l�X���x�s���      ������q
�q�����׻T,��"����;�Tnۺ=� ��I�9:Ǌ:���:� ;J!;â0;=;;̒A;�oE;|�G;ӍH;��H;�I;9I;ZI; I;�I;oI;��H;=�H;x�H;�H;�H;��H;��H;Z�H;1�H;Z�H;��H;��H;�H;�H;x�H;=�H;��H;oI;�I; I;ZI;9I;�I;��H;ӍH;|�G;�oE;̒A;=;;â0;J!;� ;���::Ǌ:�I�9=� �Tnۺ�;�"���T,����׻q����q
���      �����8����_�k�ɆO�4/�VB�\�׻����@��Q����'�>:g3�:�;�a;��/;=;;J�A;��E;ɾG;��H;�	I;gI;I;�I;�I;�I;� I;��H;;�H;��H;��H;��H;�H;c�H;)�H;c�H;�H;��H;��H;��H;;�H;��H;� I;�I;�I;�I;I;gI;�	I;��H;ɾG;��E;J�A;=;;��/;�a;�;g3�:'�>:���Q���@����\�׻VB�4/�ɆO�_�k����8��      F��	}�<�ݼ��˼"d��-��
�}�&�G������һ�������"/�i:�ճ:"�;�a;â0;�<;��B;�HF;uH;,�H;�I;yI;I;8I;Y	I;�I;�H;/�H;T�H;�H;#�H;�H;r�H;5�H;r�H;�H;#�H;�H;T�H;/�H;�H;�I;Y	I;8I;I;yI;�I;,�H;uH;�HF;��B;�<;â0;�a;"�;�ճ:i:�"/���������һ���&�G�
�}�-��"d����˼<�ݼ	}�      F�B�MR?��5���&��3��J��߮Ҽ0F����c=�J?�c.����/��qk����9�ճ:�;J!;l3;��=;��C;*�F;cH;��H;�I;I;�I;#I;�I;�I;C�H;��H;��H;|�H;?�H;|�H;3�H;|�H;?�H;|�H;��H;��H;C�H;�I;�I;#I;�I;I;�I;��H;cH;*�F;��C;��=;l3;J!;�;�ճ:���9�qk���/�c.��J?�c=���0F��߮Ҽ�J���3���&��5�MR?�      &��"W��撐�!�����j�Q`I���&����Pϼ�,���T[����I��;��qk�i:g3�:� ; &;�6;� @;C1E;�G;��H;�I;�I;OI;I;�	I;:I;t�H;��H;�H;��H;^�H;��H;D�H;��H;^�H;��H;�H;��H;t�H;:I;�	I;I;OI;�I;�I;��H;�G;C1E;� @;�6; &;� ;g3�:i:�qk�;��I�����T[��,��Pϼ�����&�Q`I���j�!���撐�"W��      �J���D��ͽ���$�������L�(��.��;��&�k����I����/��"/�'�>:���:�A;v�,;��:;=�B;�wF;�;H;��H;	I;�I;�I;AI;�I;�I;��H;s�H;4�H;n�H;��H;k�H;��H;n�H;4�H;s�H;��H;�I;�I;AI;�I;�I;	I;��H;�;H;�wF;=�B;��:;v�,;�A;���:'�>:�"/���/��I����&�k�;��.��(����L����$������ͽ�Dὼ��      K�:��*7���,�+�~�	�j��~���W����j�?�/��J���I��&�k���c.������:Ǌ:�m�:';mq3;1�>;8�D;t�G;R�H;I;. I;�I;�I;�	I;�I;_�H;��H;��H;��H;��H;^�H;��H;��H;��H;��H;_�H;�I;�	I;�I;�I;. I;I;R�H;t�G;8�D;1�>;mq3;';�m�::Ǌ:����c.����&�k��I���J��?�/���j�W��~���j��~�	�+���,��*7�      ^���p��
��)�l���M���,�Tl�K9ݽ�A���{���5��J��;���T[�J?������Q���I�9�:��;9*;4�9;ijB;چF;�MH;��H;I;�I;�I;!I;I;@I;^�H;��H;��H;��H;i�H;��H;��H;��H;^�H;@I;I;!I;�I;�I;I;��H;�MH;چF;ijB;4�9;9*;��;�:�I�9�Q������J?��T[�;���J����5��{��A��K9ݽTl���,���M�)�l�
���p��      +m־G�Ѿ�>ľ����̗����{���I�+����V���{�?�/�.���,��c=���һ�@�=� ���k:B�:#a;��3;@i?;v1E;��G;o�H;7I;wI;�I;�I;%I;�I;��H;��H;��H;��H;V�H;��H;��H;��H;��H;�I;%I;�I;�I;wI;7I;o�H;��G;v1E;@i?;��3;#a;B�:��k:=� ��@���һc=��,��.��?�/��{��V�����+���I���{�̗�������>ľG�Ѿ      =\����l5��z ��E۾�ճ��]��q�Z�F?#����A����j�(��Pϼ��������Tnۺi3�9�2�:o�;y�,;��;;B�C;�G;Q�H;�
I;� I;�I;FI;.
I;�I;> I;�H;�H;��H;!�H;��H;�H;�H;> I;�I;.
I;FI;�I;� I;�
I;Q�H;�G;B�C;��;;y�,;o�;�2�:i3�9Tnۺ��������Pϼ(����j��A�����F?#�q�Z��]���ճ��E۾�z �l5����      <�b��>]���M���6�����$���>ľq��q�Z�+�K9ݽW����L����0F��&�G�\�׻�;�u�Ǌ:�h;5O$;�7;x�A;IF;9BH;��H;�I;mI;wI;I;-I;�I;�H;��H;��H;�H;��H;��H;�H;�I;-I;I;wI;mI;�I;��H;9BH;IF;x�A;�7;5O$;�h;Ǌ:u칹;�\�׻&�G�0F�������L�W��K9ݽ+�q�Z�q���>ľ�$�������6���M��>]�      �o��벗����-�y�s�R���)�iv��>ľ�]����I�Tl�~��������&�߮Ҽ
�}�VB�"���������!:=)�:Vy;�3;ki?;�[E;��G;��H;tI;�I;�I;�I;|I;�I;�H;��H;c�H;��H;c�H;��H;�H;�I;|I;�I;�I;�I;tI;��H;��G;�[E;ki?;�3;Vy;=)�:��!:����"���VB�
�}�߮Ҽ��&����~���Tl���I��]���>ľiv���)�s�R�-�y����벗�      �˿�<ƿjL��:1��蟉��>]���)��$���ճ���{���,�j��$��Q`I��J��-��4/�T,��˻ ��!69	3�:�;o.;0-=;n`D;�G;n�H;�I;? I;`I;SI;�I;�I;��H;��H;�H;d�H;�H;��H;��H;�I;�I;SI;`I;? I;�I;n�H;�G;n`D;0-=;o.;�;	3�:�!69˻ �T,��4/�-���J��Q`I�$��j�齞�,���{��ճ��$����)��>]�蟉�:1��jL���<ƿ      ����2���K[忭˿�T��蟉�s�R�����E۾̗����M�~�	������j��3�"d��ɆO���׻c�/��
�����:��	;$*;k;;�iC;�&G;�H;�I;
!I;�I;�I;�	I;�I;� I;I�H;��H;��H;��H;I�H;� I;�I;�	I;�I;�I;
!I;�I;�H;�&G;�iC;k;;$*;��	;���:�
��c�/���׻ɆO�"d���3���j����~�	���M�̗���E۾���s�R�蟉��T���˿K[�2���      O�0��o����˿:1��-�y���6��z �����)�l�+��ͽ!�����&���˼_�k�q���l�X��� �ϳ�:o�;(&;�9;��B;�F;�|H;�I;e!I;5I;�I;�
I;qI;EI;��H;"�H;��H;"�H;��H;EI;qI;�
I;�I;5I;e!I;�I;�|H;�F;��B;�9;(&;o�;ϳ�:�� �l�X�q���_�k���˼��&�!����ͽ+�)�l������z ���6�-�y�:1���˿���o�0��      ��*��g&��#�o�K[�jL�������M�l5��>ľ
����,��D�撐��5�<�ݼ���q
���x��wk�}�b:�j�:#;ږ7;��A;�F;�cH;�I;\!I;I;oI;AI;�I;�I; �H;x�H;��H;x�H; �H;�I;�I;AI;oI;I;\!I;�I;�cH;�F;��A;ږ7;#;�j�:}�b:�wk���x��q
���<�ݼ�5�撐��Dὤ�,�
���>ľl5���M����jL��K[�o��#��g&�      ��8��4��g&�0��2����<ƿ벗��>]����G�Ѿ�p���*7����"W��MR?�	}鼀8����s������6�G:���: !;&�6;'kA;�XF;�SH;s�H;!I;�I;�I;�I;FI;�I;e�H;��H;�H;��H;e�H;�I;FI;�I;�I;�I;!I;s�H;�SH;�XF;'kA;&�6; !;���:6�G:���s������8��	}�MR?�"W�����*7��p��G�Ѿ����>]�벗��<ƿ2���0���g&��4�      ���$������꿥�ſ�ޞ�3s��2�/����� j���nHͽ������'�B<ͼ��n������Q^�0.�車:�V;�R%;~n8;��A;mCF;�H;��H;��H;��H;L�H;>�H;C�H;��H;��H;��H;+�H;��H;��H;��H;C�H;>�H;L�H;��H;��H;��H;�H;mCF;��A;~n8;�R%;�V;車:0.��Q^�������n�B<ͼ��'�����nHͽ�� j���/����2�3s��ޞ���ſ������$�      $��������~�����cm�L�-�����Fh��Ide�-�̪ɽ�v��#�$���ɼ�mj�o����X�9��lĆ:�w;i�%;L�8;~B;zQF;H;4�H;U�H;�H;p�H;B�H;5�H;��H;��H;��H;$�H;��H;��H;��H;5�H;B�H;p�H;�H;U�H;4�H;H;zQF;~B;L�8;i�%;�w;lĆ:9���X�o����mj���ɼ#�$��v��̪ɽ-�Ide�Fh������L�-�cm����~���忖����      ������{���ԿBw�����/�\��"����b��M0X�}���;����w����������]�X��VF�3��nȒ:0�;^�';׎9;1oB;�yF;� H;��H;7�H;�H;��H;F�H;:�H;��H;��H;��H;�H;��H;��H;��H;:�H;F�H;��H;�H;7�H;��H;� H;�yF;1oB;׎9;^�';0�;nȒ:3��VF�X�黼�]����������w��;��}��M0X�b������"�/�\����Bw���Կ{�𿖏�      ������Կp���ޞ�RF�]�C�$E��;�I��sD�|�"��]�c�y��֯���J�P�ѻ]�)���K����:P�
;M*;��:;�C;�F;�7H;Z�H;��H;w�H;��H;>�H;9�H;��H;��H;��H;��H;��H;��H;��H;9�H;>�H;��H;w�H;��H;Z�H;�7H;�F;�C;��:;M*;P�
;���:��K�]�)�P�ѻ��J��֯�y�]�c�"��|�sD��I���;$E�]�C�RF��ޞ�p���Կ��      ��ſ~��Bw���ޞ�|���3�W�,�%�����^ɰ��|x�\{+�ű����J��  �Ҷ��n�1�f����+�
9p�:�;4�-;��<;��C;�G;�SH;Q�H;��H;��H;��H;V�H;2�H;��H;��H;��H;��H;��H;��H;��H;2�H;V�H;��H;��H;��H;Q�H;�SH;�G;��C;��<;4�-;�;p�:
9�+�f���n�1�Ҷ���  ��J���ű�\{+��|x�^ɰ�����,�%�3�W�|����ޞ�Bw��~��      �ޞ�������RF�3�W�M�-���4Kɾ�G����O�z��ƽ����Ȅ-���ۼㄼL4�[ǐ�-ж��Z:m��:�;ʕ1;
c>;{�D;�[G;KrH;��H;i�H;e�H;'�H;u�H;(�H;h�H;��H;|�H;��H;|�H;��H;h�H;(�H;u�H;'�H;e�H;i�H;��H;KrH;�[G;{�D;
c>;ʕ1;�;m��:�Z:-ж�[ǐ�L4�ㄼ��ۼȄ-�����ƽz����O��G��4Kɾ��M�-�3�W�RF�������      3s�cm�/�\�]�C�,�%����TҾa����i��C(����UP����[�x������Y�l���X���<���k:���:)� ;�5;ZQ@;otE;�G;9�H;L�H;��H;�H;I�H;l�H;$�H;b�H;s�H;W�H;��H;W�H;s�H;b�H;$�H;l�H;I�H;�H;��H;L�H;9�H;�G;otE;ZQ@;�5;)� ;���:��k:��<��X�l����Y����x���[�UP����콡C(���i�a���TҾ��,�%�]�C�/�\�cm�      �2�L�-��"�$E�����4Kɾa��w�s�.�5�y�k㻽�v��z0��;��+��-�*�S����6�YjS��K�:��	;��(;5�9;�.B;CF;YH;ԪH;��H;��H;��H;w�H;��H;�H;/�H;C�H;<�H;Y�H;<�H;C�H;/�H;�H;��H;w�H;��H;��H;��H;ԪH;YH;CF;�.B;5�9;��(;��	;�K�:YjS��6�S���-�*��+���;�z0��v��k㻽y�.�5�w�s�a��4Kɾ����$E��"�L�-�      /�����������;^ɰ��G����i�.�5��	�ĪɽR����J�p���沼��]�J���V
x��
��}k:4��:v;��/;�,=;��C;M�F;#HH;��H;'�H;��H;#�H;��H;��H;��H;�H;�H;�H;#�H;�H;�H;�H;��H;��H;��H;#�H;��H;'�H;��H;#HH;M�F;��C;�,=;��/;v;4��:}k:�
��V
x�J�����]��沼p���J�R���Īɽ�	�.�5���i��G��^ɰ��;��徨���      ��Fh��b���I���|x���O��C(�y�Īɽ����JDX�D��'<ͼㄼ�X!�t��iX��K����:�x;7�#;#H6;HQ@;�OE;��G;��H;��H;1�H;��H;��H;��H;v�H;��H;��H;��H;��H;��H;��H;��H;��H;��H;v�H;��H;��H;��H;1�H;��H;��H;��G;�OE;HQ@;#H6;7�#;�x;���:�K�iX�t���X!�ㄼ'<ͼD��JDX�����Īɽy��C(���O��|x��I��b��Fh��       j�Ide�M0X�sD�\{+�z�����k㻽R���JDX������ۼо����;�>ۻ�X���y�:<":H��:��;��-;��;;�B;�yF;�H;��H;{�H;&�H;��H;��H;��H;m�H;��H;��H;��H;��H;z�H;��H;��H;��H;��H;m�H;��H;��H;��H;&�H;{�H;��H;�H;�yF;�B;��;;��-;��;H��::<":��y��X�>ۻ��;�о����ۼ���JDX�R���k㻽���z��\{+�sD�M0X�Ide�      ��-�}��|�ű�ƽUP���v���J�D����ۼ��v�J������+���sѺ!
9eL�:�;�$;#�5;�?;��D;j[G;eH;��H;��H;��H;��H;!�H;��H;T�H;n�H;Y�H;T�H;a�H;7�H;a�H;T�H;Y�H;n�H;T�H;��H;!�H;��H;��H;��H;��H;eH;j[G;��D;�?;#�5;�$;�;eL�:!
9�sѺ�+������v�J�����ۼD���J��v��UP��ƽű�|�}��-�      nHͽ̪ɽ�;��"����������[�z0�p��'<ͼо��v�J���k��+��(����:�`�:|�;
�/;�K<; C;9lF;��G;�H;
�H;�H;�H;A�H;T�H;��H;%�H;/�H;�H;�H;�H;��H;�H;�H;�H;/�H;%�H;��H;T�H;A�H;�H;�H;
�H;�H;��G;9lF; C;�K<;
�/;|�;�`�:���:�(�+�k����v�J�о��'<ͼp��z0���[�������"���;��̪ɽ      �����v����w�]�c��J�Ȅ-�x��;缈沼ㄼ��;�����k��66�k��J<Q:գ�:�h;M*;��8;��@;�OE;�tG;DhH;��H;��H;�H;"�H;��H;y�H;��H;��H;��H;��H;��H;��H;��H;��H;��H;��H;��H;��H;��H;y�H;��H;"�H;�H;��H;��H;DhH;�tG;�OE;��@;��8;M*;�h;գ�:J<Q:k��66�k��������;�ㄼ�沼�;�x�Ȅ-��J�]�c���w��v��      ��'�#�$����y��  ���ۼ����+����]��X!�>ۻ�+��+�k���>:[��:?�;Z�%;�5;��>;�'D;�F;� H;8�H;[�H;��H;��H;��H;��H;k�H;��H;��H;��H;��H;g�H;J�H;m�H;J�H;g�H;��H;��H;��H;��H;k�H;��H;��H;��H;��H;[�H;8�H;� H;�F;�'D;��>;�5;Z�%;?�;[��:�>:k��+��+��>ۻ�X!���]��+�������ۼ�  �y����#�$�      B<ͼ��ɼ�����֯�Ҷ��ㄼ��Y�-�*�J���t���X��sѺ�(�J<Q:[��:��
;u�#;��3;�b=;#C;3CF;�G;�H;��H;�H;8�H;��H;W�H;!�H;d�H;��H;b�H;5�H;O�H;	�H;��H;�H;��H;	�H;O�H;5�H;b�H;��H;d�H;!�H;W�H;��H;8�H;�H;��H;�H;�G;3CF;#C;�b=;��3;u�#;��
;[��:J<Q:�(��sѺ�X�t��J���-�*���Y�ㄼҶ���֯�������ɼ      ��n��mj���]���J�n�1�L4�l��S���V
x�iX���y�!
9���:գ�:?�;u�#;v�2;�<;�oB;7�E;��G;�dH;��H;8�H;��H;��H;��H;��H;9�H;F�H;7�H;�H;��H;��H;��H;��H;��H;��H;��H;��H;��H;�H;7�H;F�H;9�H;��H;��H;��H;��H;8�H;��H;�dH;��G;7�E;�oB;�<;v�2;u�#;?�;գ�:���:!
9��y�iX�V
x�S���l��L4�n�1���J���]��mj�      ����o���X��P�ѻf���[ǐ��X��6��
���K�:<":eL�:�`�:�h;Z�%;��3;�<;X/B;��E;�[G;�GH;M�H;��H;a�H;�H;7�H;=�H;��H;�H;�H;��H;��H;��H;]�H;O�H;K�H;'�H;K�H;O�H;]�H;��H;��H;��H;�H;�H;��H;=�H;7�H;�H;a�H;��H;M�H;�GH;�[G;��E;X/B;�<;��3;Z�%;�h;�`�:eL�::<":�K��
���6��X�[ǐ�f���P�ѻX��o���      �Q^��X�VF�]�)��+�-ж���<�YjS�}k:���:H��:�;|�;M*;�5;�b=;�oB;��E;�IG;\7H;s�H;��H;�H;,�H;��H;��H;��H;��H;��H;��H;��H;t�H;P�H;��H;��H;��H;��H;��H;��H;��H;P�H;t�H;��H;��H;��H;��H;��H;��H;��H;,�H;�H;��H;s�H;\7H;�IG;��E;�oB;�b=;�5;M*;|�;�;H��:���:}k:YjS���<�-ж��+�]�)�VF��X�      0.�9��3�깩�K�
9�Z:��k:�K�:4��:�x;��;�$;
�/;��8;��>;#C;7�E;�[G;\7H;̤H;�H;&�H;��H;5�H;��H;P�H;��H;��H;��H;y�H;5�H;�H;��H;��H;��H;��H;t�H;��H;��H;��H;��H;�H;5�H;y�H;��H;��H;��H;P�H;��H;5�H;��H;&�H;�H;̤H;\7H;�[G;7�E;#C;��>;��8;
�/;�$;��;�x;4��:�K�:��k:�Z:
9��K�3��9��      車:lĆ:nȒ:���:p�:m��:���:��	;v;7�#;��-;#�5;�K<;��@;�'D;3CF;��G;�GH;s�H;�H;��H;O�H;��H;\�H;"�H;��H;��H;��H;[�H;�H;��H;��H;m�H;[�H;)�H;�H;�H;�H;)�H;[�H;m�H;��H;��H;�H;[�H;��H;��H;��H;"�H;\�H;��H;O�H;��H;�H;s�H;�GH;��G;3CF;�'D;��@;�K<;#�5;��-;7�#;v;��	;���:m��:p�:���:nȒ:lĆ:      �V;�w;0�;P�
;�;�;)� ;��(;��/;#H6;��;;�?; C;�OE;�F;�G;�dH;M�H;��H;&�H;O�H;��H;0�H;��H;e�H;~�H;��H;a�H;��H;��H;��H;A�H;�H;�H;��H;��H;��H;��H;��H;�H;�H;A�H;��H;��H;��H;a�H;��H;~�H;e�H;��H;0�H;��H;O�H;&�H;��H;M�H;�dH;�G;�F;�OE; C;�?;��;;#H6;��/;��(;)� ;�;�;P�
;0�;�w;      �R%;i�%;^�';M*;4�-;ʕ1;�5;5�9;�,=;HQ@;�B;��D;9lF;�tG;� H;�H;��H;��H;�H;��H;��H;0�H;�H;a�H;��H;r�H;4�H;��H;��H;��H;�H;��H;��H;��H;|�H;e�H;L�H;e�H;|�H;��H;��H;��H;�H;��H;��H;��H;4�H;r�H;��H;a�H;�H;0�H;��H;��H;�H;��H;��H;�H;� H;�tG;9lF;��D;�B;HQ@;�,=;5�9;�5;ʕ1;4�-;M*;^�';i�%;      ~n8;L�8;׎9;��:;��<;
c>;ZQ@;�.B;��C;�OE;�yF;j[G;��G;DhH;8�H;��H;8�H;a�H;,�H;5�H;\�H;��H;a�H;j�H;i�H;D�H;��H;��H;e�H;	�H;��H;��H;Y�H;(�H;!�H;�H;��H;�H;!�H;(�H;Y�H;��H;��H;	�H;e�H;��H;��H;D�H;i�H;j�H;a�H;��H;\�H;5�H;,�H;a�H;8�H;��H;8�H;DhH;��G;j[G;�yF;�OE;��C;�.B;ZQ@;
c>;��<;��:;׎9;L�8;      ��A;~B;1oB;�C;��C;{�D;otE;CF;M�F;��G;�H;eH;�H;��H;[�H;�H;��H;�H;��H;��H;"�H;e�H;��H;i�H;-�H;��H;��H;h�H;��H;��H;r�H;@�H;
�H;��H;��H;��H;��H;��H;��H;��H;
�H;@�H;r�H;��H;��H;h�H;��H;��H;-�H;i�H;��H;e�H;"�H;��H;��H;�H;��H;�H;[�H;��H;�H;eH;�H;��G;M�F;CF;otE;{�D;��C;�C;1oB;~B;      mCF;zQF;�yF;�F;�G;�[G;�G;YH;#HH;��H;��H;��H;
�H;��H;��H;8�H;��H;7�H;��H;P�H;��H;~�H;r�H;D�H;��H;��H;_�H;��H;��H;`�H;�H;��H;��H;��H;o�H;\�H;n�H;\�H;o�H;��H;��H;��H;�H;`�H;��H;��H;_�H;��H;��H;D�H;r�H;~�H;��H;P�H;��H;7�H;��H;8�H;��H;��H;
�H;��H;��H;��H;#HH;YH;�G;�[G;�G;�F;�yF;zQF;      �H;H;� H;�7H;�SH;KrH;9�H;ԪH;��H;��H;{�H;��H;�H;�H;��H;��H;��H;=�H;��H;��H;��H;��H;4�H;��H;��H;_�H;��H;��H;H�H;�H;��H;��H;b�H;C�H;(�H;�H;�H;�H;(�H;C�H;b�H;��H;��H;�H;H�H;��H;��H;_�H;��H;��H;4�H;��H;��H;��H;��H;=�H;��H;��H;��H;�H;�H;��H;{�H;��H;��H;ԪH;9�H;KrH;�SH;�7H;� H;H;      ��H;4�H;��H;Z�H;Q�H;��H;L�H;��H;'�H;1�H;&�H;��H;�H;"�H;��H;W�H;��H;��H;��H;��H;��H;a�H;��H;��H;h�H;��H;��H;W�H;�H;��H;u�H;F�H; �H;��H;��H;��H;��H;��H;��H;��H; �H;F�H;u�H;��H;�H;W�H;��H;��H;h�H;��H;��H;a�H;��H;��H;��H;��H;��H;W�H;��H;"�H;�H;��H;&�H;1�H;'�H;��H;L�H;��H;Q�H;Z�H;��H;4�H;      ��H;U�H;7�H;��H;��H;i�H;��H;��H;��H;��H;��H;��H;A�H;��H;��H;!�H;9�H;�H;��H;��H;[�H;��H;��H;e�H;��H;��H;H�H;�H;��H;k�H;7�H;��H;��H;��H;��H;��H;�H;��H;��H;��H;��H;��H;7�H;k�H;��H;�H;H�H;��H;��H;e�H;��H;��H;[�H;��H;��H;�H;9�H;!�H;��H;��H;A�H;��H;��H;��H;��H;��H;��H;i�H;��H;��H;7�H;U�H;      ��H;�H;�H;w�H;��H;e�H;�H;��H;#�H;��H;��H;!�H;T�H;y�H;k�H;d�H;F�H;�H;��H;y�H;�H;��H;��H;	�H;��H;`�H;�H;��H;k�H;-�H;��H;��H;��H;��H;c�H;K�H;A�H;K�H;c�H;��H;��H;��H;��H;-�H;k�H;��H;�H;`�H;��H;	�H;��H;��H;�H;y�H;��H;�H;F�H;d�H;k�H;y�H;T�H;!�H;��H;��H;#�H;��H;�H;e�H;��H;w�H;�H;�H;      L�H;p�H;��H;��H;��H;'�H;I�H;w�H;��H;��H;��H;��H;��H;��H;��H;��H;7�H;��H;��H;5�H;��H;��H;�H;��H;r�H;�H;��H;u�H;7�H;��H;��H;��H;w�H;?�H;�H;'�H;(�H;'�H;�H;?�H;w�H;��H;��H;��H;7�H;u�H;��H;�H;r�H;��H;�H;��H;��H;5�H;��H;��H;7�H;��H;��H;��H;��H;��H;��H;��H;��H;w�H;I�H;'�H;��H;��H;��H;p�H;      >�H;B�H;F�H;>�H;V�H;u�H;l�H;��H;��H;v�H;m�H;T�H;%�H;��H;��H;b�H;�H;��H;t�H;�H;��H;A�H;��H;��H;@�H;��H;��H;F�H;��H;��H;��H;_�H;A�H;�H;��H;��H;��H;��H;��H;�H;A�H;_�H;��H;��H;��H;F�H;��H;��H;@�H;��H;��H;A�H;��H;�H;t�H;��H;�H;b�H;��H;��H;%�H;T�H;m�H;v�H;��H;��H;l�H;u�H;V�H;>�H;F�H;B�H;      C�H;5�H;:�H;9�H;2�H;(�H;$�H;�H;��H;��H;��H;n�H;/�H;��H;��H;5�H;��H;��H;P�H;��H;m�H;�H;��H;Y�H;
�H;��H;b�H; �H;��H;��H;w�H;A�H;��H;��H;��H;��H;��H;��H;��H;��H;��H;A�H;w�H;��H;��H; �H;b�H;��H;
�H;Y�H;��H;�H;m�H;��H;P�H;��H;��H;5�H;��H;��H;/�H;n�H;��H;��H;��H;�H;$�H;(�H;2�H;9�H;:�H;5�H;      ��H;��H;��H;��H;��H;h�H;b�H;/�H;�H;��H;��H;Y�H;�H;��H;��H;O�H;��H;]�H;��H;��H;[�H;�H;��H;(�H;��H;��H;C�H;��H;��H;��H;?�H;�H;��H;��H;��H;��H;��H;��H;��H;��H;��H;�H;?�H;��H;��H;��H;C�H;��H;��H;(�H;��H;�H;[�H;��H;��H;]�H;��H;O�H;��H;��H;�H;Y�H;��H;��H;�H;/�H;b�H;h�H;��H;��H;��H;��H;      ��H;��H;��H;��H;��H;��H;s�H;C�H;�H;��H;��H;T�H;�H;��H;g�H;	�H;��H;O�H;��H;��H;)�H;��H;|�H;!�H;��H;o�H;(�H;��H;��H;c�H;�H;��H;��H;��H;��H;��H;��H;��H;��H;��H;��H;��H;�H;c�H;��H;��H;(�H;o�H;��H;!�H;|�H;��H;)�H;��H;��H;O�H;��H;	�H;g�H;��H;�H;T�H;��H;��H;�H;C�H;s�H;��H;��H;��H;��H;��H;      ��H;��H;��H;��H;��H;|�H;W�H;<�H;�H;��H;��H;a�H;�H;��H;J�H;��H;��H;K�H;��H;��H;�H;��H;e�H;�H;��H;\�H;�H;��H;��H;K�H;'�H;��H;��H;��H;��H;��H;��H;��H;��H;��H;��H;��H;'�H;K�H;��H;��H;�H;\�H;��H;�H;e�H;��H;�H;��H;��H;K�H;��H;��H;J�H;��H;�H;a�H;��H;��H;�H;<�H;W�H;|�H;��H;��H;��H;��H;      +�H;$�H;�H;��H;��H;��H;��H;Y�H;#�H;��H;z�H;7�H;��H;��H;m�H;�H;��H;'�H;��H;t�H;�H;��H;L�H;��H;��H;n�H;�H;��H;�H;A�H;(�H;��H;��H;��H;��H;��H;~�H;��H;��H;��H;��H;��H;(�H;A�H;�H;��H;�H;n�H;��H;��H;L�H;��H;�H;t�H;��H;'�H;��H;�H;m�H;��H;��H;7�H;z�H;��H;#�H;Y�H;��H;��H;��H;��H;�H;$�H;      ��H;��H;��H;��H;��H;|�H;W�H;<�H;�H;��H;��H;a�H;�H;��H;J�H;��H;��H;K�H;��H;��H;�H;��H;e�H;�H;��H;\�H;�H;��H;��H;K�H;'�H;��H;��H;��H;��H;��H;��H;��H;��H;��H;��H;��H;'�H;K�H;��H;��H;�H;\�H;��H;�H;e�H;��H;�H;��H;��H;K�H;��H;��H;J�H;��H;�H;a�H;��H;��H;�H;<�H;W�H;|�H;��H;��H;��H;��H;      ��H;��H;��H;��H;��H;��H;s�H;C�H;�H;��H;��H;T�H;�H;��H;g�H;	�H;��H;O�H;��H;��H;)�H;��H;|�H;!�H;��H;o�H;(�H;��H;��H;c�H;�H;��H;��H;��H;��H;��H;��H;��H;��H;��H;��H;��H;�H;c�H;��H;��H;(�H;o�H;��H;!�H;|�H;��H;)�H;��H;��H;O�H;��H;	�H;g�H;��H;�H;T�H;��H;��H;�H;C�H;s�H;��H;��H;��H;��H;��H;      ��H;��H;��H;��H;��H;h�H;b�H;/�H;�H;��H;��H;Y�H;�H;��H;��H;O�H;��H;]�H;��H;��H;[�H;�H;��H;(�H;��H;��H;C�H;��H;��H;��H;?�H;�H;��H;��H;��H;��H;��H;��H;��H;��H;��H;�H;?�H;��H;��H;��H;C�H;��H;��H;(�H;��H;�H;[�H;��H;��H;]�H;��H;O�H;��H;��H;�H;Y�H;��H;��H;�H;/�H;b�H;h�H;��H;��H;��H;��H;      C�H;5�H;:�H;9�H;2�H;(�H;$�H;�H;��H;��H;��H;n�H;/�H;��H;��H;5�H;��H;��H;P�H;��H;m�H;�H;��H;Y�H;
�H;��H;b�H; �H;��H;��H;w�H;A�H;��H;��H;��H;��H;��H;��H;��H;��H;��H;A�H;w�H;��H;��H; �H;b�H;��H;
�H;Y�H;��H;�H;m�H;��H;P�H;��H;��H;5�H;��H;��H;/�H;n�H;��H;��H;��H;�H;$�H;(�H;2�H;9�H;:�H;5�H;      >�H;B�H;F�H;>�H;V�H;u�H;l�H;��H;��H;v�H;m�H;T�H;%�H;��H;��H;b�H;�H;��H;t�H;�H;��H;A�H;��H;��H;@�H;��H;��H;F�H;��H;��H;��H;_�H;A�H;�H;��H;��H;��H;��H;��H;�H;A�H;_�H;��H;��H;��H;F�H;��H;��H;@�H;��H;��H;A�H;��H;�H;t�H;��H;�H;b�H;��H;��H;%�H;T�H;m�H;v�H;��H;��H;l�H;u�H;V�H;>�H;F�H;B�H;      L�H;p�H;��H;��H;��H;'�H;I�H;w�H;��H;��H;��H;��H;��H;��H;��H;��H;7�H;��H;��H;5�H;��H;��H;�H;��H;r�H;�H;��H;u�H;7�H;��H;��H;��H;w�H;?�H;�H;'�H;(�H;'�H;�H;?�H;w�H;��H;��H;��H;7�H;u�H;��H;�H;r�H;��H;�H;��H;��H;5�H;��H;��H;7�H;��H;��H;��H;��H;��H;��H;��H;��H;w�H;I�H;'�H;��H;��H;��H;p�H;      ��H;�H;�H;w�H;��H;e�H;�H;��H;#�H;��H;��H;!�H;T�H;y�H;k�H;d�H;F�H;�H;��H;y�H;�H;��H;��H;	�H;��H;`�H;�H;��H;k�H;-�H;��H;��H;��H;��H;c�H;K�H;A�H;K�H;c�H;��H;��H;��H;��H;-�H;k�H;��H;�H;`�H;��H;	�H;��H;��H;�H;y�H;��H;�H;F�H;d�H;k�H;y�H;T�H;!�H;��H;��H;#�H;��H;�H;e�H;��H;w�H;�H;�H;      ��H;U�H;7�H;��H;��H;i�H;��H;��H;��H;��H;��H;��H;A�H;��H;��H;!�H;9�H;�H;��H;��H;[�H;��H;��H;e�H;��H;��H;H�H;�H;��H;k�H;7�H;��H;��H;��H;��H;��H;�H;��H;��H;��H;��H;��H;7�H;k�H;��H;�H;H�H;��H;��H;e�H;��H;��H;[�H;��H;��H;�H;9�H;!�H;��H;��H;A�H;��H;��H;��H;��H;��H;��H;i�H;��H;��H;7�H;U�H;      ��H;4�H;��H;Z�H;Q�H;��H;L�H;��H;'�H;1�H;&�H;��H;�H;"�H;��H;W�H;��H;��H;��H;��H;��H;a�H;��H;��H;h�H;��H;��H;W�H;�H;��H;u�H;F�H; �H;��H;��H;��H;��H;��H;��H;��H; �H;F�H;u�H;��H;�H;W�H;��H;��H;h�H;��H;��H;a�H;��H;��H;��H;��H;��H;W�H;��H;"�H;�H;��H;&�H;1�H;'�H;��H;L�H;��H;Q�H;Z�H;��H;4�H;      �H;H;� H;�7H;�SH;KrH;9�H;ԪH;��H;��H;{�H;��H;�H;�H;��H;��H;��H;=�H;��H;��H;��H;��H;4�H;��H;��H;_�H;��H;��H;H�H;�H;��H;��H;b�H;C�H;(�H;�H;�H;�H;(�H;C�H;b�H;��H;��H;�H;H�H;��H;��H;_�H;��H;��H;4�H;��H;��H;��H;��H;=�H;��H;��H;��H;�H;�H;��H;{�H;��H;��H;ԪH;9�H;KrH;�SH;�7H;� H;H;      mCF;zQF;�yF;�F;�G;�[G;�G;YH;#HH;��H;��H;��H;
�H;��H;��H;8�H;��H;7�H;��H;P�H;��H;~�H;r�H;D�H;��H;��H;_�H;��H;��H;`�H;�H;��H;��H;��H;o�H;\�H;n�H;\�H;o�H;��H;��H;��H;�H;`�H;��H;��H;_�H;��H;��H;D�H;r�H;~�H;��H;P�H;��H;7�H;��H;8�H;��H;��H;
�H;��H;��H;��H;#HH;YH;�G;�[G;�G;�F;�yF;zQF;      ��A;~B;1oB;�C;��C;{�D;otE;CF;M�F;��G;�H;eH;�H;��H;[�H;�H;��H;�H;��H;��H;"�H;e�H;��H;i�H;-�H;��H;��H;h�H;��H;��H;r�H;@�H;
�H;��H;��H;��H;��H;��H;��H;��H;
�H;@�H;r�H;��H;��H;h�H;��H;��H;-�H;i�H;��H;e�H;"�H;��H;��H;�H;��H;�H;[�H;��H;�H;eH;�H;��G;M�F;CF;otE;{�D;��C;�C;1oB;~B;      ~n8;L�8;׎9;��:;��<;
c>;ZQ@;�.B;��C;�OE;�yF;j[G;��G;DhH;8�H;��H;8�H;a�H;,�H;5�H;\�H;��H;a�H;j�H;i�H;D�H;��H;��H;e�H;	�H;��H;��H;Y�H;(�H;!�H;�H;��H;�H;!�H;(�H;Y�H;��H;��H;	�H;e�H;��H;��H;D�H;i�H;j�H;a�H;��H;\�H;5�H;,�H;a�H;8�H;��H;8�H;DhH;��G;j[G;�yF;�OE;��C;�.B;ZQ@;
c>;��<;��:;׎9;L�8;      �R%;i�%;^�';M*;4�-;ʕ1;�5;5�9;�,=;HQ@;�B;��D;9lF;�tG;� H;�H;��H;��H;�H;��H;��H;0�H;�H;a�H;��H;r�H;4�H;��H;��H;��H;�H;��H;��H;��H;|�H;e�H;L�H;e�H;|�H;��H;��H;��H;�H;��H;��H;��H;4�H;r�H;��H;a�H;�H;0�H;��H;��H;�H;��H;��H;�H;� H;�tG;9lF;��D;�B;HQ@;�,=;5�9;�5;ʕ1;4�-;M*;^�';i�%;      �V;�w;0�;P�
;�;�;)� ;��(;��/;#H6;��;;�?; C;�OE;�F;�G;�dH;M�H;��H;&�H;O�H;��H;0�H;��H;e�H;~�H;��H;a�H;��H;��H;��H;A�H;�H;�H;��H;��H;��H;��H;��H;�H;�H;A�H;��H;��H;��H;a�H;��H;~�H;e�H;��H;0�H;��H;O�H;&�H;��H;M�H;�dH;�G;�F;�OE; C;�?;��;;#H6;��/;��(;)� ;�;�;P�
;0�;�w;      車:lĆ:nȒ:���:p�:m��:���:��	;v;7�#;��-;#�5;�K<;��@;�'D;3CF;��G;�GH;s�H;�H;��H;O�H;��H;\�H;"�H;��H;��H;��H;[�H;�H;��H;��H;m�H;[�H;)�H;�H;�H;�H;)�H;[�H;m�H;��H;��H;�H;[�H;��H;��H;��H;"�H;\�H;��H;O�H;��H;�H;s�H;�GH;��G;3CF;�'D;��@;�K<;#�5;��-;7�#;v;��	;���:m��:p�:���:nȒ:lĆ:      0.�9��3�깩�K�
9�Z:��k:�K�:4��:�x;��;�$;
�/;��8;��>;#C;7�E;�[G;\7H;̤H;�H;&�H;��H;5�H;��H;P�H;��H;��H;��H;y�H;5�H;�H;��H;��H;��H;��H;t�H;��H;��H;��H;��H;�H;5�H;y�H;��H;��H;��H;P�H;��H;5�H;��H;&�H;�H;̤H;\7H;�[G;7�E;#C;��>;��8;
�/;�$;��;�x;4��:�K�:��k:�Z:
9��K�3��9��      �Q^��X�VF�]�)��+�-ж���<�YjS�}k:���:H��:�;|�;M*;�5;�b=;�oB;��E;�IG;\7H;s�H;��H;�H;,�H;��H;��H;��H;��H;��H;��H;��H;t�H;P�H;��H;��H;��H;��H;��H;��H;��H;P�H;t�H;��H;��H;��H;��H;��H;��H;��H;,�H;�H;��H;s�H;\7H;�IG;��E;�oB;�b=;�5;M*;|�;�;H��:���:}k:YjS���<�-ж��+�]�)�VF��X�      ����o���X��P�ѻf���[ǐ��X��6��
���K�:<":eL�:�`�:�h;Z�%;��3;�<;X/B;��E;�[G;�GH;M�H;��H;a�H;�H;7�H;=�H;��H;�H;�H;��H;��H;��H;]�H;O�H;K�H;'�H;K�H;O�H;]�H;��H;��H;��H;�H;�H;��H;=�H;7�H;�H;a�H;��H;M�H;�GH;�[G;��E;X/B;�<;��3;Z�%;�h;�`�:eL�::<":�K��
���6��X�[ǐ�f���P�ѻX��o���      ��n��mj���]���J�n�1�L4�l��S���V
x�iX���y�!
9���:գ�:?�;u�#;v�2;�<;�oB;7�E;��G;�dH;��H;8�H;��H;��H;��H;��H;9�H;F�H;7�H;�H;��H;��H;��H;��H;��H;��H;��H;��H;��H;�H;7�H;F�H;9�H;��H;��H;��H;��H;8�H;��H;�dH;��G;7�E;�oB;�<;v�2;u�#;?�;գ�:���:!
9��y�iX�V
x�S���l��L4�n�1���J���]��mj�      B<ͼ��ɼ�����֯�Ҷ��ㄼ��Y�-�*�J���t���X��sѺ�(�J<Q:[��:��
;u�#;��3;�b=;#C;3CF;�G;�H;��H;�H;8�H;��H;W�H;!�H;d�H;��H;b�H;5�H;O�H;	�H;��H;�H;��H;	�H;O�H;5�H;b�H;��H;d�H;!�H;W�H;��H;8�H;�H;��H;�H;�G;3CF;#C;�b=;��3;u�#;��
;[��:J<Q:�(��sѺ�X�t��J���-�*���Y�ㄼҶ���֯�������ɼ      ��'�#�$����y��  ���ۼ����+����]��X!�>ۻ�+��+�k���>:[��:?�;Z�%;�5;��>;�'D;�F;� H;8�H;[�H;��H;��H;��H;��H;k�H;��H;��H;��H;��H;g�H;J�H;m�H;J�H;g�H;��H;��H;��H;��H;k�H;��H;��H;��H;��H;[�H;8�H;� H;�F;�'D;��>;�5;Z�%;?�;[��:�>:k��+��+��>ۻ�X!���]��+�������ۼ�  �y����#�$�      �����v����w�]�c��J�Ȅ-�x��;缈沼ㄼ��;�����k��66�k��J<Q:գ�:�h;M*;��8;��@;�OE;�tG;DhH;��H;��H;�H;"�H;��H;y�H;��H;��H;��H;��H;��H;��H;��H;��H;��H;��H;��H;��H;��H;y�H;��H;"�H;�H;��H;��H;DhH;�tG;�OE;��@;��8;M*;�h;գ�:J<Q:k��66�k��������;�ㄼ�沼�;�x�Ȅ-��J�]�c���w��v��      nHͽ̪ɽ�;��"����������[�z0�p��'<ͼо��v�J���k��+��(����:�`�:|�;
�/;�K<; C;9lF;��G;�H;
�H;�H;�H;A�H;T�H;��H;%�H;/�H;�H;�H;�H;��H;�H;�H;�H;/�H;%�H;��H;T�H;A�H;�H;�H;
�H;�H;��G;9lF; C;�K<;
�/;|�;�`�:���:�(�+�k����v�J�о��'<ͼp��z0���[�������"���;��̪ɽ      ��-�}��|�ű�ƽUP���v���J�D����ۼ��v�J������+���sѺ!
9eL�:�;�$;#�5;�?;��D;j[G;eH;��H;��H;��H;��H;!�H;��H;T�H;n�H;Y�H;T�H;a�H;7�H;a�H;T�H;Y�H;n�H;T�H;��H;!�H;��H;��H;��H;��H;eH;j[G;��D;�?;#�5;�$;�;eL�:!
9�sѺ�+������v�J�����ۼD���J��v��UP��ƽű�|�}��-�       j�Ide�M0X�sD�\{+�z�����k㻽R���JDX������ۼо����;�>ۻ�X���y�:<":H��:��;��-;��;;�B;�yF;�H;��H;{�H;&�H;��H;��H;��H;m�H;��H;��H;��H;��H;z�H;��H;��H;��H;��H;m�H;��H;��H;��H;&�H;{�H;��H;�H;�yF;�B;��;;��-;��;H��::<":��y��X�>ۻ��;�о����ۼ���JDX�R���k㻽���z��\{+�sD�M0X�Ide�      ��Fh��b���I���|x���O��C(�y�Īɽ����JDX�D��'<ͼㄼ�X!�t��iX��K����:�x;7�#;#H6;HQ@;�OE;��G;��H;��H;1�H;��H;��H;��H;v�H;��H;��H;��H;��H;��H;��H;��H;��H;��H;v�H;��H;��H;��H;1�H;��H;��H;��G;�OE;HQ@;#H6;7�#;�x;���:�K�iX�t���X!�ㄼ'<ͼD��JDX�����Īɽy��C(���O��|x��I��b��Fh��      /�����������;^ɰ��G����i�.�5��	�ĪɽR����J�p���沼��]�J���V
x��
��}k:4��:v;��/;�,=;��C;M�F;#HH;��H;'�H;��H;#�H;��H;��H;��H;�H;�H;�H;#�H;�H;�H;�H;��H;��H;��H;#�H;��H;'�H;��H;#HH;M�F;��C;�,=;��/;v;4��:}k:�
��V
x�J�����]��沼p���J�R���Īɽ�	�.�5���i��G��^ɰ��;��徨���      �2�L�-��"�$E�����4Kɾa��w�s�.�5�y�k㻽�v��z0��;��+��-�*�S����6�YjS��K�:��	;��(;5�9;�.B;CF;YH;ԪH;��H;��H;��H;w�H;��H;�H;/�H;C�H;<�H;Y�H;<�H;C�H;/�H;�H;��H;w�H;��H;��H;��H;ԪH;YH;CF;�.B;5�9;��(;��	;�K�:YjS��6�S���-�*��+���;�z0��v��k㻽y�.�5�w�s�a��4Kɾ����$E��"�L�-�      3s�cm�/�\�]�C�,�%����TҾa����i��C(����UP����[�x������Y�l���X���<���k:���:)� ;�5;ZQ@;otE;�G;9�H;L�H;��H;�H;I�H;l�H;$�H;b�H;s�H;W�H;��H;W�H;s�H;b�H;$�H;l�H;I�H;�H;��H;L�H;9�H;�G;otE;ZQ@;�5;)� ;���:��k:��<��X�l����Y����x���[�UP����콡C(���i�a���TҾ��,�%�]�C�/�\�cm�      �ޞ�������RF�3�W�M�-���4Kɾ�G����O�z��ƽ����Ȅ-���ۼㄼL4�[ǐ�-ж��Z:m��:�;ʕ1;
c>;{�D;�[G;KrH;��H;i�H;e�H;'�H;u�H;(�H;h�H;��H;|�H;��H;|�H;��H;h�H;(�H;u�H;'�H;e�H;i�H;��H;KrH;�[G;{�D;
c>;ʕ1;�;m��:�Z:-ж�[ǐ�L4�ㄼ��ۼȄ-�����ƽz����O��G��4Kɾ��M�-�3�W�RF�������      ��ſ~��Bw���ޞ�|���3�W�,�%�����^ɰ��|x�\{+�ű����J��  �Ҷ��n�1�f����+�
9p�:�;4�-;��<;��C;�G;�SH;Q�H;��H;��H;��H;V�H;2�H;��H;��H;��H;��H;��H;��H;��H;2�H;V�H;��H;��H;��H;Q�H;�SH;�G;��C;��<;4�-;�;p�:
9�+�f���n�1�Ҷ���  ��J���ű�\{+��|x�^ɰ�����,�%�3�W�|����ޞ�Bw��~��      ������Կp���ޞ�RF�]�C�$E��;�I��sD�|�"��]�c�y��֯���J�P�ѻ]�)���K����:P�
;M*;��:;�C;�F;�7H;Z�H;��H;w�H;��H;>�H;9�H;��H;��H;��H;��H;��H;��H;��H;9�H;>�H;��H;w�H;��H;Z�H;�7H;�F;�C;��:;M*;P�
;���:��K�]�)�P�ѻ��J��֯�y�]�c�"��|�sD��I���;$E�]�C�RF��ޞ�p���Կ��      ������{���ԿBw�����/�\��"����b��M0X�}���;����w����������]�X��VF�3��nȒ:0�;^�';׎9;1oB;�yF;� H;��H;7�H;�H;��H;F�H;:�H;��H;��H;��H;�H;��H;��H;��H;:�H;F�H;��H;�H;7�H;��H;� H;�yF;1oB;׎9;^�';0�;nȒ:3��VF�X�黼�]����������w��;��}��M0X�b������"�/�\����Bw���Կ{�𿖏�      $��������~�����cm�L�-�����Fh��Ide�-�̪ɽ�v��#�$���ɼ�mj�o����X�9��lĆ:�w;i�%;L�8;~B;zQF;H;4�H;U�H;�H;p�H;B�H;5�H;��H;��H;��H;$�H;��H;��H;��H;5�H;B�H;p�H;�H;U�H;4�H;H;zQF;~B;L�8;i�%;�w;lĆ:9���X�o����mj���ɼ#�$��v��̪ɽ-�Ide�Fh������L�-�cm����~���忖����      Vܿ%�ֿ�aǿ2^��&���Io���7����iþ�(���-=��` ��@����_�&]�&p����I�r�ѻ��)�"�R�[�:��
;*;C�:;�B;UHF;=�G;�kH;3�H;��H;h�H;��H;��H;o�H;��H;(�H;��H;(�H;��H;o�H;��H;��H;h�H;��H;3�H;�kH;=�G;UHF;�B;C�:;*;��
;[�:"�R���)�r�ѻ��I�&p��&]���_��@���` ��-=��(���iþ����7�Io�&���2^���aǿ%�ֿ      %�ֿ5pѿ֊¿������PXi�Õ3��
�GD��;l��1�9�j.���R��\� �\x��1�E��ͻ��$�� ����:��;��*;[�:;-�B;3TF;��G;ZmH;ϠH;ܶH;��H;��H;��H;�H;��H;<�H;��H;<�H;��H;�H;��H;��H;��H;ܶH;ϠH;ZmH;��G;3TF;-�B;[�:;��*;��;���:� ���$��ͻ1�E�\x�� �\��R��j.��1�9�;l��GD���
�Õ3�PXi�������֊¿5pѿ      �aǿ֊¿���������s"Y��f'�����)o���.}��k/�m��ڟ�<Q�%#�ע��(;�P������l�7���:I�;�,;��;;�C;RvF;/�G;�qH;[�H;��H;<�H;�H;�H;��H;��H;j�H;��H;j�H;��H;��H;�H;�H;<�H;��H;[�H;�qH;/�G;RvF;�C;��;;�,;I�;��:l�7����P����(;�ע�%#�<Q�ڟ�m���k/��.}�)o�������f'�s"Y����������֊¿      2^������b���Io���@���޾����&ce�"����ڽ绒��f@������R���O*�mG�����r<^9Ѳ�:[;�c.;&�<;ԏC;F�F;��G;�xH;äH;7�H;I�H;��H;��H;��H;�H;��H;6�H;��H;�H;��H;��H;��H;I�H;7�H;äH;�xH;��G;F�F;ԏC;&�<;�c.;[;Ѳ�:r<^9���mG���O*��R�������f@�绒���ڽ"��&ce������޾���@�Io�b�������      &����������Io��!J�@�#��\��HD������jPH�����b��C��t +�u�ټ%��������������:���:��;�X1;3>;�/D;��F;�H;r�H;��H;)�H;��H;��H;)�H;��H;p�H;��H;~�H;��H;p�H;��H;)�H;��H;��H;)�H;��H;r�H;�H;��F;�/D;3>;�X1;��;���:��:����������%��u�ټt +�C���b�����jPH�����HD���\��@�#��!J�Io��������      Io�PXi�s"Y���@�@�#��
��о�A�� �i���(�i��gr����_��5��ɺ�o�`��<����d�A�\�L�X:NO�:6`;#�4;�?;��D;�7G;�/H;ȊH;��H;��H;.�H;��H;��H;�H;��H;-�H;��H;-�H;��H;�H;��H;��H;.�H;��H;��H;ȊH;�/H;�7G;��D;�?;#�4;6`;NO�:L�X:A�\���d��<��o�`��ɺ��5���_�gr��i����(� �i��A���о�
�@�#���@�s"Y�PXi�      ��7�Õ3��f'���\���о�����.}��-=�o
�y�ĽO��:����������7�@GĻ+�$�S�����:�z;�C&;D+8;EIA;0�E;��G;�KH;�H;��H;R�H;�H;(�H;��H;��H;@�H;��H;5�H;��H;@�H;��H;��H;(�H;�H;R�H;��H;�H;�KH;��G;0�E;EIA;D+8;�C&;�z;���:S��+�$�@GĻ�7���������:�O��y�Ľo
��-=��.}������о�\����f'�Õ3�      ���
������޾HD���A���.}��D�[t���ڽ�!��\����P�ļ�
v�F�����Jɺ�N�9���:h';�-;ӊ;;��B;�HF;��G;?eH;ʜH;�H;M�H;��H;��H;��H;{�H;��H;�H;��H;�H;��H;{�H;��H;��H;��H;M�H;�H;ʜH;?eH;��G;�HF;��B;ӊ;;�-;h';���:�N�9�Jɺ��F���
v�P�ļ���\��!����ڽ[t��D��.}��A��HD���޾�����
�      �iþGD��)o���������� �i��-=�[t����R��Tys�m +����s񗼗(;�H�ѻt@�Ї!��1j:�O�:3�;�C3;}�>;CED;��F;�H;_{H;��H;��H;V�H;�H;�H;��H;9�H;R�H;��H;�H;��H;R�H;9�H;��H;�H;�H;V�H;��H;��H;_{H;�H;��F;CED;}�>;�C3;3�;�O�:�1j:Ї!�t@�H�ѻ�(;�s����m +�Tys��R����[t��-=� �i���������)o��GD��      �(��;l���.}�&ce�jPH���(�o
���ڽ�R����{�4�6�� �$p��\�`�ר�-��JҺ�C^9_��:=�;�}(;t�8;IA;5{E;FiG;�<H;i�H;��H;H�H;�H;N�H;��H;��H;��H;��H;�H;i�H;�H;��H;��H;��H;��H;N�H;�H;H�H;��H;i�H;�<H;FiG;5{E;IA;t�8;�}(;=�;_��:�C^9JҺ-��ר�\�`�$p��� �4�6���{��R����ڽo
���(�jPH�&ce��.}�;l��      �-=�1�9��k/�"�����i��y�Ľ�!��Tys�4�6�#��ɺ��vz����c^��̃$������r:���:6�;�X1;>H=;iwC;VvF;R�G;/eH;m�H;��H;��H;��H;u�H;�H;��H;��H;��H;��H;��H;��H;��H;��H;��H;�H;u�H;��H;��H;��H;m�H;/eH;R�G;VvF;iwC;>H=;�X1;6�;���:��r:���̃$�c^������vz��ɺ�#�4�6�Tys��!��y�Ľi���"���k/�1�9�      �` �j.��m��ڽ�b��gr��O��\�m +�� ��ɺ�=��O*�bͻQ6R��ǅ���:���:ڃ;�);6t8;��@;�)E;�7G;s#H;o�H;c�H;�H;I�H;��H;��H;��H;�H;m�H;�H; �H;>�H; �H;�H;m�H;�H;��H;��H;��H;I�H;�H;c�H;o�H;s#H;�7G;�)E;��@;6t8;�);ڃ;���:��:�ǅ�Q6R�bͻ�O*�=��ɺ�� �m +�\�O��gr���b����ڽm��j.��      �@���R��ڟ�绒�C����_�:�������$p���vz��O*�5ֻgk������09�:_0;�� ;�C3;��=;�C;kF;��G;�[H;H;o�H;%�H;a�H;��H;��H;��H;�H;&�H;��H;n�H;��H;n�H;��H;&�H;�H;��H;��H;��H;a�H;%�H;o�H;H;�[H;��G;kF;�C;��=;�C3;�� ;_0;�:��09���gk�5ֻ�O*��vz�$p����輙��:���_�C��绒�ڟ��R��      ��_�\�<Q��f@�t +��5�����P�ļs�\�`����bͻgk��Iɺ
7��:�O�:x�;%d.;��:;Z�A;c{E;�MG;p&H;/�H;�H;��H;��H;I�H;m�H;|�H;R�H;�H;��H;*�H;��H;�H;��H;*�H;��H;�H;R�H;|�H;m�H;I�H;��H;��H;�H;/�H;p&H;�MG;c{E;Z�A;��:;%d.;x�;�O�:�:
7��Iɺgk�bͻ���\�`�s�P�ļ�����5�t +��f@�<Q�\�      &]� �%#�����u�ټ�ɺ������
v��(;�ר�c^��Q6R����
7����:���:N�;k�*;+8;� @;��D;��F;'�G; eH;��H;��H;ľH;��H;�H;��H;A�H;��H;��H;��H;��H;B�H;u�H;B�H;��H;��H;��H;��H;A�H;��H;�H;��H;ľH;��H;��H; eH;'�G;��F;��D;� @;+8;k�*;N�;���:���:
7����Q6R�c^��ר��(;��
v������ɺ�u�ټ����%#� �      &p��\x��ע��R��%��o�`��7�F��H�ѻ-��̃$��ǅ���09�:���:�; ~(;�Y6;��>;�C;%HF;�G;DH;s�H;�H;θH;2�H;K�H;2�H;�H;��H;��H;��H;,�H;�H;��H;��H;��H;�H;,�H;��H;��H;��H;�H;2�H;K�H;2�H;θH;�H;s�H;DH;�G;%HF;�C;��>;�Y6; ~(;�;���:�:��09�ǅ�̃$�-��H�ѻF���7�o�`�%���R��ע�\x��      ��I�1�E��(;��O*�����<��@GĻ��t@�JҺ���:�:�O�:N�; ~(;R�5;>;pC;j�E;�bG;k#H;"{H;^�H;H�H;��H;��H;Y�H;��H;:�H;w�H;��H;h�H;��H;Y�H;��H;�H;��H;Y�H;��H;h�H;��H;w�H;:�H;��H;Y�H;��H;��H;H�H;^�H;"{H;k#H;�bG;j�E;pC;>;R�5; ~(;N�;�O�:�:��:���JҺt@���@GĻ�<������O*��(;�1�E�      r�ѻ�ͻP���mG�������d�+�$��JɺЇ!��C^9��r:���:_0;x�;k�*;�Y6;>;n�B;��E;8G;�H;+mH;@�H;m�H;μH;��H;��H;��H;g�H;�H;��H;��H;�H;�H;��H;�H;<�H;�H;��H;�H;�H;��H;��H;�H;g�H;��H;��H;��H;μH;m�H;@�H;+mH;�H;8G;��E;n�B;>;�Y6;k�*;x�;_0;���:��r:�C^9Ї!��Jɺ+�$���d����mG��P����ͻ      ��)���$�����������A�\�S���N�9�1j:_��:���:ڃ;�� ;%d.;+8;��>;pC;��E;�(G;��G;=cH;��H;��H;��H;��H;T�H;��H;��H;��H;��H;��H;a�H;��H;w�H;�H;I�H;b�H;I�H;�H;w�H;��H;a�H;��H;��H;��H;��H;��H;T�H;��H;��H;��H;��H;=cH;��G;�(G;��E;pC;��>;+8;%d.;�� ;ڃ;���:_��:�1j:�N�9S��A�\�������������$�      "�R�� �l�7�r<^9��:L�X:���:���:�O�:=�;6�;�);�C3;��:;� @;�C;j�E;8G;��G;�_H;��H;>�H;?�H;��H;d�H;Q�H;h�H;w�H;��H;��H;��H;$�H;��H;��H;@�H;{�H;{�H;{�H;@�H;��H;��H;$�H;��H;��H;��H;w�H;h�H;Q�H;d�H;��H;?�H;>�H;��H;�_H;��G;8G;j�E;�C;� @;��:;�C3;�);6�;=�;�O�:���:���:L�X:��:r<^9l�7�� �      [�:���:��:Ѳ�:���:NO�:�z;h';3�;�}(;�X1;6t8;��=;Z�A;��D;%HF;�bG;�H;=cH;��H;m�H;��H;R�H;�H;��H;Y�H;d�H;��H;<�H;��H;��H;��H;l�H;��H;X�H;��H;��H;��H;X�H;��H;l�H;��H;��H;��H;<�H;��H;d�H;Y�H;��H;�H;R�H;��H;m�H;��H;=cH;�H;�bG;%HF;��D;Z�A;��=;6t8;�X1;�}(;3�;h';�z;NO�:���:Ѳ�:��:���:      ��
;��;I�;[;��;6`;�C&;�-;�C3;t�8;>H=;��@;�C;c{E;��F;�G;k#H;+mH;��H;>�H;��H;��H;Y�H;9�H;��H;��H;��H;��H;~�H;�H;4�H;�H;��H;1�H;r�H;��H;��H;��H;r�H;1�H;��H;�H;4�H;�H;~�H;��H;��H;��H;��H;9�H;Y�H;��H;��H;>�H;��H;+mH;k#H;�G;��F;c{E;�C;��@;>H=;t�8;�C3;�-;�C&;6`;��;[;I�;��;      *;��*;�,;�c.;�X1;#�4;D+8;ӊ;;}�>;IA;iwC;�)E;kF;�MG;'�G;DH;"{H;@�H;��H;?�H;R�H;Y�H;��H;�H;�H;w�H;"�H;�H;��H;��H;��H;��H;��H;L�H;��H;��H;��H;��H;��H;L�H;��H;��H;��H;��H;��H;�H;"�H;w�H;�H;�H;��H;Y�H;R�H;?�H;��H;@�H;"{H;DH;'�G;�MG;kF;�)E;iwC;IA;}�>;ӊ;;D+8;#�4;�X1;�c.;�,;��*;      C�:;[�:;��;;&�<;3>;�?;EIA;��B;CED;5{E;VvF;�7G;��G;p&H; eH;s�H;^�H;m�H;��H;��H;�H;9�H;�H;��H;5�H;��H;��H;G�H;��H;~�H;(�H;��H;,�H;l�H;��H;��H;��H;��H;��H;l�H;,�H;��H;(�H;~�H;��H;G�H;��H;��H;5�H;��H;�H;9�H;�H;��H;��H;m�H;^�H;s�H; eH;p&H;��G;�7G;VvF;5{E;CED;��B;EIA;�?;3>;&�<;��;;[�:;      �B;-�B;�C;ԏC;�/D;��D;0�E;�HF;��F;FiG;R�G;s#H;�[H;/�H;��H;�H;H�H;μH;��H;d�H;��H;��H;�H;5�H;��H;��H;�H;T�H;8�H;�H;��H;��H;=�H;��H;��H;��H;��H;��H;��H;��H;=�H;��H;��H;�H;8�H;T�H;�H;��H;��H;5�H;�H;��H;��H;d�H;��H;μH;H�H;�H;��H;/�H;�[H;s#H;R�G;FiG;��F;�HF;0�E;��D;�/D;ԏC;�C;-�B;      UHF;3TF;RvF;F�F;��F;�7G;��G;��G;�H;�<H;/eH;o�H;H;�H;��H;θH;��H;��H;T�H;Q�H;Y�H;��H;w�H;��H;��H;	�H;9�H;�H;��H;R�H;��H;.�H;C�H;}�H;��H;��H;��H;��H;��H;}�H;C�H;.�H;��H;R�H;��H;�H;9�H;	�H;��H;��H;w�H;��H;Y�H;Q�H;T�H;��H;��H;θH;��H;�H;H;o�H;/eH;�<H;�H;��G;��G;�7G;��F;F�F;RvF;3TF;      =�G;��G;/�G;��G;�H;�/H;�KH;?eH;_{H;i�H;m�H;c�H;o�H;��H;ľH;2�H;��H;��H;��H;h�H;d�H;��H;"�H;��H;�H;9�H;�H;��H;[�H;��H;��H;<�H;\�H;�H;��H;��H;��H;��H;��H;�H;\�H;<�H;��H;��H;[�H;��H;�H;9�H;�H;��H;"�H;��H;d�H;h�H;��H;��H;��H;2�H;ľH;��H;o�H;c�H;m�H;i�H;_{H;?eH;�KH;�/H;�H;��G;/�G;��G;      �kH;ZmH;�qH;�xH;r�H;ȊH;�H;ʜH;��H;��H;��H;�H;%�H;��H;��H;K�H;Y�H;��H;��H;w�H;��H;��H;�H;G�H;T�H;�H;��H;B�H;��H;��H;�H;B�H;k�H;l�H;��H;��H;��H;��H;��H;l�H;k�H;B�H;�H;��H;��H;B�H;��H;�H;T�H;G�H;�H;��H;��H;w�H;��H;��H;Y�H;K�H;��H;��H;%�H;�H;��H;��H;��H;ʜH;�H;ȊH;r�H;�xH;�qH;ZmH;      3�H;ϠH;[�H;äH;��H;��H;��H;�H;��H;H�H;��H;I�H;a�H;I�H;�H;2�H;��H;g�H;��H;��H;<�H;~�H;��H;��H;8�H;��H;[�H;��H;��H;�H;6�H;S�H;j�H;k�H;j�H;u�H;u�H;u�H;j�H;k�H;j�H;S�H;6�H;�H;��H;��H;[�H;��H;8�H;��H;��H;~�H;<�H;��H;��H;g�H;��H;2�H;�H;I�H;a�H;I�H;��H;H�H;��H;�H;��H;��H;��H;äH;[�H;ϠH;      ��H;ܶH;��H;7�H;)�H;��H;R�H;M�H;V�H;�H;��H;��H;��H;m�H;��H;�H;:�H;�H;��H;��H;��H;�H;��H;~�H;�H;R�H;��H;��H;�H;+�H;J�H;I�H;X�H;h�H;O�H;a�H;{�H;a�H;O�H;h�H;X�H;I�H;J�H;+�H;�H;��H;��H;R�H;�H;~�H;��H;�H;��H;��H;��H;�H;:�H;�H;��H;m�H;��H;��H;��H;�H;V�H;M�H;R�H;��H;)�H;7�H;��H;ܶH;      h�H;��H;<�H;I�H;��H;.�H;�H;��H;�H;N�H;u�H;��H;��H;|�H;A�H;��H;w�H;��H;��H;��H;��H;4�H;��H;(�H;��H;��H;��H;�H;6�H;J�H;a�H;T�H;E�H;E�H;c�H;U�H;6�H;U�H;c�H;E�H;E�H;T�H;a�H;J�H;6�H;�H;��H;��H;��H;(�H;��H;4�H;��H;��H;��H;��H;w�H;��H;A�H;|�H;��H;��H;u�H;N�H;�H;��H;�H;.�H;��H;I�H;<�H;��H;      ��H;��H;�H;��H;��H;��H;(�H;��H;�H;��H;�H;��H;��H;R�H;��H;��H;��H;��H;a�H;$�H;��H;�H;��H;��H;��H;.�H;<�H;B�H;S�H;I�H;T�H;Z�H;C�H;=�H;O�H;4�H;+�H;4�H;O�H;=�H;C�H;Z�H;T�H;I�H;S�H;B�H;<�H;.�H;��H;��H;��H;�H;��H;$�H;a�H;��H;��H;��H;��H;R�H;��H;��H;�H;��H;�H;��H;(�H;��H;��H;��H;�H;��H;      ��H;��H;�H;��H;)�H;��H;��H;��H;��H;��H;��H;�H;�H;�H;��H;��H;h�H;�H;��H;��H;l�H;��H;��H;,�H;=�H;C�H;\�H;k�H;j�H;X�H;E�H;C�H;G�H;C�H;"�H;#�H;S�H;#�H;"�H;C�H;G�H;C�H;E�H;X�H;j�H;k�H;\�H;C�H;=�H;,�H;��H;��H;l�H;��H;��H;�H;h�H;��H;��H;�H;�H;�H;��H;��H;��H;��H;��H;��H;)�H;��H;�H;��H;      o�H;�H;��H;��H;��H;�H;��H;{�H;9�H;��H;��H;m�H;&�H;��H;��H;,�H;��H;�H;w�H;��H;��H;1�H;L�H;l�H;��H;}�H;�H;l�H;k�H;h�H;E�H;=�H;C�H;-�H;�H;#�H;)�H;#�H;�H;-�H;C�H;=�H;E�H;h�H;k�H;l�H;�H;}�H;��H;l�H;L�H;1�H;��H;��H;w�H;�H;��H;,�H;��H;��H;&�H;m�H;��H;��H;9�H;{�H;��H;�H;��H;��H;��H;�H;      ��H;��H;��H;�H;p�H;��H;@�H;��H;R�H;��H;��H;�H;��H;*�H;��H;�H;Y�H;��H;�H;@�H;X�H;r�H;��H;��H;��H;��H;��H;��H;j�H;O�H;c�H;O�H;"�H;�H;'�H;�H;�H;�H;'�H;�H;"�H;O�H;c�H;O�H;j�H;��H;��H;��H;��H;��H;��H;r�H;X�H;@�H;�H;��H;Y�H;�H;��H;*�H;��H;�H;��H;��H;R�H;��H;@�H;��H;p�H;�H;��H;��H;      (�H;<�H;j�H;��H;��H;-�H;��H;�H;��H;�H;��H; �H;n�H;��H;B�H;��H;��H;�H;I�H;{�H;��H;��H;��H;��H;��H;��H;��H;��H;u�H;a�H;U�H;4�H;#�H;#�H;�H;�H;�H;�H;�H;#�H;#�H;4�H;U�H;a�H;u�H;��H;��H;��H;��H;��H;��H;��H;��H;{�H;I�H;�H;��H;��H;B�H;��H;n�H; �H;��H;�H;��H;�H;��H;-�H;��H;��H;j�H;<�H;      ��H;��H;��H;6�H;~�H;��H;5�H;��H;�H;i�H;��H;>�H;��H;�H;u�H;��H;�H;<�H;b�H;{�H;��H;��H;��H;��H;��H;��H;��H;��H;u�H;{�H;6�H;+�H;S�H;)�H;�H;�H;�H;�H;�H;)�H;S�H;+�H;6�H;{�H;u�H;��H;��H;��H;��H;��H;��H;��H;��H;{�H;b�H;<�H;�H;��H;u�H;�H;��H;>�H;��H;i�H;�H;��H;5�H;��H;~�H;6�H;��H;��H;      (�H;<�H;j�H;��H;��H;-�H;��H;�H;��H;�H;��H; �H;n�H;��H;B�H;��H;��H;�H;I�H;{�H;��H;��H;��H;��H;��H;��H;��H;��H;u�H;a�H;U�H;4�H;#�H;#�H;�H;�H;�H;�H;�H;#�H;#�H;4�H;U�H;a�H;u�H;��H;��H;��H;��H;��H;��H;��H;��H;{�H;I�H;�H;��H;��H;B�H;��H;n�H; �H;��H;�H;��H;�H;��H;-�H;��H;��H;j�H;<�H;      ��H;��H;��H;�H;p�H;��H;@�H;��H;R�H;��H;��H;�H;��H;*�H;��H;�H;Y�H;��H;�H;@�H;X�H;r�H;��H;��H;��H;��H;��H;��H;j�H;O�H;c�H;O�H;"�H;�H;'�H;�H;�H;�H;'�H;�H;"�H;O�H;c�H;O�H;j�H;��H;��H;��H;��H;��H;��H;r�H;X�H;@�H;�H;��H;Y�H;�H;��H;*�H;��H;�H;��H;��H;R�H;��H;@�H;��H;p�H;�H;��H;��H;      o�H;�H;��H;��H;��H;�H;��H;{�H;9�H;��H;��H;m�H;&�H;��H;��H;,�H;��H;�H;w�H;��H;��H;1�H;L�H;l�H;��H;}�H;�H;l�H;k�H;h�H;E�H;=�H;C�H;-�H;�H;#�H;)�H;#�H;�H;-�H;C�H;=�H;E�H;h�H;k�H;l�H;�H;}�H;��H;l�H;L�H;1�H;��H;��H;w�H;�H;��H;,�H;��H;��H;&�H;m�H;��H;��H;9�H;{�H;��H;�H;��H;��H;��H;�H;      ��H;��H;�H;��H;)�H;��H;��H;��H;��H;��H;��H;�H;�H;�H;��H;��H;h�H;�H;��H;��H;l�H;��H;��H;,�H;=�H;C�H;\�H;k�H;j�H;X�H;E�H;C�H;G�H;C�H;"�H;#�H;S�H;#�H;"�H;C�H;G�H;C�H;E�H;X�H;j�H;k�H;\�H;C�H;=�H;,�H;��H;��H;l�H;��H;��H;�H;h�H;��H;��H;�H;�H;�H;��H;��H;��H;��H;��H;��H;)�H;��H;�H;��H;      ��H;��H;�H;��H;��H;��H;(�H;��H;�H;��H;�H;��H;��H;R�H;��H;��H;��H;��H;a�H;$�H;��H;�H;��H;��H;��H;.�H;<�H;B�H;S�H;I�H;T�H;Z�H;C�H;=�H;O�H;4�H;+�H;4�H;O�H;=�H;C�H;Z�H;T�H;I�H;S�H;B�H;<�H;.�H;��H;��H;��H;�H;��H;$�H;a�H;��H;��H;��H;��H;R�H;��H;��H;�H;��H;�H;��H;(�H;��H;��H;��H;�H;��H;      h�H;��H;<�H;I�H;��H;.�H;�H;��H;�H;N�H;u�H;��H;��H;|�H;A�H;��H;w�H;��H;��H;��H;��H;4�H;��H;(�H;��H;��H;��H;�H;6�H;J�H;a�H;T�H;E�H;E�H;c�H;U�H;6�H;U�H;c�H;E�H;E�H;T�H;a�H;J�H;6�H;�H;��H;��H;��H;(�H;��H;4�H;��H;��H;��H;��H;w�H;��H;A�H;|�H;��H;��H;u�H;N�H;�H;��H;�H;.�H;��H;I�H;<�H;��H;      ��H;ܶH;��H;7�H;)�H;��H;R�H;M�H;V�H;�H;��H;��H;��H;m�H;��H;�H;:�H;�H;��H;��H;��H;�H;��H;~�H;�H;R�H;��H;��H;�H;+�H;J�H;I�H;X�H;h�H;O�H;a�H;{�H;a�H;O�H;h�H;X�H;I�H;J�H;+�H;�H;��H;��H;R�H;�H;~�H;��H;�H;��H;��H;��H;�H;:�H;�H;��H;m�H;��H;��H;��H;�H;V�H;M�H;R�H;��H;)�H;7�H;��H;ܶH;      3�H;ϠH;[�H;äH;��H;��H;��H;�H;��H;H�H;��H;I�H;a�H;I�H;�H;2�H;��H;g�H;��H;��H;<�H;~�H;��H;��H;8�H;��H;[�H;��H;��H;�H;6�H;S�H;j�H;k�H;j�H;u�H;u�H;u�H;j�H;k�H;j�H;S�H;6�H;�H;��H;��H;[�H;��H;8�H;��H;��H;~�H;<�H;��H;��H;g�H;��H;2�H;�H;I�H;a�H;I�H;��H;H�H;��H;�H;��H;��H;��H;äH;[�H;ϠH;      �kH;ZmH;�qH;�xH;r�H;ȊH;�H;ʜH;��H;��H;��H;�H;%�H;��H;��H;K�H;Y�H;��H;��H;w�H;��H;��H;�H;G�H;T�H;�H;��H;B�H;��H;��H;�H;B�H;k�H;l�H;��H;��H;��H;��H;��H;l�H;k�H;B�H;�H;��H;��H;B�H;��H;�H;T�H;G�H;�H;��H;��H;w�H;��H;��H;Y�H;K�H;��H;��H;%�H;�H;��H;��H;��H;ʜH;�H;ȊH;r�H;�xH;�qH;ZmH;      =�G;��G;/�G;��G;�H;�/H;�KH;?eH;_{H;i�H;m�H;c�H;o�H;��H;ľH;2�H;��H;��H;��H;h�H;d�H;��H;"�H;��H;�H;9�H;�H;��H;[�H;��H;��H;<�H;\�H;�H;��H;��H;��H;��H;��H;�H;\�H;<�H;��H;��H;[�H;��H;�H;9�H;�H;��H;"�H;��H;d�H;h�H;��H;��H;��H;2�H;ľH;��H;o�H;c�H;m�H;i�H;_{H;?eH;�KH;�/H;�H;��G;/�G;��G;      UHF;3TF;RvF;F�F;��F;�7G;��G;��G;�H;�<H;/eH;o�H;H;�H;��H;θH;��H;��H;T�H;Q�H;Y�H;��H;w�H;��H;��H;	�H;9�H;�H;��H;R�H;��H;.�H;C�H;}�H;��H;��H;��H;��H;��H;}�H;C�H;.�H;��H;R�H;��H;�H;9�H;	�H;��H;��H;w�H;��H;Y�H;Q�H;T�H;��H;��H;θH;��H;�H;H;o�H;/eH;�<H;�H;��G;��G;�7G;��F;F�F;RvF;3TF;      �B;-�B;�C;ԏC;�/D;��D;0�E;�HF;��F;FiG;R�G;s#H;�[H;/�H;��H;�H;H�H;μH;��H;d�H;��H;��H;�H;5�H;��H;��H;�H;T�H;8�H;�H;��H;��H;=�H;��H;��H;��H;��H;��H;��H;��H;=�H;��H;��H;�H;8�H;T�H;�H;��H;��H;5�H;�H;��H;��H;d�H;��H;μH;H�H;�H;��H;/�H;�[H;s#H;R�G;FiG;��F;�HF;0�E;��D;�/D;ԏC;�C;-�B;      C�:;[�:;��;;&�<;3>;�?;EIA;��B;CED;5{E;VvF;�7G;��G;p&H; eH;s�H;^�H;m�H;��H;��H;�H;9�H;�H;��H;5�H;��H;��H;G�H;��H;~�H;(�H;��H;,�H;l�H;��H;��H;��H;��H;��H;l�H;,�H;��H;(�H;~�H;��H;G�H;��H;��H;5�H;��H;�H;9�H;�H;��H;��H;m�H;^�H;s�H; eH;p&H;��G;�7G;VvF;5{E;CED;��B;EIA;�?;3>;&�<;��;;[�:;      *;��*;�,;�c.;�X1;#�4;D+8;ӊ;;}�>;IA;iwC;�)E;kF;�MG;'�G;DH;"{H;@�H;��H;?�H;R�H;Y�H;��H;�H;�H;w�H;"�H;�H;��H;��H;��H;��H;��H;L�H;��H;��H;��H;��H;��H;L�H;��H;��H;��H;��H;��H;�H;"�H;w�H;�H;�H;��H;Y�H;R�H;?�H;��H;@�H;"{H;DH;'�G;�MG;kF;�)E;iwC;IA;}�>;ӊ;;D+8;#�4;�X1;�c.;�,;��*;      ��
;��;I�;[;��;6`;�C&;�-;�C3;t�8;>H=;��@;�C;c{E;��F;�G;k#H;+mH;��H;>�H;��H;��H;Y�H;9�H;��H;��H;��H;��H;~�H;�H;4�H;�H;��H;1�H;r�H;��H;��H;��H;r�H;1�H;��H;�H;4�H;�H;~�H;��H;��H;��H;��H;9�H;Y�H;��H;��H;>�H;��H;+mH;k#H;�G;��F;c{E;�C;��@;>H=;t�8;�C3;�-;�C&;6`;��;[;I�;��;      [�:���:��:Ѳ�:���:NO�:�z;h';3�;�}(;�X1;6t8;��=;Z�A;��D;%HF;�bG;�H;=cH;��H;m�H;��H;R�H;�H;��H;Y�H;d�H;��H;<�H;��H;��H;��H;l�H;��H;X�H;��H;��H;��H;X�H;��H;l�H;��H;��H;��H;<�H;��H;d�H;Y�H;��H;�H;R�H;��H;m�H;��H;=cH;�H;�bG;%HF;��D;Z�A;��=;6t8;�X1;�}(;3�;h';�z;NO�:���:Ѳ�:��:���:      "�R�� �l�7�r<^9��:L�X:���:���:�O�:=�;6�;�);�C3;��:;� @;�C;j�E;8G;��G;�_H;��H;>�H;?�H;��H;d�H;Q�H;h�H;w�H;��H;��H;��H;$�H;��H;��H;@�H;{�H;{�H;{�H;@�H;��H;��H;$�H;��H;��H;��H;w�H;h�H;Q�H;d�H;��H;?�H;>�H;��H;�_H;��G;8G;j�E;�C;� @;��:;�C3;�);6�;=�;�O�:���:���:L�X:��:r<^9l�7�� �      ��)���$�����������A�\�S���N�9�1j:_��:���:ڃ;�� ;%d.;+8;��>;pC;��E;�(G;��G;=cH;��H;��H;��H;��H;T�H;��H;��H;��H;��H;��H;a�H;��H;w�H;�H;I�H;b�H;I�H;�H;w�H;��H;a�H;��H;��H;��H;��H;��H;T�H;��H;��H;��H;��H;=cH;��G;�(G;��E;pC;��>;+8;%d.;�� ;ڃ;���:_��:�1j:�N�9S��A�\�������������$�      r�ѻ�ͻP���mG�������d�+�$��JɺЇ!��C^9��r:���:_0;x�;k�*;�Y6;>;n�B;��E;8G;�H;+mH;@�H;m�H;μH;��H;��H;��H;g�H;�H;��H;��H;�H;�H;��H;�H;<�H;�H;��H;�H;�H;��H;��H;�H;g�H;��H;��H;��H;μH;m�H;@�H;+mH;�H;8G;��E;n�B;>;�Y6;k�*;x�;_0;���:��r:�C^9Ї!��Jɺ+�$���d����mG��P����ͻ      ��I�1�E��(;��O*�����<��@GĻ��t@�JҺ���:�:�O�:N�; ~(;R�5;>;pC;j�E;�bG;k#H;"{H;^�H;H�H;��H;��H;Y�H;��H;:�H;w�H;��H;h�H;��H;Y�H;��H;�H;��H;Y�H;��H;h�H;��H;w�H;:�H;��H;Y�H;��H;��H;H�H;^�H;"{H;k#H;�bG;j�E;pC;>;R�5; ~(;N�;�O�:�:��:���JҺt@���@GĻ�<������O*��(;�1�E�      &p��\x��ע��R��%��o�`��7�F��H�ѻ-��̃$��ǅ���09�:���:�; ~(;�Y6;��>;�C;%HF;�G;DH;s�H;�H;θH;2�H;K�H;2�H;�H;��H;��H;��H;,�H;�H;��H;��H;��H;�H;,�H;��H;��H;��H;�H;2�H;K�H;2�H;θH;�H;s�H;DH;�G;%HF;�C;��>;�Y6; ~(;�;���:�:��09�ǅ�̃$�-��H�ѻF���7�o�`�%���R��ע�\x��      &]� �%#�����u�ټ�ɺ������
v��(;�ר�c^��Q6R����
7����:���:N�;k�*;+8;� @;��D;��F;'�G; eH;��H;��H;ľH;��H;�H;��H;A�H;��H;��H;��H;��H;B�H;u�H;B�H;��H;��H;��H;��H;A�H;��H;�H;��H;ľH;��H;��H; eH;'�G;��F;��D;� @;+8;k�*;N�;���:���:
7����Q6R�c^��ר��(;��
v������ɺ�u�ټ����%#� �      ��_�\�<Q��f@�t +��5�����P�ļs�\�`����bͻgk��Iɺ
7��:�O�:x�;%d.;��:;Z�A;c{E;�MG;p&H;/�H;�H;��H;��H;I�H;m�H;|�H;R�H;�H;��H;*�H;��H;�H;��H;*�H;��H;�H;R�H;|�H;m�H;I�H;��H;��H;�H;/�H;p&H;�MG;c{E;Z�A;��:;%d.;x�;�O�:�:
7��Iɺgk�bͻ���\�`�s�P�ļ�����5�t +��f@�<Q�\�      �@���R��ڟ�绒�C����_�:�������$p���vz��O*�5ֻgk������09�:_0;�� ;�C3;��=;�C;kF;��G;�[H;H;o�H;%�H;a�H;��H;��H;��H;�H;&�H;��H;n�H;��H;n�H;��H;&�H;�H;��H;��H;��H;a�H;%�H;o�H;H;�[H;��G;kF;�C;��=;�C3;�� ;_0;�:��09���gk�5ֻ�O*��vz�$p����輙��:���_�C��绒�ڟ��R��      �` �j.��m��ڽ�b��gr��O��\�m +�� ��ɺ�=��O*�bͻQ6R��ǅ���:���:ڃ;�);6t8;��@;�)E;�7G;s#H;o�H;c�H;�H;I�H;��H;��H;��H;�H;m�H;�H; �H;>�H; �H;�H;m�H;�H;��H;��H;��H;I�H;�H;c�H;o�H;s#H;�7G;�)E;��@;6t8;�);ڃ;���:��:�ǅ�Q6R�bͻ�O*�=��ɺ�� �m +�\�O��gr���b����ڽm��j.��      �-=�1�9��k/�"�����i��y�Ľ�!��Tys�4�6�#��ɺ��vz����c^��̃$������r:���:6�;�X1;>H=;iwC;VvF;R�G;/eH;m�H;��H;��H;��H;u�H;�H;��H;��H;��H;��H;��H;��H;��H;��H;��H;�H;u�H;��H;��H;��H;m�H;/eH;R�G;VvF;iwC;>H=;�X1;6�;���:��r:���̃$�c^������vz��ɺ�#�4�6�Tys��!��y�Ľi���"���k/�1�9�      �(��;l���.}�&ce�jPH���(�o
���ڽ�R����{�4�6�� �$p��\�`�ר�-��JҺ�C^9_��:=�;�}(;t�8;IA;5{E;FiG;�<H;i�H;��H;H�H;�H;N�H;��H;��H;��H;��H;�H;i�H;�H;��H;��H;��H;��H;N�H;�H;H�H;��H;i�H;�<H;FiG;5{E;IA;t�8;�}(;=�;_��:�C^9JҺ-��ר�\�`�$p��� �4�6���{��R����ڽo
���(�jPH�&ce��.}�;l��      �iþGD��)o���������� �i��-=�[t����R��Tys�m +����s񗼗(;�H�ѻt@�Ї!��1j:�O�:3�;�C3;}�>;CED;��F;�H;_{H;��H;��H;V�H;�H;�H;��H;9�H;R�H;��H;�H;��H;R�H;9�H;��H;�H;�H;V�H;��H;��H;_{H;�H;��F;CED;}�>;�C3;3�;�O�:�1j:Ї!�t@�H�ѻ�(;�s����m +�Tys��R����[t��-=� �i���������)o��GD��      ���
������޾HD���A���.}��D�[t���ڽ�!��\����P�ļ�
v�F�����Jɺ�N�9���:h';�-;ӊ;;��B;�HF;��G;?eH;ʜH;�H;M�H;��H;��H;��H;{�H;��H;�H;��H;�H;��H;{�H;��H;��H;��H;M�H;�H;ʜH;?eH;��G;�HF;��B;ӊ;;�-;h';���:�N�9�Jɺ��F���
v�P�ļ���\��!����ڽ[t��D��.}��A��HD���޾�����
�      ��7�Õ3��f'���\���о�����.}��-=�o
�y�ĽO��:����������7�@GĻ+�$�S�����:�z;�C&;D+8;EIA;0�E;��G;�KH;�H;��H;R�H;�H;(�H;��H;��H;@�H;��H;5�H;��H;@�H;��H;��H;(�H;�H;R�H;��H;�H;�KH;��G;0�E;EIA;D+8;�C&;�z;���:S��+�$�@GĻ�7���������:�O��y�Ľo
��-=��.}������о�\����f'�Õ3�      Io�PXi�s"Y���@�@�#��
��о�A�� �i���(�i��gr����_��5��ɺ�o�`��<����d�A�\�L�X:NO�:6`;#�4;�?;��D;�7G;�/H;ȊH;��H;��H;.�H;��H;��H;�H;��H;-�H;��H;-�H;��H;�H;��H;��H;.�H;��H;��H;ȊH;�/H;�7G;��D;�?;#�4;6`;NO�:L�X:A�\���d��<��o�`��ɺ��5���_�gr��i����(� �i��A���о�
�@�#���@�s"Y�PXi�      &����������Io��!J�@�#��\��HD������jPH�����b��C��t +�u�ټ%��������������:���:��;�X1;3>;�/D;��F;�H;r�H;��H;)�H;��H;��H;)�H;��H;p�H;��H;~�H;��H;p�H;��H;)�H;��H;��H;)�H;��H;r�H;�H;��F;�/D;3>;�X1;��;���:��:����������%��u�ټt +�C���b�����jPH�����HD���\��@�#��!J�Io��������      2^������b���Io���@���޾����&ce�"����ڽ绒��f@������R���O*�mG�����r<^9Ѳ�:[;�c.;&�<;ԏC;F�F;��G;�xH;äH;7�H;I�H;��H;��H;��H;�H;��H;6�H;��H;�H;��H;��H;��H;I�H;7�H;äH;�xH;��G;F�F;ԏC;&�<;�c.;[;Ѳ�:r<^9���mG���O*��R�������f@�绒���ڽ"��&ce������޾���@�Io�b�������      �aǿ֊¿���������s"Y��f'�����)o���.}��k/�m��ڟ�<Q�%#�ע��(;�P������l�7���:I�;�,;��;;�C;RvF;/�G;�qH;[�H;��H;<�H;�H;�H;��H;��H;j�H;��H;j�H;��H;��H;�H;�H;<�H;��H;[�H;�qH;/�G;RvF;�C;��;;�,;I�;��:l�7����P����(;�ע�%#�<Q�ڟ�m���k/��.}�)o�������f'�s"Y����������֊¿      %�ֿ5pѿ֊¿������PXi�Õ3��
�GD��;l��1�9�j.���R��\� �\x��1�E��ͻ��$�� ����:��;��*;[�:;-�B;3TF;��G;ZmH;ϠH;ܶH;��H;��H;��H;�H;��H;<�H;��H;<�H;��H;�H;��H;��H;��H;ܶH;ϠH;ZmH;��G;3TF;-�B;[�:;��*;��;���:� ���$��ͻ1�E�\x�� �\��R��j.��1�9�;l��GD���
�Õ3�PXi�������֊¿5pѿ      �?��ph��1v��� ��$�X��O/�#y�-�;Ѱ��j+X�����ѽ����Gn;�>�＿����B(�暩���� �e9��:^;Y.;��<;�VC;?ZF;�G;4/H;tiH;X�H;s�H;��H;E�H;��H;~�H;��H;��H;��H;~�H;��H;E�H;��H;s�H;X�H;tiH;4/H;�G;?ZF;�VC;��<;Y.;^;��: �e9���暩��B(�����>��Gn;�������ѽ��j+X�Ѱ��-�;#y��O/�$�X�� ��1v��ph��      ph��"���V�����y�EvS�aM+��v� 9ɾ�����T�]��[ν����`\8�����x���%�\��������9A,�:��;�.;M�<; nC;�cF;�G;�0H;!jH;ǋH;ѣH;��H;��H;��H;��H;��H;��H;��H;��H;��H;��H;��H;ѣH;ǋH;!jH;�0H;�G;�cF; nC;M�<;�.;��;A,�:��9���\����%��x�����`\8������[ν]��T����� 9ɾ�v�aM+�EvS���y�V���"���      1v��V���L ��M�h�%E�I��R���i㼾n���nH�È�a�ý�Ȅ��s/��o༼#�����4J���к��9"f�:Ml;�0;P\=; �C;5�F;��G;Q5H;^lH;G�H;ϤH;��H;�H;b�H;��H;#�H; �H;#�H;��H;b�H;�H;��H;ϤH;G�H;^lH;Q5H;��G;5�F; �C;P\=;�0;Ml;"f�:��9�к4J������#���o��s/��Ȅ�a�ýÈ��nH�n��i㼾R���I��%E�M�h�L ��V���      � ����y�M�h�ބN��O/����-�߾�A���*|�ؕ6�a}��㳽KSt�(�!�Wrμ(F{��_�Y��h����:���:VZ;2;�N>;�D;��F;��G;J<H;�oH;��H;t�H;��H;��H;��H;��H;��H;�H;��H;��H;��H;��H;��H;t�H;��H;�oH;J<H;��G;��F;�D;�N>;2;VZ;���:�:h���Y���_�(F{�Wrμ(�!�KSt��㳽a}�ؕ6��*|��A��-�߾����O/�ބN�M�h���y�      $�X�EvS�%E��O/��S�1W����������4S\�� �q�&�����Y�h��������]�}���T�b��Y���Y:~~�:�_;��4;�?;|�D;�F;/�G;5EH;tH;�H;��H;��H;3�H;��H;D�H;7�H;�H;7�H;D�H;��H;3�H;��H;��H;�H;tH;5EH;/�G;�F;|�D;�?;��4;�_;~~�:��Y:�Y�T�b�}�����]�����h����Y�&���q�� �4S\���������1W���S��O/�%E�EvS�      �O/�aM+�I�����1W�� 9ɾ0���Mw�� :�Y��_�ý�L��Dn;�>���bv���E<��˻)�-����x�:^;%;�7;��@;V4E;�!G;,�G;hOH;0zH;��H;��H;��H;��H;�H;2�H;�H;��H;�H;2�H;�H;��H;��H;��H;��H;0zH;hOH;,�G;�!G;V4E;��@;�7;%;^;�x�:��)�-��˻�E<�bv��>���Dn;��L��_�ýY��� :��Mw�0�� 9ɾ1W�����I��aM+�      #y��v�R���-�߾����0��1����nH���(Ὁu��r�d�O�Prμ="�����	��3���k89u:�:��;+;�{:;�6B;)�E;EaG;�H;ZH;��H;L�H;ĮH;�H;e�H;e�H;*�H;��H;��H;��H;*�H;e�H;e�H;�H;ĮH;L�H;��H;ZH;�H;EaG;)�E;�6B;�{:;+;��;u:�:�k893��	�����="��PrμO�r�d��u��(����nH�1���0������-�߾R����v�      -�; 9ɾi㼾�A�������Mw��nH�����Z��㳽����Z\8�P#�������]N�J��.�b�ZJx�v5:��:��;8�0;u\=;u�C;�ZF;�G;)H;eH;��H;F�H;g�H;��H;6�H;��H;P�H;��H;��H;��H;P�H;��H;6�H;��H;g�H;F�H;��H;eH;)H;�G;�ZF;u�C;u\=;8�0;��;��:v5:ZJx�.�b�J���]N�����P#��Z\8������㳽�Z񽞯��nH��Mw������A��i㼾 9ɾ      Ѱ������n���*|�4S\�� :����Z�U$������K�c���Oļ����������y&�1��N.�:/^;��#;G6;��?;,�D;��F;��G;)?H;�oH;�H;��H;9�H;q�H;J�H;��H;��H;��H;��H;��H;��H;��H;J�H;q�H;9�H;��H;�H;�oH;)?H;��G;��F;,�D;��?;G6;��#;/^;N.�:1��y&������������Oļc���K����U$���Z���� :�4S\��*|�n������      j+X��T��nH�ؕ6�� �Y��(��㳽����mR����ټ�����E<��?ݻbd\�c ��":�c�:7�;y�,;��:;�6B;̱E;�KG;iH;�RH;�zH;��H;
�H;9�H;_�H;n�H;+�H;��H;�H;��H;�H;��H;+�H;n�H;_�H;9�H;
�H;��H;�zH;�RH;iH;�KG;̱E;�6B;��:;y�,;7�;�c�:":c ��bd\��?ݻ�E<������ټ���mR�����㳽(�Y��� �ؕ6��nH��T�      ��]�È�a}�q�_�ý�u�������K����o�Wv���&R���f^����>@���:�A;�";��4;��>;�D;��F;,�G; )H;�cH;��H;5�H;��H;N�H;M�H;��H;��H;<�H;(�H;��H;(�H;<�H;��H;��H;M�H;N�H;��H;5�H;��H;�cH; )H;,�G;��F;�D;��>;��4;�";�A;��:>@���f^�����&R�Wv���o����K������u��_�ýq�a}�È�]�      ��ѽ�[νa�ý�㳽&����L��r�d�Z\8�c���ټWv����Y��_����z��]���Y:?��:�l;r-;Q�:;��A;qnE;�!G;��G;�FH;�rH;�H;��H;�H;J�H;5�H;��H;��H;��H;B�H;�H;B�H;��H;��H;��H;5�H;J�H;�H;��H;�H;�rH;�FH;��G;�!G;qnE;��A;Q�:;r-;�l;?��:��Y:]�z������_���Y�Wv���ټc��Z\8�r�d��L��&����㳽a�ý�[ν      ���������Ȅ�KSt���Y�Dn;�O�P#���Oļ�����&R��_������N3�0�Y�,2:�:8�;@?&;(G6;�W?;�D;fwF;�G;c H;�]H;��H;�H;�H;a�H;#�H;�H;��H;'�H;��H;i�H;$�H;i�H;��H;'�H;��H;�H;#�H;a�H;�H;�H;��H;�]H;c H;�G;fwF;�D;�W?;(G6;@?&;8�;�:,2:0�Y��N3������_��&R������OļP#��O�Dn;���Y�KSt��Ȅ�����      Gn;�`\8��s/�(�!�h��>���Prμ��������E<�������N3��Ix�_�9��:T^;� ;~2;��<;.�B;�E;e4G;1�G;^EH;�pH;��H;h�H;ϳH;k�H;��H;��H;�H;��H;1�H;��H;�H;��H;1�H;��H;�H;��H;��H;k�H;ϳH;h�H;��H;�pH;^EH;1�G;e4G;�E;.�B;��<;~2;� ;T^;��:_�9�Ix��N3�������E<��������Prμ>���h��(�!��s/�`\8�      >�Ｘ���o�Wrμ����bv��="���]N�����?ݻf^��z��0�Y�_�9��:���:B�;��.;�{:;2>A;��D;`�F;ߵG;
)H;D`H;5�H;��H;�H;R�H;5�H;R�H;t�H;�H;.�H;k�H;��H;��H;��H;k�H;.�H;�H;t�H;R�H;5�H;R�H;�H;��H;5�H;D`H;
)H;ߵG;`�F;��D;2>A;�{:;��.;B�;���:��:_�90�Y�z��f^���?ݻ����]N�="��bv������Wrμ�o༸��      �����x���#��(F{���]��E<����J�뻲���bd\���]�,2:��:���:�Z;��,;/�8;` @;0D;�ZF;PzG;
H;iOH;=uH;�H;[�H;�H;B�H;z�H;��H;��H;��H;��H;��H;��H;��H;��H;��H;��H;��H;��H;��H;z�H;B�H;�H;[�H;�H;=uH;iOH;
H;PzG;�ZF;0D;` @;/�8;��,;�Z;���:��:,2:]���bd\�����J�뻛���E<���]�(F{��#���x��      �B(��%�����_�}����˻	��.�b�y&�c ��>@���Y:�:T^;B�;��,;Z_8;��?;��C;�F;FG;t�G;?H;FjH;#�H; �H;
�H;k�H;��H;~�H;��H;/�H;��H;��H;��H;��H;��H;��H;��H;��H;��H;/�H;��H;~�H;��H;k�H;
�H; �H;#�H;FjH;?H;t�G;FG;�F;��C;��?;Z_8;��,;B�;T^;�:��Y:>@�c ��y&�.�b�	���˻}����_�����%�      暩�\���4J��Y��T�b�)�-�3��ZJx�1��":��:?��:8�;� ;��.;/�8;��?;1�C;�E;e"G;�G;1H;aH;gH;��H;��H;��H;��H;s�H;(�H;I�H;J�H;��H;(�H;��H;G�H;��H;G�H;��H;(�H;��H;J�H;I�H;(�H;s�H;��H;��H;��H;��H;gH;aH;1H;�G;e"G;�E;1�C;��?;/�8;��.;� ;8�;?��:��:":1��ZJx�3��)�-�T�b�Y��4J��\���      �����뺸кh����Y����k89v5:N.�:�c�:�A;�l;@?&;~2;�{:;` @;��C;�E;�G;�G;}'H;ZH;�yH;W�H;��H;��H;{�H;��H;��H;l�H;��H;
�H;[�H;<�H;W�H;
�H;��H;
�H;W�H;<�H;[�H;
�H;��H;l�H;��H;��H;{�H;��H;��H;W�H;�yH;ZH;}'H;�G;�G;�E;��C;` @;�{:;~2;@?&;�l;�A;�c�:N.�:v5:�k89���Y�h����к���       �e9��9��9�:��Y:�x�:u:�:��:/^;7�;�";r-;(G6;��<;2>A;0D;�F;e"G;�G;$H;~VH;�uH;��H;X�H;b�H;��H;!�H;��H;��H;E�H;��H;��H;��H;6�H;�H;��H;�H;��H;�H;6�H;��H;��H;��H;E�H;��H;��H;!�H;��H;b�H;X�H;��H;�uH;~VH;$H;�G;e"G;�F;0D;2>A;��<;(G6;r-;�";7�;/^;��:u:�:�x�:��Y:�:��9��9      ��:A,�:"f�:���:~~�:^;��;��;��#;y�,;��4;Q�:;�W?;.�B;��D;�ZF;FG;�G;}'H;~VH;�tH;��H;.�H;�H;<�H;	�H;��H;��H;��H;��H;��H;��H;��H;��H;��H;^�H;b�H;^�H;��H;��H;��H;��H;��H;��H;��H;��H;��H;	�H;<�H;�H;.�H;��H;�tH;~VH;}'H;�G;FG;�ZF;��D;.�B;�W?;Q�:;��4;y�,;��#;��;��;^;~~�:���:"f�:A,�:      ^;��;Ml;VZ;�_;%;+;8�0;G6;��:;��>;��A;�D;�E;`�F;PzG;t�G;1H;ZH;�uH;��H;g�H;ܫH;߷H;��H;e�H;��H;��H;��H;��H;H�H;G�H;��H;��H;p�H;��H;��H;��H;p�H;��H;��H;G�H;H�H;��H;��H;��H;��H;e�H;��H;߷H;ܫH;g�H;��H;�uH;ZH;1H;t�G;PzG;`�F;�E;�D;��A;��>;��:;G6;8�0;+;%;�_;VZ;Ml;��;      Y.;�.;�0;2;��4;�7;�{:;u\=;��?;�6B;�D;qnE;fwF;e4G;ߵG;
H;?H;aH;�yH;��H;.�H;ܫH;`�H;��H;�H;��H;��H;�H;)�H;��H;��H;h�H;c�H;O�H;��H;(�H;P�H;(�H;��H;O�H;c�H;h�H;��H;��H;)�H;�H;��H;��H;�H;��H;`�H;ܫH;.�H;��H;�yH;aH;?H;
H;ߵG;e4G;fwF;qnE;�D;�6B;��?;u\=;�{:;�7;��4;2;�0;�.;      ��<;M�<;P\=;�N>;�?;��@;�6B;u�C;,�D;̱E;��F;�!G;�G;1�G;
)H;iOH;FjH;gH;W�H;X�H;�H;߷H;��H;H�H;H�H;E�H;W�H;��H;,�H;A�H;�H;�H;�H;��H;H�H;��H;��H;��H;H�H;��H;�H;�H;�H;A�H;,�H;��H;W�H;E�H;H�H;H�H;��H;߷H;�H;X�H;W�H;gH;FjH;iOH;
)H;1�G;�G;�!G;��F;̱E;,�D;u�C;�6B;��@;�?;�N>;P\=;M�<;      �VC; nC; �C;�D;|�D;V4E;)�E;�ZF;��F;�KG;,�G;��G;c H;^EH;D`H;=uH;#�H;��H;��H;b�H;<�H;��H;�H;H�H;�H;�H;O�H;��H;��H;��H;��H;��H;��H;=�H;��H;��H;��H;��H;��H;=�H;��H;��H;��H;��H;��H;��H;O�H;�H;�H;H�H;�H;��H;<�H;b�H;��H;��H;#�H;=uH;D`H;^EH;c H;��G;,�G;�KG;��F;�ZF;)�E;V4E;|�D;�D; �C; nC;      ?ZF;�cF;5�F;��F;�F;�!G;EaG;�G;��G;iH; )H;�FH;�]H;�pH;5�H;�H; �H;��H;��H;��H;	�H;e�H;��H;E�H;�H;5�H;��H;��H;t�H;��H;��H;��H;,�H;~�H;��H;�H;�H;�H;��H;~�H;,�H;��H;��H;��H;t�H;��H;��H;5�H;�H;E�H;��H;e�H;	�H;��H;��H;��H; �H;�H;5�H;�pH;�]H;�FH; )H;iH;��G;�G;EaG;�!G;�F;��F;5�F;�cF;      �G;�G;��G;��G;/�G;,�G;�H;)H;)?H;�RH;�cH;�rH;��H;��H;��H;[�H;
�H;��H;{�H;!�H;��H;��H;��H;W�H;O�H;��H;��H;J�H;��H;��H;j�H; �H;}�H;��H;�H;:�H;Y�H;:�H;�H;��H;}�H; �H;j�H;��H;��H;J�H;��H;��H;O�H;W�H;��H;��H;��H;!�H;{�H;��H;
�H;[�H;��H;��H;��H;�rH;�cH;�RH;)?H;)H;�H;,�G;/�G;��G;��G;�G;      4/H;�0H;Q5H;J<H;5EH;hOH;ZH;eH;�oH;�zH;��H;�H;�H;h�H;�H;�H;k�H;��H;��H;��H;��H;��H;�H;��H;��H;��H;J�H;��H;e�H;S�H;�H;i�H;��H;�H;E�H;[�H;L�H;[�H;E�H;�H;��H;i�H;�H;S�H;e�H;��H;J�H;��H;��H;��H;�H;��H;��H;��H;��H;��H;k�H;�H;�H;h�H;�H;�H;��H;�zH;�oH;eH;ZH;hOH;5EH;J<H;Q5H;�0H;      tiH;!jH;^lH;�oH;tH;0zH;��H;��H;�H;��H;5�H;��H;�H;ϳH;R�H;B�H;��H;s�H;��H;��H;��H;��H;)�H;,�H;��H;t�H;��H;e�H;[�H;��H;Y�H;��H;��H;5�H;e�H;o�H;b�H;o�H;e�H;5�H;��H;��H;Y�H;��H;[�H;e�H;��H;t�H;��H;,�H;)�H;��H;��H;��H;��H;s�H;��H;B�H;R�H;ϳH;�H;��H;5�H;��H;�H;��H;��H;0zH;tH;�oH;^lH;!jH;      X�H;ǋH;G�H;��H;�H;��H;L�H;F�H;��H;
�H;��H;�H;a�H;k�H;5�H;z�H;~�H;(�H;l�H;E�H;��H;��H;��H;A�H;��H;��H;��H;S�H;��H;J�H;��H;��H;6�H;]�H;h�H;��H;��H;��H;h�H;]�H;6�H;��H;��H;J�H;��H;S�H;��H;��H;��H;A�H;��H;��H;��H;E�H;l�H;(�H;~�H;z�H;5�H;k�H;a�H;�H;��H;
�H;��H;F�H;L�H;��H;�H;��H;G�H;ǋH;      s�H;ѣH;ϤH;t�H;��H;��H;ĮH;g�H;9�H;9�H;N�H;J�H;#�H;��H;R�H;��H;��H;I�H;��H;��H;��H;H�H;��H;�H;��H;��H;j�H;�H;Y�H;��H;��H;)�H;a�H;o�H;��H;��H;��H;��H;��H;o�H;a�H;)�H;��H;��H;Y�H;�H;j�H;��H;��H;�H;��H;H�H;��H;��H;��H;I�H;��H;��H;R�H;��H;#�H;J�H;N�H;9�H;9�H;g�H;ĮH;��H;��H;t�H;ϤH;ѣH;      ��H;��H;��H;��H;��H;��H;�H;��H;q�H;_�H;M�H;5�H;�H;��H;t�H;��H;/�H;J�H;
�H;��H;��H;G�H;h�H;�H;��H;��H; �H;i�H;��H;��H;)�H;A�H;k�H;��H;��H;��H;��H;��H;��H;��H;k�H;A�H;)�H;��H;��H;i�H; �H;��H;��H;�H;h�H;G�H;��H;��H;
�H;J�H;/�H;��H;t�H;��H;�H;5�H;M�H;_�H;q�H;��H;�H;��H;��H;��H;��H;��H;      E�H;��H;�H;��H;3�H;��H;e�H;6�H;J�H;n�H;��H;��H;��H;�H;�H;��H;��H;��H;[�H;��H;��H;��H;c�H;�H;��H;,�H;}�H;��H;��H;6�H;a�H;k�H;{�H;��H;��H;��H;��H;��H;��H;��H;{�H;k�H;a�H;6�H;��H;��H;}�H;,�H;��H;�H;c�H;��H;��H;��H;[�H;��H;��H;��H;�H;�H;��H;��H;��H;n�H;J�H;6�H;e�H;��H;3�H;��H;�H;��H;      ��H;��H;b�H;��H;��H;�H;e�H;��H;��H;+�H;��H;��H;'�H;��H;.�H;��H;��H;(�H;<�H;6�H;��H;��H;O�H;��H;=�H;~�H;��H;�H;5�H;]�H;o�H;��H;��H;��H;��H;��H;��H;��H;��H;��H;��H;��H;o�H;]�H;5�H;�H;��H;~�H;=�H;��H;O�H;��H;��H;6�H;<�H;(�H;��H;��H;.�H;��H;'�H;��H;��H;+�H;��H;��H;e�H;�H;��H;��H;b�H;��H;      ~�H;��H;��H;��H;D�H;2�H;*�H;P�H;��H;��H;<�H;��H;��H;1�H;k�H;��H;��H;��H;W�H;�H;��H;p�H;��H;H�H;��H;��H;�H;E�H;e�H;h�H;��H;��H;��H;��H;��H;��H;��H;��H;��H;��H;��H;��H;��H;h�H;e�H;E�H;�H;��H;��H;H�H;��H;p�H;��H;�H;W�H;��H;��H;��H;k�H;1�H;��H;��H;<�H;��H;��H;P�H;*�H;2�H;D�H;��H;��H;��H;      ��H;��H;#�H;��H;7�H;�H;��H;��H;��H;�H;(�H;B�H;i�H;��H;��H;��H;��H;G�H;
�H;��H;^�H;��H;(�H;��H;��H;�H;:�H;[�H;o�H;��H;��H;��H;��H;��H;��H;��H;��H;��H;��H;��H;��H;��H;��H;��H;o�H;[�H;:�H;�H;��H;��H;(�H;��H;^�H;��H;
�H;G�H;��H;��H;��H;��H;i�H;B�H;(�H;�H;��H;��H;��H;�H;7�H;��H;#�H;��H;      ��H;��H; �H;�H;�H;��H;��H;��H;��H;��H;��H;�H;$�H;�H;��H;��H;��H;��H;��H;�H;b�H;��H;P�H;��H;��H;�H;Y�H;L�H;b�H;��H;��H;��H;��H;��H;��H;��H;��H;��H;��H;��H;��H;��H;��H;��H;b�H;L�H;Y�H;�H;��H;��H;P�H;��H;b�H;�H;��H;��H;��H;��H;��H;�H;$�H;�H;��H;��H;��H;��H;��H;��H;�H;�H; �H;��H;      ��H;��H;#�H;��H;7�H;�H;��H;��H;��H;�H;(�H;B�H;i�H;��H;��H;��H;��H;G�H;
�H;��H;^�H;��H;(�H;��H;��H;�H;:�H;[�H;o�H;��H;��H;��H;��H;��H;��H;��H;��H;��H;��H;��H;��H;��H;��H;��H;o�H;[�H;:�H;�H;��H;��H;(�H;��H;^�H;��H;
�H;G�H;��H;��H;��H;��H;i�H;B�H;(�H;�H;��H;��H;��H;�H;7�H;��H;#�H;��H;      ~�H;��H;��H;��H;D�H;2�H;*�H;P�H;��H;��H;<�H;��H;��H;1�H;k�H;��H;��H;��H;W�H;�H;��H;p�H;��H;H�H;��H;��H;�H;E�H;e�H;h�H;��H;��H;��H;��H;��H;��H;��H;��H;��H;��H;��H;��H;��H;h�H;e�H;E�H;�H;��H;��H;H�H;��H;p�H;��H;�H;W�H;��H;��H;��H;k�H;1�H;��H;��H;<�H;��H;��H;P�H;*�H;2�H;D�H;��H;��H;��H;      ��H;��H;b�H;��H;��H;�H;e�H;��H;��H;+�H;��H;��H;'�H;��H;.�H;��H;��H;(�H;<�H;6�H;��H;��H;O�H;��H;=�H;~�H;��H;�H;5�H;]�H;o�H;��H;��H;��H;��H;��H;��H;��H;��H;��H;��H;��H;o�H;]�H;5�H;�H;��H;~�H;=�H;��H;O�H;��H;��H;6�H;<�H;(�H;��H;��H;.�H;��H;'�H;��H;��H;+�H;��H;��H;e�H;�H;��H;��H;b�H;��H;      E�H;��H;�H;��H;3�H;��H;e�H;6�H;J�H;n�H;��H;��H;��H;�H;�H;��H;��H;��H;[�H;��H;��H;��H;c�H;�H;��H;,�H;}�H;��H;��H;6�H;a�H;k�H;{�H;��H;��H;��H;��H;��H;��H;��H;{�H;k�H;a�H;6�H;��H;��H;}�H;,�H;��H;�H;c�H;��H;��H;��H;[�H;��H;��H;��H;�H;�H;��H;��H;��H;n�H;J�H;6�H;e�H;��H;3�H;��H;�H;��H;      ��H;��H;��H;��H;��H;��H;�H;��H;q�H;_�H;M�H;5�H;�H;��H;t�H;��H;/�H;J�H;
�H;��H;��H;G�H;h�H;�H;��H;��H; �H;i�H;��H;��H;)�H;A�H;k�H;��H;��H;��H;��H;��H;��H;��H;k�H;A�H;)�H;��H;��H;i�H; �H;��H;��H;�H;h�H;G�H;��H;��H;
�H;J�H;/�H;��H;t�H;��H;�H;5�H;M�H;_�H;q�H;��H;�H;��H;��H;��H;��H;��H;      s�H;ѣH;ϤH;t�H;��H;��H;ĮH;g�H;9�H;9�H;N�H;J�H;#�H;��H;R�H;��H;��H;I�H;��H;��H;��H;H�H;��H;�H;��H;��H;j�H;�H;Y�H;��H;��H;)�H;a�H;o�H;��H;��H;��H;��H;��H;o�H;a�H;)�H;��H;��H;Y�H;�H;j�H;��H;��H;�H;��H;H�H;��H;��H;��H;I�H;��H;��H;R�H;��H;#�H;J�H;N�H;9�H;9�H;g�H;ĮH;��H;��H;t�H;ϤH;ѣH;      X�H;ǋH;G�H;��H;�H;��H;L�H;F�H;��H;
�H;��H;�H;a�H;k�H;5�H;z�H;~�H;(�H;l�H;E�H;��H;��H;��H;A�H;��H;��H;��H;S�H;��H;J�H;��H;��H;6�H;]�H;h�H;��H;��H;��H;h�H;]�H;6�H;��H;��H;J�H;��H;S�H;��H;��H;��H;A�H;��H;��H;��H;E�H;l�H;(�H;~�H;z�H;5�H;k�H;a�H;�H;��H;
�H;��H;F�H;L�H;��H;�H;��H;G�H;ǋH;      tiH;!jH;^lH;�oH;tH;0zH;��H;��H;�H;��H;5�H;��H;�H;ϳH;R�H;B�H;��H;s�H;��H;��H;��H;��H;)�H;,�H;��H;t�H;��H;e�H;[�H;��H;Y�H;��H;��H;5�H;e�H;o�H;b�H;o�H;e�H;5�H;��H;��H;Y�H;��H;[�H;e�H;��H;t�H;��H;,�H;)�H;��H;��H;��H;��H;s�H;��H;B�H;R�H;ϳH;�H;��H;5�H;��H;�H;��H;��H;0zH;tH;�oH;^lH;!jH;      4/H;�0H;Q5H;J<H;5EH;hOH;ZH;eH;�oH;�zH;��H;�H;�H;h�H;�H;�H;k�H;��H;��H;��H;��H;��H;�H;��H;��H;��H;J�H;��H;e�H;S�H;�H;i�H;��H;�H;E�H;[�H;L�H;[�H;E�H;�H;��H;i�H;�H;S�H;e�H;��H;J�H;��H;��H;��H;�H;��H;��H;��H;��H;��H;k�H;�H;�H;h�H;�H;�H;��H;�zH;�oH;eH;ZH;hOH;5EH;J<H;Q5H;�0H;      �G;�G;��G;��G;/�G;,�G;�H;)H;)?H;�RH;�cH;�rH;��H;��H;��H;[�H;
�H;��H;{�H;!�H;��H;��H;��H;W�H;O�H;��H;��H;J�H;��H;��H;j�H; �H;}�H;��H;�H;:�H;Y�H;:�H;�H;��H;}�H; �H;j�H;��H;��H;J�H;��H;��H;O�H;W�H;��H;��H;��H;!�H;{�H;��H;
�H;[�H;��H;��H;��H;�rH;�cH;�RH;)?H;)H;�H;,�G;/�G;��G;��G;�G;      ?ZF;�cF;5�F;��F;�F;�!G;EaG;�G;��G;iH; )H;�FH;�]H;�pH;5�H;�H; �H;��H;��H;��H;	�H;e�H;��H;E�H;�H;5�H;��H;��H;t�H;��H;��H;��H;,�H;~�H;��H;�H;�H;�H;��H;~�H;,�H;��H;��H;��H;t�H;��H;��H;5�H;�H;E�H;��H;e�H;	�H;��H;��H;��H; �H;�H;5�H;�pH;�]H;�FH; )H;iH;��G;�G;EaG;�!G;�F;��F;5�F;�cF;      �VC; nC; �C;�D;|�D;V4E;)�E;�ZF;��F;�KG;,�G;��G;c H;^EH;D`H;=uH;#�H;��H;��H;b�H;<�H;��H;�H;H�H;�H;�H;O�H;��H;��H;��H;��H;��H;��H;=�H;��H;��H;��H;��H;��H;=�H;��H;��H;��H;��H;��H;��H;O�H;�H;�H;H�H;�H;��H;<�H;b�H;��H;��H;#�H;=uH;D`H;^EH;c H;��G;,�G;�KG;��F;�ZF;)�E;V4E;|�D;�D; �C; nC;      ��<;M�<;P\=;�N>;�?;��@;�6B;u�C;,�D;̱E;��F;�!G;�G;1�G;
)H;iOH;FjH;gH;W�H;X�H;�H;߷H;��H;H�H;H�H;E�H;W�H;��H;,�H;A�H;�H;�H;�H;��H;H�H;��H;��H;��H;H�H;��H;�H;�H;�H;A�H;,�H;��H;W�H;E�H;H�H;H�H;��H;߷H;�H;X�H;W�H;gH;FjH;iOH;
)H;1�G;�G;�!G;��F;̱E;,�D;u�C;�6B;��@;�?;�N>;P\=;M�<;      Y.;�.;�0;2;��4;�7;�{:;u\=;��?;�6B;�D;qnE;fwF;e4G;ߵG;
H;?H;aH;�yH;��H;.�H;ܫH;`�H;��H;�H;��H;��H;�H;)�H;��H;��H;h�H;c�H;O�H;��H;(�H;P�H;(�H;��H;O�H;c�H;h�H;��H;��H;)�H;�H;��H;��H;�H;��H;`�H;ܫH;.�H;��H;�yH;aH;?H;
H;ߵG;e4G;fwF;qnE;�D;�6B;��?;u\=;�{:;�7;��4;2;�0;�.;      ^;��;Ml;VZ;�_;%;+;8�0;G6;��:;��>;��A;�D;�E;`�F;PzG;t�G;1H;ZH;�uH;��H;g�H;ܫH;߷H;��H;e�H;��H;��H;��H;��H;H�H;G�H;��H;��H;p�H;��H;��H;��H;p�H;��H;��H;G�H;H�H;��H;��H;��H;��H;e�H;��H;߷H;ܫH;g�H;��H;�uH;ZH;1H;t�G;PzG;`�F;�E;�D;��A;��>;��:;G6;8�0;+;%;�_;VZ;Ml;��;      ��:A,�:"f�:���:~~�:^;��;��;��#;y�,;��4;Q�:;�W?;.�B;��D;�ZF;FG;�G;}'H;~VH;�tH;��H;.�H;�H;<�H;	�H;��H;��H;��H;��H;��H;��H;��H;��H;��H;^�H;b�H;^�H;��H;��H;��H;��H;��H;��H;��H;��H;��H;	�H;<�H;�H;.�H;��H;�tH;~VH;}'H;�G;FG;�ZF;��D;.�B;�W?;Q�:;��4;y�,;��#;��;��;^;~~�:���:"f�:A,�:       �e9��9��9�:��Y:�x�:u:�:��:/^;7�;�";r-;(G6;��<;2>A;0D;�F;e"G;�G;$H;~VH;�uH;��H;X�H;b�H;��H;!�H;��H;��H;E�H;��H;��H;��H;6�H;�H;��H;�H;��H;�H;6�H;��H;��H;��H;E�H;��H;��H;!�H;��H;b�H;X�H;��H;�uH;~VH;$H;�G;e"G;�F;0D;2>A;��<;(G6;r-;�";7�;/^;��:u:�:�x�:��Y:�:��9��9      �����뺸кh����Y����k89v5:N.�:�c�:�A;�l;@?&;~2;�{:;` @;��C;�E;�G;�G;}'H;ZH;�yH;W�H;��H;��H;{�H;��H;��H;l�H;��H;
�H;[�H;<�H;W�H;
�H;��H;
�H;W�H;<�H;[�H;
�H;��H;l�H;��H;��H;{�H;��H;��H;W�H;�yH;ZH;}'H;�G;�G;�E;��C;` @;�{:;~2;@?&;�l;�A;�c�:N.�:v5:�k89���Y�h����к���      暩�\���4J��Y��T�b�)�-�3��ZJx�1��":��:?��:8�;� ;��.;/�8;��?;1�C;�E;e"G;�G;1H;aH;gH;��H;��H;��H;��H;s�H;(�H;I�H;J�H;��H;(�H;��H;G�H;��H;G�H;��H;(�H;��H;J�H;I�H;(�H;s�H;��H;��H;��H;��H;gH;aH;1H;�G;e"G;�E;1�C;��?;/�8;��.;� ;8�;?��:��:":1��ZJx�3��)�-�T�b�Y��4J��\���      �B(��%�����_�}����˻	��.�b�y&�c ��>@���Y:�:T^;B�;��,;Z_8;��?;��C;�F;FG;t�G;?H;FjH;#�H; �H;
�H;k�H;��H;~�H;��H;/�H;��H;��H;��H;��H;��H;��H;��H;��H;��H;/�H;��H;~�H;��H;k�H;
�H; �H;#�H;FjH;?H;t�G;FG;�F;��C;��?;Z_8;��,;B�;T^;�:��Y:>@�c ��y&�.�b�	���˻}����_�����%�      �����x���#��(F{���]��E<����J�뻲���bd\���]�,2:��:���:�Z;��,;/�8;` @;0D;�ZF;PzG;
H;iOH;=uH;�H;[�H;�H;B�H;z�H;��H;��H;��H;��H;��H;��H;��H;��H;��H;��H;��H;��H;��H;z�H;B�H;�H;[�H;�H;=uH;iOH;
H;PzG;�ZF;0D;` @;/�8;��,;�Z;���:��:,2:]���bd\�����J�뻛���E<���]�(F{��#���x��      >�Ｘ���o�Wrμ����bv��="���]N�����?ݻf^��z��0�Y�_�9��:���:B�;��.;�{:;2>A;��D;`�F;ߵG;
)H;D`H;5�H;��H;�H;R�H;5�H;R�H;t�H;�H;.�H;k�H;��H;��H;��H;k�H;.�H;�H;t�H;R�H;5�H;R�H;�H;��H;5�H;D`H;
)H;ߵG;`�F;��D;2>A;�{:;��.;B�;���:��:_�90�Y�z��f^���?ݻ����]N�="��bv������Wrμ�o༸��      Gn;�`\8��s/�(�!�h��>���Prμ��������E<�������N3��Ix�_�9��:T^;� ;~2;��<;.�B;�E;e4G;1�G;^EH;�pH;��H;h�H;ϳH;k�H;��H;��H;�H;��H;1�H;��H;�H;��H;1�H;��H;�H;��H;��H;k�H;ϳH;h�H;��H;�pH;^EH;1�G;e4G;�E;.�B;��<;~2;� ;T^;��:_�9�Ix��N3�������E<��������Prμ>���h��(�!��s/�`\8�      ���������Ȅ�KSt���Y�Dn;�O�P#���Oļ�����&R��_������N3�0�Y�,2:�:8�;@?&;(G6;�W?;�D;fwF;�G;c H;�]H;��H;�H;�H;a�H;#�H;�H;��H;'�H;��H;i�H;$�H;i�H;��H;'�H;��H;�H;#�H;a�H;�H;�H;��H;�]H;c H;�G;fwF;�D;�W?;(G6;@?&;8�;�:,2:0�Y��N3������_��&R������OļP#��O�Dn;���Y�KSt��Ȅ�����      ��ѽ�[νa�ý�㳽&����L��r�d�Z\8�c���ټWv����Y��_����z��]���Y:?��:�l;r-;Q�:;��A;qnE;�!G;��G;�FH;�rH;�H;��H;�H;J�H;5�H;��H;��H;��H;B�H;�H;B�H;��H;��H;��H;5�H;J�H;�H;��H;�H;�rH;�FH;��G;�!G;qnE;��A;Q�:;r-;�l;?��:��Y:]�z������_���Y�Wv���ټc��Z\8�r�d��L��&����㳽a�ý�[ν      ��]�È�a}�q�_�ý�u�������K����o�Wv���&R���f^����>@���:�A;�";��4;��>;�D;��F;,�G; )H;�cH;��H;5�H;��H;N�H;M�H;��H;��H;<�H;(�H;��H;(�H;<�H;��H;��H;M�H;N�H;��H;5�H;��H;�cH; )H;,�G;��F;�D;��>;��4;�";�A;��:>@���f^�����&R�Wv���o����K������u��_�ýq�a}�È�]�      j+X��T��nH�ؕ6�� �Y��(��㳽����mR����ټ�����E<��?ݻbd\�c ��":�c�:7�;y�,;��:;�6B;̱E;�KG;iH;�RH;�zH;��H;
�H;9�H;_�H;n�H;+�H;��H;�H;��H;�H;��H;+�H;n�H;_�H;9�H;
�H;��H;�zH;�RH;iH;�KG;̱E;�6B;��:;y�,;7�;�c�:":c ��bd\��?ݻ�E<������ټ���mR�����㳽(�Y��� �ؕ6��nH��T�      Ѱ������n���*|�4S\�� :����Z�U$������K�c���Oļ����������y&�1��N.�:/^;��#;G6;��?;,�D;��F;��G;)?H;�oH;�H;��H;9�H;q�H;J�H;��H;��H;��H;��H;��H;��H;��H;J�H;q�H;9�H;��H;�H;�oH;)?H;��G;��F;,�D;��?;G6;��#;/^;N.�:1��y&������������Oļc���K����U$���Z���� :�4S\��*|�n������      -�; 9ɾi㼾�A�������Mw��nH�����Z��㳽����Z\8�P#�������]N�J��.�b�ZJx�v5:��:��;8�0;u\=;u�C;�ZF;�G;)H;eH;��H;F�H;g�H;��H;6�H;��H;P�H;��H;��H;��H;P�H;��H;6�H;��H;g�H;F�H;��H;eH;)H;�G;�ZF;u�C;u\=;8�0;��;��:v5:ZJx�.�b�J���]N�����P#��Z\8������㳽�Z񽞯��nH��Mw������A��i㼾 9ɾ      #y��v�R���-�߾����0��1����nH���(Ὁu��r�d�O�Prμ="�����	��3���k89u:�:��;+;�{:;�6B;)�E;EaG;�H;ZH;��H;L�H;ĮH;�H;e�H;e�H;*�H;��H;��H;��H;*�H;e�H;e�H;�H;ĮH;L�H;��H;ZH;�H;EaG;)�E;�6B;�{:;+;��;u:�:�k893��	�����="��PrμO�r�d��u��(����nH�1���0������-�߾R����v�      �O/�aM+�I�����1W�� 9ɾ0���Mw�� :�Y��_�ý�L��Dn;�>���bv���E<��˻)�-����x�:^;%;�7;��@;V4E;�!G;,�G;hOH;0zH;��H;��H;��H;��H;�H;2�H;�H;��H;�H;2�H;�H;��H;��H;��H;��H;0zH;hOH;,�G;�!G;V4E;��@;�7;%;^;�x�:��)�-��˻�E<�bv��>���Dn;��L��_�ýY��� :��Mw�0�� 9ɾ1W�����I��aM+�      $�X�EvS�%E��O/��S�1W����������4S\�� �q�&�����Y�h��������]�}���T�b��Y���Y:~~�:�_;��4;�?;|�D;�F;/�G;5EH;tH;�H;��H;��H;3�H;��H;D�H;7�H;�H;7�H;D�H;��H;3�H;��H;��H;�H;tH;5EH;/�G;�F;|�D;�?;��4;�_;~~�:��Y:�Y�T�b�}�����]�����h����Y�&���q�� �4S\���������1W���S��O/�%E�EvS�      � ����y�M�h�ބN��O/����-�߾�A���*|�ؕ6�a}��㳽KSt�(�!�Wrμ(F{��_�Y��h����:���:VZ;2;�N>;�D;��F;��G;J<H;�oH;��H;t�H;��H;��H;��H;��H;��H;�H;��H;��H;��H;��H;��H;t�H;��H;�oH;J<H;��G;��F;�D;�N>;2;VZ;���:�:h���Y���_�(F{�Wrμ(�!�KSt��㳽a}�ؕ6��*|��A��-�߾����O/�ބN�M�h���y�      1v��V���L ��M�h�%E�I��R���i㼾n���nH�È�a�ý�Ȅ��s/��o༼#�����4J���к��9"f�:Ml;�0;P\=; �C;5�F;��G;Q5H;^lH;G�H;ϤH;��H;�H;b�H;��H;#�H; �H;#�H;��H;b�H;�H;��H;ϤH;G�H;^lH;Q5H;��G;5�F; �C;P\=;�0;Ml;"f�:��9�к4J������#���o��s/��Ȅ�a�ýÈ��nH�n��i㼾R���I��%E�M�h�L ��V���      ph��"���V�����y�EvS�aM+��v� 9ɾ�����T�]��[ν����`\8�����x���%�\��������9A,�:��;�.;M�<; nC;�cF;�G;�0H;!jH;ǋH;ѣH;��H;��H;��H;��H;��H;��H;��H;��H;��H;��H;��H;ѣH;ǋH;!jH;�0H;�G;�cF; nC;M�<;�.;��;A,�:��9���\����%��x�����`\8������[ν]��T����� 9ɾ�v�aM+�EvS���y�V���"���      .Eb�I]�tN�ߛ7����e� �{�˾��	�j��!,�J���0��m���,˼��x�E���1��b���P�:e�:2;��1;n+>;��C;�vF;�G;��G;>H;�gH;Z�H;v�H;8�H;�H;��H;(�H;��H;(�H;��H;�H;8�H;v�H;Z�H;�gH;>H;��G;�G;�vF;��C;n+>;��1;2;e�:P�:b����1��E����x�,˼��m�0��J����!,�	�j���{�˾e� ����ߛ7�tN�I]�      I]�N�W��TI�v3��D�������Ǿb���ȟf� )� ��W;���Fi��k�x�Ǽ�[t�8�	�(Ȅ�tX��Ο:���:%�;�I2;�Y>;pD;�~F;[�G;+H;�>H;�hH;�H;�H;q�H;7�H;��H;S�H;��H;S�H;��H;7�H;q�H;�H;�H;�hH;�>H;+H;[�G;�~F;pD;�Y>;�I2;%�;���:Ο:tX��(Ȅ�8�	��[t�x�Ǽ�k��Fi�W;�� �� )�ȟf�b�����Ǿ�����D�v3��TI�N�W�      tN��TI���;��'��k���i���f󐾖Z��K ��s�&����&^����"����g����Ѩu�S!���1<:��:m
;�f3;-�>;�AD;ՕF;�G;�H;UAH;~jH;\�H;ߟH;(�H;ԻH;k�H;��H;B�H;��H;k�H;ԻH;(�H;ߟH;\�H;~jH;UAH;�H;�G;ՕF;�AD;-�>;�f3;m
;��:�1<:S!��Ѩu������g��"�����&^�&����s潎K ��Z�f�i������k��'���;��TI�      ߛ7�v3��'����e� ��{Ծ
���6���]�F�����ӽ���;�L�1v�x뮼-T�ǘ��PV�r�=�1(i:_��:!z ;�#5;�?;2�D;�F;�G;�H;�EH;�mH;��H;}�H;j�H;ۼH;4�H;O�H;��H;O�H;4�H;ۼH;j�H;}�H;��H;�mH;�EH;�H;�G;�F;2�D;�?;�#5;!z ;_��:1(i:r�=��PV�ǘ�-T�x뮼1v�;�L�����ӽ���]�F�6���
����{Ծe� �����'�v3�      ����D��k�e� �<�ݾS���C͓�ȟf��>/�x��~'��n섽/�6�Rt��v��?�:�Tʻ�.�ݷ��s�:1; �$;�X7;��@;	E;:�F;P�G;�H;EKH;�qH;��H;ɣH;�H;�H;.�H;D�H;��H;D�H;.�H;�H;�H;ɣH;��H;�qH;EKH;�H;P�G;:�F;	E;��@;�X7; �$;1;�s�:ݷ��.�Tʻ?�:��v��Rt�/�6�n섽~'��x���>/�ȟf�C͓�S���<�ݾe� ��k��D�      e� ������쾻{ԾS���b���9�x�rSC��^�ͻ޽%���Q�e����ѼG������R������Ԥ8��:�X;��);5�9;-�A;��E;�G;2�G;s H;DRH;�vH;v�H;��H;:�H;��H;r�H;u�H;��H;u�H;r�H;��H;:�H;��H;v�H;�vH;DRH;s H;2�G;�G;��E;-�A;5�9;��);�X;��:�Ԥ8����R�����G���Ѽ��Q�e�%���ͻ޽�^�rSC�9�x�b���S����{Ծ�쾃���      {�˾��Ǿi���
���C͓�9�x�ؘJ��K �H��� �������?���t뮼�[�����3|��W��;�:u~�:';�
/;�f<;�C;� F;�MG;��G;9,H;sZH;�|H;ǖH;©H;��H;��H;��H;��H;��H;��H;��H;��H;��H;©H;ǖH;�|H;sZH;9,H;��G;�MG;� F;�C;�f<;�
/;';u~�:;�:�W��3|������[�t뮼����?���� ��H����K �ؘJ�9�x�C͓�
���i�����Ǿ      ��b���f�6���ȟf�rSC��K �Gn����Ž����Z��k��|ռX��Ey-����x.�z���O�:�*�:��;o4;s�>;)D;�vF;I�G;��G;�8H;\cH;w�H;��H;[�H;e�H;��H;��H;K�H;f�H;K�H;��H;��H;e�H;[�H;��H;w�H;\cH;�8H;��G;I�G;�vF;)D;s�>;o4;��;�*�:�O�:z��x.����Ey-�X���|ռ�k��Z������ŽGn���K �rSC�ȟf�6���f�b���      	�j�ȟf��Z�]�F��>/��^�H�����Ž- ���Fi�kQ+�Ot�PT��H�W�����1��jȺ�U�9�O�:	Y;��(;T�8;1A;�E;!�F;|�G;�H;�EH;�lH;��H;��H;8�H;d�H;��H;��H;��H;��H;��H;��H;��H;d�H;8�H;��H;��H;�lH;�EH;�H;|�G;!�F;�E;1A;T�8;��(;	Y;�O�:�U�9jȺ�1�����H�W�PT��Ot�kQ+��Fi�- ����ŽH����^��>/�]�F��Z�ȟf�      �!,� )��K ����x��ͻ޽ ������Fi���0�����跼z�x�����.��c�(�����)i:���:��;�0;��<;�C;��E;)<G;
�G;�#H;jSH;�vH;�H;�H;E�H;t�H;4�H;��H;��H;n�H;��H;��H;4�H;t�H;E�H;�H;�H;�vH;jSH;�#H;
�G;)<G;��E;�C;��<;�0;��;���:�)i:���c�(��.�����z�x��跼�����0��Fi���� ��ͻ޽x������K � )�      J��� ��s��ӽ~'��%�������Z�kQ+�����"��G����0���׻͕b��W���V�9�:�_;�)';/Y7;G#@;S�D;�F;+�G;��G;@7H;aH;��H;Y�H;��H;l�H;��H;��H;z�H;A�H;.�H;A�H;z�H;��H;��H;l�H;��H;Y�H;��H;aH;@7H;��G;+�G;�F;S�D;G#@;/Y7;�)';�_;�:�V�9�W��͕b���׻��0�G���"�����kQ+��Z����%���~'���ӽ�s� ��      0��W;��&������n섽Q�e���?��k�Ot��跼G��ee7�����Ǆ��0�K�t�^t�:�*�:�
;�1;��<;��B;N�E;G;�G;iH;vIH;`nH;��H;��H;�H;��H;��H;�H;��H; �H;��H; �H;��H;�H;��H;��H;�H;��H;��H;`nH;vIH;iH;�G;G;N�E;��B;��<;�1;�
;�*�:^t�:K�t��0��Ǆ����ee7�G���跼Ot�k���?�Q�e�n섽���&���W;��      m��Fi��&^�;�L�/�6������|ռPT��z�x���0��������1���ڷ�wm`:��:��;��*;}�8;G�@;d�D;��F;}G;��G;�0H;�ZH;m{H;��H;֧H;�H;��H;��H;|�H;��H;��H;d�H;��H;��H;|�H;��H;��H;�H;֧H;��H;m{H;�ZH;�0H;��G;}G;��F;d�D;G�@;}�8;��*;��;��:wm`:�ڷ�1��������껣�0�z�x�PT���|ռ����/�6�;�L��&^��Fi�      ���k���1v�Rt��Ѽt뮼X��H�W������׻�Ǆ�1�����3<:v��::Y;�s%;<$5;�Y>;-`C;��E;N)G;u�G;"H;GH;lkH;�H;��H;��H;ȻH;��H;��H;��H;g�H;^�H;�H;^�H;g�H;��H;��H;��H;ȻH;��H;��H;�H;lkH;GH;"H;u�G;N)G;��E;-`C;�Y>;<$5;�s%;:Y;v��:�3<:���1���Ǆ���׻���H�W�X��t뮼�ѼRt�1v����k�      ,˼x�Ǽ�"��x뮼�v��G���[�Ey-�����.��͕b��0㺋ڷ��3<:L�:^\;��!;1J2;�f<;/B;QBE;J�F;a�G; �G;�3H;�[H;{H;��H;��H;P�H;��H;5�H;��H;B�H;A�H;��H;��H;��H;A�H;B�H;��H;5�H;��H;P�H;��H;��H;{H;�[H;�3H; �G;a�G;J�F;QBE;/B;�f<;1J2;��!;^\;L�:�3<:�ڷ��0�͕b��.�����Ey-��[�G���v��x뮼�"��x�Ǽ      ��x��[t���g�-T�?�:������������1��c�(��W��K�t�wm`:v��:^\;pz ;�0;�;;9<A;?�D;�vF;�bG;d�G;� H;�LH;�nH;o�H;~�H;��H;��H;Z�H;��H;H�H;_�H;��H;��H;�H;��H;��H;_�H;H�H;��H;Z�H;��H;��H;~�H;o�H;�nH;�LH;� H;d�G;�bG;�vF;?�D;9<A;�;;�0;pz ;^\;v��:wm`:K�t��W��c�(��1������������?�:�-T���g��[t�      E��8�	����ǘ�Tʻ�R��3|�x.�jȺ����V�9^t�:��::Y;��!;�0;-�:;�@;4BD;�1F;�7G;��G;�H;j?H;*cH;�H;m�H;:�H;<�H;>�H;��H;��H;��H;[�H;��H;��H;s�H;��H;��H;[�H;��H;��H;��H;>�H;<�H;:�H;m�H;�H;*cH;j?H;�H;��G;�7G;�1F;4BD;�@;-�:;�0;��!;:Y;��:^t�:�V�9���jȺx.�3|��R��Tʻǘ����8�	�      �1��(Ȅ�Ѩu��PV��.�����W��z��U�9�)i:�:�*�:��;�s%;1J2;�;;�@;�D;/F;>G;��G;�H;�4H;�YH;5wH;7�H;�H;	�H;�H;H�H;^�H;�H;�H;�H;*�H;E�H;��H;E�H;*�H;�H;�H;�H;^�H;H�H;�H;	�H;�H;7�H;5wH;�YH;�4H;�H;��G;>G;/F;�D;�@;�;;1J2;�s%;��;�*�:�:�)i:�U�9z���W������.��PV�Ѩu�(Ȅ�      b���tX��S!��r�=�ݷ��Ԥ8;�:�O�:�O�:���:�_;�
;��*;<$5;�f<;9<A;4BD;/F;�G;��G;q�G;�,H;RH;UpH;�H;��H;r�H;�H;)�H;��H;��H;��H;?�H;��H;��H;{�H;��H;{�H;��H;��H;?�H;��H;��H;��H;)�H;�H;r�H;��H;�H;UpH;RH;�,H;q�G;��G;�G;/F;4BD;9<A;�f<;<$5;��*;�
;�_;���:�O�:�O�:;�:�Ԥ8ݷ�r�=�S!��tX��      P�:Ο:�1<:1(i:�s�:��:u~�:�*�:	Y;��;�)';�1;}�8;�Y>;/B;?�D;�1F;>G;��G;%�G;�(H;�MH;qkH;C�H;c�H;u�H;��H;�H;t�H;��H;$�H;�H;�H;D�H;��H;��H;��H;��H;��H;D�H;�H;�H;$�H;��H;t�H;�H;��H;u�H;c�H;C�H;qkH;�MH;�(H;%�G;��G;>G;�1F;?�D;/B;�Y>;}�8;�1;�)';��;	Y;�*�:u~�:��:�s�:1(i:�1<:Ο:      e�:���:��:_��:1;�X;';��;��(;�0;/Y7;��<;G�@;-`C;QBE;�vF;�7G;��G;q�G;�(H;�KH;�hH;.�H;O�H;��H;��H;��H;N�H;�H;��H;��H;A�H;��H;��H;��H;��H;��H;��H;��H;��H;��H;A�H;��H;��H;�H;N�H;��H;��H;��H;O�H;.�H;�hH;�KH;�(H;q�G;��G;�7G;�vF;QBE;-`C;G�@;��<;/Y7;�0;��(;��;';�X;1;_��:��:���:      2;%�;m
;!z ; �$;��);�
/;o4;T�8;��<;G#@;��B;d�D;��E;J�F;�bG;��G;�H;�,H;�MH;�hH;B�H;��H;��H;ͰH;��H;��H;��H;2�H;��H;^�H;�H;0�H;��H;��H;P�H;��H;P�H;��H;��H;0�H;�H;^�H;��H;2�H;��H;��H;��H;ͰH;��H;��H;B�H;�hH;�MH;�,H;�H;��G;�bG;J�F;��E;d�D;��B;G#@;��<;T�8;o4;�
/;��); �$;!z ;m
;%�;      ��1;�I2;�f3;�#5;�X7;5�9;�f<;s�>;1A;�C;S�D;N�E;��F;N)G;a�G;d�G;�H;�4H;RH;qkH;.�H;��H;�H;ɯH;�H;U�H;L�H; �H;��H;��H;u�H;��H;o�H;��H;��H;�H;\�H;�H;��H;��H;o�H;��H;u�H;��H;��H; �H;L�H;U�H;�H;ɯH;�H;��H;.�H;qkH;RH;�4H;�H;d�G;a�G;N)G;��F;N�E;S�D;�C;1A;s�>;�f<;5�9;�X7;�#5;�f3;�I2;      n+>;�Y>;-�>;�?;��@;-�A;�C;)D;�E;��E;�F;G;}G;u�G; �G;� H;j?H;�YH;UpH;C�H;O�H;��H;ɯH;�H;��H;��H;5�H;��H;��H;��H;O�H; �H;��H;��H;H�H;��H;��H;��H;H�H;��H;��H; �H;O�H;��H;��H;��H;5�H;��H;��H;�H;ɯH;��H;O�H;C�H;UpH;�YH;j?H;� H; �G;u�G;}G;G;�F;��E;�E;)D;�C;-�A;��@;�?;-�>;�Y>;      ��C;pD;�AD;2�D;	E;��E;� F;�vF;!�F;)<G;+�G;�G;��G;"H;�3H;�LH;*cH;5wH;�H;c�H;��H;ͰH;�H;��H;<�H;��H;��H;^�H;c�H;��H;��H;f�H;��H;?�H;��H;C�H;L�H;C�H;��H;?�H;��H;f�H;��H;��H;c�H;^�H;��H;��H;<�H;��H;�H;ͰH;��H;c�H;�H;5wH;*cH;�LH;�3H;"H;��G;�G;+�G;)<G;!�F;�vF;� F;��E;	E;2�D;�AD;pD;      �vF;�~F;ՕF;�F;:�F;�G;�MG;I�G;|�G;
�G;��G;iH;�0H;GH;�[H;�nH;�H;7�H;��H;u�H;��H;��H;U�H;��H;��H;W�H;$�H;�H;��H;��H;�H;S�H;6�H;��H;m�H;��H;��H;��H;m�H;��H;6�H;S�H;�H;��H;��H;�H;$�H;W�H;��H;��H;U�H;��H;��H;u�H;��H;7�H;�H;�nH;�[H;GH;�0H;iH;��G;
�G;|�G;I�G;�MG;�G;:�F;�F;ՕF;�~F;      �G;[�G;�G;�G;P�G;2�G;��G;��G;�H;�#H;@7H;vIH;�ZH;lkH;{H;o�H;m�H;�H;r�H;��H;��H;��H;L�H;5�H;��H;$�H;�H;h�H;J�H;��H;7�H;�H;��H;��H;��H;�H;�H;�H;��H;��H;��H;�H;7�H;��H;J�H;h�H;�H;$�H;��H;5�H;L�H;��H;��H;��H;r�H;�H;m�H;o�H;{H;lkH;�ZH;vIH;@7H;�#H;�H;��G;��G;2�G;P�G;�G;�G;[�G;      ��G;+H;�H;�H;�H;s H;9,H;�8H;�EH;jSH;aH;`nH;m{H;�H;��H;~�H;:�H;	�H;�H;�H;N�H;��H; �H;��H;^�H;�H;h�H;\�H;��H;�H;�H;��H;z�H;��H;�H;^�H;g�H;^�H;�H;��H;z�H;��H;�H;�H;��H;\�H;h�H;�H;^�H;��H; �H;��H;N�H;�H;�H;	�H;:�H;~�H;��H;�H;m{H;`nH;aH;jSH;�EH;�8H;9,H;s H;�H;�H;�H;+H;      >H;�>H;UAH;�EH;EKH;DRH;sZH;\cH;�lH;�vH;��H;��H;��H;��H;��H;��H;<�H;�H;)�H;t�H;�H;2�H;��H;��H;c�H;��H;J�H;��H;#�H;��H;��H;k�H;��H;5�H;p�H;��H;��H;��H;p�H;5�H;��H;k�H;��H;��H;#�H;��H;J�H;��H;c�H;��H;��H;2�H;�H;t�H;)�H;�H;<�H;��H;��H;��H;��H;��H;��H;�vH;�lH;\cH;sZH;DRH;EKH;�EH;UAH;�>H;      �gH;�hH;~jH;�mH;�qH;�vH;�|H;w�H;��H;�H;Y�H;��H;֧H;��H;P�H;��H;>�H;H�H;��H;��H;��H;��H;��H;��H;��H;��H;��H;�H;��H;��H;t�H;��H;$�H;y�H;��H;��H;��H;��H;��H;y�H;$�H;��H;t�H;��H;��H;�H;��H;��H;��H;��H;��H;��H;��H;��H;��H;H�H;>�H;��H;P�H;��H;֧H;��H;Y�H;�H;��H;w�H;�|H;�vH;�qH;�mH;~jH;�hH;      Z�H;�H;\�H;��H;��H;v�H;ǖH;��H;��H;�H;��H;�H;�H;ȻH;��H;Z�H;��H;^�H;��H;$�H;��H;^�H;u�H;O�H;��H;�H;7�H;�H;��H;t�H;��H;.�H;��H;��H;��H;��H;��H;��H;��H;��H;��H;.�H;��H;t�H;��H;�H;7�H;�H;��H;O�H;u�H;^�H;��H;$�H;��H;^�H;��H;Z�H;��H;ȻH;�H;�H;��H;�H;��H;��H;ǖH;v�H;��H;��H;\�H;�H;      v�H;�H;ߟH;}�H;ɣH;��H;©H;[�H;8�H;E�H;l�H;��H;��H;��H;5�H;��H;��H;�H;��H;�H;A�H;�H;��H; �H;f�H;S�H;�H;��H;k�H;��H;.�H;z�H;��H;��H;��H;�H;�H;�H;��H;��H;��H;z�H;.�H;��H;k�H;��H;�H;S�H;f�H; �H;��H;�H;A�H;�H;��H;�H;��H;��H;5�H;��H;��H;��H;l�H;E�H;8�H;[�H;©H;��H;ɣH;}�H;ߟH;�H;      8�H;q�H;(�H;j�H;�H;:�H;��H;e�H;d�H;t�H;��H;��H;��H;��H;��H;H�H;��H;�H;?�H;�H;��H;0�H;o�H;��H;��H;6�H;��H;z�H;��H;$�H;��H;��H;��H;��H;�H;�H;�H;�H;�H;��H;��H;��H;��H;$�H;��H;z�H;��H;6�H;��H;��H;o�H;0�H;��H;�H;?�H;�H;��H;H�H;��H;��H;��H;��H;��H;t�H;d�H;e�H;��H;:�H;�H;j�H;(�H;q�H;      �H;7�H;ԻH;ۼH;�H;��H;��H;��H;��H;4�H;��H;�H;|�H;��H;B�H;_�H;[�H;�H;��H;D�H;��H;��H;��H;��H;?�H;��H;��H;��H;5�H;y�H;��H;��H;��H; �H;-�H;8�H;�H;8�H;-�H; �H;��H;��H;��H;y�H;5�H;��H;��H;��H;?�H;��H;��H;��H;��H;D�H;��H;�H;[�H;_�H;B�H;��H;|�H;�H;��H;4�H;��H;��H;��H;��H;�H;ۼH;ԻH;7�H;      ��H;��H;k�H;4�H;.�H;r�H;��H;��H;��H;��H;z�H;��H;��H;g�H;A�H;��H;��H;*�H;��H;��H;��H;��H;��H;H�H;��H;m�H;��H;�H;p�H;��H;��H;��H;�H;-�H;�H;-�H;J�H;-�H;�H;-�H;�H;��H;��H;��H;p�H;�H;��H;m�H;��H;H�H;��H;��H;��H;��H;��H;*�H;��H;��H;A�H;g�H;��H;��H;z�H;��H;��H;��H;��H;r�H;.�H;4�H;k�H;��H;      (�H;S�H;��H;O�H;D�H;u�H;��H;K�H;��H;��H;A�H; �H;��H;^�H;��H;��H;��H;E�H;{�H;��H;��H;P�H;�H;��H;C�H;��H;�H;^�H;��H;��H;��H;�H;�H;8�H;-�H;$�H;6�H;$�H;-�H;8�H;�H;�H;��H;��H;��H;^�H;�H;��H;C�H;��H;�H;P�H;��H;��H;{�H;E�H;��H;��H;��H;^�H;��H; �H;A�H;��H;��H;K�H;��H;u�H;D�H;O�H;��H;S�H;      ��H;��H;B�H;��H;��H;��H;��H;f�H;��H;n�H;.�H;��H;d�H;�H;��H;�H;s�H;��H;��H;��H;��H;��H;\�H;��H;L�H;��H;�H;g�H;��H;��H;��H;�H;�H;�H;J�H;6�H;#�H;6�H;J�H;�H;�H;�H;��H;��H;��H;g�H;�H;��H;L�H;��H;\�H;��H;��H;��H;��H;��H;s�H;�H;��H;�H;d�H;��H;.�H;n�H;��H;f�H;��H;��H;��H;��H;B�H;��H;      (�H;S�H;��H;O�H;D�H;u�H;��H;K�H;��H;��H;A�H; �H;��H;^�H;��H;��H;��H;E�H;{�H;��H;��H;P�H;�H;��H;C�H;��H;�H;^�H;��H;��H;��H;�H;�H;8�H;-�H;$�H;6�H;$�H;-�H;8�H;�H;�H;��H;��H;��H;^�H;�H;��H;C�H;��H;�H;P�H;��H;��H;{�H;E�H;��H;��H;��H;^�H;��H; �H;A�H;��H;��H;K�H;��H;u�H;D�H;O�H;��H;S�H;      ��H;��H;k�H;4�H;.�H;r�H;��H;��H;��H;��H;z�H;��H;��H;g�H;A�H;��H;��H;*�H;��H;��H;��H;��H;��H;H�H;��H;m�H;��H;�H;p�H;��H;��H;��H;�H;-�H;�H;-�H;J�H;-�H;�H;-�H;�H;��H;��H;��H;p�H;�H;��H;m�H;��H;H�H;��H;��H;��H;��H;��H;*�H;��H;��H;A�H;g�H;��H;��H;z�H;��H;��H;��H;��H;r�H;.�H;4�H;k�H;��H;      �H;7�H;ԻH;ۼH;�H;��H;��H;��H;��H;4�H;��H;�H;|�H;��H;B�H;_�H;[�H;�H;��H;D�H;��H;��H;��H;��H;?�H;��H;��H;��H;5�H;y�H;��H;��H;��H; �H;-�H;8�H;�H;8�H;-�H; �H;��H;��H;��H;y�H;5�H;��H;��H;��H;?�H;��H;��H;��H;��H;D�H;��H;�H;[�H;_�H;B�H;��H;|�H;�H;��H;4�H;��H;��H;��H;��H;�H;ۼH;ԻH;7�H;      8�H;q�H;(�H;j�H;�H;:�H;��H;e�H;d�H;t�H;��H;��H;��H;��H;��H;H�H;��H;�H;?�H;�H;��H;0�H;o�H;��H;��H;6�H;��H;z�H;��H;$�H;��H;��H;��H;��H;�H;�H;�H;�H;�H;��H;��H;��H;��H;$�H;��H;z�H;��H;6�H;��H;��H;o�H;0�H;��H;�H;?�H;�H;��H;H�H;��H;��H;��H;��H;��H;t�H;d�H;e�H;��H;:�H;�H;j�H;(�H;q�H;      v�H;�H;ߟH;}�H;ɣH;��H;©H;[�H;8�H;E�H;l�H;��H;��H;��H;5�H;��H;��H;�H;��H;�H;A�H;�H;��H; �H;f�H;S�H;�H;��H;k�H;��H;.�H;z�H;��H;��H;��H;�H;�H;�H;��H;��H;��H;z�H;.�H;��H;k�H;��H;�H;S�H;f�H; �H;��H;�H;A�H;�H;��H;�H;��H;��H;5�H;��H;��H;��H;l�H;E�H;8�H;[�H;©H;��H;ɣH;}�H;ߟH;�H;      Z�H;�H;\�H;��H;��H;v�H;ǖH;��H;��H;�H;��H;�H;�H;ȻH;��H;Z�H;��H;^�H;��H;$�H;��H;^�H;u�H;O�H;��H;�H;7�H;�H;��H;t�H;��H;.�H;��H;��H;��H;��H;��H;��H;��H;��H;��H;.�H;��H;t�H;��H;�H;7�H;�H;��H;O�H;u�H;^�H;��H;$�H;��H;^�H;��H;Z�H;��H;ȻH;�H;�H;��H;�H;��H;��H;ǖH;v�H;��H;��H;\�H;�H;      �gH;�hH;~jH;�mH;�qH;�vH;�|H;w�H;��H;�H;Y�H;��H;֧H;��H;P�H;��H;>�H;H�H;��H;��H;��H;��H;��H;��H;��H;��H;��H;�H;��H;��H;t�H;��H;$�H;y�H;��H;��H;��H;��H;��H;y�H;$�H;��H;t�H;��H;��H;�H;��H;��H;��H;��H;��H;��H;��H;��H;��H;H�H;>�H;��H;P�H;��H;֧H;��H;Y�H;�H;��H;w�H;�|H;�vH;�qH;�mH;~jH;�hH;      >H;�>H;UAH;�EH;EKH;DRH;sZH;\cH;�lH;�vH;��H;��H;��H;��H;��H;��H;<�H;�H;)�H;t�H;�H;2�H;��H;��H;c�H;��H;J�H;��H;#�H;��H;��H;k�H;��H;5�H;p�H;��H;��H;��H;p�H;5�H;��H;k�H;��H;��H;#�H;��H;J�H;��H;c�H;��H;��H;2�H;�H;t�H;)�H;�H;<�H;��H;��H;��H;��H;��H;��H;�vH;�lH;\cH;sZH;DRH;EKH;�EH;UAH;�>H;      ��G;+H;�H;�H;�H;s H;9,H;�8H;�EH;jSH;aH;`nH;m{H;�H;��H;~�H;:�H;	�H;�H;�H;N�H;��H; �H;��H;^�H;�H;h�H;\�H;��H;�H;�H;��H;z�H;��H;�H;^�H;g�H;^�H;�H;��H;z�H;��H;�H;�H;��H;\�H;h�H;�H;^�H;��H; �H;��H;N�H;�H;�H;	�H;:�H;~�H;��H;�H;m{H;`nH;aH;jSH;�EH;�8H;9,H;s H;�H;�H;�H;+H;      �G;[�G;�G;�G;P�G;2�G;��G;��G;�H;�#H;@7H;vIH;�ZH;lkH;{H;o�H;m�H;�H;r�H;��H;��H;��H;L�H;5�H;��H;$�H;�H;h�H;J�H;��H;7�H;�H;��H;��H;��H;�H;�H;�H;��H;��H;��H;�H;7�H;��H;J�H;h�H;�H;$�H;��H;5�H;L�H;��H;��H;��H;r�H;�H;m�H;o�H;{H;lkH;�ZH;vIH;@7H;�#H;�H;��G;��G;2�G;P�G;�G;�G;[�G;      �vF;�~F;ՕF;�F;:�F;�G;�MG;I�G;|�G;
�G;��G;iH;�0H;GH;�[H;�nH;�H;7�H;��H;u�H;��H;��H;U�H;��H;��H;W�H;$�H;�H;��H;��H;�H;S�H;6�H;��H;m�H;��H;��H;��H;m�H;��H;6�H;S�H;�H;��H;��H;�H;$�H;W�H;��H;��H;U�H;��H;��H;u�H;��H;7�H;�H;�nH;�[H;GH;�0H;iH;��G;
�G;|�G;I�G;�MG;�G;:�F;�F;ՕF;�~F;      ��C;pD;�AD;2�D;	E;��E;� F;�vF;!�F;)<G;+�G;�G;��G;"H;�3H;�LH;*cH;5wH;�H;c�H;��H;ͰH;�H;��H;<�H;��H;��H;^�H;c�H;��H;��H;f�H;��H;?�H;��H;C�H;L�H;C�H;��H;?�H;��H;f�H;��H;��H;c�H;^�H;��H;��H;<�H;��H;�H;ͰH;��H;c�H;�H;5wH;*cH;�LH;�3H;"H;��G;�G;+�G;)<G;!�F;�vF;� F;��E;	E;2�D;�AD;pD;      n+>;�Y>;-�>;�?;��@;-�A;�C;)D;�E;��E;�F;G;}G;u�G; �G;� H;j?H;�YH;UpH;C�H;O�H;��H;ɯH;�H;��H;��H;5�H;��H;��H;��H;O�H; �H;��H;��H;H�H;��H;��H;��H;H�H;��H;��H; �H;O�H;��H;��H;��H;5�H;��H;��H;�H;ɯH;��H;O�H;C�H;UpH;�YH;j?H;� H; �G;u�G;}G;G;�F;��E;�E;)D;�C;-�A;��@;�?;-�>;�Y>;      ��1;�I2;�f3;�#5;�X7;5�9;�f<;s�>;1A;�C;S�D;N�E;��F;N)G;a�G;d�G;�H;�4H;RH;qkH;.�H;��H;�H;ɯH;�H;U�H;L�H; �H;��H;��H;u�H;��H;o�H;��H;��H;�H;\�H;�H;��H;��H;o�H;��H;u�H;��H;��H; �H;L�H;U�H;�H;ɯH;�H;��H;.�H;qkH;RH;�4H;�H;d�G;a�G;N)G;��F;N�E;S�D;�C;1A;s�>;�f<;5�9;�X7;�#5;�f3;�I2;      2;%�;m
;!z ; �$;��);�
/;o4;T�8;��<;G#@;��B;d�D;��E;J�F;�bG;��G;�H;�,H;�MH;�hH;B�H;��H;��H;ͰH;��H;��H;��H;2�H;��H;^�H;�H;0�H;��H;��H;P�H;��H;P�H;��H;��H;0�H;�H;^�H;��H;2�H;��H;��H;��H;ͰH;��H;��H;B�H;�hH;�MH;�,H;�H;��G;�bG;J�F;��E;d�D;��B;G#@;��<;T�8;o4;�
/;��); �$;!z ;m
;%�;      e�:���:��:_��:1;�X;';��;��(;�0;/Y7;��<;G�@;-`C;QBE;�vF;�7G;��G;q�G;�(H;�KH;�hH;.�H;O�H;��H;��H;��H;N�H;�H;��H;��H;A�H;��H;��H;��H;��H;��H;��H;��H;��H;��H;A�H;��H;��H;�H;N�H;��H;��H;��H;O�H;.�H;�hH;�KH;�(H;q�G;��G;�7G;�vF;QBE;-`C;G�@;��<;/Y7;�0;��(;��;';�X;1;_��:��:���:      P�:Ο:�1<:1(i:�s�:��:u~�:�*�:	Y;��;�)';�1;}�8;�Y>;/B;?�D;�1F;>G;��G;%�G;�(H;�MH;qkH;C�H;c�H;u�H;��H;�H;t�H;��H;$�H;�H;�H;D�H;��H;��H;��H;��H;��H;D�H;�H;�H;$�H;��H;t�H;�H;��H;u�H;c�H;C�H;qkH;�MH;�(H;%�G;��G;>G;�1F;?�D;/B;�Y>;}�8;�1;�)';��;	Y;�*�:u~�:��:�s�:1(i:�1<:Ο:      b���tX��S!��r�=�ݷ��Ԥ8;�:�O�:�O�:���:�_;�
;��*;<$5;�f<;9<A;4BD;/F;�G;��G;q�G;�,H;RH;UpH;�H;��H;r�H;�H;)�H;��H;��H;��H;?�H;��H;��H;{�H;��H;{�H;��H;��H;?�H;��H;��H;��H;)�H;�H;r�H;��H;�H;UpH;RH;�,H;q�G;��G;�G;/F;4BD;9<A;�f<;<$5;��*;�
;�_;���:�O�:�O�:;�:�Ԥ8ݷ�r�=�S!��tX��      �1��(Ȅ�Ѩu��PV��.�����W��z��U�9�)i:�:�*�:��;�s%;1J2;�;;�@;�D;/F;>G;��G;�H;�4H;�YH;5wH;7�H;�H;	�H;�H;H�H;^�H;�H;�H;�H;*�H;E�H;��H;E�H;*�H;�H;�H;�H;^�H;H�H;�H;	�H;�H;7�H;5wH;�YH;�4H;�H;��G;>G;/F;�D;�@;�;;1J2;�s%;��;�*�:�:�)i:�U�9z���W������.��PV�Ѩu�(Ȅ�      E��8�	����ǘ�Tʻ�R��3|�x.�jȺ����V�9^t�:��::Y;��!;�0;-�:;�@;4BD;�1F;�7G;��G;�H;j?H;*cH;�H;m�H;:�H;<�H;>�H;��H;��H;��H;[�H;��H;��H;s�H;��H;��H;[�H;��H;��H;��H;>�H;<�H;:�H;m�H;�H;*cH;j?H;�H;��G;�7G;�1F;4BD;�@;-�:;�0;��!;:Y;��:^t�:�V�9���jȺx.�3|��R��Tʻǘ����8�	�      ��x��[t���g�-T�?�:������������1��c�(��W��K�t�wm`:v��:^\;pz ;�0;�;;9<A;?�D;�vF;�bG;d�G;� H;�LH;�nH;o�H;~�H;��H;��H;Z�H;��H;H�H;_�H;��H;��H;�H;��H;��H;_�H;H�H;��H;Z�H;��H;��H;~�H;o�H;�nH;�LH;� H;d�G;�bG;�vF;?�D;9<A;�;;�0;pz ;^\;v��:wm`:K�t��W��c�(��1������������?�:�-T���g��[t�      ,˼x�Ǽ�"��x뮼�v��G���[�Ey-�����.��͕b��0㺋ڷ��3<:L�:^\;��!;1J2;�f<;/B;QBE;J�F;a�G; �G;�3H;�[H;{H;��H;��H;P�H;��H;5�H;��H;B�H;A�H;��H;��H;��H;A�H;B�H;��H;5�H;��H;P�H;��H;��H;{H;�[H;�3H; �G;a�G;J�F;QBE;/B;�f<;1J2;��!;^\;L�:�3<:�ڷ��0�͕b��.�����Ey-��[�G���v��x뮼�"��x�Ǽ      ���k���1v�Rt��Ѽt뮼X��H�W������׻�Ǆ�1�����3<:v��::Y;�s%;<$5;�Y>;-`C;��E;N)G;u�G;"H;GH;lkH;�H;��H;��H;ȻH;��H;��H;��H;g�H;^�H;�H;^�H;g�H;��H;��H;��H;ȻH;��H;��H;�H;lkH;GH;"H;u�G;N)G;��E;-`C;�Y>;<$5;�s%;:Y;v��:�3<:���1���Ǆ���׻���H�W�X��t뮼�ѼRt�1v����k�      m��Fi��&^�;�L�/�6������|ռPT��z�x���0��������1���ڷ�wm`:��:��;��*;}�8;G�@;d�D;��F;}G;��G;�0H;�ZH;m{H;��H;֧H;�H;��H;��H;|�H;��H;��H;d�H;��H;��H;|�H;��H;��H;�H;֧H;��H;m{H;�ZH;�0H;��G;}G;��F;d�D;G�@;}�8;��*;��;��:wm`:�ڷ�1��������껣�0�z�x�PT���|ռ����/�6�;�L��&^��Fi�      0��W;��&������n섽Q�e���?��k�Ot��跼G��ee7�����Ǆ��0�K�t�^t�:�*�:�
;�1;��<;��B;N�E;G;�G;iH;vIH;`nH;��H;��H;�H;��H;��H;�H;��H; �H;��H; �H;��H;�H;��H;��H;�H;��H;��H;`nH;vIH;iH;�G;G;N�E;��B;��<;�1;�
;�*�:^t�:K�t��0��Ǆ����ee7�G���跼Ot�k���?�Q�e�n섽���&���W;��      J��� ��s��ӽ~'��%�������Z�kQ+�����"��G����0���׻͕b��W���V�9�:�_;�)';/Y7;G#@;S�D;�F;+�G;��G;@7H;aH;��H;Y�H;��H;l�H;��H;��H;z�H;A�H;.�H;A�H;z�H;��H;��H;l�H;��H;Y�H;��H;aH;@7H;��G;+�G;�F;S�D;G#@;/Y7;�)';�_;�:�V�9�W��͕b���׻��0�G���"�����kQ+��Z����%���~'���ӽ�s� ��      �!,� )��K ����x��ͻ޽ ������Fi���0�����跼z�x�����.��c�(�����)i:���:��;�0;��<;�C;��E;)<G;
�G;�#H;jSH;�vH;�H;�H;E�H;t�H;4�H;��H;��H;n�H;��H;��H;4�H;t�H;E�H;�H;�H;�vH;jSH;�#H;
�G;)<G;��E;�C;��<;�0;��;���:�)i:���c�(��.�����z�x��跼�����0��Fi���� ��ͻ޽x������K � )�      	�j�ȟf��Z�]�F��>/��^�H�����Ž- ���Fi�kQ+�Ot�PT��H�W�����1��jȺ�U�9�O�:	Y;��(;T�8;1A;�E;!�F;|�G;�H;�EH;�lH;��H;��H;8�H;d�H;��H;��H;��H;��H;��H;��H;��H;d�H;8�H;��H;��H;�lH;�EH;�H;|�G;!�F;�E;1A;T�8;��(;	Y;�O�:�U�9jȺ�1�����H�W�PT��Ot�kQ+��Fi�- ����ŽH����^��>/�]�F��Z�ȟf�      ��b���f�6���ȟf�rSC��K �Gn����Ž����Z��k��|ռX��Ey-����x.�z���O�:�*�:��;o4;s�>;)D;�vF;I�G;��G;�8H;\cH;w�H;��H;[�H;e�H;��H;��H;K�H;f�H;K�H;��H;��H;e�H;[�H;��H;w�H;\cH;�8H;��G;I�G;�vF;)D;s�>;o4;��;�*�:�O�:z��x.����Ey-�X���|ռ�k��Z������ŽGn���K �rSC�ȟf�6���f�b���      {�˾��Ǿi���
���C͓�9�x�ؘJ��K �H��� �������?���t뮼�[�����3|��W��;�:u~�:';�
/;�f<;�C;� F;�MG;��G;9,H;sZH;�|H;ǖH;©H;��H;��H;��H;��H;��H;��H;��H;��H;��H;©H;ǖH;�|H;sZH;9,H;��G;�MG;� F;�C;�f<;�
/;';u~�:;�:�W��3|������[�t뮼����?���� ��H����K �ؘJ�9�x�C͓�
���i�����Ǿ      e� ������쾻{ԾS���b���9�x�rSC��^�ͻ޽%���Q�e����ѼG������R������Ԥ8��:�X;��);5�9;-�A;��E;�G;2�G;s H;DRH;�vH;v�H;��H;:�H;��H;r�H;u�H;��H;u�H;r�H;��H;:�H;��H;v�H;�vH;DRH;s H;2�G;�G;��E;-�A;5�9;��);�X;��:�Ԥ8����R�����G���Ѽ��Q�e�%���ͻ޽�^�rSC�9�x�b���S����{Ծ�쾃���      ����D��k�e� �<�ݾS���C͓�ȟf��>/�x��~'��n섽/�6�Rt��v��?�:�Tʻ�.�ݷ��s�:1; �$;�X7;��@;	E;:�F;P�G;�H;EKH;�qH;��H;ɣH;�H;�H;.�H;D�H;��H;D�H;.�H;�H;�H;ɣH;��H;�qH;EKH;�H;P�G;:�F;	E;��@;�X7; �$;1;�s�:ݷ��.�Tʻ?�:��v��Rt�/�6�n섽~'��x���>/�ȟf�C͓�S���<�ݾe� ��k��D�      ߛ7�v3��'����e� ��{Ծ
���6���]�F�����ӽ���;�L�1v�x뮼-T�ǘ��PV�r�=�1(i:_��:!z ;�#5;�?;2�D;�F;�G;�H;�EH;�mH;��H;}�H;j�H;ۼH;4�H;O�H;��H;O�H;4�H;ۼH;j�H;}�H;��H;�mH;�EH;�H;�G;�F;2�D;�?;�#5;!z ;_��:1(i:r�=��PV�ǘ�-T�x뮼1v�;�L�����ӽ���]�F�6���
����{Ծe� �����'�v3�      tN��TI���;��'��k���i���f󐾖Z��K ��s�&����&^����"����g����Ѩu�S!���1<:��:m
;�f3;-�>;�AD;ՕF;�G;�H;UAH;~jH;\�H;ߟH;(�H;ԻH;k�H;��H;B�H;��H;k�H;ԻH;(�H;ߟH;\�H;~jH;UAH;�H;�G;ՕF;�AD;-�>;�f3;m
;��:�1<:S!��Ѩu������g��"�����&^�&����s潎K ��Z�f�i������k��'���;��TI�      I]�N�W��TI�v3��D�������Ǿb���ȟf� )� ��W;���Fi��k�x�Ǽ�[t�8�	�(Ȅ�tX��Ο:���:%�;�I2;�Y>;pD;�~F;[�G;+H;�>H;�hH;�H;�H;q�H;7�H;��H;S�H;��H;S�H;��H;7�H;q�H;�H;�H;�hH;�>H;+H;[�G;�~F;pD;�Y>;�I2;%�;���:Ο:tX��(Ȅ�8�	��[t�x�Ǽ�k��Fi�W;�� �� )�ȟf�b�����Ǿ�����D�v3��TI�N�W�      �$��� ���������þ�*��
Dx�}�=����\Pν鰒��&K�xc����;�V�s���D^���S��v[:���:�d;��4;�_?;�lD;��F;puG;M�G;�H;�NH;�rH;�H;��H;��H;�H;q�H;E�H;q�H;�H;��H;��H;�H;�rH;�NH;�H;M�G;puG;��F;�lD;�_?;��4;�d;���:�v[:��S��D^�s��;�V����xc��&K�鰒�\Pν���}�=�
Dx��*���þ��������� �      �� �k��>��=���������0���s���:�N9���ʽZ����G��8��-��z5S�w���/X���D��Ad:�A�:� ;x�4;�?;"~D;p�F;3xG;��G;�H;NOH;HsH;:�H;�H;�H;W�H;��H;U�H;��H;W�H;�H;�H;:�H;HsH;NOH;�H;��G;3xG;p�F;"~D;�?;x�4;� ;�A�:�Ad:��D��/X�w��z5S��-���8���G�Z����ʽN9���:��s��0��������=��>��k��      ���>��&�
�����fYؾ���ȥ����f���0�C[�*8������ȟ>�|���#Ȥ�Y6H�,�ܻ�qF�1��3�}:���:�";��5;6�?;��D;��F;/�G;��G;s"H;�QH;�tH;y�H;�H;��H;�H;�H;��H;�H;�H;��H;�H;y�H;�tH;�QH;s"H;��G;/�G;��F;��D;6�?;��5;�";���:3�}:1���qF�,�ܻY6H�#Ȥ�|���ȟ>�����*8��C[���0���f�ȥ�����fYؾ����&�
�>��      ��=������I��þ�R��&���QS��Q"��s�����}��0���d���x�6��ƻ(}*����^�:�w;�%;Rl7;�@;�D;�F;��G;��G;3'H;UH;�wH;�H;f�H;±H;ۺH;�H;��H;�H;ۺH;±H;f�H;�H;�wH;UH;3'H;��G;��G;�F;�D;�@;Rl7;�%;�w;^�:���(}*��ƻx�6�d����켟0���}�����s��Q"�QS�&����R���þIᾁ���=��      ����fYؾ�þ�ê�f쏾jk���:�e�R�ؽ�����c�:y���Ҽݫ��� �B�(����'7��:�
;c�(;�^9;��A;�[E;��F;�G;��G;�-H;�YH;{H;�H;i�H;u�H;6�H;�H;��H;�H;6�H;u�H;i�H;�H;{H;�YH;�-H;��G;�G;��F;�[E;��A;�^9;c�(;�
;��:��'7(��B�� �ݫ����Ҽ:y��c�����R�ؽe���:�jk�f쏾�ê��þfYؾ��      �þ��������R��f쏾�s��H����������������D�vc�g����f�3,�����P����9/��:5;�i-;��;;��B;+�E;�G;��G;��G;�5H;�_H;�H;{�H;�H;q�H;ɽH;r�H;��H;r�H;ɽH;q�H;�H;{�H;�H;�_H;�5H;��G;��G;�G;+�E;��B;��;;�i-;5;/��:��9�P�����3,��f�g���vc���D���������������H��s�f쏾�R���������      �*���0��ȥ��&���jk��H��#%�B[�ZPν�s��0�f�/%�d��`���G�=�n?ػgFL��D�`�R:B�:��;�2;�=;��C;�/F;�FG;�G;WH;?H;�fH;��H;V�H;ͫH;��H;��H;�H;��H;�H;��H;��H;ͫH;V�H;��H;�fH;?H;WH;�G;�FG;�/F;��C;�=;�2;��;B�:`�R:�D�gFL�n?ػG�=�`���d��/%�0�f��s��ZPνB[��#%��H�jk�&���ȥ���0��      
Dx��s���f�QS���:����B[��7ս�榽��}�u�;��8�)�����r����G������Ҭ����:��;}$;,�6;f�?;3�D;�F;�oG;��G;H;XIH;dnH;i�H;��H;�H;Z�H;��H;��H;G�H;��H;��H;Z�H;�H;��H;i�H;dnH;XIH;H;��G;�oG;�F;3�D;f�?;,�6;}$;��;���:�Ҭ����G�������r�)����8�u�;���}��榽�7սB[������:�QS���f��s�      }�=���:���0��Q"�e�����ZPν�榽%����G�����Ҽ���E:�
�ܻ�D^�ϸ��ih:���:O;�{,;�:;��A;~hE;��F;\�G;��G;�'H;eTH;�vH;��H;L�H;��H;�H;��H;��H;3�H;��H;��H;�H;��H;L�H;��H;�vH;eTH;�'H;��G;\�G;��F;~hE;��A;�:;�{,;O;���:ih:ϸ���D^�
�ܻE:������Ҽ����G�%���榽ZPν����e��Q"���0���:�      ���N9�C[��s�R�ؽ���s����}���G��K��	c��!�V�%,��*�����,����:?��:� ;Ƃ3;0>;�C;"F;#8G;l�G;�H;7H;�_H;,H;�H; �H;g�H;�H;m�H;��H;3�H;��H;m�H;�H;g�H; �H;�H;,H;�_H;7H;�H;l�G;#8G;"F;�C;0>;Ƃ3;� ;?��:��:,������*��%,�!�V�	c��K�����G���}��s����R�ؽ�s�C[�N9�      \Pν��ʽ*8�������������0�f�u�;���K��Ȥ���f���$ߵ�?o5�5�D�L�-:���:X>;G+;_9;�A;��D;[�F;�uG;�G;IH;�FH;�kH;�H;��H;�H;H�H;�H;��H;"�H;F�H;"�H;��H;�H;H�H;�H;��H;�H;�kH;�FH;IH;�G;�uG;[�F;��D;�A;_9;G+;X>;���:L�-:5�D�?o5�$ߵ�����f�Ȥ�K����u�;�0�f������������*8����ʽ      鰒�Z��������}��c���D�/%��8���Ҽ	c����f�����ƻZ/X�u���9f�:ȏ;F";�3;�>;�XC;��E;G;'�G;��G;�+H;/VH;9wH;��H;W�H;�H;.�H;�H;Q�H;`�H;N�H;`�H;Q�H;�H;.�H;�H;W�H;��H;9wH;/VH;�+H;��G;'�G;G;��E;�XC;�>;�3;F";ȏ;f�:9u���Z/X��ƻ�����f�	c����Ҽ�8�/%���D��c���}�����Z��      �&K���G�ȟ>��0�:y�vc�d��)������!�V����ƻgod���º�P(7�3�:���:�;]P.;9�:;ayA;y�D;�F;�mG;t�G;!H;�?H;MeH;��H;R�H;ժH;��H;�H;	�H;��H;��H;V�H;��H;��H;	�H;�H;��H;ժH;R�H;��H;MeH;�?H;!H;t�G;�mG;�F;y�D;ayA;9�:;]P.;�;���:�3�:�P(7��ºgod��ƻ��!�V����)���d��vc�:y��0�ȟ>���G�      xc��8�|����켕�Ҽg���`�����r�E:�%,�$ߵ�Z/X���º̬�E�}:> �:v;��);�l7;i�?;�C;KF;�(G;E�G;�G;2)H;�RH;�sH;��H;��H;�H;ͼH;��H;��H;+�H;��H;l�H;��H;+�H;��H;��H;ͼH;�H;��H;��H;�sH;�RH;2)H;�G;E�G;�(G;KF;�C;i�?;�l7;��);v;> �:E�}:̬���ºZ/X�$ߵ�%,�E:���r�`���g�����Ҽ��|����8�      ����-��#Ȥ�d���ݫ���f�G�=����
�ܻ�*��?o5�u����P(7E�}:�m�:��;>&;��4;B�=;�B;+�E;S�F;ˀG;$�G;cH;�@H;�dH;d�H;��H;x�H;��H;��H;;�H;��H;��H;��H;l�H;��H;��H;��H;;�H;��H;��H;x�H;��H;d�H;�dH;�@H;cH;$�G;ˀG;S�F;+�E;�B;B�=;��4;>&;��;�m�:E�}:�P(7u���?o5��*��
�ܻ���G�=��f�ݫ��d���#Ȥ��-��      ;�V�z5S�Y6H�x�6�� �3,�n?ػG���D^����5�D�9�3�:> �:��;]%;��3;p�<;�B;�
E;>�F;�WG;8�G;t�G;�/H;wVH;�uH;�H;��H;ܰH;��H;��H;��H;j�H;��H;��H;Q�H;��H;��H;j�H;��H;��H;��H;ܰH;��H;�H;�uH;wVH;�/H;t�G;8�G;�WG;>�F;�
E;�B;p�<;��3;]%;��;> �:�3�:95�D�����D^�G��n?ػ3,�� �x�6�Y6H�z5S�      s��w��,�ܻ�ƻB󩻝��gFL����ϸ��,��L�-:f�:���:v;>&;��3;�8<;_�A;%�D;�YF;Z4G;3�G;�G;� H;`IH;VjH;ńH;ٙH;��H;��H;�H;��H;��H;��H;��H;v�H;�H;v�H;��H;��H;��H;��H;�H;��H;��H;ٙH;ńH;VjH;`IH;� H;�G;3�G;Z4G;�YF;%�D;_�A;�8<;��3;>&;v;���:f�:L�-:,��ϸ�����gFL����B��ƻ,�ܻw��      �D^��/X��qF�(}*�(���P���D��Ҭ�ih:��:���:ȏ;�;��);��4;p�<;_�A;f�D;�8F;
G;��G;w�G;jH;C>H;�`H;5|H;��H;��H;��H;��H;��H;|�H;��H;4�H;��H;8�H;��H;8�H;��H;4�H;��H;|�H;��H;��H;��H;��H;��H;5|H;�`H;C>H;jH;w�G;��G;
G;�8F;f�D;_�A;p�<;��4;��);�;ȏ;���:��:ih:�Ҭ��D��P��(��(}*��qF��/X�      ��S���D�1�������'7��9`�R:���:���:?��:X>;F";]P.;�l7;B�=;�B;%�D;�8F;XG;R�G;��G;�H;�5H;�XH;uH;=�H;�H;�H;�H;��H;9�H;��H;-�H;M�H;q�H;��H;�H;��H;q�H;M�H;-�H;��H;9�H;��H;�H;�H;�H;=�H;uH;�XH;�5H;�H;��G;R�G;XG;�8F;%�D;�B;B�=;�l7;]P.;F";X>;?��:���:���:`�R:��9��'7���1����D�      �v[:�Ad:3�}:^�:��:/��:B�:��;O;� ;G+;�3;9�:;i�?;�B;�
E;�YF;
G;R�G;��G;nH;�0H;�RH;�oH;�H;f�H; �H;��H;��H;��H;�H;��H;��H;5�H;�H;(�H;q�H;(�H;�H;5�H;��H;��H;�H;��H;��H;��H; �H;f�H;�H;�oH;�RH;�0H;nH;��G;R�G;
G;�YF;�
E;�B;i�?;9�:;�3;G+;� ;O;��;B�:/��:��:^�:3�}:�Ad:      ���:�A�:���:�w;�
;5;��;}$;�{,;Ƃ3;_9;�>;ayA;�C;+�E;>�F;Z4G;��G;��G;nH;�.H;PH;&lH;i�H;��H;��H;��H;�H;��H;)�H;r�H;��H;��H;��H;y�H;W�H;��H;W�H;y�H;��H;��H;��H;r�H;)�H;��H;�H;��H;��H;��H;i�H;&lH;PH;�.H;nH;��G;��G;Z4G;>�F;+�E;�C;ayA;�>;_9;Ƃ3;�{,;}$;��;5;�
;�w;���:�A�:      �d;� ;�";�%;c�(;�i-;�2;,�6;�:;0>;�A;�XC;y�D;KF;S�F;�WG;3�G;w�G;�H;�0H;PH;�jH;��H;��H;V�H;E�H;�H;��H;��H;�H;��H;��H;��H;�H;��H;j�H;��H;j�H;��H;�H;��H;��H;��H;�H;��H;��H;�H;E�H;V�H;��H;��H;�jH;PH;�0H;�H;w�G;3�G;�WG;S�F;KF;y�D;�XC;�A;0>;�:;,�6;�2;�i-;c�(;�%;�";� ;      ��4;x�4;��5;Rl7;�^9;��;;�=;f�?;��A;�C;��D;��E;�F;�(G;ˀG;8�G;�G;jH;�5H;�RH;&lH;��H;˓H;#�H;گH;g�H;<�H;H�H;��H;��H;(�H;��H;C�H;��H;��H;m�H;��H;m�H;��H;��H;C�H;��H;(�H;��H;��H;H�H;<�H;g�H;گH;#�H;˓H;��H;&lH;�RH;�5H;jH;�G;8�G;ˀG;�(G;�F;��E;��D;�C;��A;f�?;�=;��;;�^9;Rl7;��5;x�4;      �_?;�?;6�?;�@;��A;��B;��C;3�D;~hE;"F;[�F;G;�mG;E�G;$�G;t�G;� H;C>H;�XH;�oH;i�H;��H;#�H;\�H;��H;;�H;X�H;�H;��H;��H;g�H;��H;��H;��H;��H;E�H;^�H;E�H;��H;��H;��H;��H;g�H;��H;��H;�H;X�H;;�H;��H;\�H;#�H;��H;i�H;�oH;�XH;C>H;� H;t�G;$�G;E�G;�mG;G;[�F;"F;~hE;3�D;��C;��B;��A;�@;6�?;�?;      �lD;"~D;��D;�D;�[E;+�E;�/F;�F;��F;#8G;�uG;'�G;t�G;�G;cH;�/H;`IH;�`H;uH;�H;��H;V�H;گH;��H;�H;��H;}�H;#�H;��H;�H;n�H;N�H;��H;��H;��H;��H;6�H;��H;��H;��H;��H;N�H;n�H;�H;��H;#�H;}�H;��H;�H;��H;گH;V�H;��H;�H;uH;�`H;`IH;�/H;cH;�G;t�G;'�G;�uG;#8G;��F;�F;�/F;+�E;�[E;�D;��D;"~D;      ��F;p�F;��F;�F;��F;�G;�FG;�oG;\�G;l�G;�G;��G;!H;2)H;�@H;wVH;VjH;5|H;=�H;f�H;��H;E�H;g�H;;�H;��H;E�H;��H;��H;��H;�H;�H;��H;��H;��H;B�H;��H;��H;��H;B�H;��H;��H;��H;�H;�H;��H;��H;��H;E�H;��H;;�H;g�H;E�H;��H;f�H;=�H;5|H;VjH;wVH;�@H;2)H;!H;��G;�G;l�G;\�G;�oG;�FG;�G;��F;�F;��F;p�F;      puG;3xG;/�G;��G;�G;��G;�G;��G;��G;�H;IH;�+H;�?H;�RH;�dH;�uH;ńH;��H;�H; �H;��H;�H;<�H;X�H;}�H;��H;t�H;l�H;��H;��H;n�H;��H;��H;L�H;��H;-�H;.�H;-�H;��H;L�H;��H;��H;n�H;��H;��H;l�H;t�H;��H;}�H;X�H;<�H;�H;��H; �H;�H;��H;ńH;�uH;�dH;�RH;�?H;�+H;IH;�H;��G;��G;�G;��G;�G;��G;/�G;3xG;      M�G;��G;��G;��G;��G;��G;WH;H;�'H;7H;�FH;/VH;MeH;�sH;d�H;�H;ٙH;��H;�H;��H;�H;��H;H�H;�H;#�H;��H;l�H;��H;��H;p�H;��H;��H;c�H;��H;U�H;��H;��H;��H;U�H;��H;c�H;��H;��H;p�H;��H;��H;l�H;��H;#�H;�H;H�H;��H;�H;��H;�H;��H;ٙH;�H;d�H;�sH;MeH;/VH;�FH;7H;�'H;H;WH;��G;��G;��G;��G;��G;      �H;�H;s"H;3'H;�-H;�5H;?H;XIH;eTH;�_H;�kH;9wH;��H;��H;��H;��H;��H;��H;�H;��H;��H;��H;��H;��H;��H;��H;��H;��H;>�H;��H;��H;X�H;��H;y�H;��H;��H;��H;��H;��H;y�H;��H;X�H;��H;��H;>�H;��H;��H;��H;��H;��H;��H;��H;��H;��H;�H;��H;��H;��H;��H;��H;��H;9wH;�kH;�_H;eTH;XIH;?H;�5H;�-H;3'H;s"H;�H;      �NH;NOH;�QH;UH;�YH;�_H;�fH;dnH;�vH;,H;�H;��H;R�H;��H;x�H;ܰH;��H;��H;��H;��H;)�H;�H;��H;��H;�H;�H;��H;p�H;��H;��H;V�H;��H;q�H;��H;�H;%�H;?�H;%�H;�H;��H;q�H;��H;V�H;��H;��H;p�H;��H;�H;�H;��H;��H;�H;)�H;��H;��H;��H;��H;ܰH;x�H;��H;R�H;��H;�H;,H;�vH;dnH;�fH;�_H;�YH;UH;�QH;NOH;      �rH;HsH;�tH;�wH;{H;�H;��H;i�H;��H;�H;��H;W�H;ժH;�H;��H;��H;�H;��H;9�H;�H;r�H;��H;(�H;g�H;n�H;�H;n�H;��H;��H;V�H;��H;q�H;��H;�H;_�H;l�H;d�H;l�H;_�H;�H;��H;q�H;��H;V�H;��H;��H;n�H;�H;n�H;g�H;(�H;��H;r�H;�H;9�H;��H;�H;��H;��H;�H;ժH;W�H;��H;�H;��H;i�H;��H;�H;{H;�wH;�tH;HsH;      �H;:�H;y�H;�H;�H;{�H;V�H;��H;L�H; �H;�H;�H;��H;ͼH;��H;��H;��H;|�H;��H;��H;��H;��H;��H;��H;N�H;��H;��H;��H;X�H;��H;q�H;��H;�H;_�H;��H;��H;��H;��H;��H;_�H;�H;��H;q�H;��H;X�H;��H;��H;��H;N�H;��H;��H;��H;��H;��H;��H;|�H;��H;��H;��H;ͼH;��H;�H;�H; �H;L�H;��H;V�H;{�H;�H;�H;y�H;:�H;      ��H;�H;�H;f�H;i�H;�H;ͫH;�H;��H;g�H;H�H;.�H;�H;��H;;�H;��H;��H;��H;-�H;��H;��H;��H;C�H;��H;��H;��H;��H;c�H;��H;q�H;��H;�H;X�H;��H;��H;��H;��H;��H;��H;��H;X�H;�H;��H;q�H;��H;c�H;��H;��H;��H;��H;C�H;��H;��H;��H;-�H;��H;��H;��H;;�H;��H;�H;.�H;H�H;g�H;��H;�H;ͫH;�H;i�H;f�H;�H;�H;      ��H;�H;��H;±H;u�H;q�H;��H;Z�H;�H;�H;�H;�H;	�H;��H;��H;j�H;��H;4�H;M�H;5�H;��H;�H;��H;��H;��H;��H;L�H;��H;y�H;��H;�H;_�H;��H;��H;��H;��H;��H;��H;��H;��H;��H;_�H;�H;��H;y�H;��H;L�H;��H;��H;��H;��H;�H;��H;5�H;M�H;4�H;��H;j�H;��H;��H;	�H;�H;�H;�H;�H;Z�H;��H;q�H;u�H;±H;��H;�H;      �H;W�H;�H;ۺH;6�H;ɽH;��H;��H;��H;m�H;��H;Q�H;��H;+�H;��H;��H;��H;��H;q�H;�H;y�H;��H;��H;��H;��H;B�H;��H;U�H;��H;�H;_�H;��H;��H;��H;��H;��H;��H;��H;��H;��H;��H;��H;_�H;�H;��H;U�H;��H;B�H;��H;��H;��H;��H;y�H;�H;q�H;��H;��H;��H;��H;+�H;��H;Q�H;��H;m�H;��H;��H;��H;ɽH;6�H;ۺH;�H;W�H;      q�H;��H;�H;�H;�H;r�H;�H;��H;��H;��H;"�H;`�H;��H;��H;��H;��H;v�H;8�H;��H;(�H;W�H;j�H;m�H;E�H;��H;��H;-�H;��H;��H;%�H;l�H;��H;��H;��H;��H;��H;��H;��H;��H;��H;��H;��H;l�H;%�H;��H;��H;-�H;��H;��H;E�H;m�H;j�H;W�H;(�H;��H;8�H;v�H;��H;��H;��H;��H;`�H;"�H;��H;��H;��H;�H;r�H;�H;�H;�H;��H;      E�H;U�H;��H;��H;��H;��H;��H;G�H;3�H;3�H;F�H;N�H;V�H;l�H;l�H;Q�H;�H;��H;�H;q�H;��H;��H;��H;^�H;6�H;��H;.�H;��H;��H;?�H;d�H;��H;��H;��H;��H;��H;��H;��H;��H;��H;��H;��H;d�H;?�H;��H;��H;.�H;��H;6�H;^�H;��H;��H;��H;q�H;�H;��H;�H;Q�H;l�H;l�H;V�H;N�H;F�H;3�H;3�H;G�H;��H;��H;��H;��H;��H;U�H;      q�H;��H;�H;�H;�H;r�H;�H;��H;��H;��H;"�H;`�H;��H;��H;��H;��H;v�H;8�H;��H;(�H;W�H;j�H;m�H;E�H;��H;��H;-�H;��H;��H;%�H;l�H;��H;��H;��H;��H;��H;��H;��H;��H;��H;��H;��H;l�H;%�H;��H;��H;-�H;��H;��H;E�H;m�H;j�H;W�H;(�H;��H;8�H;v�H;��H;��H;��H;��H;`�H;"�H;��H;��H;��H;�H;r�H;�H;�H;�H;��H;      �H;W�H;�H;ۺH;6�H;ɽH;��H;��H;��H;m�H;��H;Q�H;��H;+�H;��H;��H;��H;��H;q�H;�H;y�H;��H;��H;��H;��H;B�H;��H;U�H;��H;�H;_�H;��H;��H;��H;��H;��H;��H;��H;��H;��H;��H;��H;_�H;�H;��H;U�H;��H;B�H;��H;��H;��H;��H;y�H;�H;q�H;��H;��H;��H;��H;+�H;��H;Q�H;��H;m�H;��H;��H;��H;ɽH;6�H;ۺH;�H;W�H;      ��H;�H;��H;±H;u�H;q�H;��H;Z�H;�H;�H;�H;�H;	�H;��H;��H;j�H;��H;4�H;M�H;5�H;��H;�H;��H;��H;��H;��H;L�H;��H;y�H;��H;�H;_�H;��H;��H;��H;��H;��H;��H;��H;��H;��H;_�H;�H;��H;y�H;��H;L�H;��H;��H;��H;��H;�H;��H;5�H;M�H;4�H;��H;j�H;��H;��H;	�H;�H;�H;�H;�H;Z�H;��H;q�H;u�H;±H;��H;�H;      ��H;�H;�H;f�H;i�H;�H;ͫH;�H;��H;g�H;H�H;.�H;�H;��H;;�H;��H;��H;��H;-�H;��H;��H;��H;C�H;��H;��H;��H;��H;c�H;��H;q�H;��H;�H;X�H;��H;��H;��H;��H;��H;��H;��H;X�H;�H;��H;q�H;��H;c�H;��H;��H;��H;��H;C�H;��H;��H;��H;-�H;��H;��H;��H;;�H;��H;�H;.�H;H�H;g�H;��H;�H;ͫH;�H;i�H;f�H;�H;�H;      �H;:�H;y�H;�H;�H;{�H;V�H;��H;L�H; �H;�H;�H;��H;ͼH;��H;��H;��H;|�H;��H;��H;��H;��H;��H;��H;N�H;��H;��H;��H;X�H;��H;q�H;��H;�H;_�H;��H;��H;��H;��H;��H;_�H;�H;��H;q�H;��H;X�H;��H;��H;��H;N�H;��H;��H;��H;��H;��H;��H;|�H;��H;��H;��H;ͼH;��H;�H;�H; �H;L�H;��H;V�H;{�H;�H;�H;y�H;:�H;      �rH;HsH;�tH;�wH;{H;�H;��H;i�H;��H;�H;��H;W�H;ժH;�H;��H;��H;�H;��H;9�H;�H;r�H;��H;(�H;g�H;n�H;�H;n�H;��H;��H;V�H;��H;q�H;��H;�H;_�H;l�H;d�H;l�H;_�H;�H;��H;q�H;��H;V�H;��H;��H;n�H;�H;n�H;g�H;(�H;��H;r�H;�H;9�H;��H;�H;��H;��H;�H;ժH;W�H;��H;�H;��H;i�H;��H;�H;{H;�wH;�tH;HsH;      �NH;NOH;�QH;UH;�YH;�_H;�fH;dnH;�vH;,H;�H;��H;R�H;��H;x�H;ܰH;��H;��H;��H;��H;)�H;�H;��H;��H;�H;�H;��H;p�H;��H;��H;V�H;��H;q�H;��H;�H;%�H;?�H;%�H;�H;��H;q�H;��H;V�H;��H;��H;p�H;��H;�H;�H;��H;��H;�H;)�H;��H;��H;��H;��H;ܰH;x�H;��H;R�H;��H;�H;,H;�vH;dnH;�fH;�_H;�YH;UH;�QH;NOH;      �H;�H;s"H;3'H;�-H;�5H;?H;XIH;eTH;�_H;�kH;9wH;��H;��H;��H;��H;��H;��H;�H;��H;��H;��H;��H;��H;��H;��H;��H;��H;>�H;��H;��H;X�H;��H;y�H;��H;��H;��H;��H;��H;y�H;��H;X�H;��H;��H;>�H;��H;��H;��H;��H;��H;��H;��H;��H;��H;�H;��H;��H;��H;��H;��H;��H;9wH;�kH;�_H;eTH;XIH;?H;�5H;�-H;3'H;s"H;�H;      M�G;��G;��G;��G;��G;��G;WH;H;�'H;7H;�FH;/VH;MeH;�sH;d�H;�H;ٙH;��H;�H;��H;�H;��H;H�H;�H;#�H;��H;l�H;��H;��H;p�H;��H;��H;c�H;��H;U�H;��H;��H;��H;U�H;��H;c�H;��H;��H;p�H;��H;��H;l�H;��H;#�H;�H;H�H;��H;�H;��H;�H;��H;ٙH;�H;d�H;�sH;MeH;/VH;�FH;7H;�'H;H;WH;��G;��G;��G;��G;��G;      puG;3xG;/�G;��G;�G;��G;�G;��G;��G;�H;IH;�+H;�?H;�RH;�dH;�uH;ńH;��H;�H; �H;��H;�H;<�H;X�H;}�H;��H;t�H;l�H;��H;��H;n�H;��H;��H;L�H;��H;-�H;.�H;-�H;��H;L�H;��H;��H;n�H;��H;��H;l�H;t�H;��H;}�H;X�H;<�H;�H;��H; �H;�H;��H;ńH;�uH;�dH;�RH;�?H;�+H;IH;�H;��G;��G;�G;��G;�G;��G;/�G;3xG;      ��F;p�F;��F;�F;��F;�G;�FG;�oG;\�G;l�G;�G;��G;!H;2)H;�@H;wVH;VjH;5|H;=�H;f�H;��H;E�H;g�H;;�H;��H;E�H;��H;��H;��H;�H;�H;��H;��H;��H;B�H;��H;��H;��H;B�H;��H;��H;��H;�H;�H;��H;��H;��H;E�H;��H;;�H;g�H;E�H;��H;f�H;=�H;5|H;VjH;wVH;�@H;2)H;!H;��G;�G;l�G;\�G;�oG;�FG;�G;��F;�F;��F;p�F;      �lD;"~D;��D;�D;�[E;+�E;�/F;�F;��F;#8G;�uG;'�G;t�G;�G;cH;�/H;`IH;�`H;uH;�H;��H;V�H;گH;��H;�H;��H;}�H;#�H;��H;�H;n�H;N�H;��H;��H;��H;��H;6�H;��H;��H;��H;��H;N�H;n�H;�H;��H;#�H;}�H;��H;�H;��H;گH;V�H;��H;�H;uH;�`H;`IH;�/H;cH;�G;t�G;'�G;�uG;#8G;��F;�F;�/F;+�E;�[E;�D;��D;"~D;      �_?;�?;6�?;�@;��A;��B;��C;3�D;~hE;"F;[�F;G;�mG;E�G;$�G;t�G;� H;C>H;�XH;�oH;i�H;��H;#�H;\�H;��H;;�H;X�H;�H;��H;��H;g�H;��H;��H;��H;��H;E�H;^�H;E�H;��H;��H;��H;��H;g�H;��H;��H;�H;X�H;;�H;��H;\�H;#�H;��H;i�H;�oH;�XH;C>H;� H;t�G;$�G;E�G;�mG;G;[�F;"F;~hE;3�D;��C;��B;��A;�@;6�?;�?;      ��4;x�4;��5;Rl7;�^9;��;;�=;f�?;��A;�C;��D;��E;�F;�(G;ˀG;8�G;�G;jH;�5H;�RH;&lH;��H;˓H;#�H;گH;g�H;<�H;H�H;��H;��H;(�H;��H;C�H;��H;��H;m�H;��H;m�H;��H;��H;C�H;��H;(�H;��H;��H;H�H;<�H;g�H;گH;#�H;˓H;��H;&lH;�RH;�5H;jH;�G;8�G;ˀG;�(G;�F;��E;��D;�C;��A;f�?;�=;��;;�^9;Rl7;��5;x�4;      �d;� ;�";�%;c�(;�i-;�2;,�6;�:;0>;�A;�XC;y�D;KF;S�F;�WG;3�G;w�G;�H;�0H;PH;�jH;��H;��H;V�H;E�H;�H;��H;��H;�H;��H;��H;��H;�H;��H;j�H;��H;j�H;��H;�H;��H;��H;��H;�H;��H;��H;�H;E�H;V�H;��H;��H;�jH;PH;�0H;�H;w�G;3�G;�WG;S�F;KF;y�D;�XC;�A;0>;�:;,�6;�2;�i-;c�(;�%;�";� ;      ���:�A�:���:�w;�
;5;��;}$;�{,;Ƃ3;_9;�>;ayA;�C;+�E;>�F;Z4G;��G;��G;nH;�.H;PH;&lH;i�H;��H;��H;��H;�H;��H;)�H;r�H;��H;��H;��H;y�H;W�H;��H;W�H;y�H;��H;��H;��H;r�H;)�H;��H;�H;��H;��H;��H;i�H;&lH;PH;�.H;nH;��G;��G;Z4G;>�F;+�E;�C;ayA;�>;_9;Ƃ3;�{,;}$;��;5;�
;�w;���:�A�:      �v[:�Ad:3�}:^�:��:/��:B�:��;O;� ;G+;�3;9�:;i�?;�B;�
E;�YF;
G;R�G;��G;nH;�0H;�RH;�oH;�H;f�H; �H;��H;��H;��H;�H;��H;��H;5�H;�H;(�H;q�H;(�H;�H;5�H;��H;��H;�H;��H;��H;��H; �H;f�H;�H;�oH;�RH;�0H;nH;��G;R�G;
G;�YF;�
E;�B;i�?;9�:;�3;G+;� ;O;��;B�:/��:��:^�:3�}:�Ad:      ��S���D�1�������'7��9`�R:���:���:?��:X>;F";]P.;�l7;B�=;�B;%�D;�8F;XG;R�G;��G;�H;�5H;�XH;uH;=�H;�H;�H;�H;��H;9�H;��H;-�H;M�H;q�H;��H;�H;��H;q�H;M�H;-�H;��H;9�H;��H;�H;�H;�H;=�H;uH;�XH;�5H;�H;��G;R�G;XG;�8F;%�D;�B;B�=;�l7;]P.;F";X>;?��:���:���:`�R:��9��'7���1����D�      �D^��/X��qF�(}*�(���P���D��Ҭ�ih:��:���:ȏ;�;��);��4;p�<;_�A;f�D;�8F;
G;��G;w�G;jH;C>H;�`H;5|H;��H;��H;��H;��H;��H;|�H;��H;4�H;��H;8�H;��H;8�H;��H;4�H;��H;|�H;��H;��H;��H;��H;��H;5|H;�`H;C>H;jH;w�G;��G;
G;�8F;f�D;_�A;p�<;��4;��);�;ȏ;���:��:ih:�Ҭ��D��P��(��(}*��qF��/X�      s��w��,�ܻ�ƻB󩻝��gFL����ϸ��,��L�-:f�:���:v;>&;��3;�8<;_�A;%�D;�YF;Z4G;3�G;�G;� H;`IH;VjH;ńH;ٙH;��H;��H;�H;��H;��H;��H;��H;v�H;�H;v�H;��H;��H;��H;��H;�H;��H;��H;ٙH;ńH;VjH;`IH;� H;�G;3�G;Z4G;�YF;%�D;_�A;�8<;��3;>&;v;���:f�:L�-:,��ϸ�����gFL����B��ƻ,�ܻw��      ;�V�z5S�Y6H�x�6�� �3,�n?ػG���D^����5�D�9�3�:> �:��;]%;��3;p�<;�B;�
E;>�F;�WG;8�G;t�G;�/H;wVH;�uH;�H;��H;ܰH;��H;��H;��H;j�H;��H;��H;Q�H;��H;��H;j�H;��H;��H;��H;ܰH;��H;�H;�uH;wVH;�/H;t�G;8�G;�WG;>�F;�
E;�B;p�<;��3;]%;��;> �:�3�:95�D�����D^�G��n?ػ3,�� �x�6�Y6H�z5S�      ����-��#Ȥ�d���ݫ���f�G�=����
�ܻ�*��?o5�u����P(7E�}:�m�:��;>&;��4;B�=;�B;+�E;S�F;ˀG;$�G;cH;�@H;�dH;d�H;��H;x�H;��H;��H;;�H;��H;��H;��H;l�H;��H;��H;��H;;�H;��H;��H;x�H;��H;d�H;�dH;�@H;cH;$�G;ˀG;S�F;+�E;�B;B�=;��4;>&;��;�m�:E�}:�P(7u���?o5��*��
�ܻ���G�=��f�ݫ��d���#Ȥ��-��      xc��8�|����켕�Ҽg���`�����r�E:�%,�$ߵ�Z/X���º̬�E�}:> �:v;��);�l7;i�?;�C;KF;�(G;E�G;�G;2)H;�RH;�sH;��H;��H;�H;ͼH;��H;��H;+�H;��H;l�H;��H;+�H;��H;��H;ͼH;�H;��H;��H;�sH;�RH;2)H;�G;E�G;�(G;KF;�C;i�?;�l7;��);v;> �:E�}:̬���ºZ/X�$ߵ�%,�E:���r�`���g�����Ҽ��|����8�      �&K���G�ȟ>��0�:y�vc�d��)������!�V����ƻgod���º�P(7�3�:���:�;]P.;9�:;ayA;y�D;�F;�mG;t�G;!H;�?H;MeH;��H;R�H;ժH;��H;�H;	�H;��H;��H;V�H;��H;��H;	�H;�H;��H;ժH;R�H;��H;MeH;�?H;!H;t�G;�mG;�F;y�D;ayA;9�:;]P.;�;���:�3�:�P(7��ºgod��ƻ��!�V����)���d��vc�:y��0�ȟ>���G�      鰒�Z��������}��c���D�/%��8���Ҽ	c����f�����ƻZ/X�u���9f�:ȏ;F";�3;�>;�XC;��E;G;'�G;��G;�+H;/VH;9wH;��H;W�H;�H;.�H;�H;Q�H;`�H;N�H;`�H;Q�H;�H;.�H;�H;W�H;��H;9wH;/VH;�+H;��G;'�G;G;��E;�XC;�>;�3;F";ȏ;f�:9u���Z/X��ƻ�����f�	c����Ҽ�8�/%���D��c���}�����Z��      \Pν��ʽ*8�������������0�f�u�;���K��Ȥ���f���$ߵ�?o5�5�D�L�-:���:X>;G+;_9;�A;��D;[�F;�uG;�G;IH;�FH;�kH;�H;��H;�H;H�H;�H;��H;"�H;F�H;"�H;��H;�H;H�H;�H;��H;�H;�kH;�FH;IH;�G;�uG;[�F;��D;�A;_9;G+;X>;���:L�-:5�D�?o5�$ߵ�����f�Ȥ�K����u�;�0�f������������*8����ʽ      ���N9�C[��s�R�ؽ���s����}���G��K��	c��!�V�%,��*�����,����:?��:� ;Ƃ3;0>;�C;"F;#8G;l�G;�H;7H;�_H;,H;�H; �H;g�H;�H;m�H;��H;3�H;��H;m�H;�H;g�H; �H;�H;,H;�_H;7H;�H;l�G;#8G;"F;�C;0>;Ƃ3;� ;?��:��:,������*��%,�!�V�	c��K�����G���}��s����R�ؽ�s�C[�N9�      }�=���:���0��Q"�e�����ZPν�榽%����G�����Ҽ���E:�
�ܻ�D^�ϸ��ih:���:O;�{,;�:;��A;~hE;��F;\�G;��G;�'H;eTH;�vH;��H;L�H;��H;�H;��H;��H;3�H;��H;��H;�H;��H;L�H;��H;�vH;eTH;�'H;��G;\�G;��F;~hE;��A;�:;�{,;O;���:ih:ϸ���D^�
�ܻE:������Ҽ����G�%���榽ZPν����e��Q"���0���:�      
Dx��s���f�QS���:����B[��7ս�榽��}�u�;��8�)�����r����G������Ҭ����:��;}$;,�6;f�?;3�D;�F;�oG;��G;H;XIH;dnH;i�H;��H;�H;Z�H;��H;��H;G�H;��H;��H;Z�H;�H;��H;i�H;dnH;XIH;H;��G;�oG;�F;3�D;f�?;,�6;}$;��;���:�Ҭ����G�������r�)����8�u�;���}��榽�7սB[������:�QS���f��s�      �*���0��ȥ��&���jk��H��#%�B[�ZPν�s��0�f�/%�d��`���G�=�n?ػgFL��D�`�R:B�:��;�2;�=;��C;�/F;�FG;�G;WH;?H;�fH;��H;V�H;ͫH;��H;��H;�H;��H;�H;��H;��H;ͫH;V�H;��H;�fH;?H;WH;�G;�FG;�/F;��C;�=;�2;��;B�:`�R:�D�gFL�n?ػG�=�`���d��/%�0�f��s��ZPνB[��#%��H�jk�&���ȥ���0��      �þ��������R��f쏾�s��H����������������D�vc�g����f�3,�����P����9/��:5;�i-;��;;��B;+�E;�G;��G;��G;�5H;�_H;�H;{�H;�H;q�H;ɽH;r�H;��H;r�H;ɽH;q�H;�H;{�H;�H;�_H;�5H;��G;��G;�G;+�E;��B;��;;�i-;5;/��:��9�P�����3,��f�g���vc���D���������������H��s�f쏾�R���������      ����fYؾ�þ�ê�f쏾jk���:�e�R�ؽ�����c�:y���Ҽݫ��� �B�(����'7��:�
;c�(;�^9;��A;�[E;��F;�G;��G;�-H;�YH;{H;�H;i�H;u�H;6�H;�H;��H;�H;6�H;u�H;i�H;�H;{H;�YH;�-H;��G;�G;��F;�[E;��A;�^9;c�(;�
;��:��'7(��B�� �ݫ����Ҽ:y��c�����R�ؽe���:�jk�f쏾�ê��þfYؾ��      ��=������I��þ�R��&���QS��Q"��s�����}��0���d���x�6��ƻ(}*����^�:�w;�%;Rl7;�@;�D;�F;��G;��G;3'H;UH;�wH;�H;f�H;±H;ۺH;�H;��H;�H;ۺH;±H;f�H;�H;�wH;UH;3'H;��G;��G;�F;�D;�@;Rl7;�%;�w;^�:���(}*��ƻx�6�d����켟0���}�����s��Q"�QS�&����R���þIᾁ���=��      ���>��&�
�����fYؾ���ȥ����f���0�C[�*8������ȟ>�|���#Ȥ�Y6H�,�ܻ�qF�1��3�}:���:�";��5;6�?;��D;��F;/�G;��G;s"H;�QH;�tH;y�H;�H;��H;�H;�H;��H;�H;�H;��H;�H;y�H;�tH;�QH;s"H;��G;/�G;��F;��D;6�?;��5;�";���:3�}:1���qF�,�ܻY6H�#Ȥ�|���ȟ>�����*8��C[���0���f�ȥ�����fYؾ����&�
�>��      �� �k��>��=���������0���s���:�N9���ʽZ����G��8��-��z5S�w���/X���D��Ad:�A�:� ;x�4;�?;"~D;p�F;3xG;��G;�H;NOH;HsH;:�H;�H;�H;W�H;��H;U�H;��H;W�H;�H;�H;:�H;HsH;NOH;�H;��G;3xG;p�F;"~D;�?;x�4;� ;�A�:�Ad:��D��/X�w��z5S��-���8���G�Z����ʽN9���:��s��0��������=��>��k��      3F�/h��ǰ�3Vھ�������~���S��#��o��S��R₽�6�-���<y��FB��Eֻ_A?��	�Y�:���:�";�36;�@;��D;�F;�mG;%�G;>H;9?H;fH;w�H;P�H;��H;��H;�H;�H;�H;��H;��H;P�H;w�H;fH;9?H;>H;%�G;�mG;�F;��D;�@;�36;�";���:Y�:�	�_A?��EֻFB�<y��-����6�R₽S���o���#��S��~��������3Vھǰ�/h��      /h���b���쾅*־�v������)�� �O�6� ��r�r���؀��3����ݜ��>��ѻ��9�����n�:�$ ;�L#;˃6;�@@;B�D;�F;<pG;��G;TH;@H;�fH;�H;��H;�H;=�H;�H;��H;�H;=�H;�H;��H;�H;�fH;@H;TH;��G;<pG;�F;B�D;�@@;˃6;�L#;�$ ;�n�:�����9��ѻ�>�ݜ�����3��؀��r���r�6� � �O��)������v���*־�쾼b��      ǰ�쾐�޾5ʾ/;���:����v��E�A'���L����u�X�+�bW缨A��s�4�n�Ļ�8)��j��W�:�;�%;kk7;f�@;A�D;4�F;wG;��G;uH;cBH;YhH;B�H;��H;ƩH;�H;��H;��H;��H;�H;ƩH;��H;B�H;YhH;cBH;uH;��G;wG;4�F;A�D;f�@;kk7;�%;�;W�:�j���8)�n�Ļs�4��A��bW�X�+���u�L����A'��E���v��:��/;��5ʾ��޾��      3Vھ�*־5ʾT��������M���9b��5���}�սn���Xc�ݟ���ռ�I��$�$�4T���Z�*_����:��;��';��8;]QA;�8E;��F;�G;%�G;�H;-FH;?kH;u�H;Z�H;�H;�H;��H;t�H;��H;�H;�H;Z�H;u�H;?kH;-FH;�H;%�G;�G;��F;�8E;]QA;��8;��';��;��:*_���Z�4T��$�$��I����ռݟ��Xc�n��}�ս���5��9b��M������T���5ʾ�*־      ���v��/;������:P���r�U�H�6� ��~��@������Q�K�<��վ���s�G��`񕻀ܺ�2u9�%�:��;��+;��:;"B;��E;,�F;��G;�G;mH;[KH;'oH;j�H;��H;ŬH;_�H;��H;��H;��H;_�H;ŬH;��H;j�H;'oH;[KH;mH;�G;��G;,�F;��E;"B;��:;��+;��;�%�:�2u9�ܺ`�G����s��վ�<�Q�K�����@���~��6� �U�H��r�:P������/;���v��      ��������:���M���r� �O��",�<�
��gٽKĥ�|�u�K1�(����Τ�m�P��Z�r.o�lp���:Ӵ�:{P;��/;��<;F
C;e�E;� G;^�G;5�G;�$H;�QH;�sH;$�H;f�H;��H;*�H;{�H;&�H;{�H;*�H;��H;f�H;$�H;�sH;�QH;�$H;5�G;^�G;� G;e�E;F
C;��<;��/;{P;Ӵ�:�:lp��r.o��Z�m�P��Τ�(���K1�|�u�Kĥ��gٽ<�
��",� �O��r��M���:�����      �~���)����v��9b�U�H��",�0Z���S��X^��e�N�{����μ�I���%+�ۚ����.������i~:���:�l;@�3;��>;�C;�OF;�EG;{�G;"�G;�.H;'YH;�yH;p�H;��H;��H;E�H;J�H;��H;J�H;E�H;��H;��H;p�H;�yH;'YH;�.H;"�G;{�G;�EG;�OF;�C;��>;@�3;�l;���:�i~:������.�ۚ���%+��I����μ{��e�N�X^��S����0Z��",�U�H��9b���v��)��      �S� �O��E��5�6� �<�
���|9��l���Xc���(����߈��Z�[����oݎ�ܺ?99���:��	;�c';��7;��@;��D;.�F;aiG;��G;�H;�9H;faH;�H;/�H;O�H;g�H;��H;Y�H;��H;Y�H;��H;g�H;O�H;/�H;�H;faH;�9H;�H;��G;aiG;.�F;��D;��@;��7;�c';��	;���:?99ܺoݎ����Z�[�߈�������(��Xc�l��|9����<�
�6� ��5��E� �O�      �#�6� �A'����~���gٽS��l���j��3�ji��վ�T����(�Q�Ļ,A?���B�4�@:[�:�P;v�.;P�;;�sB;[�E;��F;l�G;'�G;H;�EH;JjH;��H;H�H;.�H;��H;0�H;��H;�H;��H;0�H;��H;.�H;H�H;��H;JjH;�EH;H;'�G;l�G;��F;[�E;�sB;P�;;v�.;�P;[�:4�@:��B�,A?�Q�Ļ�(�T����վ�ji��3��j�l��S���gٽ�~����A'�6� �      �o���r���}�ս@��Kĥ�X^���Xc��3���	���˼t]��FB��Z򻆜��EӺ&��8�:z�;QM#;�<5;x?;��C;�?F;J9G;,�G;M�G;c&H;�QH;�sH;ۍH;��H;H�H;кH;��H;��H;a�H;��H;��H;кH;H�H;��H;ۍH;�sH;�QH;c&H;M�G;,�G;J9G;�?F;��C;x?;�<5;QM#;z�;�:&��8EӺ�����Z�FB�t]����˼��	��3��Xc�X^��Kĥ�@��}�ս���r�      S���r��L��n������|�u�e�N���(�ji���˼�A��b�P�=s��|������\:~�:�;�m-;E�:;N�A;�+E;��F;lnG;,�G;�H;�6H;j^H;/}H;�H;&�H;��H;/�H;��H;Y�H;��H;Y�H;��H;/�H;��H;&�H;�H;/}H;j^H;�6H;�H;,�G;lnG;��F;�+E;N�A;E�:;�m-;�;~�:�\:����|��=s�b�P��A����˼ji���(�e�N�|�u�����n��L���r��      R₽�؀���u��Xc�Q�K�K1�{�����վ�t]��b�P�m��	T��h�9��o�g2�9�%�:��	;�%;��5;�>;��C;F;� G;ݙG;�G;oH;�GH;�jH;ʆH;r�H;��H;̸H;��H;l�H;��H;��H;��H;l�H;��H;̸H;��H;r�H;ʆH;�jH;�GH;oH;�G;ݙG;� G;F;��C;�>;��5;�%;��	;�%�:g2�9�o�h�9�	T��m��b�P�t]���վ����{��K1�Q�K��Xc���u��؀�      �6��3�X�+�ݟ�<�(�����μ߈��T���FB�=s�	T����D��{���8u90q�:���:�X;`t0;S�;;1B;C9E;.�F;9gG;�G;<�G;�/H;�WH;SwH;G�H;��H;#�H;�H;��H;2�H;I�H;S�H;I�H;2�H;��H;�H;#�H;��H;G�H;SwH;�WH;�/H;<�G;�G;9gG;.�F;C9E;1B;S�;;`t0;�X;���:0q�:�8u9�{����D�	T��=s�FB�T���߈����μ(���<�ݟ�X�+��3�      -������bW缑�ռ�վ��Τ��I��Z�[��(��Z�h�9��{���99�W�:�W�:�P;�,;�8;�@@;YAD;�?F;�+G;ÛG;��G;�H;�CH;GgH;W�H;y�H;��H;�H;=�H;:�H;��H;��H;��H;��H;��H;:�H;=�H;�H;��H;y�H;W�H;GgH;�CH;�H;��G;ÛG;�+G;�?F;YAD;�@@;�8;�,;�P;�W�:�W�:�99�{��h�9���Z��(�Z�[��I���Τ��վ���ռbW缧��      <y��ݜ��A���I����s�m�P��%+����Q�Ļ����|��o��8u9�W�:8+�:�;]);8�6;װ>;�OC;��E;9�F;�wG;`�G;� H;�0H;@WH;)vH;ԎH;8�H;#�H;��H;4�H;^�H;��H;�H;��H;�H;��H;^�H;4�H;��H;#�H;8�H;ԎH;)vH;@WH;�0H;� H;`�G;�wG;9�F;��E;�OC;װ>;8�6;]);�;8+�:�W�:�8u9�o�|�����Q�Ļ����%+�m�P���s��I���A��ݜ�      FB��>�s�4�$�$�G���Z�ۚ��oݎ�,A?�EӺ����g2�90q�:�W�:�;D�';�<5;֜=;Z�B;jFE;��F;�TG;Y�G;�G;�H;�GH;9iH;�H;��H;f�H;T�H;f�H;��H;[�H;'�H;5�H;��H;5�H;'�H;[�H;��H;f�H;T�H;f�H;��H;�H;9iH;�GH;�H;�G;Y�G;�TG;��F;jFE;Z�B;֜=;�<5;D�';�;�W�:0q�:g2�9����EӺ,A?�oݎ�ۚ���Z�G��$�$�s�4��>�      �Eֻ�ѻn�Ļ4T��`�r.o���.�ܺ��B�&��8�\:�%�:���:�P;]);�<5;K:=;x"B;��D;!uF;+6G;��G;��G;�H;�9H;9]H;�yH;�H;��H;�H;'�H;��H;u�H;6�H;��H;B�H;��H;B�H;��H;6�H;u�H;��H;'�H;�H;��H;�H;�yH;9]H;�9H;�H;��G;��G;+6G;!uF;��D;x"B;K:=;�<5;]);�P;���:�%�:�\:&��8��B�ܺ��.�r.o�`�4T��n�Ļ�ѻ      _A?���9��8)��Z��ܺlp������?994�@:�:~�:��	;�X;�,;8�6;֜=;x"B;�D;�WF;!G;��G;S�G;�H; .H;�RH;�pH;�H;ԜH;��H;׸H;��H;��H;��H;��H;��H;0�H;��H;0�H;��H;��H;��H;��H;��H;׸H;��H;ԜH;�H;�pH;�RH; .H;�H;S�G;��G;!G;�WF;�D;x"B;֜=;8�6;�,;�X;��	;~�:�:4�@:?99����lp���ܺ�Z��8)���9�      �	�����j��*_���2u9�:�i~:���:[�:z�;�;�%;`t0;�8;װ>;Z�B;��D;�WF;sG;��G;��G;��G;%H;-JH;�hH;�H;��H;T�H;��H;�H;x�H;��H;��H;H�H;��H;��H;h�H;��H;��H;H�H;��H;��H;x�H;�H;��H;T�H;��H;�H;�hH;-JH;%H;��G;��G;��G;sG;�WF;��D;Z�B;װ>;�8;`t0;�%;�;z�;[�:���:�i~:�:�2u9*_���j�����      Y�:�n�:W�:��:�%�:Ӵ�:���:��	;�P;QM#;�m-;��5;S�;;�@@;�OC;jFE;!uF;!G;��G;�G;F�G;wH;7DH;�bH;d|H;��H;ӢH;��H;ۻH;��H;��H;B�H;i�H;e�H;]�H;��H;��H;��H;]�H;e�H;i�H;B�H;��H;��H;ۻH;��H;ӢH;��H;d|H;�bH;7DH;wH;F�G;�G;��G;!G;!uF;jFE;�OC;�@@;S�;;��5;�m-;QM#;�P;��	;���:Ӵ�:�%�:��:W�:�n�:      ���:�$ ;�;��;��;{P;�l;�c';v�.;�<5;E�:;�>;1B;YAD;��E;��F;+6G;��G;��G;F�G;�H;AH;/_H;lxH;��H;<�H;m�H;��H;b�H;��H;��H;F�H;��H;S�H;�H;��H;Z�H;��H;�H;S�H;��H;F�H;��H;��H;b�H;��H;m�H;<�H;��H;lxH;/_H;AH;�H;F�G;��G;��G;+6G;��F;��E;YAD;1B;�>;E�:;�<5;v�.;�c';�l;{P;��;��;�;�$ ;      �";�L#;�%;��';��+;��/;@�3;��7;P�;;x?;N�A;��C;C9E;�?F;9�F;�TG;��G;S�G;��G;wH;AH;�]H;hvH;9�H;��H;��H;��H;D�H;�H;7�H;1�H;��H;��H;��H;w�H;U�H;��H;U�H;w�H;��H;��H;��H;1�H;7�H;�H;D�H;��H;��H;��H;9�H;hvH;�]H;AH;wH;��G;S�G;��G;�TG;9�F;�?F;C9E;��C;N�A;x?;P�;;��7;@�3;��/;��+;��';�%;�L#;      �36;˃6;kk7;��8;��:;��<;��>;��@;�sB;��C;�+E;F;.�F;�+G;�wG;Y�G;��G;�H;%H;7DH;/_H;hvH;N�H;P�H;h�H;��H;��H;��H;��H;�H;=�H;Q�H;��H;m�H;��H;{�H;��H;{�H;��H;m�H;��H;Q�H;=�H;�H;��H;��H;��H;��H;h�H;P�H;N�H;hvH;/_H;7DH;%H;�H;��G;Y�G;�wG;�+G;.�F;F;�+E;��C;�sB;��@;��>;��<;��:;��8;kk7;˃6;      �@;�@@;f�@;]QA;"B;F
C;�C;��D;[�E;�?F;��F;� G;9gG;ÛG;`�G;�G;�H; .H;-JH;�bH;lxH;9�H;P�H;ۨH;#�H;��H;��H;��H;!�H;[�H;��H;[�H;K�H;��H;��H;i�H;��H;i�H;��H;��H;K�H;[�H;��H;[�H;!�H;��H;��H;��H;#�H;ۨH;P�H;9�H;lxH;�bH;-JH; .H;�H;�G;`�G;ÛG;9gG;� G;��F;�?F;[�E;��D;�C;F
C;"B;]QA;f�@;�@@;      ��D;B�D;A�D;�8E;��E;e�E;�OF;.�F;��F;J9G;lnG;ݙG;�G;��G;� H;�H;�9H;�RH;�hH;d|H;��H;��H;h�H;#�H;U�H;��H;@�H;}�H;��H;9�H;��H;�H;��H;��H;��H;-�H;q�H;-�H;��H;��H;��H;�H;��H;9�H;��H;}�H;@�H;��H;U�H;#�H;h�H;��H;��H;d|H;�hH;�RH;�9H;�H;� H;��G;�G;ݙG;lnG;J9G;��F;.�F;�OF;e�E;��E;�8E;A�D;B�D;      �F;�F;4�F;��F;,�F;� G;�EG;aiG;l�G;,�G;,�G;�G;<�G;�H;�0H;�GH;9]H;�pH;�H;��H;<�H;��H;��H;��H;��H;�H;/�H;k�H;��H;��H;��H;��H;��H;��H;��H;��H;�H;��H;��H;��H;��H;��H;��H;��H;��H;k�H;/�H;�H;��H;��H;��H;��H;<�H;��H;�H;�pH;9]H;�GH;�0H;�H;<�G;�G;,�G;,�G;l�G;aiG;�EG;� G;,�F;��F;4�F;�F;      �mG;<pG;wG;�G;��G;^�G;{�G;��G;'�G;M�G;�H;oH;�/H;�CH;@WH;9iH;�yH;�H;��H;ӢH;m�H;��H;��H;��H;@�H;/�H;N�H;��H;h�H;��H;X�H;��H;��H;��H;;�H;��H;��H;��H;;�H;��H;��H;��H;X�H;��H;h�H;��H;N�H;/�H;@�H;��H;��H;��H;m�H;ӢH;��H;�H;�yH;9iH;@WH;�CH;�/H;oH;�H;M�G;'�G;��G;{�G;^�G;��G;�G;wG;<pG;      %�G;��G;��G;%�G;�G;5�G;"�G;�H;H;c&H;�6H;�GH;�WH;GgH;)vH;�H;�H;ԜH;T�H;��H;��H;D�H;��H;��H;}�H;k�H;��H;G�H;��H;K�H;��H;��H;��H;j�H;��H;
�H; �H;
�H;��H;j�H;��H;��H;��H;K�H;��H;G�H;��H;k�H;}�H;��H;��H;D�H;��H;��H;T�H;ԜH;�H;�H;)vH;GgH;�WH;�GH;�6H;c&H;H;�H;"�G;5�G;�G;%�G;��G;��G;      >H;TH;uH;�H;mH;�$H;�.H;�9H;�EH;�QH;j^H;�jH;SwH;W�H;ԎH;��H;��H;��H;��H;ۻH;b�H;�H;��H;!�H;��H;��H;h�H;��H;,�H;��H;��H;��H;b�H;��H;L�H;�H;��H;�H;L�H;��H;b�H;��H;��H;��H;,�H;��H;h�H;��H;��H;!�H;��H;�H;b�H;ۻH;��H;��H;��H;��H;ԎH;W�H;SwH;�jH;j^H;�QH;�EH;�9H;�.H;�$H;mH;�H;uH;TH;      9?H;@H;cBH;-FH;[KH;�QH;'YH;faH;JjH;�sH;/}H;ʆH;G�H;y�H;8�H;f�H;�H;׸H;�H;��H;��H;7�H;�H;[�H;9�H;��H;��H;K�H;��H;��H;��H;m�H;�H;T�H;��H;��H;��H;��H;��H;T�H;�H;m�H;��H;��H;��H;K�H;��H;��H;9�H;[�H;�H;7�H;��H;��H;�H;׸H;�H;f�H;8�H;y�H;G�H;ʆH;/}H;�sH;JjH;faH;'YH;�QH;[KH;-FH;cBH;@H;      fH;�fH;YhH;?kH;'oH;�sH;�yH;�H;��H;ۍH;�H;r�H;��H;��H;#�H;T�H;'�H;��H;x�H;��H;��H;1�H;=�H;��H;��H;��H;X�H;��H;��H;��H;t�H;�H;h�H;��H;��H;�H;0�H;�H;��H;��H;h�H;�H;t�H;��H;��H;��H;X�H;��H;��H;��H;=�H;1�H;��H;��H;x�H;��H;'�H;T�H;#�H;��H;��H;r�H;�H;ۍH;��H;�H;�yH;�sH;'oH;?kH;YhH;�fH;      w�H;�H;B�H;u�H;j�H;$�H;p�H;/�H;H�H;��H;&�H;��H;#�H;�H;��H;f�H;��H;��H;��H;B�H;F�H;��H;Q�H;[�H;�H;��H;��H;��H;��H;m�H;�H;y�H;��H; �H;,�H;J�H;I�H;J�H;,�H; �H;��H;y�H;�H;m�H;��H;��H;��H;��H;�H;[�H;Q�H;��H;F�H;B�H;��H;��H;��H;f�H;��H;�H;#�H;��H;&�H;��H;H�H;/�H;p�H;$�H;j�H;u�H;B�H;�H;      P�H;��H;��H;Z�H;��H;f�H;��H;O�H;.�H;H�H;��H;̸H;�H;=�H;4�H;��H;u�H;��H;��H;i�H;��H;��H;��H;K�H;��H;��H;��H;��H;b�H;�H;h�H;��H;	�H;9�H;X�H;�H;��H;�H;X�H;9�H;	�H;��H;h�H;�H;b�H;��H;��H;��H;��H;K�H;��H;��H;��H;i�H;��H;��H;u�H;��H;4�H;=�H;�H;̸H;��H;H�H;.�H;O�H;��H;f�H;��H;Z�H;��H;��H;      ��H;�H;ƩH;�H;ŬH;��H;��H;g�H;��H;кH;/�H;��H;��H;:�H;^�H;[�H;6�H;��H;H�H;e�H;S�H;��H;m�H;��H;��H;��H;��H;j�H;��H;T�H;��H; �H;9�H;u�H;��H;��H;��H;��H;��H;u�H;9�H; �H;��H;T�H;��H;j�H;��H;��H;��H;��H;m�H;��H;S�H;e�H;H�H;��H;6�H;[�H;^�H;:�H;��H;��H;/�H;кH;��H;g�H;��H;��H;ŬH;�H;ƩH;�H;      ��H;=�H;�H;�H;_�H;*�H;E�H;��H;0�H;��H;��H;l�H;2�H;��H;��H;'�H;��H;��H;��H;]�H;�H;w�H;��H;��H;��H;��H;;�H;��H;L�H;��H;��H;,�H;X�H;��H;��H;��H;��H;��H;��H;��H;X�H;,�H;��H;��H;L�H;��H;;�H;��H;��H;��H;��H;w�H;�H;]�H;��H;��H;��H;'�H;��H;��H;2�H;l�H;��H;��H;0�H;��H;E�H;*�H;_�H;�H;�H;=�H;      �H;�H;��H;��H;��H;{�H;J�H;Y�H;��H;��H;Y�H;��H;I�H;��H;�H;5�H;B�H;0�H;��H;��H;��H;U�H;{�H;i�H;-�H;��H;��H;
�H;�H;��H;�H;J�H;�H;��H;��H;��H;��H;��H;��H;��H;�H;J�H;�H;��H;�H;
�H;��H;��H;-�H;i�H;{�H;U�H;��H;��H;��H;0�H;B�H;5�H;�H;��H;I�H;��H;Y�H;��H;��H;Y�H;J�H;{�H;��H;��H;��H;�H;      �H;��H;��H;t�H;��H;&�H;��H;��H;�H;a�H;��H;��H;S�H;��H;��H;��H;��H;��H;h�H;��H;Z�H;��H;��H;��H;q�H;�H;��H; �H;��H;��H;0�H;I�H;��H;��H;��H;��H;��H;��H;��H;��H;��H;I�H;0�H;��H;��H; �H;��H;�H;q�H;��H;��H;��H;Z�H;��H;h�H;��H;��H;��H;��H;��H;S�H;��H;��H;a�H;�H;��H;��H;&�H;��H;t�H;��H;��H;      �H;�H;��H;��H;��H;{�H;J�H;Y�H;��H;��H;Y�H;��H;I�H;��H;�H;5�H;B�H;0�H;��H;��H;��H;U�H;{�H;i�H;-�H;��H;��H;
�H;�H;��H;�H;J�H;�H;��H;��H;��H;��H;��H;��H;��H;�H;J�H;�H;��H;�H;
�H;��H;��H;-�H;i�H;{�H;U�H;��H;��H;��H;0�H;B�H;5�H;�H;��H;I�H;��H;Y�H;��H;��H;Y�H;J�H;{�H;��H;��H;��H;�H;      ��H;=�H;�H;�H;_�H;*�H;E�H;��H;0�H;��H;��H;l�H;2�H;��H;��H;'�H;��H;��H;��H;]�H;�H;w�H;��H;��H;��H;��H;;�H;��H;L�H;��H;��H;,�H;X�H;��H;��H;��H;��H;��H;��H;��H;X�H;,�H;��H;��H;L�H;��H;;�H;��H;��H;��H;��H;w�H;�H;]�H;��H;��H;��H;'�H;��H;��H;2�H;l�H;��H;��H;0�H;��H;E�H;*�H;_�H;�H;�H;=�H;      ��H;�H;ƩH;�H;ŬH;��H;��H;g�H;��H;кH;/�H;��H;��H;:�H;^�H;[�H;6�H;��H;H�H;e�H;S�H;��H;m�H;��H;��H;��H;��H;j�H;��H;T�H;��H; �H;9�H;u�H;��H;��H;��H;��H;��H;u�H;9�H; �H;��H;T�H;��H;j�H;��H;��H;��H;��H;m�H;��H;S�H;e�H;H�H;��H;6�H;[�H;^�H;:�H;��H;��H;/�H;кH;��H;g�H;��H;��H;ŬH;�H;ƩH;�H;      P�H;��H;��H;Z�H;��H;f�H;��H;O�H;.�H;H�H;��H;̸H;�H;=�H;4�H;��H;u�H;��H;��H;i�H;��H;��H;��H;K�H;��H;��H;��H;��H;b�H;�H;h�H;��H;	�H;9�H;X�H;�H;��H;�H;X�H;9�H;	�H;��H;h�H;�H;b�H;��H;��H;��H;��H;K�H;��H;��H;��H;i�H;��H;��H;u�H;��H;4�H;=�H;�H;̸H;��H;H�H;.�H;O�H;��H;f�H;��H;Z�H;��H;��H;      w�H;�H;B�H;u�H;j�H;$�H;p�H;/�H;H�H;��H;&�H;��H;#�H;�H;��H;f�H;��H;��H;��H;B�H;F�H;��H;Q�H;[�H;�H;��H;��H;��H;��H;m�H;�H;y�H;��H; �H;,�H;J�H;I�H;J�H;,�H; �H;��H;y�H;�H;m�H;��H;��H;��H;��H;�H;[�H;Q�H;��H;F�H;B�H;��H;��H;��H;f�H;��H;�H;#�H;��H;&�H;��H;H�H;/�H;p�H;$�H;j�H;u�H;B�H;�H;      fH;�fH;YhH;?kH;'oH;�sH;�yH;�H;��H;ۍH;�H;r�H;��H;��H;#�H;T�H;'�H;��H;x�H;��H;��H;1�H;=�H;��H;��H;��H;X�H;��H;��H;��H;t�H;�H;h�H;��H;��H;�H;0�H;�H;��H;��H;h�H;�H;t�H;��H;��H;��H;X�H;��H;��H;��H;=�H;1�H;��H;��H;x�H;��H;'�H;T�H;#�H;��H;��H;r�H;�H;ۍH;��H;�H;�yH;�sH;'oH;?kH;YhH;�fH;      9?H;@H;cBH;-FH;[KH;�QH;'YH;faH;JjH;�sH;/}H;ʆH;G�H;y�H;8�H;f�H;�H;׸H;�H;��H;��H;7�H;�H;[�H;9�H;��H;��H;K�H;��H;��H;��H;m�H;�H;T�H;��H;��H;��H;��H;��H;T�H;�H;m�H;��H;��H;��H;K�H;��H;��H;9�H;[�H;�H;7�H;��H;��H;�H;׸H;�H;f�H;8�H;y�H;G�H;ʆH;/}H;�sH;JjH;faH;'YH;�QH;[KH;-FH;cBH;@H;      >H;TH;uH;�H;mH;�$H;�.H;�9H;�EH;�QH;j^H;�jH;SwH;W�H;ԎH;��H;��H;��H;��H;ۻH;b�H;�H;��H;!�H;��H;��H;h�H;��H;,�H;��H;��H;��H;b�H;��H;L�H;�H;��H;�H;L�H;��H;b�H;��H;��H;��H;,�H;��H;h�H;��H;��H;!�H;��H;�H;b�H;ۻH;��H;��H;��H;��H;ԎH;W�H;SwH;�jH;j^H;�QH;�EH;�9H;�.H;�$H;mH;�H;uH;TH;      %�G;��G;��G;%�G;�G;5�G;"�G;�H;H;c&H;�6H;�GH;�WH;GgH;)vH;�H;�H;ԜH;T�H;��H;��H;D�H;��H;��H;}�H;k�H;��H;G�H;��H;K�H;��H;��H;��H;j�H;��H;
�H; �H;
�H;��H;j�H;��H;��H;��H;K�H;��H;G�H;��H;k�H;}�H;��H;��H;D�H;��H;��H;T�H;ԜH;�H;�H;)vH;GgH;�WH;�GH;�6H;c&H;H;�H;"�G;5�G;�G;%�G;��G;��G;      �mG;<pG;wG;�G;��G;^�G;{�G;��G;'�G;M�G;�H;oH;�/H;�CH;@WH;9iH;�yH;�H;��H;ӢH;m�H;��H;��H;��H;@�H;/�H;N�H;��H;h�H;��H;X�H;��H;��H;��H;;�H;��H;��H;��H;;�H;��H;��H;��H;X�H;��H;h�H;��H;N�H;/�H;@�H;��H;��H;��H;m�H;ӢH;��H;�H;�yH;9iH;@WH;�CH;�/H;oH;�H;M�G;'�G;��G;{�G;^�G;��G;�G;wG;<pG;      �F;�F;4�F;��F;,�F;� G;�EG;aiG;l�G;,�G;,�G;�G;<�G;�H;�0H;�GH;9]H;�pH;�H;��H;<�H;��H;��H;��H;��H;�H;/�H;k�H;��H;��H;��H;��H;��H;��H;��H;��H;�H;��H;��H;��H;��H;��H;��H;��H;��H;k�H;/�H;�H;��H;��H;��H;��H;<�H;��H;�H;�pH;9]H;�GH;�0H;�H;<�G;�G;,�G;,�G;l�G;aiG;�EG;� G;,�F;��F;4�F;�F;      ��D;B�D;A�D;�8E;��E;e�E;�OF;.�F;��F;J9G;lnG;ݙG;�G;��G;� H;�H;�9H;�RH;�hH;d|H;��H;��H;h�H;#�H;U�H;��H;@�H;}�H;��H;9�H;��H;�H;��H;��H;��H;-�H;q�H;-�H;��H;��H;��H;�H;��H;9�H;��H;}�H;@�H;��H;U�H;#�H;h�H;��H;��H;d|H;�hH;�RH;�9H;�H;� H;��G;�G;ݙG;lnG;J9G;��F;.�F;�OF;e�E;��E;�8E;A�D;B�D;      �@;�@@;f�@;]QA;"B;F
C;�C;��D;[�E;�?F;��F;� G;9gG;ÛG;`�G;�G;�H; .H;-JH;�bH;lxH;9�H;P�H;ۨH;#�H;��H;��H;��H;!�H;[�H;��H;[�H;K�H;��H;��H;i�H;��H;i�H;��H;��H;K�H;[�H;��H;[�H;!�H;��H;��H;��H;#�H;ۨH;P�H;9�H;lxH;�bH;-JH; .H;�H;�G;`�G;ÛG;9gG;� G;��F;�?F;[�E;��D;�C;F
C;"B;]QA;f�@;�@@;      �36;˃6;kk7;��8;��:;��<;��>;��@;�sB;��C;�+E;F;.�F;�+G;�wG;Y�G;��G;�H;%H;7DH;/_H;hvH;N�H;P�H;h�H;��H;��H;��H;��H;�H;=�H;Q�H;��H;m�H;��H;{�H;��H;{�H;��H;m�H;��H;Q�H;=�H;�H;��H;��H;��H;��H;h�H;P�H;N�H;hvH;/_H;7DH;%H;�H;��G;Y�G;�wG;�+G;.�F;F;�+E;��C;�sB;��@;��>;��<;��:;��8;kk7;˃6;      �";�L#;�%;��';��+;��/;@�3;��7;P�;;x?;N�A;��C;C9E;�?F;9�F;�TG;��G;S�G;��G;wH;AH;�]H;hvH;9�H;��H;��H;��H;D�H;�H;7�H;1�H;��H;��H;��H;w�H;U�H;��H;U�H;w�H;��H;��H;��H;1�H;7�H;�H;D�H;��H;��H;��H;9�H;hvH;�]H;AH;wH;��G;S�G;��G;�TG;9�F;�?F;C9E;��C;N�A;x?;P�;;��7;@�3;��/;��+;��';�%;�L#;      ���:�$ ;�;��;��;{P;�l;�c';v�.;�<5;E�:;�>;1B;YAD;��E;��F;+6G;��G;��G;F�G;�H;AH;/_H;lxH;��H;<�H;m�H;��H;b�H;��H;��H;F�H;��H;S�H;�H;��H;Z�H;��H;�H;S�H;��H;F�H;��H;��H;b�H;��H;m�H;<�H;��H;lxH;/_H;AH;�H;F�G;��G;��G;+6G;��F;��E;YAD;1B;�>;E�:;�<5;v�.;�c';�l;{P;��;��;�;�$ ;      Y�:�n�:W�:��:�%�:Ӵ�:���:��	;�P;QM#;�m-;��5;S�;;�@@;�OC;jFE;!uF;!G;��G;�G;F�G;wH;7DH;�bH;d|H;��H;ӢH;��H;ۻH;��H;��H;B�H;i�H;e�H;]�H;��H;��H;��H;]�H;e�H;i�H;B�H;��H;��H;ۻH;��H;ӢH;��H;d|H;�bH;7DH;wH;F�G;�G;��G;!G;!uF;jFE;�OC;�@@;S�;;��5;�m-;QM#;�P;��	;���:Ӵ�:�%�:��:W�:�n�:      �	�����j��*_���2u9�:�i~:���:[�:z�;�;�%;`t0;�8;װ>;Z�B;��D;�WF;sG;��G;��G;��G;%H;-JH;�hH;�H;��H;T�H;��H;�H;x�H;��H;��H;H�H;��H;��H;h�H;��H;��H;H�H;��H;��H;x�H;�H;��H;T�H;��H;�H;�hH;-JH;%H;��G;��G;��G;sG;�WF;��D;Z�B;װ>;�8;`t0;�%;�;z�;[�:���:�i~:�:�2u9*_���j�����      _A?���9��8)��Z��ܺlp������?994�@:�:~�:��	;�X;�,;8�6;֜=;x"B;�D;�WF;!G;��G;S�G;�H; .H;�RH;�pH;�H;ԜH;��H;׸H;��H;��H;��H;��H;��H;0�H;��H;0�H;��H;��H;��H;��H;��H;׸H;��H;ԜH;�H;�pH;�RH; .H;�H;S�G;��G;!G;�WF;�D;x"B;֜=;8�6;�,;�X;��	;~�:�:4�@:?99����lp���ܺ�Z��8)���9�      �Eֻ�ѻn�Ļ4T��`�r.o���.�ܺ��B�&��8�\:�%�:���:�P;]);�<5;K:=;x"B;��D;!uF;+6G;��G;��G;�H;�9H;9]H;�yH;�H;��H;�H;'�H;��H;u�H;6�H;��H;B�H;��H;B�H;��H;6�H;u�H;��H;'�H;�H;��H;�H;�yH;9]H;�9H;�H;��G;��G;+6G;!uF;��D;x"B;K:=;�<5;]);�P;���:�%�:�\:&��8��B�ܺ��.�r.o�`�4T��n�Ļ�ѻ      FB��>�s�4�$�$�G���Z�ۚ��oݎ�,A?�EӺ����g2�90q�:�W�:�;D�';�<5;֜=;Z�B;jFE;��F;�TG;Y�G;�G;�H;�GH;9iH;�H;��H;f�H;T�H;f�H;��H;[�H;'�H;5�H;��H;5�H;'�H;[�H;��H;f�H;T�H;f�H;��H;�H;9iH;�GH;�H;�G;Y�G;�TG;��F;jFE;Z�B;֜=;�<5;D�';�;�W�:0q�:g2�9����EӺ,A?�oݎ�ۚ���Z�G��$�$�s�4��>�      <y��ݜ��A���I����s�m�P��%+����Q�Ļ����|��o��8u9�W�:8+�:�;]);8�6;װ>;�OC;��E;9�F;�wG;`�G;� H;�0H;@WH;)vH;ԎH;8�H;#�H;��H;4�H;^�H;��H;�H;��H;�H;��H;^�H;4�H;��H;#�H;8�H;ԎH;)vH;@WH;�0H;� H;`�G;�wG;9�F;��E;�OC;װ>;8�6;]);�;8+�:�W�:�8u9�o�|�����Q�Ļ����%+�m�P���s��I���A��ݜ�      -������bW缑�ռ�վ��Τ��I��Z�[��(��Z�h�9��{���99�W�:�W�:�P;�,;�8;�@@;YAD;�?F;�+G;ÛG;��G;�H;�CH;GgH;W�H;y�H;��H;�H;=�H;:�H;��H;��H;��H;��H;��H;:�H;=�H;�H;��H;y�H;W�H;GgH;�CH;�H;��G;ÛG;�+G;�?F;YAD;�@@;�8;�,;�P;�W�:�W�:�99�{��h�9���Z��(�Z�[��I���Τ��վ���ռbW缧��      �6��3�X�+�ݟ�<�(�����μ߈��T���FB�=s�	T����D��{���8u90q�:���:�X;`t0;S�;;1B;C9E;.�F;9gG;�G;<�G;�/H;�WH;SwH;G�H;��H;#�H;�H;��H;2�H;I�H;S�H;I�H;2�H;��H;�H;#�H;��H;G�H;SwH;�WH;�/H;<�G;�G;9gG;.�F;C9E;1B;S�;;`t0;�X;���:0q�:�8u9�{����D�	T��=s�FB�T���߈����μ(���<�ݟ�X�+��3�      R₽�؀���u��Xc�Q�K�K1�{�����վ�t]��b�P�m��	T��h�9��o�g2�9�%�:��	;�%;��5;�>;��C;F;� G;ݙG;�G;oH;�GH;�jH;ʆH;r�H;��H;̸H;��H;l�H;��H;��H;��H;l�H;��H;̸H;��H;r�H;ʆH;�jH;�GH;oH;�G;ݙG;� G;F;��C;�>;��5;�%;��	;�%�:g2�9�o�h�9�	T��m��b�P�t]���վ����{��K1�Q�K��Xc���u��؀�      S���r��L��n������|�u�e�N���(�ji���˼�A��b�P�=s��|������\:~�:�;�m-;E�:;N�A;�+E;��F;lnG;,�G;�H;�6H;j^H;/}H;�H;&�H;��H;/�H;��H;Y�H;��H;Y�H;��H;/�H;��H;&�H;�H;/}H;j^H;�6H;�H;,�G;lnG;��F;�+E;N�A;E�:;�m-;�;~�:�\:����|��=s�b�P��A����˼ji���(�e�N�|�u�����n��L���r��      �o���r���}�ս@��Kĥ�X^���Xc��3���	���˼t]��FB��Z򻆜��EӺ&��8�:z�;QM#;�<5;x?;��C;�?F;J9G;,�G;M�G;c&H;�QH;�sH;ۍH;��H;H�H;кH;��H;��H;a�H;��H;��H;кH;H�H;��H;ۍH;�sH;�QH;c&H;M�G;,�G;J9G;�?F;��C;x?;�<5;QM#;z�;�:&��8EӺ�����Z�FB�t]����˼��	��3��Xc�X^��Kĥ�@��}�ս���r�      �#�6� �A'����~���gٽS��l���j��3�ji��վ�T����(�Q�Ļ,A?���B�4�@:[�:�P;v�.;P�;;�sB;[�E;��F;l�G;'�G;H;�EH;JjH;��H;H�H;.�H;��H;0�H;��H;�H;��H;0�H;��H;.�H;H�H;��H;JjH;�EH;H;'�G;l�G;��F;[�E;�sB;P�;;v�.;�P;[�:4�@:��B�,A?�Q�Ļ�(�T����վ�ji��3��j�l��S���gٽ�~����A'�6� �      �S� �O��E��5�6� �<�
���|9��l���Xc���(����߈��Z�[����oݎ�ܺ?99���:��	;�c';��7;��@;��D;.�F;aiG;��G;�H;�9H;faH;�H;/�H;O�H;g�H;��H;Y�H;��H;Y�H;��H;g�H;O�H;/�H;�H;faH;�9H;�H;��G;aiG;.�F;��D;��@;��7;�c';��	;���:?99ܺoݎ����Z�[�߈�������(��Xc�l��|9����<�
�6� ��5��E� �O�      �~���)����v��9b�U�H��",�0Z���S��X^��e�N�{����μ�I���%+�ۚ����.������i~:���:�l;@�3;��>;�C;�OF;�EG;{�G;"�G;�.H;'YH;�yH;p�H;��H;��H;E�H;J�H;��H;J�H;E�H;��H;��H;p�H;�yH;'YH;�.H;"�G;{�G;�EG;�OF;�C;��>;@�3;�l;���:�i~:������.�ۚ���%+��I����μ{��e�N�X^��S����0Z��",�U�H��9b���v��)��      ��������:���M���r� �O��",�<�
��gٽKĥ�|�u�K1�(����Τ�m�P��Z�r.o�lp���:Ӵ�:{P;��/;��<;F
C;e�E;� G;^�G;5�G;�$H;�QH;�sH;$�H;f�H;��H;*�H;{�H;&�H;{�H;*�H;��H;f�H;$�H;�sH;�QH;�$H;5�G;^�G;� G;e�E;F
C;��<;��/;{P;Ӵ�:�:lp��r.o��Z�m�P��Τ�(���K1�|�u�Kĥ��gٽ<�
��",� �O��r��M���:�����      ���v��/;������:P���r�U�H�6� ��~��@������Q�K�<��վ���s�G��`񕻀ܺ�2u9�%�:��;��+;��:;"B;��E;,�F;��G;�G;mH;[KH;'oH;j�H;��H;ŬH;_�H;��H;��H;��H;_�H;ŬH;��H;j�H;'oH;[KH;mH;�G;��G;,�F;��E;"B;��:;��+;��;�%�:�2u9�ܺ`�G����s��վ�<�Q�K�����@���~��6� �U�H��r�:P������/;���v��      3Vھ�*־5ʾT��������M���9b��5���}�սn���Xc�ݟ���ռ�I��$�$�4T���Z�*_����:��;��';��8;]QA;�8E;��F;�G;%�G;�H;-FH;?kH;u�H;Z�H;�H;�H;��H;t�H;��H;�H;�H;Z�H;u�H;?kH;-FH;�H;%�G;�G;��F;�8E;]QA;��8;��';��;��:*_���Z�4T��$�$��I����ռݟ��Xc�n��}�ս���5��9b��M������T���5ʾ�*־      ǰ�쾐�޾5ʾ/;���:����v��E�A'���L����u�X�+�bW缨A��s�4�n�Ļ�8)��j��W�:�;�%;kk7;f�@;A�D;4�F;wG;��G;uH;cBH;YhH;B�H;��H;ƩH;�H;��H;��H;��H;�H;ƩH;��H;B�H;YhH;cBH;uH;��G;wG;4�F;A�D;f�@;kk7;�%;�;W�:�j���8)�n�Ļs�4��A��bW�X�+���u�L����A'��E���v��:��/;��5ʾ��޾��      /h���b���쾅*־�v������)�� �O�6� ��r�r���؀��3����ݜ��>��ѻ��9�����n�:�$ ;�L#;˃6;�@@;B�D;�F;<pG;��G;TH;@H;�fH;�H;��H;�H;=�H;�H;��H;�H;=�H;�H;��H;�H;�fH;@H;TH;��G;<pG;�F;B�D;�@@;˃6;�L#;�$ ;�n�:�����9��ѻ�>�ݜ�����3��؀��r���r�6� � �O��)������v���*־�쾼b��      ����]�0_ݾ��ɾK*��Ы���zx��G�0,�U�뽘b�� @{�|�/�\���䙼�J;��ͻ��4�-WṺ��:�;]�#;��6;UZ@;��D;��F;�kG;��G;{H;�9H;�aH;�H;M�H;U�H;�H;�H;��H;�H;�H;U�H;M�H;�H;�aH;�9H;{H;��G;�kG;��F;��D;UZ@;��6;]�#;�;���:-WṬ�4��ͻ�J;��䙼\��|�/� @{��b��U��0,��G��zx�Ы��K*����ɾ0_ݾ�]�      �]����:پZ�žI�������8t�I�C�����罽���`w�-�l���_����7��Rɻ�K/�yƹb��:O/;f$;)7;~@;��D;��F;nG;-�G;gH;�:H;�bH;��H;��H;��H;5�H;L�H;B�H;L�H;5�H;��H;��H;��H;�bH;�:H;gH;-�G;nG;��F;��D;~@;)7;f$;O/;b��:yƹ�K/��Rɻ��7��_��l��-�`w����������I�C��8t����I���Z�ž�:پ��      0_ݾ�:پ�V;�*���Ƥ�3a����g�g$:��Z�?ݽkƣ�Al�:.%��߼=��n9.�����#V� 2p��@�:�w;�'&;��7;~�@;O
E;F�F;�tG;Z�G;�
H;=H;|dH;��H;��H;s�H;ձH;ݷH;عH;ݷH;ձH;s�H;��H;��H;|dH;=H;�
H;Z�G;�tG;F�F;O
E;~�@;��7;�'&;�w;�@�: 2p�#V�����n9.�=���߼:.%�Al�kƣ�?ݽ�Z�g$:���g�3a���Ƥ��*���V;�:پ      ��ɾZ�ž�*��Sת�Ы��	�����T��J+��a2̽ss���yZ����μ>y�����!Ϩ�,,����6���:��
;��(;�M9;C�A;�ME;��F;�~G;�G;�H;�@H;agH;�H;`�H;��H;��H;ǸH;��H;ǸH;��H;��H;`�H;�H;agH;�@H;�H;�G;�~G;��F;�ME;C�A;�M9;��(;��
;���:���6,,�!Ϩ����>y��μ����yZ�ss��a2̽��J+���T�	���Ы��Sת��*��Z�ž      K*��I����Ƥ�Ы���/���c��G=����z�gж��ɇ� �C�����!��);k�{&�}-��G�˺LX�9	��:�8;hh,;8	;;?PB;��E; G;�G;�G;�H;2FH;|kH;/�H;��H;��H;d�H;&�H;��H;&�H;d�H;��H;��H;/�H;|kH;2FH;�H;�G;�G; G;��E;?PB;8	;;hh,;�8;	��:LX�9G�˺}-��{&�);k��!����� �C��ɇ�gж��z����G=��c��/��Ы���Ƥ�I���      Ы�����3a��	����c�J�C�Z#���$vϽ����Al�8g*�T��v
���I�X��q\c��쀺0t,:g��:u�;D_0;��<;�0C;2�E;�"G;}�G;B�G;GH;�LH;epH;׊H;��H;�H;T�H;��H;��H;��H;T�H;�H;��H;׊H;epH;�LH;GH;B�G;}�G;�"G;2�E;�0C;��<;D_0;u�;g��:0t,:�쀺q\c�X�軞I�v
��T��8g*�Al�����$vϽ��Z#�J�C��c�	���3a�����      �zx��8t���g���T��G=�Z#��5�?ݽ�b������G������Ǽ?y���$�'����$�%vƹ棆:6&�:2� ;�~4;��>;�D;[F;�EG;��G;:�G;7)H;�TH;%vH;%�H;
�H;��H;��H;��H;M�H;��H;��H;��H;
�H;%�H;%vH;�TH;7)H;:�G;��G;�EG;[F;�D;��>;�~4;2� ;6&�:棆:%vƹ�$�'����$�?y����Ǽ���G������b��?ݽ�5�Z#��G=���T���g��8t�      �G�I�C�g$:��J+�����?ݽ4���I���yZ�Ơ"�k�鼣���T�Y� ��L��j�˺�m9�ض:�;�_(;}8;��@;��D;'�F;�gG;��G;� H;e4H; ]H;�|H;�H;ۥH;y�H;�H;ɿH;X�H;ɿH;�H;y�H;ۥH;�H;�|H; ]H;e4H;� H;��G;�gG;'�F;��D;��@;}8;�_(;�;�ض:�m9j�˺�L��Y� �T�����k��Ơ"��yZ�I��4���?ݽ�����J+�g$:�I�C�      0,����Z���z�$vϽ�b��I��.]a�-�D� ��!��)�{��!�g���i�4��P(�<nQ:L�:��;H�/;:'<;A�B;=�E;)�F;φG;��G;hH;o@H;=fH;y�H;\�H;�H;��H;��H;�H;u�H;�H;��H;��H;�H;\�H;y�H;=fH;o@H;hH;��G;φG;)�F;=�E;A�B;:'<;H�/;��;L�:<nQ:�P(�i�4�g����!�)�{��!��D� �-�.]a�I���b��$vϽ�z���Z���      U�뽱��?ݽa2̽gж����������yZ�-�����`ļ-O���J;�6��&�|�_�ºAM@9;��:��;Tf$;��5;)N?;�D;�KF;?:G;ߣG;#�G;� H;MH;�oH;��H;��H;K�H;�H;f�H;��H;��H;��H;f�H;�H;K�H;��H;��H;�oH;MH;� H;#�G;ߣG;?:G;�KF;�D;)N?;��5;Tf$;��;;��:AM@9_�º&�|�6�軃J;�-O���`ļ���-��yZ���������gж�a2̽?ݽ���      �b������kƣ�ss���ɇ�Al�G�Ơ"�D� ��`ļ6���I��C��ۙ��Vuƹ��k:��:��;�=.;|	;;*�A;-AE;��F;NlG;��G;��G;�1H;ZH;�yH;�H;��H;��H;{�H;O�H;�H;3�H;�H;O�H;{�H;��H;��H;�H;�yH;ZH;�1H;��G;��G;NlG;��F;-AE;*�A;|	;;�=.;��;��:��k:Vuƹ��ۙ��C��I�6���`ļD� �Ơ"�G�Al��ɇ�ss��kƣ�����       @{�`w�Al��yZ� �C�8g*����k���!��-O���I�|��Ψ�3K/�b$T��P:���:3�;6(&;]#6;%?;��C;�"F;9#G;^�G;��G;�H;XBH;gH;��H;��H;��H;�H;�H;?�H;��H;��H;��H;?�H;�H;�H;��H;��H;��H;gH;XBH;�H;��G;^�G;9#G;�"F;��C;%?;]#6;6(&;3�;���:�P:b$T�3K/��Ψ�|��I�-O���!��k�鼇��8g*� �C��yZ�Al�`w�      |�/�-�:.%�������T���Ǽ����)�{��J;��C��Ψ�
O:�����vZ�9L��:;�;�-1;k'<;$5B;%NE;Z�F;jeG;�G;h�G;"*H;
SH;�sH;F�H;�H;@�H;i�H;��H;�H;�H;=�H;�H;�H;��H;i�H;@�H;�H;F�H;�sH;
SH;"*H;h�G;�G;jeG;Z�F;%NE;$5B;k'<;�-1;�;;L��:vZ�9����
O:��Ψ��C��J;�)�{�������ǼT��������:.%�-�      \��l�鼟߼μ�!��v
��?y��T��!�6�軉ۙ�3K/�����hm9pA�:���:Ž;��,;,N9;�~@;^D;
LF;�-G;�G;��G;�H;�>H;CcH;;�H;��H;+�H;��H;��H;��H;��H;��H;��H;��H;��H;��H;��H;��H;+�H;��H;;�H;CcH;�>H;�H;��G;�G;�-G;
LF;^D;�~@;,N9;��,;Ž;���:pA�:hm9����3K/��ۙ�6���!�T�?y��v
���!��μ�߼l��      �䙼�_��=��>y��);k��I��$�Y� �g���&�|��b$T�vZ�9pA�:���:��;��);�7;=�>; tC;_�E;1�F;$uG;O�G;��G;/+H;�RH;�rH;��H;��H;/�H;�H;��H;S�H;��H;�H;��H;�H;��H;S�H;��H;�H;/�H;��H;��H;�rH;�RH;/+H;��G;O�G;$uG;1�F;_�E; tC;=�>;�7;��);��;���:pA�:vZ�9b$T��&�|�g���Y� ��$��I�);k�>y��=���_��      �J;���7�n9.����{&�X��'����L��i�4�_�ºVuƹ�P:L��:���:��;,�(;-�5;#�=;�B;�ZE;��F;TG;ߨG;��G;�H;�BH;9eH;�H;��H;�H;��H;�H;��H;o�H;�H;Q�H;9�H;Q�H;�H;o�H;��H;�H;��H;�H;��H;�H;9eH;�BH;�H;��G;ߨG;TG;��F;�ZE;�B;#�=;-�5;,�(;��;���:L��:�P:Vuƹ_�ºi�4��L��'���X��{&����n9.���7�      �ͻ�Rɻ����!Ϩ�}-��q\c��$�j�˺�P(�AM@9��k:���:;Ž;��);-�5;��=;uPB;�
E;5F;d7G;y�G;{�G;�H;�4H;�XH;gvH;��H;ѠH;�H;��H;��H;l�H;<�H;��H;��H;9�H;��H;��H;<�H;l�H;��H;��H;�H;ѠH;��H;gvH;�XH;�4H;�H;{�G;y�G;d7G;5F;�
E;uPB;��=;-�5;��);Ž;;���:��k:AM@9�P(�j�˺�$�q\c�}-��!Ϩ������Rɻ      ��4��K/�#V�,,�G�˺�쀺%vƹ�m9<nQ:;��:��:3�;�;��,;�7;#�=;uPB;�D;�bF;]#G;�G;�G;�G;�(H;�MH;�lH;��H;�H;E�H;-�H;-�H;��H;��H;��H;��H;��H;'�H;��H;��H;��H;��H;��H;-�H;-�H;E�H;�H;��H;�lH;�MH;�(H;�G;�G;�G;]#G;�bF;�D;uPB;#�=;�7;��,;�;3�;��:;��:<nQ:�m9%vƹ�쀺G�˺,,�#V��K/�      -W�yƹ 2p����6LX�90t,:棆:�ض:L�:��;��;6(&;�-1;,N9;=�>;�B;�
E;�bF;+G;eG;�G;��G;�H;EH;�dH;�~H;ٓH;�H;ҲH;��H;'�H;��H;��H;g�H; �H;Z�H;��H;Z�H; �H;g�H;��H;��H;'�H;��H;ҲH;�H;ٓH;�~H;�dH;EH;�H;��G;�G;eG;+G;�bF;�
E;�B;=�>;,N9;�-1;6(&;��;��;L�:�ض:棆:0t,:LX�9���6 2p�yƹ      ���:b��:�@�:���:	��:g��:6&�:�;��;Tf$;�=.;]#6;k'<;�~@; tC;�ZE;5F;]#G;eG;�G;K�G;�H;?H;�^H;yH;y�H;<�H;ѮH;J�H;��H;��H;d�H;��H;��H;��H;�H;{�H;�H;��H;��H;��H;d�H;��H;��H;J�H;ѮH;<�H;y�H;yH;�^H;?H;�H;K�G;�G;eG;]#G;5F;�ZE; tC;�~@;k'<;]#6;�=.;Tf$;��;�;6&�:g��:	��:���:�@�:b��:      �;O/;�w;��
;�8;u�;2� ;�_(;H�/;��5;|	;;%?;$5B;^D;_�E;��F;d7G;�G;�G;K�G;�H;�;H;�ZH;
uH;��H;p�H;U�H;T�H;��H;��H;��H;}�H;�H;��H;��H;��H;��H;��H;��H;��H;�H;}�H;��H;��H;��H;T�H;U�H;p�H;��H;
uH;�ZH;�;H;�H;K�G;�G;�G;d7G;��F;_�E;^D;$5B;%?;|	;;��5;H�/;�_(;2� ;u�;�8;��
;�w;O/;      ]�#;f$;�'&;��(;hh,;D_0;�~4;}8;:'<;)N?;*�A;��C;%NE;
LF;1�F;TG;y�G;�G;��G;�H;�;H;�YH;sH;�H;��H;��H;�H;�H;��H;)�H;Q�H;F�H;e�H;��H;��H;��H;%�H;��H;��H;��H;e�H;F�H;Q�H;)�H;��H;�H;�H;��H;��H;�H;sH;�YH;�;H;�H;��G;�G;y�G;TG;1�F;
LF;%NE;��C;*�A;)N?;:'<;}8;�~4;D_0;hh,;��(;�'&;f$;      ��6;)7;��7;�M9;8	;;��<;��>;��@;A�B;�D;-AE;�"F;Z�F;�-G;$uG;ߨG;{�G;�G;�H;?H;�ZH;sH;V�H;r�H;�H;?�H;�H;;�H;�H;4�H;d�H;��H;U�H;>�H;G�H;�H;@�H;�H;G�H;>�H;U�H;��H;d�H;4�H;�H;;�H;�H;?�H;�H;r�H;V�H;sH;�ZH;?H;�H;�G;{�G;ߨG;$uG;�-G;Z�F;�"F;-AE;�D;A�B;��@;��>;��<;8	;;�M9;��7;)7;      UZ@;~@;~�@;C�A;?PB;�0C;�D;��D;=�E;�KF;��F;9#G;jeG;�G;O�G;��G;�H;�(H;EH;�^H;
uH;�H;r�H;|�H;W�H;/�H;@�H;��H;c�H;��H;�H;��H;��H;x�H;t�H;
�H;Q�H;
�H;t�H;x�H;��H;��H;�H;��H;c�H;��H;@�H;/�H;W�H;|�H;r�H;�H;
uH;�^H;EH;�(H;�H;��G;O�G;�G;jeG;9#G;��F;�KF;=�E;��D;�D;�0C;?PB;C�A;~�@;~@;      ��D;��D;O
E;�ME;��E;2�E;[F;'�F;)�F;?:G;NlG;^�G;�G;��G;��G;�H;�4H;�MH;�dH;yH;��H;��H;�H;W�H;��H;��H;=�H;��H;�H;��H;c�H;��H;b�H;��H;��H;��H;�H;��H;��H;��H;b�H;��H;c�H;��H;�H;��H;=�H;��H;��H;W�H;�H;��H;��H;yH;�dH;�MH;�4H;�H;��G;��G;�G;^�G;NlG;?:G;)�F;'�F;[F;2�E;��E;�ME;O
E;��D;      ��F;��F;F�F;��F; G;�"G;�EG;�gG;φG;ߣG;��G;��G;h�G;�H;/+H;�BH;�XH;�lH;�~H;y�H;p�H;��H;?�H;/�H;��H;�H;G�H;��H;#�H;)�H;k�H;�H;��H;��H;e�H;��H;��H;��H;e�H;��H;��H;�H;k�H;)�H;#�H;��H;G�H;�H;��H;/�H;?�H;��H;p�H;y�H;�~H;�lH;�XH;�BH;/+H;�H;h�G;��G;��G;ߣG;φG;�gG;�EG;�"G; G;��F;F�F;��F;      �kG;nG;�tG;�~G;�G;}�G;��G;��G;��G;#�G;��G;�H;"*H;�>H;�RH;9eH;gvH;��H;ٓH;<�H;U�H;�H;�H;@�H;=�H;G�H;e�H;��H;��H;5�H;*�H;t�H;��H;x�H;�H;d�H;��H;d�H;�H;x�H;��H;t�H;*�H;5�H;��H;��H;e�H;G�H;=�H;@�H;�H;�H;U�H;<�H;ٓH;��H;gvH;9eH;�RH;�>H;"*H;�H;��G;#�G;��G;��G;��G;}�G;�G;�~G;�tG;nG;      ��G;-�G;Z�G;�G;�G;B�G;:�G;� H;hH;� H;�1H;XBH;
SH;CcH;�rH;�H;��H;�H;�H;ѮH;T�H;�H;;�H;��H;��H;��H;��H;��H;�H;��H;q�H;��H;��H;B�H;��H;��H;#�H;��H;��H;B�H;��H;��H;q�H;��H;�H;��H;��H;��H;��H;��H;;�H;�H;T�H;ѮH;�H;�H;��H;�H;�rH;CcH;
SH;XBH;�1H;� H;hH;� H;:�G;B�G;�G;�G;Z�G;-�G;      {H;gH;�
H;�H;�H;GH;7)H;e4H;o@H;MH;ZH;gH;�sH;;�H;��H;��H;ѠH;E�H;ҲH;J�H;��H;��H;�H;c�H;�H;#�H;��H;�H;��H;V�H;�H;��H;@�H;��H;�H;V�H;b�H;V�H;�H;��H;@�H;��H;�H;V�H;��H;�H;��H;#�H;�H;c�H;�H;��H;��H;J�H;ҲH;E�H;ѠH;��H;��H;;�H;�sH;gH;ZH;MH;o@H;e4H;7)H;GH;�H;�H;�
H;gH;      �9H;�:H;=H;�@H;2FH;�LH;�TH; ]H;=fH;�oH;�yH;��H;F�H;��H;��H;�H;�H;-�H;��H;��H;��H;)�H;4�H;��H;��H;)�H;5�H;��H;V�H;��H;w�H;1�H;��H;8�H;��H;��H;��H;��H;��H;8�H;��H;1�H;w�H;��H;V�H;��H;5�H;)�H;��H;��H;4�H;)�H;��H;��H;��H;-�H;�H;�H;��H;��H;F�H;��H;�yH;�oH;=fH; ]H;�TH;�LH;2FH;�@H;=H;�:H;      �aH;�bH;|dH;agH;|kH;epH;%vH;�|H;y�H;��H;�H;��H;�H;+�H;/�H;��H;��H;-�H;'�H;��H;��H;Q�H;d�H;�H;c�H;k�H;*�H;q�H;�H;w�H;H�H;��H;2�H;��H;��H;��H;�H;��H;��H;��H;2�H;��H;H�H;w�H;�H;q�H;*�H;k�H;c�H;�H;d�H;Q�H;��H;��H;'�H;-�H;��H;��H;/�H;+�H;�H;��H;�H;��H;y�H;�|H;%vH;epH;|kH;agH;|dH;�bH;      �H;��H;��H;�H;/�H;׊H;%�H;�H;\�H;��H;��H;��H;@�H;��H;�H;�H;��H;��H;��H;d�H;}�H;F�H;��H;��H;��H;�H;t�H;��H;��H;1�H;��H;B�H;��H;��H;�H;C�H;5�H;C�H;�H;��H;��H;B�H;��H;1�H;��H;��H;t�H;�H;��H;��H;��H;F�H;}�H;d�H;��H;��H;��H;�H;�H;��H;@�H;��H;��H;��H;\�H;�H;%�H;׊H;/�H;�H;��H;��H;      M�H;��H;��H;`�H;��H;��H;
�H;ۥH;�H;K�H;��H;�H;i�H;��H;��H;��H;l�H;��H;��H;��H;�H;e�H;U�H;��H;b�H;��H;��H;��H;@�H;��H;2�H;��H;�H;�H;V�H;l�H;6�H;l�H;V�H;�H;�H;��H;2�H;��H;@�H;��H;��H;��H;b�H;��H;U�H;e�H;�H;��H;��H;��H;l�H;��H;��H;��H;i�H;�H;��H;K�H;�H;ۥH;
�H;��H;��H;`�H;��H;��H;      U�H;��H;s�H;��H;��H;�H;��H;y�H;��H;�H;{�H;�H;��H;��H;S�H;o�H;<�H;��H;g�H;��H;��H;��H;>�H;x�H;��H;��H;x�H;B�H;��H;8�H;��H;��H;�H;M�H;m�H;y�H;��H;y�H;m�H;M�H;�H;��H;��H;8�H;��H;B�H;x�H;��H;��H;x�H;>�H;��H;��H;��H;g�H;��H;<�H;o�H;S�H;��H;��H;�H;{�H;�H;��H;y�H;��H;�H;��H;��H;s�H;��H;      �H;5�H;ձH;��H;d�H;T�H;��H;�H;��H;f�H;O�H;?�H;�H;��H;��H;�H;��H;��H; �H;��H;��H;��H;G�H;t�H;��H;e�H;�H;��H;�H;��H;��H;�H;V�H;m�H;u�H;��H;��H;��H;u�H;m�H;V�H;�H;��H;��H;�H;��H;�H;e�H;��H;t�H;G�H;��H;��H;��H; �H;��H;��H;�H;��H;��H;�H;?�H;O�H;f�H;��H;�H;��H;T�H;d�H;��H;ձH;5�H;      �H;L�H;ݷH;ǸH;&�H;��H;��H;ɿH;�H;��H;�H;��H;�H;��H;�H;Q�H;��H;��H;Z�H;�H;��H;��H;�H;
�H;��H;��H;d�H;��H;V�H;��H;��H;C�H;l�H;y�H;��H;��H;��H;��H;��H;y�H;l�H;C�H;��H;��H;V�H;��H;d�H;��H;��H;
�H;�H;��H;��H;�H;Z�H;��H;��H;Q�H;�H;��H;�H;��H;�H;��H;�H;ɿH;��H;��H;&�H;ǸH;ݷH;L�H;      ��H;B�H;عH;��H;��H;��H;M�H;X�H;u�H;��H;3�H;��H;=�H;��H;��H;9�H;9�H;'�H;��H;{�H;��H;%�H;@�H;Q�H;�H;��H;��H;#�H;b�H;��H;�H;5�H;6�H;��H;��H;��H;��H;��H;��H;��H;6�H;5�H;�H;��H;b�H;#�H;��H;��H;�H;Q�H;@�H;%�H;��H;{�H;��H;'�H;9�H;9�H;��H;��H;=�H;��H;3�H;��H;u�H;X�H;M�H;��H;��H;��H;عH;B�H;      �H;L�H;ݷH;ǸH;&�H;��H;��H;ɿH;�H;��H;�H;��H;�H;��H;�H;Q�H;��H;��H;Z�H;�H;��H;��H;�H;
�H;��H;��H;d�H;��H;V�H;��H;��H;C�H;l�H;y�H;��H;��H;��H;��H;��H;y�H;l�H;C�H;��H;��H;V�H;��H;d�H;��H;��H;
�H;�H;��H;��H;�H;Z�H;��H;��H;Q�H;�H;��H;�H;��H;�H;��H;�H;ɿH;��H;��H;&�H;ǸH;ݷH;L�H;      �H;5�H;ձH;��H;d�H;T�H;��H;�H;��H;f�H;O�H;?�H;�H;��H;��H;�H;��H;��H; �H;��H;��H;��H;G�H;t�H;��H;e�H;�H;��H;�H;��H;��H;�H;V�H;m�H;u�H;��H;��H;��H;u�H;m�H;V�H;�H;��H;��H;�H;��H;�H;e�H;��H;t�H;G�H;��H;��H;��H; �H;��H;��H;�H;��H;��H;�H;?�H;O�H;f�H;��H;�H;��H;T�H;d�H;��H;ձH;5�H;      U�H;��H;s�H;��H;��H;�H;��H;y�H;��H;�H;{�H;�H;��H;��H;S�H;o�H;<�H;��H;g�H;��H;��H;��H;>�H;x�H;��H;��H;x�H;B�H;��H;8�H;��H;��H;�H;M�H;m�H;y�H;��H;y�H;m�H;M�H;�H;��H;��H;8�H;��H;B�H;x�H;��H;��H;x�H;>�H;��H;��H;��H;g�H;��H;<�H;o�H;S�H;��H;��H;�H;{�H;�H;��H;y�H;��H;�H;��H;��H;s�H;��H;      M�H;��H;��H;`�H;��H;��H;
�H;ۥH;�H;K�H;��H;�H;i�H;��H;��H;��H;l�H;��H;��H;��H;�H;e�H;U�H;��H;b�H;��H;��H;��H;@�H;��H;2�H;��H;�H;�H;V�H;l�H;6�H;l�H;V�H;�H;�H;��H;2�H;��H;@�H;��H;��H;��H;b�H;��H;U�H;e�H;�H;��H;��H;��H;l�H;��H;��H;��H;i�H;�H;��H;K�H;�H;ۥH;
�H;��H;��H;`�H;��H;��H;      �H;��H;��H;�H;/�H;׊H;%�H;�H;\�H;��H;��H;��H;@�H;��H;�H;�H;��H;��H;��H;d�H;}�H;F�H;��H;��H;��H;�H;t�H;��H;��H;1�H;��H;B�H;��H;��H;�H;C�H;5�H;C�H;�H;��H;��H;B�H;��H;1�H;��H;��H;t�H;�H;��H;��H;��H;F�H;}�H;d�H;��H;��H;��H;�H;�H;��H;@�H;��H;��H;��H;\�H;�H;%�H;׊H;/�H;�H;��H;��H;      �aH;�bH;|dH;agH;|kH;epH;%vH;�|H;y�H;��H;�H;��H;�H;+�H;/�H;��H;��H;-�H;'�H;��H;��H;Q�H;d�H;�H;c�H;k�H;*�H;q�H;�H;w�H;H�H;��H;2�H;��H;��H;��H;�H;��H;��H;��H;2�H;��H;H�H;w�H;�H;q�H;*�H;k�H;c�H;�H;d�H;Q�H;��H;��H;'�H;-�H;��H;��H;/�H;+�H;�H;��H;�H;��H;y�H;�|H;%vH;epH;|kH;agH;|dH;�bH;      �9H;�:H;=H;�@H;2FH;�LH;�TH; ]H;=fH;�oH;�yH;��H;F�H;��H;��H;�H;�H;-�H;��H;��H;��H;)�H;4�H;��H;��H;)�H;5�H;��H;V�H;��H;w�H;1�H;��H;8�H;��H;��H;��H;��H;��H;8�H;��H;1�H;w�H;��H;V�H;��H;5�H;)�H;��H;��H;4�H;)�H;��H;��H;��H;-�H;�H;�H;��H;��H;F�H;��H;�yH;�oH;=fH; ]H;�TH;�LH;2FH;�@H;=H;�:H;      {H;gH;�
H;�H;�H;GH;7)H;e4H;o@H;MH;ZH;gH;�sH;;�H;��H;��H;ѠH;E�H;ҲH;J�H;��H;��H;�H;c�H;�H;#�H;��H;�H;��H;V�H;�H;��H;@�H;��H;�H;V�H;b�H;V�H;�H;��H;@�H;��H;�H;V�H;��H;�H;��H;#�H;�H;c�H;�H;��H;��H;J�H;ҲH;E�H;ѠH;��H;��H;;�H;�sH;gH;ZH;MH;o@H;e4H;7)H;GH;�H;�H;�
H;gH;      ��G;-�G;Z�G;�G;�G;B�G;:�G;� H;hH;� H;�1H;XBH;
SH;CcH;�rH;�H;��H;�H;�H;ѮH;T�H;�H;;�H;��H;��H;��H;��H;��H;�H;��H;q�H;��H;��H;B�H;��H;��H;#�H;��H;��H;B�H;��H;��H;q�H;��H;�H;��H;��H;��H;��H;��H;;�H;�H;T�H;ѮH;�H;�H;��H;�H;�rH;CcH;
SH;XBH;�1H;� H;hH;� H;:�G;B�G;�G;�G;Z�G;-�G;      �kG;nG;�tG;�~G;�G;}�G;��G;��G;��G;#�G;��G;�H;"*H;�>H;�RH;9eH;gvH;��H;ٓH;<�H;U�H;�H;�H;@�H;=�H;G�H;e�H;��H;��H;5�H;*�H;t�H;��H;x�H;�H;d�H;��H;d�H;�H;x�H;��H;t�H;*�H;5�H;��H;��H;e�H;G�H;=�H;@�H;�H;�H;U�H;<�H;ٓH;��H;gvH;9eH;�RH;�>H;"*H;�H;��G;#�G;��G;��G;��G;}�G;�G;�~G;�tG;nG;      ��F;��F;F�F;��F; G;�"G;�EG;�gG;φG;ߣG;��G;��G;h�G;�H;/+H;�BH;�XH;�lH;�~H;y�H;p�H;��H;?�H;/�H;��H;�H;G�H;��H;#�H;)�H;k�H;�H;��H;��H;e�H;��H;��H;��H;e�H;��H;��H;�H;k�H;)�H;#�H;��H;G�H;�H;��H;/�H;?�H;��H;p�H;y�H;�~H;�lH;�XH;�BH;/+H;�H;h�G;��G;��G;ߣG;φG;�gG;�EG;�"G; G;��F;F�F;��F;      ��D;��D;O
E;�ME;��E;2�E;[F;'�F;)�F;?:G;NlG;^�G;�G;��G;��G;�H;�4H;�MH;�dH;yH;��H;��H;�H;W�H;��H;��H;=�H;��H;�H;��H;c�H;��H;b�H;��H;��H;��H;�H;��H;��H;��H;b�H;��H;c�H;��H;�H;��H;=�H;��H;��H;W�H;�H;��H;��H;yH;�dH;�MH;�4H;�H;��G;��G;�G;^�G;NlG;?:G;)�F;'�F;[F;2�E;��E;�ME;O
E;��D;      UZ@;~@;~�@;C�A;?PB;�0C;�D;��D;=�E;�KF;��F;9#G;jeG;�G;O�G;��G;�H;�(H;EH;�^H;
uH;�H;r�H;|�H;W�H;/�H;@�H;��H;c�H;��H;�H;��H;��H;x�H;t�H;
�H;Q�H;
�H;t�H;x�H;��H;��H;�H;��H;c�H;��H;@�H;/�H;W�H;|�H;r�H;�H;
uH;�^H;EH;�(H;�H;��G;O�G;�G;jeG;9#G;��F;�KF;=�E;��D;�D;�0C;?PB;C�A;~�@;~@;      ��6;)7;��7;�M9;8	;;��<;��>;��@;A�B;�D;-AE;�"F;Z�F;�-G;$uG;ߨG;{�G;�G;�H;?H;�ZH;sH;V�H;r�H;�H;?�H;�H;;�H;�H;4�H;d�H;��H;U�H;>�H;G�H;�H;@�H;�H;G�H;>�H;U�H;��H;d�H;4�H;�H;;�H;�H;?�H;�H;r�H;V�H;sH;�ZH;?H;�H;�G;{�G;ߨG;$uG;�-G;Z�F;�"F;-AE;�D;A�B;��@;��>;��<;8	;;�M9;��7;)7;      ]�#;f$;�'&;��(;hh,;D_0;�~4;}8;:'<;)N?;*�A;��C;%NE;
LF;1�F;TG;y�G;�G;��G;�H;�;H;�YH;sH;�H;��H;��H;�H;�H;��H;)�H;Q�H;F�H;e�H;��H;��H;��H;%�H;��H;��H;��H;e�H;F�H;Q�H;)�H;��H;�H;�H;��H;��H;�H;sH;�YH;�;H;�H;��G;�G;y�G;TG;1�F;
LF;%NE;��C;*�A;)N?;:'<;}8;�~4;D_0;hh,;��(;�'&;f$;      �;O/;�w;��
;�8;u�;2� ;�_(;H�/;��5;|	;;%?;$5B;^D;_�E;��F;d7G;�G;�G;K�G;�H;�;H;�ZH;
uH;��H;p�H;U�H;T�H;��H;��H;��H;}�H;�H;��H;��H;��H;��H;��H;��H;��H;�H;}�H;��H;��H;��H;T�H;U�H;p�H;��H;
uH;�ZH;�;H;�H;K�G;�G;�G;d7G;��F;_�E;^D;$5B;%?;|	;;��5;H�/;�_(;2� ;u�;�8;��
;�w;O/;      ���:b��:�@�:���:	��:g��:6&�:�;��;Tf$;�=.;]#6;k'<;�~@; tC;�ZE;5F;]#G;eG;�G;K�G;�H;?H;�^H;yH;y�H;<�H;ѮH;J�H;��H;��H;d�H;��H;��H;��H;�H;{�H;�H;��H;��H;��H;d�H;��H;��H;J�H;ѮH;<�H;y�H;yH;�^H;?H;�H;K�G;�G;eG;]#G;5F;�ZE; tC;�~@;k'<;]#6;�=.;Tf$;��;�;6&�:g��:	��:���:�@�:b��:      -W�yƹ 2p����6LX�90t,:棆:�ض:L�:��;��;6(&;�-1;,N9;=�>;�B;�
E;�bF;+G;eG;�G;��G;�H;EH;�dH;�~H;ٓH;�H;ҲH;��H;'�H;��H;��H;g�H; �H;Z�H;��H;Z�H; �H;g�H;��H;��H;'�H;��H;ҲH;�H;ٓH;�~H;�dH;EH;�H;��G;�G;eG;+G;�bF;�
E;�B;=�>;,N9;�-1;6(&;��;��;L�:�ض:棆:0t,:LX�9���6 2p�yƹ      ��4��K/�#V�,,�G�˺�쀺%vƹ�m9<nQ:;��:��:3�;�;��,;�7;#�=;uPB;�D;�bF;]#G;�G;�G;�G;�(H;�MH;�lH;��H;�H;E�H;-�H;-�H;��H;��H;��H;��H;��H;'�H;��H;��H;��H;��H;��H;-�H;-�H;E�H;�H;��H;�lH;�MH;�(H;�G;�G;�G;]#G;�bF;�D;uPB;#�=;�7;��,;�;3�;��:;��:<nQ:�m9%vƹ�쀺G�˺,,�#V��K/�      �ͻ�Rɻ����!Ϩ�}-��q\c��$�j�˺�P(�AM@9��k:���:;Ž;��);-�5;��=;uPB;�
E;5F;d7G;y�G;{�G;�H;�4H;�XH;gvH;��H;ѠH;�H;��H;��H;l�H;<�H;��H;��H;9�H;��H;��H;<�H;l�H;��H;��H;�H;ѠH;��H;gvH;�XH;�4H;�H;{�G;y�G;d7G;5F;�
E;uPB;��=;-�5;��);Ž;;���:��k:AM@9�P(�j�˺�$�q\c�}-��!Ϩ������Rɻ      �J;���7�n9.����{&�X��'����L��i�4�_�ºVuƹ�P:L��:���:��;,�(;-�5;#�=;�B;�ZE;��F;TG;ߨG;��G;�H;�BH;9eH;�H;��H;�H;��H;�H;��H;o�H;�H;Q�H;9�H;Q�H;�H;o�H;��H;�H;��H;�H;��H;�H;9eH;�BH;�H;��G;ߨG;TG;��F;�ZE;�B;#�=;-�5;,�(;��;���:L��:�P:Vuƹ_�ºi�4��L��'���X��{&����n9.���7�      �䙼�_��=��>y��);k��I��$�Y� �g���&�|��b$T�vZ�9pA�:���:��;��);�7;=�>; tC;_�E;1�F;$uG;O�G;��G;/+H;�RH;�rH;��H;��H;/�H;�H;��H;S�H;��H;�H;��H;�H;��H;S�H;��H;�H;/�H;��H;��H;�rH;�RH;/+H;��G;O�G;$uG;1�F;_�E; tC;=�>;�7;��);��;���:pA�:vZ�9b$T��&�|�g���Y� ��$��I�);k�>y��=���_��      \��l�鼟߼μ�!��v
��?y��T��!�6�軉ۙ�3K/�����hm9pA�:���:Ž;��,;,N9;�~@;^D;
LF;�-G;�G;��G;�H;�>H;CcH;;�H;��H;+�H;��H;��H;��H;��H;��H;��H;��H;��H;��H;��H;��H;+�H;��H;;�H;CcH;�>H;�H;��G;�G;�-G;
LF;^D;�~@;,N9;��,;Ž;���:pA�:hm9����3K/��ۙ�6���!�T�?y��v
���!��μ�߼l��      |�/�-�:.%�������T���Ǽ����)�{��J;��C��Ψ�
O:�����vZ�9L��:;�;�-1;k'<;$5B;%NE;Z�F;jeG;�G;h�G;"*H;
SH;�sH;F�H;�H;@�H;i�H;��H;�H;�H;=�H;�H;�H;��H;i�H;@�H;�H;F�H;�sH;
SH;"*H;h�G;�G;jeG;Z�F;%NE;$5B;k'<;�-1;�;;L��:vZ�9����
O:��Ψ��C��J;�)�{�������ǼT��������:.%�-�       @{�`w�Al��yZ� �C�8g*����k���!��-O���I�|��Ψ�3K/�b$T��P:���:3�;6(&;]#6;%?;��C;�"F;9#G;^�G;��G;�H;XBH;gH;��H;��H;��H;�H;�H;?�H;��H;��H;��H;?�H;�H;�H;��H;��H;��H;gH;XBH;�H;��G;^�G;9#G;�"F;��C;%?;]#6;6(&;3�;���:�P:b$T�3K/��Ψ�|��I�-O���!��k�鼇��8g*� �C��yZ�Al�`w�      �b������kƣ�ss���ɇ�Al�G�Ơ"�D� ��`ļ6���I��C��ۙ��Vuƹ��k:��:��;�=.;|	;;*�A;-AE;��F;NlG;��G;��G;�1H;ZH;�yH;�H;��H;��H;{�H;O�H;�H;3�H;�H;O�H;{�H;��H;��H;�H;�yH;ZH;�1H;��G;��G;NlG;��F;-AE;*�A;|	;;�=.;��;��:��k:Vuƹ��ۙ��C��I�6���`ļD� �Ơ"�G�Al��ɇ�ss��kƣ�����      U�뽱��?ݽa2̽gж����������yZ�-�����`ļ-O���J;�6��&�|�_�ºAM@9;��:��;Tf$;��5;)N?;�D;�KF;?:G;ߣG;#�G;� H;MH;�oH;��H;��H;K�H;�H;f�H;��H;��H;��H;f�H;�H;K�H;��H;��H;�oH;MH;� H;#�G;ߣG;?:G;�KF;�D;)N?;��5;Tf$;��;;��:AM@9_�º&�|�6�軃J;�-O���`ļ���-��yZ���������gж�a2̽?ݽ���      0,����Z���z�$vϽ�b��I��.]a�-�D� ��!��)�{��!�g���i�4��P(�<nQ:L�:��;H�/;:'<;A�B;=�E;)�F;φG;��G;hH;o@H;=fH;y�H;\�H;�H;��H;��H;�H;u�H;�H;��H;��H;�H;\�H;y�H;=fH;o@H;hH;��G;φG;)�F;=�E;A�B;:'<;H�/;��;L�:<nQ:�P(�i�4�g����!�)�{��!��D� �-�.]a�I���b��$vϽ�z���Z���      �G�I�C�g$:��J+�����?ݽ4���I���yZ�Ơ"�k�鼣���T�Y� ��L��j�˺�m9�ض:�;�_(;}8;��@;��D;'�F;�gG;��G;� H;e4H; ]H;�|H;�H;ۥH;y�H;�H;ɿH;X�H;ɿH;�H;y�H;ۥH;�H;�|H; ]H;e4H;� H;��G;�gG;'�F;��D;��@;}8;�_(;�;�ض:�m9j�˺�L��Y� �T�����k��Ơ"��yZ�I��4���?ݽ�����J+�g$:�I�C�      �zx��8t���g���T��G=�Z#��5�?ݽ�b������G������Ǽ?y���$�'����$�%vƹ棆:6&�:2� ;�~4;��>;�D;[F;�EG;��G;:�G;7)H;�TH;%vH;%�H;
�H;��H;��H;��H;M�H;��H;��H;��H;
�H;%�H;%vH;�TH;7)H;:�G;��G;�EG;[F;�D;��>;�~4;2� ;6&�:棆:%vƹ�$�'����$�?y����Ǽ���G������b��?ݽ�5�Z#��G=���T���g��8t�      Ы�����3a��	����c�J�C�Z#���$vϽ����Al�8g*�T��v
���I�X��q\c��쀺0t,:g��:u�;D_0;��<;�0C;2�E;�"G;}�G;B�G;GH;�LH;epH;׊H;��H;�H;T�H;��H;��H;��H;T�H;�H;��H;׊H;epH;�LH;GH;B�G;}�G;�"G;2�E;�0C;��<;D_0;u�;g��:0t,:�쀺q\c�X�軞I�v
��T��8g*�Al�����$vϽ��Z#�J�C��c�	���3a�����      K*��I����Ƥ�Ы���/���c��G=����z�gж��ɇ� �C�����!��);k�{&�}-��G�˺LX�9	��:�8;hh,;8	;;?PB;��E; G;�G;�G;�H;2FH;|kH;/�H;��H;��H;d�H;&�H;��H;&�H;d�H;��H;��H;/�H;|kH;2FH;�H;�G;�G; G;��E;?PB;8	;;hh,;�8;	��:LX�9G�˺}-��{&�);k��!����� �C��ɇ�gж��z����G=��c��/��Ы���Ƥ�I���      ��ɾZ�ž�*��Sת�Ы��	�����T��J+��a2̽ss���yZ����μ>y�����!Ϩ�,,����6���:��
;��(;�M9;C�A;�ME;��F;�~G;�G;�H;�@H;agH;�H;`�H;��H;��H;ǸH;��H;ǸH;��H;��H;`�H;�H;agH;�@H;�H;�G;�~G;��F;�ME;C�A;�M9;��(;��
;���:���6,,�!Ϩ����>y��μ����yZ�ss��a2̽��J+���T�	���Ы��Sת��*��Z�ž      0_ݾ�:پ�V;�*���Ƥ�3a����g�g$:��Z�?ݽkƣ�Al�:.%��߼=��n9.�����#V� 2p��@�:�w;�'&;��7;~�@;O
E;F�F;�tG;Z�G;�
H;=H;|dH;��H;��H;s�H;ձH;ݷH;عH;ݷH;ձH;s�H;��H;��H;|dH;=H;�
H;Z�G;�tG;F�F;O
E;~�@;��7;�'&;�w;�@�: 2p�#V�����n9.�=���߼:.%�Al�kƣ�?ݽ�Z�g$:���g�3a���Ƥ��*���V;�:پ      �]����:پZ�žI�������8t�I�C�����罽���`w�-�l���_����7��Rɻ�K/�yƹb��:O/;f$;)7;~@;��D;��F;nG;-�G;gH;�:H;�bH;��H;��H;��H;5�H;L�H;B�H;L�H;5�H;��H;��H;��H;�bH;�:H;gH;-�G;nG;��F;��D;~@;)7;f$;O/;b��:yƹ�K/��Rɻ��7��_��l��-�`w����������I�C��8t����I���Z�ž�:پ��      3F�/h��ǰ�3Vھ�������~���S��#��o��S��R₽�6�-���<y��FB��Eֻ_A?��	�Y�:���:�";�36;�@;��D;�F;�mG;%�G;>H;9?H;fH;w�H;P�H;��H;��H;�H;�H;�H;��H;��H;P�H;w�H;fH;9?H;>H;%�G;�mG;�F;��D;�@;�36;�";���:Y�:�	�_A?��EֻFB�<y��-����6�R₽S���o���#��S��~��������3Vھǰ�/h��      /h���b���쾅*־�v������)�� �O�6� ��r�r���؀��3����ݜ��>��ѻ��9�����n�:�$ ;�L#;˃6;�@@;B�D;�F;<pG;��G;TH;@H;�fH;�H;��H;�H;=�H;�H;��H;�H;=�H;�H;��H;�H;�fH;@H;TH;��G;<pG;�F;B�D;�@@;˃6;�L#;�$ ;�n�:�����9��ѻ�>�ݜ�����3��؀��r���r�6� � �O��)������v���*־�쾼b��      ǰ�쾐�޾5ʾ/;���:����v��E�A'���L����u�X�+�bW缨A��s�4�n�Ļ�8)��j��W�:�;�%;kk7;f�@;A�D;4�F;wG;��G;uH;cBH;YhH;B�H;��H;ƩH;�H;��H;��H;��H;�H;ƩH;��H;B�H;YhH;cBH;uH;��G;wG;4�F;A�D;f�@;kk7;�%;�;W�:�j���8)�n�Ļs�4��A��bW�X�+���u�L����A'��E���v��:��/;��5ʾ��޾��      3Vھ�*־5ʾT��������M���9b��5���}�սn���Xc�ݟ���ռ�I��$�$�4T���Z�(_����:��;��';��8;]QA;�8E;��F;�G;%�G;�H;-FH;?kH;u�H;Z�H;�H;�H;��H;t�H;��H;�H;�H;Z�H;u�H;?kH;-FH;�H;%�G;�G;��F;�8E;]QA;��8;��';��;��:(_���Z�4T��$�$��I����ռݟ��Xc�n��}�ս���5��9b��M������T���5ʾ�*־      ���v��/;������:P���r�U�H�6� ��~��@������Q�K�<��վ���s�G��`�ܺ�2u9�%�:��;��+;��:;"B;��E;,�F;��G;�G;mH;[KH;'oH;j�H;��H;ŬH;_�H;��H;��H;��H;_�H;ŬH;��H;j�H;'oH;[KH;mH;�G;��G;,�F;��E;"B;��:;��+;��;�%�:�2u9ܺ`�G����s��վ�<�Q�K�����@���~��6� �U�H��r�:P������/;���v��      ��������:���M���r� �O��",�<�
��gٽKĥ�|�u�K1�(����Τ�m�P��Z�r.o�lp���:Ӵ�:{P;��/;��<;F
C;e�E;� G;^�G;5�G;�$H;�QH;�sH;$�H;f�H;��H;*�H;{�H;&�H;{�H;*�H;��H;f�H;$�H;�sH;�QH;�$H;5�G;^�G;� G;e�E;F
C;��<;��/;{P;Ӵ�:�:lp��r.o��Z�m�P��Τ�(���K1�|�u�Kĥ��gٽ<�
��",� �O��r��M���:�����      �~���)����v��9b�U�H��",�0Z���S��X^��e�N�{����μ�I���%+�ۚ����.������i~:���:�l;@�3;��>;�C;�OF;�EG;{�G;"�G;�.H;'YH;�yH;p�H;��H;��H;E�H;J�H;��H;J�H;E�H;��H;��H;p�H;�yH;'YH;�.H;"�G;{�G;�EG;�OF;�C;��>;@�3;�l;���:�i~:������.�ۚ���%+��I����μ{��e�N�X^��S����0Z��",�U�H��9b���v��)��      �S� �O��E��5�6� �<�
���|9��l���Xc���(����߈��Z�[����oݎ�ܺ@99���:��	;�c';��7;��@;��D;.�F;aiG;��G;�H;�9H;faH;�H;/�H;O�H;g�H;��H;Y�H;��H;Y�H;��H;g�H;O�H;/�H;�H;faH;�9H;�H;��G;aiG;.�F;��D;��@;��7;�c';��	;���:@99ܺoݎ����Z�[�߈�������(��Xc�l��|9����<�
�6� ��5��E� �O�      �#�6� �A'����~���gٽS��l���j��3�ji��վ�T����(�Q�Ļ,A?���B�4�@:[�:�P;v�.;P�;;�sB;[�E;��F;l�G;'�G;H;�EH;JjH;��H;H�H;.�H;��H;0�H;��H;�H;��H;0�H;��H;.�H;H�H;��H;JjH;�EH;H;'�G;l�G;��F;[�E;�sB;P�;;v�.;�P;[�:4�@:��B�,A?�Q�Ļ�(�T����վ�ji��3��j�l��S���gٽ�~����A'�6� �      �o���r���}�ս@��Kĥ�X^���Xc��3���	���˼t]��FB��Z򻆜��EӺ'��8�:z�;RM#;�<5;x?;��C;�?F;J9G;,�G;M�G;c&H;�QH;�sH;ۍH;��H;H�H;кH;��H;��H;a�H;��H;��H;кH;H�H;��H;ۍH;�sH;�QH;c&H;M�G;,�G;J9G;�?F;��C;x?;�<5;RM#;z�;�:'��8EӺ�����Z�FB�t]����˼��	��3��Xc�X^��Kĥ�@��}�ս���r�      S���r��L��n������|�u�e�N���(�ji���˼�A��b�P�=s��|������\:~�:�;�m-;E�:;N�A;�+E;��F;lnG;,�G;�H;�6H;j^H;/}H;�H;&�H;��H;/�H;��H;Y�H;��H;Y�H;��H;/�H;��H;&�H;�H;/}H;j^H;�6H;�H;,�G;lnG;��F;�+E;N�A;E�:;�m-;�;~�:�\:����|��=s�b�P��A����˼ji���(�e�N�|�u�����n��L���r��      R₽�؀���u��Xc�Q�K�K1�{�����վ�t]��b�P�m��	T��h�9��o�g2�9�%�:��	;�%;��5;�>;��C;F;� G;ݙG;�G;oH;�GH;�jH;ʆH;r�H;��H;̸H;��H;l�H;��H;��H;��H;l�H;��H;̸H;��H;r�H;ʆH;�jH;�GH;oH;�G;ݙG;� G;F;��C;�>;��5;�%;��	;�%�:g2�9�o�h�9�	T��m��b�P�t]���վ����{��K1�Q�K��Xc���u��؀�      �6��3�X�+�ݟ�<�(�����μ߈��T���FB�=s�	T����D��{���8u90q�:���:�X;at0;S�;;1B;C9E;.�F;9gG;�G;<�G;�/H;�WH;SwH;G�H;��H;#�H;�H;��H;2�H;I�H;S�H;I�H;2�H;��H;�H;#�H;��H;G�H;SwH;�WH;�/H;<�G;�G;9gG;.�F;C9E;1B;S�;;at0;�X;���:0q�:�8u9�{����D�	T��=s�FB�T���߈����μ(���<�ݟ�X�+��3�      -������bW缑�ռ�վ��Τ��I��Z�[��(��Z�h�9��{���99�W�:�W�:�P;�,;�8;�@@;YAD;�?F;�+G;ÛG;��G;�H;�CH;GgH;W�H;y�H;��H;�H;=�H;:�H;��H;��H;��H;��H;��H;:�H;=�H;�H;��H;y�H;W�H;GgH;�CH;�H;��G;ÛG;�+G;�?F;YAD;�@@;�8;�,;�P;�W�:�W�:�99�{��h�9���Z��(�Z�[��I���Τ��վ���ռbW缧��      <y��ݜ��A���I����s�m�P��%+����Q�Ļ����|��o��8u9�W�:8+�:�;]);8�6;װ>;�OC;��E;9�F;�wG;`�G;� H;�0H;@WH;)vH;ԎH;8�H;#�H;��H;4�H;^�H;��H;�H;��H;�H;��H;^�H;4�H;��H;#�H;8�H;ԎH;)vH;@WH;�0H;� H;`�G;�wG;9�F;��E;�OC;װ>;8�6;]);�;8+�:�W�:�8u9�o�|�����Q�Ļ����%+�m�P���s��I���A��ݜ�      FB��>�s�4�$�$�G���Z�ۚ��oݎ�,A?�EӺ����g2�90q�:�W�:�;D�';�<5;֜=;Z�B;jFE;��F;�TG;Y�G;�G;�H;�GH;9iH;�H;��H;f�H;T�H;f�H;��H;[�H;(�H;5�H;��H;5�H;(�H;[�H;��H;f�H;T�H;f�H;��H;�H;9iH;�GH;�H;�G;Y�G;�TG;��F;jFE;Z�B;֜=;�<5;D�';�;�W�:0q�:g2�9����EӺ,A?�oݎ�ۚ���Z�G��$�$�s�4��>�      �Eֻ�ѻn�Ļ4T��`�r.o���.�ܺ��B�'��8�\:�%�:���:�P;]);�<5;K:=;x"B;��D;!uF;+6G;��G;��G;�H;�9H;9]H;�yH;�H;��H;�H;'�H;��H;u�H;6�H;��H;B�H;��H;B�H;��H;6�H;u�H;��H;'�H;�H;��H;�H;�yH;9]H;�9H;�H;��G;��G;+6G;!uF;��D;x"B;K:=;�<5;]);�P;���:�%�:�\:'��8��B�ܺ��.�r.o�`�4T��n�Ļ�ѻ      _A?���9��8)��Z�ܺlp������@994�@:�:~�:��	;�X;�,;8�6;֜=;x"B; �D;�WF;!G;��G;S�G;�H; .H;�RH;�pH;�H;ԜH;��H;׸H;��H;��H;��H;��H;��H;0�H;��H;0�H;��H;��H;��H;��H;��H;׸H;��H;ԜH;�H;�pH;�RH; .H;�H;S�G;��G;!G;�WF; �D;x"B;֜=;8�6;�,;�X;��	;~�:�:4�@:@99����lp��ܺ�Z��8)���9�      �	�����j��(_���2u9�:�i~:���:[�:z�;�;�%;at0;�8;װ>;Z�B;��D;�WF;sG;��G;��G;��G;%H;-JH;�hH;�H;��H;T�H;��H;�H;x�H;��H;��H;H�H;��H;��H;h�H;��H;��H;H�H;��H;��H;x�H;�H;��H;T�H;��H;�H;�hH;-JH;%H;��G;��G;��G;sG;�WF;��D;Z�B;װ>;�8;at0;�%;�;z�;[�:���:�i~:�:�2u9(_���j�����      Y�:�n�:W�:��:�%�:Ӵ�:���:��	;�P;RM#;�m-;��5;S�;;�@@;�OC;jFE;!uF;!G;��G;�G;F�G;wH;7DH;�bH;d|H;��H;ӢH;��H;ۻH;��H;��H;B�H;i�H;e�H;]�H;��H;��H;��H;]�H;e�H;i�H;B�H;��H;��H;ۻH;��H;ӢH;��H;d|H;�bH;7DH;wH;F�G;�G;��G;!G;!uF;jFE;�OC;�@@;S�;;��5;�m-;RM#;�P;��	;���:Ӵ�:�%�:��:W�:�n�:      ���:�$ ;�;��;��;{P;�l;�c';v�.;�<5;E�:;�>;1B;YAD;��E;��F;+6G;��G;��G;F�G;�H;AH;/_H;lxH;��H;<�H;m�H;��H;b�H;��H;��H;F�H;��H;S�H;�H;��H;Z�H;��H;�H;S�H;��H;F�H;��H;��H;b�H;��H;m�H;<�H;��H;lxH;/_H;AH;�H;F�G;��G;��G;+6G;��F;��E;YAD;1B;�>;E�:;�<5;v�.;�c';�l;{P;��;��;�;�$ ;      �";�L#;�%;��';��+;��/;@�3;��7;P�;;x?;N�A;��C;C9E;�?F;9�F;�TG;��G;S�G;��G;wH;AH;�]H;hvH;9�H;��H;��H;��H;D�H;�H;7�H;1�H;��H;��H;��H;w�H;U�H;��H;U�H;w�H;��H;��H;��H;1�H;7�H;�H;D�H;��H;��H;��H;9�H;hvH;�]H;AH;wH;��G;S�G;��G;�TG;9�F;�?F;C9E;��C;N�A;x?;P�;;��7;@�3;��/;��+;��';�%;�L#;      �36;˃6;kk7;��8;��:;��<;��>;��@;�sB;��C;�+E;F;.�F;�+G;�wG;Y�G;��G;�H;%H;7DH;/_H;hvH;N�H;P�H;h�H;��H;��H;��H;��H;�H;=�H;Q�H;��H;m�H;��H;{�H;��H;{�H;��H;m�H;��H;Q�H;=�H;�H;��H;��H;��H;��H;h�H;P�H;N�H;hvH;/_H;7DH;%H;�H;��G;Y�G;�wG;�+G;.�F;F;�+E;��C;�sB;��@;��>;��<;��:;��8;kk7;˃6;      �@;�@@;f�@;]QA;"B;F
C;�C;��D;[�E;�?F;��F;� G;9gG;ÛG;`�G;�G;�H; .H;-JH;�bH;lxH;9�H;P�H;ۨH;#�H;��H;��H;��H;!�H;[�H;��H;[�H;K�H;��H;��H;i�H;��H;i�H;��H;��H;K�H;[�H;��H;[�H;!�H;��H;��H;��H;#�H;ۨH;P�H;9�H;lxH;�bH;-JH; .H;�H;�G;`�G;ÛG;9gG;� G;��F;�?F;[�E;��D;�C;F
C;"B;]QA;f�@;�@@;      ��D;B�D;A�D;�8E;��E;e�E;�OF;.�F;��F;J9G;lnG;ݙG;�G;��G;� H;�H;�9H;�RH;�hH;d|H;��H;��H;h�H;#�H;U�H;��H;@�H;}�H;��H;9�H;��H;�H;��H;��H;��H;-�H;q�H;-�H;��H;��H;��H;�H;��H;9�H;��H;}�H;@�H;��H;U�H;#�H;h�H;��H;��H;d|H;�hH;�RH;�9H;�H;� H;��G;�G;ݙG;lnG;J9G;��F;.�F;�OF;e�E;��E;�8E;A�D;B�D;      �F;�F;4�F;��F;,�F;� G;�EG;aiG;l�G;,�G;,�G;�G;<�G;�H;�0H;�GH;9]H;�pH;�H;��H;<�H;��H;��H;��H;��H;�H;/�H;k�H;��H;��H;��H;��H;��H;��H;��H;��H;�H;��H;��H;��H;��H;��H;��H;��H;��H;k�H;/�H;�H;��H;��H;��H;��H;<�H;��H;�H;�pH;9]H;�GH;�0H;�H;<�G;�G;,�G;,�G;l�G;aiG;�EG;� G;,�F;��F;4�F;�F;      �mG;<pG;wG;�G;��G;^�G;{�G;��G;'�G;M�G;�H;oH;�/H;�CH;@WH;9iH;�yH;�H;��H;ӢH;m�H;��H;��H;��H;@�H;/�H;N�H;��H;h�H;��H;X�H;��H;��H;��H;;�H;��H;��H;��H;;�H;��H;��H;��H;X�H;��H;h�H;��H;N�H;/�H;@�H;��H;��H;��H;m�H;ӢH;��H;�H;�yH;9iH;@WH;�CH;�/H;oH;�H;M�G;'�G;��G;{�G;^�G;��G;�G;wG;<pG;      %�G;��G;��G;%�G;�G;5�G;"�G;�H;H;c&H;�6H;�GH;�WH;GgH;)vH;�H;�H;ԜH;T�H;��H;��H;D�H;��H;��H;}�H;k�H;��H;G�H;��H;K�H;��H;��H;��H;j�H;��H;�H; �H;�H;��H;j�H;��H;��H;��H;K�H;��H;G�H;��H;k�H;}�H;��H;��H;D�H;��H;��H;T�H;ԜH;�H;�H;)vH;GgH;�WH;�GH;�6H;c&H;H;�H;"�G;5�G;�G;%�G;��G;��G;      >H;TH;uH;�H;mH;�$H;�.H;�9H;�EH;�QH;j^H;�jH;SwH;W�H;ԎH;��H;��H;��H;��H;ۻH;b�H;�H;��H;!�H;��H;��H;h�H;��H;,�H;��H;��H;��H;b�H;��H;L�H;�H;��H;�H;L�H;��H;b�H;��H;��H;��H;,�H;��H;h�H;��H;��H;!�H;��H;�H;b�H;ۻH;��H;��H;��H;��H;ԎH;W�H;SwH;�jH;j^H;�QH;�EH;�9H;�.H;�$H;mH;�H;uH;TH;      9?H;@H;cBH;-FH;[KH;�QH;'YH;faH;JjH;�sH;/}H;ʆH;G�H;y�H;8�H;f�H;�H;׸H;�H;��H;��H;7�H;�H;[�H;9�H;��H;��H;K�H;��H;��H;��H;m�H;�H;T�H;��H;��H;��H;��H;��H;T�H;�H;m�H;��H;��H;��H;K�H;��H;��H;9�H;[�H;�H;7�H;��H;��H;�H;׸H;�H;f�H;8�H;y�H;G�H;ʆH;/}H;�sH;JjH;faH;'YH;�QH;[KH;-FH;cBH;@H;      fH;�fH;YhH;?kH;'oH;�sH;�yH;�H;��H;ۍH;�H;r�H;��H;��H;#�H;T�H;'�H;��H;x�H;��H;��H;1�H;=�H;��H;��H;��H;X�H;��H;��H;��H;t�H;�H;h�H;��H;��H;�H;0�H;�H;��H;��H;h�H;�H;t�H;��H;��H;��H;X�H;��H;��H;��H;=�H;1�H;��H;��H;x�H;��H;'�H;T�H;#�H;��H;��H;r�H;�H;ۍH;��H;�H;�yH;�sH;'oH;?kH;YhH;�fH;      w�H;�H;B�H;u�H;j�H;$�H;p�H;/�H;H�H;��H;&�H;��H;#�H;�H;��H;f�H;��H;��H;��H;B�H;F�H;��H;Q�H;[�H;�H;��H;��H;��H;��H;m�H;�H;y�H;��H; �H;,�H;J�H;I�H;J�H;,�H; �H;��H;y�H;�H;m�H;��H;��H;��H;��H;�H;[�H;Q�H;��H;F�H;B�H;��H;��H;��H;f�H;��H;�H;#�H;��H;&�H;��H;H�H;/�H;p�H;$�H;j�H;u�H;B�H;�H;      P�H;��H;��H;Z�H;��H;f�H;��H;O�H;.�H;H�H;��H;̸H;�H;=�H;4�H;��H;u�H;��H;��H;i�H;��H;��H;��H;K�H;��H;��H;��H;��H;b�H;�H;h�H;��H;	�H;9�H;X�H;�H;��H;�H;X�H;9�H;	�H;��H;h�H;�H;b�H;��H;��H;��H;��H;K�H;��H;��H;��H;i�H;��H;��H;u�H;��H;4�H;=�H;�H;̸H;��H;H�H;.�H;O�H;��H;f�H;��H;Z�H;��H;��H;      ��H;�H;ƩH;�H;ŬH;��H;��H;g�H;��H;кH;/�H;��H;��H;:�H;^�H;[�H;6�H;��H;H�H;e�H;S�H;��H;m�H;��H;��H;��H;��H;j�H;��H;T�H;��H; �H;9�H;u�H;��H;��H;��H;��H;��H;u�H;9�H; �H;��H;T�H;��H;j�H;��H;��H;��H;��H;m�H;��H;S�H;e�H;H�H;��H;6�H;[�H;^�H;:�H;��H;��H;/�H;кH;��H;g�H;��H;��H;ŬH;�H;ƩH;�H;      ��H;=�H;�H;�H;_�H;*�H;E�H;��H;0�H;��H;��H;l�H;2�H;��H;��H;(�H;��H;��H;��H;]�H;�H;w�H;��H;��H;��H;��H;;�H;��H;L�H;��H;��H;,�H;X�H;��H;��H;��H;��H;��H;��H;��H;X�H;,�H;��H;��H;L�H;��H;;�H;��H;��H;��H;��H;w�H;�H;]�H;��H;��H;��H;(�H;��H;��H;2�H;l�H;��H;��H;0�H;��H;E�H;*�H;_�H;�H;�H;=�H;      �H;�H;��H;��H;��H;{�H;J�H;Y�H;��H;��H;Y�H;��H;I�H;��H;�H;5�H;B�H;0�H;��H;��H;��H;U�H;{�H;i�H;-�H;��H;��H;�H;�H;��H;�H;J�H;�H;��H;��H;��H;��H;��H;��H;��H;�H;J�H;�H;��H;�H;�H;��H;��H;-�H;i�H;{�H;U�H;��H;��H;��H;0�H;B�H;5�H;�H;��H;I�H;��H;Y�H;��H;��H;Y�H;J�H;{�H;��H;��H;��H;�H;      �H;��H;��H;t�H;��H;&�H;��H;��H;�H;a�H;��H;��H;S�H;��H;��H;��H;��H;��H;h�H;��H;Z�H;��H;��H;��H;q�H;�H;��H; �H;��H;��H;0�H;I�H;��H;��H;��H;��H;��H;��H;��H;��H;��H;I�H;0�H;��H;��H; �H;��H;�H;q�H;��H;��H;��H;Z�H;��H;h�H;��H;��H;��H;��H;��H;S�H;��H;��H;a�H;�H;��H;��H;&�H;��H;t�H;��H;��H;      �H;�H;��H;��H;��H;{�H;J�H;Y�H;��H;��H;Y�H;��H;I�H;��H;�H;5�H;B�H;0�H;��H;��H;��H;U�H;{�H;i�H;-�H;��H;��H;�H;�H;��H;�H;J�H;�H;��H;��H;��H;��H;��H;��H;��H;�H;J�H;�H;��H;�H;�H;��H;��H;-�H;i�H;{�H;U�H;��H;��H;��H;0�H;B�H;5�H;�H;��H;I�H;��H;Y�H;��H;��H;Y�H;J�H;{�H;��H;��H;��H;�H;      ��H;=�H;�H;�H;_�H;*�H;E�H;��H;0�H;��H;��H;l�H;2�H;��H;��H;(�H;��H;��H;��H;]�H;�H;w�H;��H;��H;��H;��H;;�H;��H;L�H;��H;��H;,�H;X�H;��H;��H;��H;��H;��H;��H;��H;X�H;,�H;��H;��H;L�H;��H;;�H;��H;��H;��H;��H;w�H;�H;]�H;��H;��H;��H;(�H;��H;��H;2�H;l�H;��H;��H;0�H;��H;E�H;*�H;_�H;�H;�H;=�H;      ��H;�H;ƩH;�H;ŬH;��H;��H;g�H;��H;кH;/�H;��H;��H;:�H;^�H;[�H;6�H;��H;H�H;e�H;S�H;��H;m�H;��H;��H;��H;��H;j�H;��H;T�H;��H; �H;9�H;u�H;��H;��H;��H;��H;��H;u�H;9�H; �H;��H;T�H;��H;j�H;��H;��H;��H;��H;m�H;��H;S�H;e�H;H�H;��H;6�H;[�H;^�H;:�H;��H;��H;/�H;кH;��H;g�H;��H;��H;ŬH;�H;ƩH;�H;      P�H;��H;��H;Z�H;��H;f�H;��H;O�H;.�H;H�H;��H;̸H;�H;=�H;4�H;��H;u�H;��H;��H;i�H;��H;��H;��H;K�H;��H;��H;��H;��H;b�H;�H;h�H;��H;	�H;9�H;X�H;�H;��H;�H;X�H;9�H;	�H;��H;h�H;�H;b�H;��H;��H;��H;��H;K�H;��H;��H;��H;i�H;��H;��H;u�H;��H;4�H;=�H;�H;̸H;��H;H�H;.�H;O�H;��H;f�H;��H;Z�H;��H;��H;      w�H;�H;B�H;u�H;j�H;$�H;p�H;/�H;H�H;��H;&�H;��H;#�H;�H;��H;f�H;��H;��H;��H;B�H;F�H;��H;Q�H;[�H;�H;��H;��H;��H;��H;m�H;�H;y�H;��H; �H;,�H;J�H;I�H;J�H;,�H; �H;��H;y�H;�H;m�H;��H;��H;��H;��H;�H;[�H;Q�H;��H;F�H;B�H;��H;��H;��H;f�H;��H;�H;#�H;��H;&�H;��H;H�H;/�H;p�H;$�H;j�H;u�H;B�H;�H;      fH;�fH;YhH;?kH;'oH;�sH;�yH;�H;��H;ۍH;�H;r�H;��H;��H;#�H;T�H;'�H;��H;x�H;��H;��H;1�H;=�H;��H;��H;��H;X�H;��H;��H;��H;t�H;�H;h�H;��H;��H;�H;0�H;�H;��H;��H;h�H;�H;t�H;��H;��H;��H;X�H;��H;��H;��H;=�H;1�H;��H;��H;x�H;��H;'�H;T�H;#�H;��H;��H;r�H;�H;ۍH;��H;�H;�yH;�sH;'oH;?kH;YhH;�fH;      9?H;@H;cBH;-FH;[KH;�QH;'YH;faH;JjH;�sH;/}H;ʆH;G�H;y�H;8�H;f�H;�H;׸H;�H;��H;��H;7�H;�H;[�H;9�H;��H;��H;K�H;��H;��H;��H;m�H;�H;T�H;��H;��H;��H;��H;��H;T�H;�H;m�H;��H;��H;��H;K�H;��H;��H;9�H;[�H;�H;7�H;��H;��H;�H;׸H;�H;f�H;8�H;y�H;G�H;ʆH;/}H;�sH;JjH;faH;'YH;�QH;[KH;-FH;cBH;@H;      >H;TH;uH;�H;mH;�$H;�.H;�9H;�EH;�QH;j^H;�jH;SwH;W�H;ԎH;��H;��H;��H;��H;ۻH;b�H;�H;��H;!�H;��H;��H;h�H;��H;,�H;��H;��H;��H;b�H;��H;L�H;�H;��H;�H;L�H;��H;b�H;��H;��H;��H;,�H;��H;h�H;��H;��H;!�H;��H;�H;b�H;ۻH;��H;��H;��H;��H;ԎH;W�H;SwH;�jH;j^H;�QH;�EH;�9H;�.H;�$H;mH;�H;uH;TH;      %�G;��G;��G;%�G;�G;5�G;"�G;�H;H;c&H;�6H;�GH;�WH;GgH;)vH;�H;�H;ԜH;T�H;��H;��H;D�H;��H;��H;}�H;k�H;��H;G�H;��H;K�H;��H;��H;��H;j�H;��H;�H; �H;�H;��H;j�H;��H;��H;��H;K�H;��H;G�H;��H;k�H;}�H;��H;��H;D�H;��H;��H;T�H;ԜH;�H;�H;)vH;GgH;�WH;�GH;�6H;c&H;H;�H;"�G;5�G;�G;%�G;��G;��G;      �mG;<pG;wG;�G;��G;^�G;{�G;��G;'�G;M�G;�H;oH;�/H;�CH;@WH;9iH;�yH;�H;��H;ӢH;m�H;��H;��H;��H;@�H;/�H;N�H;��H;h�H;��H;X�H;��H;��H;��H;;�H;��H;��H;��H;;�H;��H;��H;��H;X�H;��H;h�H;��H;N�H;/�H;@�H;��H;��H;��H;m�H;ӢH;��H;�H;�yH;9iH;@WH;�CH;�/H;oH;�H;M�G;'�G;��G;{�G;^�G;��G;�G;wG;<pG;      �F;�F;4�F;��F;,�F;� G;�EG;aiG;l�G;,�G;,�G;�G;<�G;�H;�0H;�GH;9]H;�pH;�H;��H;<�H;��H;��H;��H;��H;�H;/�H;k�H;��H;��H;��H;��H;��H;��H;��H;��H;�H;��H;��H;��H;��H;��H;��H;��H;��H;k�H;/�H;�H;��H;��H;��H;��H;<�H;��H;�H;�pH;9]H;�GH;�0H;�H;<�G;�G;,�G;,�G;l�G;aiG;�EG;� G;,�F;��F;4�F;�F;      ��D;B�D;A�D;�8E;��E;e�E;�OF;.�F;��F;J9G;lnG;ݙG;�G;��G;� H;�H;�9H;�RH;�hH;d|H;��H;��H;h�H;#�H;U�H;��H;@�H;}�H;��H;9�H;��H;�H;��H;��H;��H;-�H;q�H;-�H;��H;��H;��H;�H;��H;9�H;��H;}�H;@�H;��H;U�H;#�H;h�H;��H;��H;d|H;�hH;�RH;�9H;�H;� H;��G;�G;ݙG;lnG;J9G;��F;.�F;�OF;e�E;��E;�8E;A�D;B�D;      �@;�@@;f�@;]QA;"B;F
C;�C;��D;[�E;�?F;��F;� G;9gG;ÛG;`�G;�G;�H; .H;-JH;�bH;lxH;9�H;P�H;ۨH;#�H;��H;��H;��H;!�H;[�H;��H;[�H;K�H;��H;��H;i�H;��H;i�H;��H;��H;K�H;[�H;��H;[�H;!�H;��H;��H;��H;#�H;ۨH;P�H;9�H;lxH;�bH;-JH; .H;�H;�G;`�G;ÛG;9gG;� G;��F;�?F;[�E;��D;�C;F
C;"B;]QA;f�@;�@@;      �36;˃6;kk7;��8;��:;��<;��>;��@;�sB;��C;�+E;F;.�F;�+G;�wG;Y�G;��G;�H;%H;7DH;/_H;hvH;N�H;P�H;h�H;��H;��H;��H;��H;�H;=�H;Q�H;��H;m�H;��H;{�H;��H;{�H;��H;m�H;��H;Q�H;=�H;�H;��H;��H;��H;��H;h�H;P�H;N�H;hvH;/_H;7DH;%H;�H;��G;Y�G;�wG;�+G;.�F;F;�+E;��C;�sB;��@;��>;��<;��:;��8;kk7;˃6;      �";�L#;�%;��';��+;��/;@�3;��7;P�;;x?;N�A;��C;C9E;�?F;9�F;�TG;��G;S�G;��G;wH;AH;�]H;hvH;9�H;��H;��H;��H;D�H;�H;7�H;1�H;��H;��H;��H;w�H;U�H;��H;U�H;w�H;��H;��H;��H;1�H;7�H;�H;D�H;��H;��H;��H;9�H;hvH;�]H;AH;wH;��G;S�G;��G;�TG;9�F;�?F;C9E;��C;N�A;x?;P�;;��7;@�3;��/;��+;��';�%;�L#;      ���:�$ ;�;��;��;{P;�l;�c';v�.;�<5;E�:;�>;1B;YAD;��E;��F;+6G;��G;��G;F�G;�H;AH;/_H;lxH;��H;<�H;m�H;��H;b�H;��H;��H;F�H;��H;S�H;�H;��H;Z�H;��H;�H;S�H;��H;F�H;��H;��H;b�H;��H;m�H;<�H;��H;lxH;/_H;AH;�H;F�G;��G;��G;+6G;��F;��E;YAD;1B;�>;E�:;�<5;v�.;�c';�l;{P;��;��;�;�$ ;      Y�:�n�:W�:��:�%�:Ӵ�:���:��	;�P;RM#;�m-;��5;S�;;�@@;�OC;jFE;!uF;!G;��G;�G;F�G;wH;7DH;�bH;d|H;��H;ӢH;��H;ۻH;��H;��H;B�H;i�H;e�H;]�H;��H;��H;��H;]�H;e�H;i�H;B�H;��H;��H;ۻH;��H;ӢH;��H;d|H;�bH;7DH;wH;F�G;�G;��G;!G;!uF;jFE;�OC;�@@;S�;;��5;�m-;RM#;�P;��	;���:Ӵ�:�%�:��:W�:�n�:      �	�����j��(_���2u9�:�i~:���:[�:z�;�;�%;at0;�8;װ>;Z�B;��D;�WF;sG;��G;��G;��G;%H;-JH;�hH;�H;��H;T�H;��H;�H;x�H;��H;��H;H�H;��H;��H;h�H;��H;��H;H�H;��H;��H;x�H;�H;��H;T�H;��H;�H;�hH;-JH;%H;��G;��G;��G;sG;�WF;��D;Z�B;װ>;�8;at0;�%;�;z�;[�:���:�i~:�:�2u9(_���j�����      _A?���9��8)��Z�ܺlp������@994�@:�:~�:��	;�X;�,;8�6;֜=;x"B; �D;�WF;!G;��G;S�G;�H; .H;�RH;�pH;�H;ԜH;��H;׸H;��H;��H;��H;��H;��H;0�H;��H;0�H;��H;��H;��H;��H;��H;׸H;��H;ԜH;�H;�pH;�RH; .H;�H;S�G;��G;!G;�WF; �D;x"B;֜=;8�6;�,;�X;��	;~�:�:4�@:@99����lp��ܺ�Z��8)���9�      �Eֻ�ѻn�Ļ4T��`�r.o���.�ܺ��B�'��8�\:�%�:���:�P;]);�<5;K:=;x"B;��D;!uF;+6G;��G;��G;�H;�9H;9]H;�yH;�H;��H;�H;'�H;��H;u�H;6�H;��H;B�H;��H;B�H;��H;6�H;u�H;��H;'�H;�H;��H;�H;�yH;9]H;�9H;�H;��G;��G;+6G;!uF;��D;x"B;K:=;�<5;]);�P;���:�%�:�\:'��8��B�ܺ��.�r.o�`�4T��n�Ļ�ѻ      FB��>�s�4�$�$�G���Z�ۚ��oݎ�,A?�EӺ����g2�90q�:�W�:�;D�';�<5;֜=;Z�B;jFE;��F;�TG;Y�G;�G;�H;�GH;9iH;�H;��H;f�H;T�H;f�H;��H;[�H;(�H;5�H;��H;5�H;(�H;[�H;��H;f�H;T�H;f�H;��H;�H;9iH;�GH;�H;�G;Y�G;�TG;��F;jFE;Z�B;֜=;�<5;D�';�;�W�:0q�:g2�9����EӺ,A?�oݎ�ۚ���Z�G��$�$�s�4��>�      <y��ݜ��A���I����s�m�P��%+����Q�Ļ����|��o��8u9�W�:8+�:�;]);8�6;װ>;�OC;��E;9�F;�wG;`�G;� H;�0H;@WH;)vH;ԎH;8�H;#�H;��H;4�H;^�H;��H;�H;��H;�H;��H;^�H;4�H;��H;#�H;8�H;ԎH;)vH;@WH;�0H;� H;`�G;�wG;9�F;��E;�OC;װ>;8�6;]);�;8+�:�W�:�8u9�o�|�����Q�Ļ����%+�m�P���s��I���A��ݜ�      -������bW缑�ռ�վ��Τ��I��Z�[��(��Z�h�9��{���99�W�:�W�:�P;�,;�8;�@@;YAD;�?F;�+G;ÛG;��G;�H;�CH;GgH;W�H;y�H;��H;�H;=�H;:�H;��H;��H;��H;��H;��H;:�H;=�H;�H;��H;y�H;W�H;GgH;�CH;�H;��G;ÛG;�+G;�?F;YAD;�@@;�8;�,;�P;�W�:�W�:�99�{��h�9���Z��(�Z�[��I���Τ��վ���ռbW缧��      �6��3�X�+�ݟ�<�(�����μ߈��T���FB�=s�	T����D��{���8u90q�:���:�X;at0;S�;;1B;C9E;.�F;9gG;�G;<�G;�/H;�WH;SwH;G�H;��H;#�H;�H;��H;2�H;I�H;S�H;I�H;2�H;��H;�H;#�H;��H;G�H;SwH;�WH;�/H;<�G;�G;9gG;.�F;C9E;1B;S�;;at0;�X;���:0q�:�8u9�{����D�	T��=s�FB�T���߈����μ(���<�ݟ�X�+��3�      R₽�؀���u��Xc�Q�K�K1�{�����վ�t]��b�P�m��	T��h�9��o�g2�9�%�:��	;�%;��5;�>;��C;F;� G;ݙG;�G;oH;�GH;�jH;ʆH;r�H;��H;̸H;��H;l�H;��H;��H;��H;l�H;��H;̸H;��H;r�H;ʆH;�jH;�GH;oH;�G;ݙG;� G;F;��C;�>;��5;�%;��	;�%�:g2�9�o�h�9�	T��m��b�P�t]���վ����{��K1�Q�K��Xc���u��؀�      S���r��L��n������|�u�e�N���(�ji���˼�A��b�P�=s��|������\:~�:�;�m-;E�:;N�A;�+E;��F;lnG;,�G;�H;�6H;j^H;/}H;�H;&�H;��H;/�H;��H;Y�H;��H;Y�H;��H;/�H;��H;&�H;�H;/}H;j^H;�6H;�H;,�G;lnG;��F;�+E;N�A;E�:;�m-;�;~�:�\:����|��=s�b�P��A����˼ji���(�e�N�|�u�����n��L���r��      �o���r���}�ս@��Kĥ�X^���Xc��3���	���˼t]��FB��Z򻆜��EӺ'��8�:z�;RM#;�<5;x?;��C;�?F;J9G;,�G;M�G;c&H;�QH;�sH;ۍH;��H;H�H;кH;��H;��H;a�H;��H;��H;кH;H�H;��H;ۍH;�sH;�QH;c&H;M�G;,�G;J9G;�?F;��C;x?;�<5;RM#;z�;�:'��8EӺ�����Z�FB�t]����˼��	��3��Xc�X^��Kĥ�@��}�ս���r�      �#�6� �A'����~���gٽS��l���j��3�ji��վ�T����(�Q�Ļ,A?���B�4�@:[�:�P;v�.;P�;;�sB;[�E;��F;l�G;'�G;H;�EH;JjH;��H;H�H;.�H;��H;0�H;��H;�H;��H;0�H;��H;.�H;H�H;��H;JjH;�EH;H;'�G;l�G;��F;[�E;�sB;P�;;v�.;�P;[�:4�@:��B�,A?�Q�Ļ�(�T����վ�ji��3��j�l��S���gٽ�~����A'�6� �      �S� �O��E��5�6� �<�
���|9��l���Xc���(����߈��Z�[����oݎ�ܺ@99���:��	;�c';��7;��@;��D;.�F;aiG;��G;�H;�9H;faH;�H;/�H;O�H;g�H;��H;Y�H;��H;Y�H;��H;g�H;O�H;/�H;�H;faH;�9H;�H;��G;aiG;.�F;��D;��@;��7;�c';��	;���:@99ܺoݎ����Z�[�߈�������(��Xc�l��|9����<�
�6� ��5��E� �O�      �~���)����v��9b�U�H��",�0Z���S��X^��e�N�{����μ�I���%+�ۚ����.������i~:���:�l;@�3;��>;�C;�OF;�EG;{�G;"�G;�.H;'YH;�yH;p�H;��H;��H;E�H;J�H;��H;J�H;E�H;��H;��H;p�H;�yH;'YH;�.H;"�G;{�G;�EG;�OF;�C;��>;@�3;�l;���:�i~:������.�ۚ���%+��I����μ{��e�N�X^��S����0Z��",�U�H��9b���v��)��      ��������:���M���r� �O��",�<�
��gٽKĥ�|�u�K1�(����Τ�m�P��Z�r.o�lp���:Ӵ�:{P;��/;��<;F
C;e�E;� G;^�G;5�G;�$H;�QH;�sH;$�H;f�H;��H;*�H;{�H;&�H;{�H;*�H;��H;f�H;$�H;�sH;�QH;�$H;5�G;^�G;� G;e�E;F
C;��<;��/;{P;Ӵ�:�:lp��r.o��Z�m�P��Τ�(���K1�|�u�Kĥ��gٽ<�
��",� �O��r��M���:�����      ���v��/;������:P���r�U�H�6� ��~��@������Q�K�<��վ���s�G��`�ܺ�2u9�%�:��;��+;��:;"B;��E;,�F;��G;�G;mH;[KH;'oH;j�H;��H;ŬH;_�H;��H;��H;��H;_�H;ŬH;��H;j�H;'oH;[KH;mH;�G;��G;,�F;��E;"B;��:;��+;��;�%�:�2u9ܺ`�G����s��վ�<�Q�K�����@���~��6� �U�H��r�:P������/;���v��      3Vھ�*־5ʾT��������M���9b��5���}�սn���Xc�ݟ���ռ�I��$�$�4T���Z�(_����:��;��';��8;]QA;�8E;��F;�G;%�G;�H;-FH;?kH;u�H;Z�H;�H;�H;��H;t�H;��H;�H;�H;Z�H;u�H;?kH;-FH;�H;%�G;�G;��F;�8E;]QA;��8;��';��;��:(_���Z�4T��$�$��I����ռݟ��Xc�n��}�ս���5��9b��M������T���5ʾ�*־      ǰ�쾐�޾5ʾ/;���:����v��E�A'���L����u�X�+�bW缨A��s�4�n�Ļ�8)��j��W�:�;�%;kk7;f�@;A�D;4�F;wG;��G;uH;cBH;YhH;B�H;��H;ƩH;�H;��H;��H;��H;�H;ƩH;��H;B�H;YhH;cBH;uH;��G;wG;4�F;A�D;f�@;kk7;�%;�;W�:�j���8)�n�Ļs�4��A��bW�X�+���u�L����A'��E���v��:��/;��5ʾ��޾��      /h���b���쾅*־�v������)�� �O�6� ��r�r���؀��3����ݜ��>��ѻ��9�����n�:�$ ;�L#;˃6;�@@;B�D;�F;<pG;��G;TH;@H;�fH;�H;��H;�H;=�H;�H;��H;�H;=�H;�H;��H;�H;�fH;@H;TH;��G;<pG;�F;B�D;�@@;˃6;�L#;�$ ;�n�:�����9��ѻ�>�ݜ�����3��؀��r���r�6� � �O��)������v���*־�쾼b��      �$��� ���������þ�*��
Dx�}�=����\Pν鰒��&K�xc����;�V�s���D^���S��v[:���:�d;��4;�_?;�lD;��F;puG;M�G;�H;�NH;�rH;�H;��H;��H;�H;q�H;E�H;q�H;�H;��H;��H;�H;�rH;�NH;�H;M�G;puG;��F;�lD;�_?;��4;�d;���:�v[:��S��D^�s��;�V����xc��&K�鰒�\Pν���}�=�
Dx��*���þ��������� �      �� �k��>��=���������0���s���:�N9���ʽZ����G��8��-��z5S�w���/X���D��Ad:�A�:� ;x�4;	�?;#~D;p�F;3xG;��G;�H;NOH;HsH;:�H;�H;�H;W�H;��H;U�H;��H;W�H;�H;�H;:�H;HsH;NOH;�H;��G;3xG;p�F;#~D;	�?;x�4;� ;�A�:�Ad:��D��/X�w��z5S��-���8���G�Z����ʽN9���:��s��0��������=��>��k��      ���>��&�
�����fYؾ���ȥ����f���0�C[�*8������ȟ>�|���#Ȥ�Y6H�,�ܻ�qF�0��4�}:���:�";��5;6�?;��D;��F;/�G;��G;s"H;�QH;�tH;y�H;�H;��H;�H;�H;��H;�H;�H;��H;�H;y�H;�tH;�QH;s"H;��G;/�G;��F;��D;6�?;��5;�";���:4�}:0���qF�,�ܻY6H�#Ȥ�|���ȟ>�����*8��C[���0���f�ȥ�����fYؾ����&�
�>��      ��=������I��þ�R��&���QS��Q"��s�����}��0���d���x�6��ƻ(}*����^�:�w;�%;Rl7;�@;�D;�F;��G;��G;3'H;UH;�wH;�H;f�H;±H;ۺH;�H;��H;�H;ۺH;±H;f�H;�H;�wH;UH;3'H;��G;��G;�F;�D;�@;Rl7;�%;�w;^�:���(}*��ƻx�6�d����켟0���}�����s��Q"�QS�&����R���þIᾁ���=��      ����fYؾ�þ�ê�f쏾jk���:�e�R�ؽ�����c�:y���Ҽݫ��� �B�(���'7��:�
;c�(;�^9;��A;�[E;��F;�G;��G;�-H;�YH;{H;�H;i�H;u�H;6�H;�H;��H;�H;6�H;u�H;i�H;�H;{H;�YH;�-H;��G;�G;��F;�[E;��A;�^9;c�(;�
;��:�'7(��B�� �ݫ����Ҽ:y��c�����R�ؽe���:�jk�f쏾�ê��þfYؾ��      �þ��������R��f쏾�s��H����������������D�vc�g����f�3,�����P����9/��:5;�i-;��;;��B;+�E;�G;��G;��G;�5H;�_H;�H;{�H;�H;q�H;ɽH;r�H;��H;r�H;ɽH;q�H;�H;{�H;�H;�_H;�5H;��G;��G;�G;+�E;��B;��;;�i-;5;/��:��9�P�����3,��f�g���vc���D���������������H��s�f쏾�R���������      �*���0��ȥ��&���jk��H��#%�B[�ZPν�s��0�f�/%�d��`���G�=�n?ػgFL��D�`�R:B�:��;�2;�=;��C;�/F;�FG;�G;WH;?H;�fH;��H;V�H;ͫH;��H;��H;�H;��H;�H;��H;��H;ͫH;V�H;��H;�fH;?H;WH;�G;�FG;�/F;��C;�=;�2;��;B�:`�R:�D�gFL�n?ػG�=�`���d��/%�0�f��s��ZPνB[��#%��H�jk�&���ȥ���0��      
Dx��s���f�QS���:����B[��7ս�榽��}�u�;��8�)�����r����G������Ҭ����:��;}$;,�6;f�?;3�D;�F;�oG;��G;H;XIH;dnH;i�H;��H;�H;Z�H;��H;��H;G�H;��H;��H;Z�H;�H;��H;i�H;dnH;XIH;H;��G;�oG;�F;3�D;f�?;,�6;}$;��;���:�Ҭ����G�������r�)����8�u�;���}��榽�7սB[������:�QS���f��s�      }�=���:���0��Q"�e�����ZPν�榽%����G�����Ҽ���E:�
�ܻ�D^�ϸ��ih:���:O;�{,;�:;��A;~hE;��F;\�G;��G;�'H;eTH;�vH;��H;L�H;��H;�H;��H;��H;3�H;��H;��H;�H;��H;L�H;��H;�vH;eTH;�'H;��G;\�G;��F;~hE;��A;�:;�{,;O;���:ih:ϸ���D^�
�ܻE:������Ҽ����G�%���榽ZPν����e��Q"���0���:�      ���N9�C[��s�R�ؽ���s����}���G��K��	c��!�V�%,��*�����+����:?��:� ;ǂ3;0>;�C;"F;#8G;l�G;�H;7H;�_H;,H;�H; �H;g�H;�H;m�H;��H;3�H;��H;m�H;�H;g�H; �H;�H;,H;�_H;7H;�H;l�G;#8G;"F;�C;0>;ǂ3;� ;?��:��:+������*��%,�!�V�	c��K�����G���}��s����R�ؽ�s�C[�N9�      \Pν��ʽ*8�������������0�f�u�;���K��Ȥ���f���$ߵ�?o5�5�D�L�-:���:X>;G+;_9;�A;��D;[�F;�uG;�G;IH;�FH;�kH;�H;��H;�H;H�H;�H;��H;"�H;F�H;"�H;��H;�H;H�H;�H;��H;�H;�kH;�FH;IH;�G;�uG;[�F;��D;�A;_9;G+;X>;���:L�-:5�D�?o5�$ߵ�����f�Ȥ�K����u�;�0�f������������*8����ʽ      鰒�Z��������}��c���D�/%��8���Ҽ	c����f�����ƻZ/X�u���年9f�:ȏ;F";�3;�>;�XC;��E;G;'�G;��G;�+H;/VH;9wH;��H;W�H;�H;.�H;�H;Q�H;`�H;N�H;`�H;Q�H;�H;.�H;�H;W�H;��H;9wH;/VH;�+H;��G;'�G;G;��E;�XC;�>;�3;F";ȏ;f�:年9u���Z/X��ƻ�����f�	c����Ҽ�8�/%���D��c���}�����Z��      �&K���G�ȟ>��0�:y�vc�d��)������!�V����ƻgod���º�P(7�3�:���:�;]P.;9�:;ayA;y�D;�F;�mG;t�G;!H;�?H;MeH;��H;R�H;ժH;��H;�H;	�H;��H;��H;V�H;��H;��H;	�H;�H;��H;ժH;R�H;��H;MeH;�?H;!H;t�G;�mG;�F;y�D;ayA;9�:;]P.;�;���:�3�:�P(7��ºgod��ƻ��!�V����)���d��vc�:y��0�ȟ>���G�      xc��8�|����켔�Ҽg���`�����r�E:�%,�$ߵ�Z/X���º̬�E�}:> �:v;��);�l7;i�?;�C;KF;�(G;E�G;�G;2)H;�RH;�sH;��H;��H;�H;ͼH;��H;��H;+�H;��H;l�H;��H;+�H;��H;��H;ͼH;�H;��H;��H;�sH;�RH;2)H;�G;E�G;�(G;KF;�C;i�?;�l7;��);v;> �:E�}:̬���ºZ/X�$ߵ�%,�E:���r�`���g�����Ҽ��|����8�      ����-��#Ȥ�d���ݫ���f�G�=����
�ܻ�*��?o5�u����P(7E�}:�m�:��;>&;��4;B�=;�B;+�E;S�F;ˀG;$�G;cH;�@H;�dH;d�H;��H;x�H;��H;��H;;�H;��H;��H;��H;l�H;��H;��H;��H;;�H;��H;��H;x�H;��H;d�H;�dH;�@H;cH;$�G;ˀG;S�F;+�E;�B;B�=;��4;>&;��;�m�:E�}:�P(7u���?o5��*��
�ܻ���G�=��f�ݫ��d���#Ȥ��-��      ;�V�z5S�Y6H�x�6�� �3,�n?ػG���D^����5�D�年9�3�:> �:��;]%;��3;p�<;�B;�
E;>�F;�WG;8�G;t�G;�/H;wVH;�uH;�H;��H;ܰH;��H;��H;��H;k�H;��H;��H;Q�H;��H;��H;k�H;��H;��H;��H;ܰH;��H;�H;�uH;wVH;�/H;t�G;8�G;�WG;>�F;�
E;�B;p�<;��3;]%;��;> �:�3�:年95�D�����D^�G��n?ػ3,�� �x�6�Y6H�z5S�      s��w��,�ܻ�ƻB󩻜��gFL����ϸ��+��L�-:f�:���:v;>&;��3;�8<;_�A;%�D;�YF;Z4G;3�G;�G;� H;`IH;VjH;ńH;ٙH;��H;��H;�H;��H;��H;��H;��H;v�H;�H;v�H;��H;��H;��H;��H;�H;��H;��H;ٙH;ńH;VjH;`IH;� H;�G;3�G;Z4G;�YF;%�D;_�A;�8<;��3;>&;v;���:f�:L�-:+��ϸ�����gFL����B��ƻ,�ܻw��      �D^��/X��qF�(}*�(���P���D��Ҭ�ih:��:���:ȏ;�;��);��4;p�<;_�A;f�D;�8F;
G;��G;w�G;jH;C>H;�`H;5|H;��H;��H;��H;��H;��H;|�H;��H;4�H;��H;8�H;��H;8�H;��H;4�H;��H;|�H;��H;��H;��H;��H;��H;5|H;�`H;C>H;jH;w�G;��G;
G;�8F;f�D;_�A;p�<;��4;��);�;ȏ;���:��:ih:�Ҭ��D��P��(��(}*��qF��/X�      ��S���D�0������'7��9`�R:���:���:?��:X>;F";]P.;�l7;B�=;�B;%�D;�8F;XG;R�G;��G;�H;�5H;�XH;uH;=�H;�H;�H;�H;��H;9�H;��H;-�H;M�H;r�H;��H;�H;��H;r�H;M�H;-�H;��H;9�H;��H;�H;�H;�H;=�H;uH;�XH;�5H;�H;��G;R�G;XG;�8F;%�D;�B;B�=;�l7;]P.;F";X>;?��:���:���:`�R:��9�'7���0����D�      �v[:�Ad:4�}:^�:��:/��:B�:��;O;� ;G+;�3;9�:;i�?;�B;�
E;�YF;
G;R�G;��G;nH;�0H;�RH;�oH;�H;f�H; �H;��H;��H;��H;�H;��H;��H;5�H;�H;(�H;q�H;(�H;�H;5�H;��H;��H;�H;��H;��H;��H; �H;f�H;�H;�oH;�RH;�0H;nH;��G;R�G;
G;�YF;�
E;�B;i�?;9�:;�3;G+;� ;O;��;B�:/��:��:^�:4�}:�Ad:      ���:�A�:���:�w;�
;5;��;}$;�{,;ǂ3;_9;�>;ayA;�C;+�E;>�F;Z4G;��G;��G;nH;�.H;PH;&lH;i�H;��H;��H;��H;�H;��H;)�H;r�H;��H;��H;��H;y�H;W�H;��H;W�H;y�H;��H;��H;��H;r�H;)�H;��H;�H;��H;��H;��H;i�H;&lH;PH;�.H;nH;��G;��G;Z4G;>�F;+�E;�C;ayA;�>;_9;ǂ3;�{,;}$;��;5;�
;�w;���:�A�:      �d;� ;�";�%;c�(;�i-;�2;,�6;�:;0>;�A;�XC;y�D;KF;S�F;�WG;3�G;w�G;�H;�0H;PH;�jH;��H;��H;V�H;E�H;�H;��H;��H;�H;��H;��H;��H;�H;��H;j�H;��H;j�H;��H;�H;��H;��H;��H;�H;��H;��H;�H;E�H;V�H;��H;��H;�jH;PH;�0H;�H;w�G;3�G;�WG;S�F;KF;y�D;�XC;�A;0>;�:;,�6;�2;�i-;c�(;�%;�";� ;      ��4;x�4;��5;Rl7;�^9;��;;�=;f�?;��A;�C;��D;��E;�F;�(G;ˀG;8�G;�G;jH;�5H;�RH;&lH;��H;˓H;#�H;گH;g�H;<�H;H�H;��H;��H;(�H;��H;C�H;��H;��H;m�H;��H;m�H;��H;��H;C�H;��H;(�H;��H;��H;H�H;<�H;g�H;گH;#�H;˓H;��H;&lH;�RH;�5H;jH;�G;8�G;ˀG;�(G;�F;��E;��D;�C;��A;f�?;�=;��;;�^9;Rl7;��5;x�4;      �_?;	�?;6�?;�@;��A;��B;��C;3�D;~hE;"F;[�F;G;�mG;E�G;$�G;t�G;� H;C>H;�XH;�oH;i�H;��H;#�H;\�H;��H;;�H;Y�H;�H;��H;��H;g�H;��H;��H;��H;��H;E�H;^�H;E�H;��H;��H;��H;��H;g�H;��H;��H;�H;Y�H;;�H;��H;\�H;#�H;��H;i�H;�oH;�XH;C>H;� H;t�G;$�G;E�G;�mG;G;[�F;"F;~hE;3�D;��C;��B;��A;�@;6�?;	�?;      �lD;#~D;��D;�D;�[E;+�E;�/F;�F;��F;#8G;�uG;'�G;t�G;�G;cH;�/H;`IH;�`H;uH;�H;��H;V�H;گH;��H;�H;��H;}�H;#�H;��H;�H;n�H;N�H;��H;��H;��H;��H;6�H;��H;��H;��H;��H;N�H;n�H;�H;��H;#�H;}�H;��H;�H;��H;گH;V�H;��H;�H;uH;�`H;`IH;�/H;cH;�G;t�G;'�G;�uG;#8G;��F;�F;�/F;+�E;�[E;�D;��D;#~D;      ��F;p�F;��F;�F;��F;�G;�FG;�oG;\�G;l�G;�G;��G;!H;2)H;�@H;wVH;VjH;5|H;=�H;f�H;��H;E�H;g�H;;�H;��H;E�H;��H;��H;��H;�H;�H;��H;��H;��H;B�H;��H;��H;��H;B�H;��H;��H;��H;�H;�H;��H;��H;��H;E�H;��H;;�H;g�H;E�H;��H;f�H;=�H;5|H;VjH;wVH;�@H;2)H;!H;��G;�G;l�G;\�G;�oG;�FG;�G;��F;�F;��F;p�F;      puG;3xG;/�G;��G;�G;��G;�G;��G;��G;�H;IH;�+H;�?H;�RH;�dH;�uH;ńH;��H;�H; �H;��H;�H;<�H;Y�H;}�H;��H;t�H;l�H;��H;��H;n�H;��H;��H;L�H;��H;-�H;.�H;-�H;��H;L�H;��H;��H;n�H;��H;��H;l�H;t�H;��H;}�H;Y�H;<�H;�H;��H; �H;�H;��H;ńH;�uH;�dH;�RH;�?H;�+H;IH;�H;��G;��G;�G;��G;�G;��G;/�G;3xG;      M�G;��G;��G;��G;��G;��G;WH;H;�'H;7H;�FH;/VH;MeH;�sH;d�H;�H;ٙH;��H;�H;��H;�H;��H;H�H;�H;#�H;��H;l�H;��H;��H;p�H;��H;��H;c�H;��H;U�H;��H;��H;��H;U�H;��H;c�H;��H;��H;p�H;��H;��H;l�H;��H;#�H;�H;H�H;��H;�H;��H;�H;��H;ٙH;�H;d�H;�sH;MeH;/VH;�FH;7H;�'H;H;WH;��G;��G;��G;��G;��G;      �H;�H;s"H;3'H;�-H;�5H;?H;XIH;eTH;�_H;�kH;9wH;��H;��H;��H;��H;��H;��H;�H;��H;��H;��H;��H;��H;��H;��H;��H;��H;>�H;��H;��H;X�H;��H;y�H;��H;��H;��H;��H;��H;y�H;��H;X�H;��H;��H;>�H;��H;��H;��H;��H;��H;��H;��H;��H;��H;�H;��H;��H;��H;��H;��H;��H;9wH;�kH;�_H;eTH;XIH;?H;�5H;�-H;3'H;s"H;�H;      �NH;NOH;�QH;UH;�YH;�_H;�fH;dnH;�vH;,H;�H;��H;R�H;��H;x�H;ܰH;��H;��H;��H;��H;)�H;�H;��H;��H;�H;�H;��H;p�H;��H;��H;V�H;��H;q�H;��H;�H;%�H;?�H;%�H;�H;��H;q�H;��H;V�H;��H;��H;p�H;��H;�H;�H;��H;��H;�H;)�H;��H;��H;��H;��H;ܰH;x�H;��H;R�H;��H;�H;,H;�vH;dnH;�fH;�_H;�YH;UH;�QH;NOH;      �rH;HsH;�tH;�wH;{H;�H;��H;i�H;��H;�H;��H;W�H;ժH;�H;��H;��H;�H;��H;9�H;�H;r�H;��H;(�H;g�H;n�H;�H;n�H;��H;��H;V�H;��H;q�H;��H;�H;_�H;l�H;d�H;l�H;_�H;�H;��H;q�H;��H;V�H;��H;��H;n�H;�H;n�H;g�H;(�H;��H;r�H;�H;9�H;��H;�H;��H;��H;�H;ժH;W�H;��H;�H;��H;i�H;��H;�H;{H;�wH;�tH;HsH;      �H;:�H;y�H;�H;�H;{�H;V�H;��H;L�H; �H;�H;�H;��H;ͼH;��H;��H;��H;|�H;��H;��H;��H;��H;��H;��H;N�H;��H;��H;��H;X�H;��H;q�H;��H;�H;_�H;��H;��H;��H;��H;��H;_�H;�H;��H;q�H;��H;X�H;��H;��H;��H;N�H;��H;��H;��H;��H;��H;��H;|�H;��H;��H;��H;ͼH;��H;�H;�H; �H;L�H;��H;V�H;{�H;�H;�H;y�H;:�H;      ��H;�H;�H;f�H;i�H;�H;ͫH;�H;��H;g�H;H�H;.�H;�H;��H;;�H;��H;��H;��H;-�H;��H;��H;��H;C�H;��H;��H;��H;��H;c�H;��H;q�H;��H;�H;X�H;��H;��H;��H;��H;��H;��H;��H;X�H;�H;��H;q�H;��H;c�H;��H;��H;��H;��H;C�H;��H;��H;��H;-�H;��H;��H;��H;;�H;��H;�H;.�H;H�H;g�H;��H;�H;ͫH;�H;i�H;f�H;�H;�H;      ��H;�H;��H;±H;u�H;q�H;��H;Z�H;�H;�H;�H;�H;	�H;��H;��H;k�H;��H;4�H;M�H;5�H;��H;�H;��H;��H;��H;��H;L�H;��H;y�H;��H;�H;_�H;��H;��H;��H;��H;��H;��H;��H;��H;��H;_�H;�H;��H;y�H;��H;L�H;��H;��H;��H;��H;�H;��H;5�H;M�H;4�H;��H;k�H;��H;��H;	�H;�H;�H;�H;�H;Z�H;��H;q�H;u�H;±H;��H;�H;      �H;W�H;�H;ۺH;6�H;ɽH;��H;��H;��H;m�H;��H;Q�H;��H;+�H;��H;��H;��H;��H;r�H;�H;y�H;��H;��H;��H;��H;B�H;��H;U�H;��H;�H;_�H;��H;��H;��H;��H;��H;��H;��H;��H;��H;��H;��H;_�H;�H;��H;U�H;��H;B�H;��H;��H;��H;��H;y�H;�H;r�H;��H;��H;��H;��H;+�H;��H;Q�H;��H;m�H;��H;��H;��H;ɽH;6�H;ۺH;�H;W�H;      q�H;��H;�H;�H;�H;r�H;�H;��H;��H;��H;"�H;`�H;��H;��H;��H;��H;v�H;8�H;��H;(�H;W�H;j�H;m�H;E�H;��H;��H;-�H;��H;��H;%�H;l�H;��H;��H;��H;��H;��H;��H;��H;��H;��H;��H;��H;l�H;%�H;��H;��H;-�H;��H;��H;E�H;m�H;j�H;W�H;(�H;��H;8�H;v�H;��H;��H;��H;��H;`�H;"�H;��H;��H;��H;�H;r�H;�H;�H;�H;��H;      E�H;U�H;��H;��H;��H;��H;��H;G�H;3�H;3�H;F�H;N�H;V�H;l�H;l�H;Q�H;�H;��H;�H;q�H;��H;��H;��H;^�H;6�H;��H;.�H;��H;��H;?�H;d�H;��H;��H;��H;��H;��H;��H;��H;��H;��H;��H;��H;d�H;?�H;��H;��H;.�H;��H;6�H;^�H;��H;��H;��H;q�H;�H;��H;�H;Q�H;l�H;l�H;V�H;N�H;F�H;3�H;3�H;G�H;��H;��H;��H;��H;��H;U�H;      q�H;��H;�H;�H;�H;r�H;�H;��H;��H;��H;"�H;`�H;��H;��H;��H;��H;v�H;8�H;��H;(�H;W�H;j�H;m�H;E�H;��H;��H;-�H;��H;��H;%�H;l�H;��H;��H;��H;��H;��H;��H;��H;��H;��H;��H;��H;l�H;%�H;��H;��H;-�H;��H;��H;E�H;m�H;j�H;W�H;(�H;��H;8�H;v�H;��H;��H;��H;��H;`�H;"�H;��H;��H;��H;�H;r�H;�H;�H;�H;��H;      �H;W�H;�H;ۺH;6�H;ɽH;��H;��H;��H;m�H;��H;Q�H;��H;+�H;��H;��H;��H;��H;r�H;�H;y�H;��H;��H;��H;��H;B�H;��H;U�H;��H;�H;_�H;��H;��H;��H;��H;��H;��H;��H;��H;��H;��H;��H;_�H;�H;��H;U�H;��H;B�H;��H;��H;��H;��H;y�H;�H;r�H;��H;��H;��H;��H;+�H;��H;Q�H;��H;m�H;��H;��H;��H;ɽH;6�H;ۺH;�H;W�H;      ��H;�H;��H;±H;u�H;q�H;��H;Z�H;�H;�H;�H;�H;	�H;��H;��H;k�H;��H;4�H;M�H;5�H;��H;�H;��H;��H;��H;��H;L�H;��H;y�H;��H;�H;_�H;��H;��H;��H;��H;��H;��H;��H;��H;��H;_�H;�H;��H;y�H;��H;L�H;��H;��H;��H;��H;�H;��H;5�H;M�H;4�H;��H;k�H;��H;��H;	�H;�H;�H;�H;�H;Z�H;��H;q�H;u�H;±H;��H;�H;      ��H;�H;�H;f�H;i�H;�H;ͫH;�H;��H;g�H;H�H;.�H;�H;��H;;�H;��H;��H;��H;-�H;��H;��H;��H;C�H;��H;��H;��H;��H;c�H;��H;q�H;��H;�H;X�H;��H;��H;��H;��H;��H;��H;��H;X�H;�H;��H;q�H;��H;c�H;��H;��H;��H;��H;C�H;��H;��H;��H;-�H;��H;��H;��H;;�H;��H;�H;.�H;H�H;g�H;��H;�H;ͫH;�H;i�H;f�H;�H;�H;      �H;:�H;y�H;�H;�H;{�H;V�H;��H;L�H; �H;�H;�H;��H;ͼH;��H;��H;��H;|�H;��H;��H;��H;��H;��H;��H;N�H;��H;��H;��H;X�H;��H;q�H;��H;�H;_�H;��H;��H;��H;��H;��H;_�H;�H;��H;q�H;��H;X�H;��H;��H;��H;N�H;��H;��H;��H;��H;��H;��H;|�H;��H;��H;��H;ͼH;��H;�H;�H; �H;L�H;��H;V�H;{�H;�H;�H;y�H;:�H;      �rH;HsH;�tH;�wH;{H;�H;��H;i�H;��H;�H;��H;W�H;ժH;�H;��H;��H;�H;��H;9�H;�H;r�H;��H;(�H;g�H;n�H;�H;n�H;��H;��H;V�H;��H;q�H;��H;�H;_�H;l�H;d�H;l�H;_�H;�H;��H;q�H;��H;V�H;��H;��H;n�H;�H;n�H;g�H;(�H;��H;r�H;�H;9�H;��H;�H;��H;��H;�H;ժH;W�H;��H;�H;��H;i�H;��H;�H;{H;�wH;�tH;HsH;      �NH;NOH;�QH;UH;�YH;�_H;�fH;dnH;�vH;,H;�H;��H;R�H;��H;x�H;ܰH;��H;��H;��H;��H;)�H;�H;��H;��H;�H;�H;��H;p�H;��H;��H;V�H;��H;q�H;��H;�H;%�H;?�H;%�H;�H;��H;q�H;��H;V�H;��H;��H;p�H;��H;�H;�H;��H;��H;�H;)�H;��H;��H;��H;��H;ܰH;x�H;��H;R�H;��H;�H;,H;�vH;dnH;�fH;�_H;�YH;UH;�QH;NOH;      �H;�H;s"H;3'H;�-H;�5H;?H;XIH;eTH;�_H;�kH;9wH;��H;��H;��H;��H;��H;��H;�H;��H;��H;��H;��H;��H;��H;��H;��H;��H;>�H;��H;��H;X�H;��H;y�H;��H;��H;��H;��H;��H;y�H;��H;X�H;��H;��H;>�H;��H;��H;��H;��H;��H;��H;��H;��H;��H;�H;��H;��H;��H;��H;��H;��H;9wH;�kH;�_H;eTH;XIH;?H;�5H;�-H;3'H;s"H;�H;      M�G;��G;��G;��G;��G;��G;WH;H;�'H;7H;�FH;/VH;MeH;�sH;d�H;�H;ٙH;��H;�H;��H;�H;��H;H�H;�H;#�H;��H;l�H;��H;��H;p�H;��H;��H;c�H;��H;U�H;��H;��H;��H;U�H;��H;c�H;��H;��H;p�H;��H;��H;l�H;��H;#�H;�H;H�H;��H;�H;��H;�H;��H;ٙH;�H;d�H;�sH;MeH;/VH;�FH;7H;�'H;H;WH;��G;��G;��G;��G;��G;      puG;3xG;/�G;��G;�G;��G;�G;��G;��G;�H;IH;�+H;�?H;�RH;�dH;�uH;ńH;��H;�H; �H;��H;�H;<�H;Y�H;}�H;��H;t�H;l�H;��H;��H;n�H;��H;��H;L�H;��H;-�H;.�H;-�H;��H;L�H;��H;��H;n�H;��H;��H;l�H;t�H;��H;}�H;Y�H;<�H;�H;��H; �H;�H;��H;ńH;�uH;�dH;�RH;�?H;�+H;IH;�H;��G;��G;�G;��G;�G;��G;/�G;3xG;      ��F;p�F;��F;�F;��F;�G;�FG;�oG;\�G;l�G;�G;��G;!H;2)H;�@H;wVH;VjH;5|H;=�H;f�H;��H;E�H;g�H;;�H;��H;E�H;��H;��H;��H;�H;�H;��H;��H;��H;B�H;��H;��H;��H;B�H;��H;��H;��H;�H;�H;��H;��H;��H;E�H;��H;;�H;g�H;E�H;��H;f�H;=�H;5|H;VjH;wVH;�@H;2)H;!H;��G;�G;l�G;\�G;�oG;�FG;�G;��F;�F;��F;p�F;      �lD;#~D;��D;�D;�[E;+�E;�/F;�F;��F;#8G;�uG;'�G;t�G;�G;cH;�/H;`IH;�`H;uH;�H;��H;V�H;گH;��H;�H;��H;}�H;#�H;��H;�H;n�H;N�H;��H;��H;��H;��H;6�H;��H;��H;��H;��H;N�H;n�H;�H;��H;#�H;}�H;��H;�H;��H;گH;V�H;��H;�H;uH;�`H;`IH;�/H;cH;�G;t�G;'�G;�uG;#8G;��F;�F;�/F;+�E;�[E;�D;��D;#~D;      �_?;	�?;6�?;�@;��A;��B;��C;3�D;~hE;"F;[�F;G;�mG;E�G;$�G;t�G;� H;C>H;�XH;�oH;i�H;��H;#�H;\�H;��H;;�H;Y�H;�H;��H;��H;g�H;��H;��H;��H;��H;E�H;^�H;E�H;��H;��H;��H;��H;g�H;��H;��H;�H;Y�H;;�H;��H;\�H;#�H;��H;i�H;�oH;�XH;C>H;� H;t�G;$�G;E�G;�mG;G;[�F;"F;~hE;3�D;��C;��B;��A;�@;6�?;	�?;      ��4;x�4;��5;Rl7;�^9;��;;�=;f�?;��A;�C;��D;��E;�F;�(G;ˀG;8�G;�G;jH;�5H;�RH;&lH;��H;˓H;#�H;گH;g�H;<�H;H�H;��H;��H;(�H;��H;C�H;��H;��H;m�H;��H;m�H;��H;��H;C�H;��H;(�H;��H;��H;H�H;<�H;g�H;گH;#�H;˓H;��H;&lH;�RH;�5H;jH;�G;8�G;ˀG;�(G;�F;��E;��D;�C;��A;f�?;�=;��;;�^9;Rl7;��5;x�4;      �d;� ;�";�%;c�(;�i-;�2;,�6;�:;0>;�A;�XC;y�D;KF;S�F;�WG;3�G;w�G;�H;�0H;PH;�jH;��H;��H;V�H;E�H;�H;��H;��H;�H;��H;��H;��H;�H;��H;j�H;��H;j�H;��H;�H;��H;��H;��H;�H;��H;��H;�H;E�H;V�H;��H;��H;�jH;PH;�0H;�H;w�G;3�G;�WG;S�F;KF;y�D;�XC;�A;0>;�:;,�6;�2;�i-;c�(;�%;�";� ;      ���:�A�:���:�w;�
;5;��;}$;�{,;ǂ3;_9;�>;ayA;�C;+�E;>�F;Z4G;��G;��G;nH;�.H;PH;&lH;i�H;��H;��H;��H;�H;��H;)�H;r�H;��H;��H;��H;y�H;W�H;��H;W�H;y�H;��H;��H;��H;r�H;)�H;��H;�H;��H;��H;��H;i�H;&lH;PH;�.H;nH;��G;��G;Z4G;>�F;+�E;�C;ayA;�>;_9;ǂ3;�{,;}$;��;5;�
;�w;���:�A�:      �v[:�Ad:4�}:^�:��:/��:B�:��;O;� ;G+;�3;9�:;i�?;�B;�
E;�YF;
G;R�G;��G;nH;�0H;�RH;�oH;�H;f�H; �H;��H;��H;��H;�H;��H;��H;5�H;�H;(�H;q�H;(�H;�H;5�H;��H;��H;�H;��H;��H;��H; �H;f�H;�H;�oH;�RH;�0H;nH;��G;R�G;
G;�YF;�
E;�B;i�?;9�:;�3;G+;� ;O;��;B�:/��:��:^�:4�}:�Ad:      ��S���D�0������'7��9`�R:���:���:?��:X>;F";]P.;�l7;B�=;�B;%�D;�8F;XG;R�G;��G;�H;�5H;�XH;uH;=�H;�H;�H;�H;��H;9�H;��H;-�H;M�H;r�H;��H;�H;��H;r�H;M�H;-�H;��H;9�H;��H;�H;�H;�H;=�H;uH;�XH;�5H;�H;��G;R�G;XG;�8F;%�D;�B;B�=;�l7;]P.;F";X>;?��:���:���:`�R:��9�'7���0����D�      �D^��/X��qF�(}*�(���P���D��Ҭ�ih:��:���:ȏ;�;��);��4;p�<;_�A;f�D;�8F;
G;��G;w�G;jH;C>H;�`H;5|H;��H;��H;��H;��H;��H;|�H;��H;4�H;��H;8�H;��H;8�H;��H;4�H;��H;|�H;��H;��H;��H;��H;��H;5|H;�`H;C>H;jH;w�G;��G;
G;�8F;f�D;_�A;p�<;��4;��);�;ȏ;���:��:ih:�Ҭ��D��P��(��(}*��qF��/X�      s��w��,�ܻ�ƻB󩻜��gFL����ϸ��+��L�-:f�:���:v;>&;��3;�8<;_�A;%�D;�YF;Z4G;3�G;�G;� H;`IH;VjH;ńH;ٙH;��H;��H;�H;��H;��H;��H;��H;v�H;�H;v�H;��H;��H;��H;��H;�H;��H;��H;ٙH;ńH;VjH;`IH;� H;�G;3�G;Z4G;�YF;%�D;_�A;�8<;��3;>&;v;���:f�:L�-:+��ϸ�����gFL����B��ƻ,�ܻw��      ;�V�z5S�Y6H�x�6�� �3,�n?ػG���D^����5�D�年9�3�:> �:��;]%;��3;p�<;�B;�
E;>�F;�WG;8�G;t�G;�/H;wVH;�uH;�H;��H;ܰH;��H;��H;��H;k�H;��H;��H;Q�H;��H;��H;k�H;��H;��H;��H;ܰH;��H;�H;�uH;wVH;�/H;t�G;8�G;�WG;>�F;�
E;�B;p�<;��3;]%;��;> �:�3�:年95�D�����D^�G��n?ػ3,�� �x�6�Y6H�z5S�      ����-��#Ȥ�d���ݫ���f�G�=����
�ܻ�*��?o5�u����P(7E�}:�m�:��;>&;��4;B�=;�B;+�E;S�F;ˀG;$�G;cH;�@H;�dH;d�H;��H;x�H;��H;��H;;�H;��H;��H;��H;l�H;��H;��H;��H;;�H;��H;��H;x�H;��H;d�H;�dH;�@H;cH;$�G;ˀG;S�F;+�E;�B;B�=;��4;>&;��;�m�:E�}:�P(7u���?o5��*��
�ܻ���G�=��f�ݫ��d���#Ȥ��-��      xc��8�|����켔�Ҽg���`�����r�E:�%,�$ߵ�Z/X���º̬�E�}:> �:v;��);�l7;i�?;�C;KF;�(G;E�G;�G;2)H;�RH;�sH;��H;��H;�H;ͼH;��H;��H;+�H;��H;l�H;��H;+�H;��H;��H;ͼH;�H;��H;��H;�sH;�RH;2)H;�G;E�G;�(G;KF;�C;i�?;�l7;��);v;> �:E�}:̬���ºZ/X�$ߵ�%,�E:���r�`���g�����Ҽ��|����8�      �&K���G�ȟ>��0�:y�vc�d��)������!�V����ƻgod���º�P(7�3�:���:�;]P.;9�:;ayA;y�D;�F;�mG;t�G;!H;�?H;MeH;��H;R�H;ժH;��H;�H;	�H;��H;��H;V�H;��H;��H;	�H;�H;��H;ժH;R�H;��H;MeH;�?H;!H;t�G;�mG;�F;y�D;ayA;9�:;]P.;�;���:�3�:�P(7��ºgod��ƻ��!�V����)���d��vc�:y��0�ȟ>���G�      鰒�Z��������}��c���D�/%��8���Ҽ	c����f�����ƻZ/X�u���年9f�:ȏ;F";�3;�>;�XC;��E;G;'�G;��G;�+H;/VH;9wH;��H;W�H;�H;.�H;�H;Q�H;`�H;N�H;`�H;Q�H;�H;.�H;�H;W�H;��H;9wH;/VH;�+H;��G;'�G;G;��E;�XC;�>;�3;F";ȏ;f�:年9u���Z/X��ƻ�����f�	c����Ҽ�8�/%���D��c���}�����Z��      \Pν��ʽ*8�������������0�f�u�;���K��Ȥ���f���$ߵ�?o5�5�D�L�-:���:X>;G+;_9;�A;��D;[�F;�uG;�G;IH;�FH;�kH;�H;��H;�H;H�H;�H;��H;"�H;F�H;"�H;��H;�H;H�H;�H;��H;�H;�kH;�FH;IH;�G;�uG;[�F;��D;�A;_9;G+;X>;���:L�-:5�D�?o5�$ߵ�����f�Ȥ�K����u�;�0�f������������*8����ʽ      ���N9�C[��s�R�ؽ���s����}���G��K��	c��!�V�%,��*�����+����:?��:� ;ǂ3;0>;�C;"F;#8G;l�G;�H;7H;�_H;,H;�H; �H;g�H;�H;m�H;��H;3�H;��H;m�H;�H;g�H; �H;�H;,H;�_H;7H;�H;l�G;#8G;"F;�C;0>;ǂ3;� ;?��:��:+������*��%,�!�V�	c��K�����G���}��s����R�ؽ�s�C[�N9�      }�=���:���0��Q"�e�����ZPν�榽%����G�����Ҽ���E:�
�ܻ�D^�ϸ��ih:���:O;�{,;�:;��A;~hE;��F;\�G;��G;�'H;eTH;�vH;��H;L�H;��H;�H;��H;��H;3�H;��H;��H;�H;��H;L�H;��H;�vH;eTH;�'H;��G;\�G;��F;~hE;��A;�:;�{,;O;���:ih:ϸ���D^�
�ܻE:������Ҽ����G�%���榽ZPν����e��Q"���0���:�      
Dx��s���f�QS���:����B[��7ս�榽��}�u�;��8�)�����r����G������Ҭ����:��;}$;,�6;f�?;3�D;�F;�oG;��G;H;XIH;dnH;i�H;��H;�H;Z�H;��H;��H;G�H;��H;��H;Z�H;�H;��H;i�H;dnH;XIH;H;��G;�oG;�F;3�D;f�?;,�6;}$;��;���:�Ҭ����G�������r�)����8�u�;���}��榽�7սB[������:�QS���f��s�      �*���0��ȥ��&���jk��H��#%�B[�ZPν�s��0�f�/%�d��`���G�=�n?ػgFL��D�`�R:B�:��;�2;�=;��C;�/F;�FG;�G;WH;?H;�fH;��H;V�H;ͫH;��H;��H;�H;��H;�H;��H;��H;ͫH;V�H;��H;�fH;?H;WH;�G;�FG;�/F;��C;�=;�2;��;B�:`�R:�D�gFL�n?ػG�=�`���d��/%�0�f��s��ZPνB[��#%��H�jk�&���ȥ���0��      �þ��������R��f쏾�s��H����������������D�vc�g����f�3,�����P����9/��:5;�i-;��;;��B;+�E;�G;��G;��G;�5H;�_H;�H;{�H;�H;q�H;ɽH;r�H;��H;r�H;ɽH;q�H;�H;{�H;�H;�_H;�5H;��G;��G;�G;+�E;��B;��;;�i-;5;/��:��9�P�����3,��f�g���vc���D���������������H��s�f쏾�R���������      ����fYؾ�þ�ê�f쏾jk���:�e�R�ؽ�����c�:y���Ҽݫ��� �B�(���'7��:�
;c�(;�^9;��A;�[E;��F;�G;��G;�-H;�YH;{H;�H;i�H;u�H;6�H;�H;��H;�H;6�H;u�H;i�H;�H;{H;�YH;�-H;��G;�G;��F;�[E;��A;�^9;c�(;�
;��:�'7(��B�� �ݫ����Ҽ:y��c�����R�ؽe���:�jk�f쏾�ê��þfYؾ��      ��=������I��þ�R��&���QS��Q"��s�����}��0���d���x�6��ƻ(}*����^�:�w;�%;Rl7;�@;�D;�F;��G;��G;3'H;UH;�wH;�H;f�H;±H;ۺH;�H;��H;�H;ۺH;±H;f�H;�H;�wH;UH;3'H;��G;��G;�F;�D;�@;Rl7;�%;�w;^�:���(}*��ƻx�6�d����켟0���}�����s��Q"�QS�&����R���þIᾁ���=��      ���>��&�
�����fYؾ���ȥ����f���0�C[�*8������ȟ>�|���#Ȥ�Y6H�,�ܻ�qF�0��4�}:���:�";��5;6�?;��D;��F;/�G;��G;s"H;�QH;�tH;y�H;�H;��H;�H;�H;��H;�H;�H;��H;�H;y�H;�tH;�QH;s"H;��G;/�G;��F;��D;6�?;��5;�";���:4�}:0���qF�,�ܻY6H�#Ȥ�|���ȟ>�����*8��C[���0���f�ȥ�����fYؾ����&�
�>��      �� �k��>��=���������0���s���:�N9���ʽZ����G��8��-��z5S�w���/X���D��Ad:�A�:� ;x�4;	�?;#~D;p�F;3xG;��G;�H;NOH;HsH;:�H;�H;�H;W�H;��H;U�H;��H;W�H;�H;�H;:�H;HsH;NOH;�H;��G;3xG;p�F;#~D;	�?;x�4;� ;�A�:�Ad:��D��/X�w��z5S��-���8���G�Z����ʽN9���:��s��0��������=��>��k��      .Eb�I]�tN�ߛ7����e� �{�˾��	�j��!,�J���0��m���,˼��x�E���1��a���Q�:e�:2;��1;n+>;��C;�vF;�G;��G;>H;�gH;Z�H;v�H;8�H;�H;��H;(�H;��H;(�H;��H;�H;8�H;v�H;Z�H;�gH;>H;��G;�G;�vF;��C;n+>;��1;2;e�:Q�:a����1��E����x�,˼��m�0��J����!,�	�j���{�˾e� ����ߛ7�tN�I]�      I]�N�W��TI�v3��D�������Ǿb���ȟf� )� ��W;���Fi��k�x�Ǽ�[t�8�	�(Ȅ�tX��Ο:���:%�;�I2;�Y>;qD;�~F;\�G;+H;�>H;�hH;�H;�H;q�H;7�H;��H;S�H;��H;S�H;��H;7�H;q�H;�H;�H;�hH;�>H;+H;\�G;�~F;qD;�Y>;�I2;%�;���:Ο:tX��(Ȅ�8�	��[t�x�Ǽ�k��Fi�W;�� �� )�ȟf�b�����Ǿ�����D�v3��TI�N�W�      tN��TI���;��'��k���i���f󐾖Z��K ��s�&����&^����"����g����Ѩu�R!���1<:��:n
;�f3;-�>;�AD;ՕF;�G;�H;UAH;jH;\�H;ߟH;(�H;ԻH;k�H;��H;B�H;��H;k�H;ԻH;(�H;ߟH;\�H;jH;UAH;�H;�G;ՕF;�AD;-�>;�f3;n
;��:�1<:R!��Ѩu������g��"�����&^�&����s潎K ��Z�f�i������k��'���;��TI�      ߛ7�v3��'����e� ��{Ծ
���6���]�F�����ӽ���;�L�1v�x뮼-T�ǘ��PV�q�=�1(i:_��:!z ;�#5;�?;2�D;�F;�G;�H;�EH;�mH;��H;}�H;j�H;ۼH;4�H;O�H;��H;O�H;4�H;ۼH;j�H;}�H;��H;�mH;�EH;�H;�G;�F;2�D;�?;�#5;!z ;_��:1(i:q�=��PV�ǘ�-T�x뮼1v�;�L�����ӽ���]�F�6���
����{Ծe� �����'�v3�      ����D��k�e� �<�ݾS���C͓�ȟf��>/�x��~'��n섽/�6�Rt��v��?�:�Tʻ�.�ݷ��s�:1; �$;�X7;��@;	E;:�F;P�G;�H;EKH;�qH;��H;ɣH;�H;�H;.�H;D�H;��H;D�H;.�H;�H;�H;ɣH;��H;�qH;EKH;�H;P�G;:�F;	E;��@;�X7; �$;1;�s�:ݷ��.�Tʻ?�:��v��Rt�/�6�n섽~'��x���>/�ȟf�C͓�S���<�ݾe� ��k��D�      e� ������쾻{ԾS���b���9�x�rSC��^�ͻ޽%���Q�e����ѼG������R�����դ8��:�X;��);5�9;-�A;��E;�G;2�G;s H;DRH;�vH;v�H;��H;:�H;��H;r�H;u�H;��H;u�H;r�H;��H;:�H;��H;v�H;�vH;DRH;s H;2�G;�G;��E;-�A;5�9;��);�X;��:դ8����R�����G���Ѽ��Q�e�%���ͻ޽�^�rSC�9�x�b���S����{Ծ�쾃���      {�˾��Ǿi���
���C͓�9�x�ؘJ��K �H��� �������?���t뮼�[�����3|��W��<�:u~�:';�
/;�f<;�C;� F;�MG;��G;9,H;sZH;�|H;ǖH;©H;��H;��H;��H;��H;��H;��H;��H;��H;��H;©H;ǖH;�|H;sZH;9,H;��G;�MG;� F;�C;�f<;�
/;';u~�:<�:�W��3|������[�t뮼����?���� ��H����K �ؘJ�9�x�C͓�
���i�����Ǿ      ��b���f�6���ȟf�rSC��K �Gn����Ž����Z��k��|ռX��Ey-����x.�y���O�:�*�:��;o4;s�>;)D;�vF;I�G;��G;�8H;\cH;x�H;��H;[�H;e�H;��H;��H;K�H;f�H;K�H;��H;��H;e�H;[�H;��H;x�H;\cH;�8H;��G;I�G;�vF;)D;s�>;o4;��;�*�:�O�:y��x.����Ey-�X���|ռ�k��Z������ŽGn���K �rSC�ȟf�6���f�b���      	�j�ȟf��Z�]�F��>/��^�H�����Ž- ���Fi�kQ+�Ot�PT��H�W�����1��jȺ�U�9�O�:	Y;��(;T�8;1A;�E;!�F;|�G;�H;�EH;�lH;��H;��H;8�H;d�H;��H;��H;��H;��H;��H;��H;��H;d�H;8�H;��H;��H;�lH;�EH;�H;|�G;!�F;�E;1A;T�8;��(;	Y;�O�:�U�9jȺ�1�����H�W�PT��Ot�kQ+��Fi�- ����ŽH����^��>/�]�F��Z�ȟf�      �!,� )��K ����x��ͻ޽ ������Fi���0�����跼z�x�����.��b�(�����)i:���:��;�0;��<;�C;��E;)<G;
�G;�#H;jSH;�vH;�H;�H;E�H;t�H;4�H;��H;��H;n�H;��H;��H;4�H;t�H;E�H;�H;�H;�vH;jSH;�#H;
�G;)<G;��E;�C;��<;�0;��;���:�)i:���b�(��.�����z�x��跼�����0��Fi���� ��ͻ޽x������K � )�      J��� ��s��ӽ~'��%�������Z�kQ+�����"��G����0���׻͕b��W���V�9�:�_;�)';/Y7;G#@;S�D;�F;+�G;��G;@7H;aH;��H;Z�H;��H;l�H;��H;��H;{�H;A�H;.�H;A�H;{�H;��H;��H;l�H;��H;Z�H;��H;aH;@7H;��G;+�G;�F;S�D;G#@;/Y7;�)';�_;�:�V�9�W��͕b���׻��0�G���"�����kQ+��Z����%���~'���ӽ�s� ��      0��W;��&������n섽Q�e���?��k�Ot��跼G��ee7�����Ǆ��0�?�t�^t�:�*�:�
;�1;��<;��B;N�E;G;�G;iH;wIH;`nH;��H;��H;�H;��H;��H;�H;��H;�H;��H;�H;��H;�H;��H;��H;�H;��H;��H;`nH;wIH;iH;�G;G;N�E;��B;��<;�1;�
;�*�:^t�:?�t��0��Ǆ����ee7�G���跼Ot�k���?�Q�e�n섽���&���W;��      m��Fi��&^�;�L�/�6������|ռPT��z�x���0��������1���ڷ�xm`:��:��;��*;}�8;G�@;d�D;��F;}G;��G;�0H;�ZH;m{H;��H;֧H;�H;��H;��H;|�H;��H;��H;d�H;��H;��H;|�H;��H;��H;�H;֧H;��H;m{H;�ZH;�0H;��G;}G;��F;d�D;G�@;}�8;��*;��;��:xm`:�ڷ�1��������껣�0�z�x�PT���|ռ����/�6�;�L��&^��Fi�      ���k���1v�Rt��Ѽt뮼X��H�W������׻�Ǆ�1�����3<:v��:;Y;�s%;<$5;�Y>;-`C;��E;O)G;u�G;"H;GH;lkH;�H;��H;��H;ȻH;��H;��H;��H;g�H;^�H;�H;^�H;g�H;��H;��H;��H;ȻH;��H;��H;�H;lkH;GH;"H;u�G;O)G;��E;-`C;�Y>;<$5;�s%;;Y;v��:�3<:���1���Ǆ���׻���H�W�X��t뮼�ѼRt�1v����k�      ,˼x�Ǽ�"��x뮼�v��G���[�Ey-�����.��͕b��0㺉ڷ��3<:L�:_\;��!;1J2;�f<;/B;QBE;J�F;a�G; �G;�3H;�[H;{H;��H;��H;P�H;��H;5�H;��H;B�H;A�H;��H;��H;��H;A�H;B�H;��H;5�H;��H;P�H;��H;��H;{H;�[H;�3H; �G;a�G;J�F;QBE;/B;�f<;1J2;��!;_\;L�:�3<:�ڷ��0�͕b��.�����Ey-��[�G���v��x뮼�"��x�Ǽ      ��x��[t���g�-T�?�:������������1��b�(��W��?�t�xm`:v��:_\;pz ;�0;�;;9<A;?�D;�vF;�bG;d�G;� H;�LH;�nH;o�H;~�H;��H;��H;Z�H;��H;H�H;_�H;��H;��H;�H;��H;��H;_�H;H�H;��H;Z�H;��H;��H;~�H;o�H;�nH;�LH;� H;d�G;�bG;�vF;?�D;9<A;�;;�0;pz ;_\;v��:xm`:?�t��W��b�(��1������������?�:�-T���g��[t�      E��8�	����ǘ�Tʻ�R��3|�x.�jȺ����V�9^t�:��:;Y;��!;�0;-�:;�@;4BD;�1F;�7G;��G;�H;k?H;*cH;�H;m�H;:�H;<�H;>�H;��H;��H;��H;[�H;��H;��H;s�H;��H;��H;[�H;��H;��H;��H;>�H;<�H;:�H;m�H;�H;*cH;k?H;�H;��G;�7G;�1F;4BD;�@;-�:;�0;��!;;Y;��:^t�:�V�9���jȺx.�3|��R��Tʻǘ����8�	�      �1��(Ȅ�Ѩu��PV��.�����W��y��U�9�)i:�:�*�:��;�s%;1J2;�;;�@;�D;/F;>G;��G;�H;�4H;�YH;5wH;7�H;�H;	�H;�H;H�H;^�H;�H;�H;�H;*�H;E�H;��H;E�H;*�H;�H;�H;�H;^�H;H�H;�H;	�H;�H;7�H;5wH;�YH;�4H;�H;��G;>G;/F;�D;�@;�;;1J2;�s%;��;�*�:�:�)i:�U�9y���W������.��PV�Ѩu�(Ȅ�      a���tX��R!��q�=�ݷ�դ8<�:�O�:�O�:���:�_;�
;��*;<$5;�f<;9<A;4BD;/F;�G;��G;q�G;�,H;RH;UpH;�H;��H;r�H;�H;)�H;��H;��H;��H;?�H;��H;��H;{�H;��H;{�H;��H;��H;?�H;��H;��H;��H;)�H;�H;r�H;��H;�H;UpH;RH;�,H;q�G;��G;�G;/F;4BD;9<A;�f<;<$5;��*;�
;�_;���:�O�:�O�:<�:դ8ݷ�q�=�R!��tX��      Q�:Ο:�1<:1(i:�s�:��:u~�:�*�:	Y;��;�)';�1;}�8;�Y>;/B;?�D;�1F;>G;��G;%�G;�(H;�MH;qkH;C�H;c�H;v�H;��H;�H;t�H;��H;$�H;�H;�H;D�H;��H;��H;��H;��H;��H;D�H;�H;�H;$�H;��H;t�H;�H;��H;v�H;c�H;C�H;qkH;�MH;�(H;%�G;��G;>G;�1F;?�D;/B;�Y>;}�8;�1;�)';��;	Y;�*�:u~�:��:�s�:1(i:�1<:Ο:      e�:���:��:_��:1;�X;';��;��(;�0;/Y7;��<;G�@;-`C;QBE;�vF;�7G;��G;q�G;�(H;�KH;�hH;.�H;O�H;��H;��H;��H;N�H;�H;��H;��H;A�H;��H;��H;��H;��H;��H;��H;��H;��H;��H;A�H;��H;��H;�H;N�H;��H;��H;��H;O�H;.�H;�hH;�KH;�(H;q�G;��G;�7G;�vF;QBE;-`C;G�@;��<;/Y7;�0;��(;��;';�X;1;_��:��:���:      2;%�;n
;!z ; �$;��);�
/;o4;T�8;��<;G#@;��B;d�D;��E;J�F;�bG;��G;�H;�,H;�MH;�hH;B�H;��H;��H;ΰH;��H;��H;��H;2�H;��H;^�H;�H;0�H;��H;��H;P�H;��H;P�H;��H;��H;0�H;�H;^�H;��H;2�H;��H;��H;��H;ΰH;��H;��H;B�H;�hH;�MH;�,H;�H;��G;�bG;J�F;��E;d�D;��B;G#@;��<;T�8;o4;�
/;��); �$;!z ;n
;%�;      ��1;�I2;�f3;�#5;�X7;5�9;�f<;s�>;1A;�C;S�D;N�E;��F;O)G;a�G;d�G;�H;�4H;RH;qkH;.�H;��H;�H;ɯH;�H;U�H;L�H; �H;��H;��H;u�H;��H;o�H;��H;��H;�H;\�H;�H;��H;��H;o�H;��H;u�H;��H;��H; �H;L�H;U�H;�H;ɯH;�H;��H;.�H;qkH;RH;�4H;�H;d�G;a�G;O)G;��F;N�E;S�D;�C;1A;s�>;�f<;5�9;�X7;�#5;�f3;�I2;      n+>;�Y>;-�>;�?;��@;-�A;�C;)D;�E;��E;�F;G;}G;u�G; �G;� H;k?H;�YH;UpH;C�H;O�H;��H;ɯH;�H;��H;��H;5�H;��H;��H;��H;O�H; �H;��H;��H;H�H;��H;��H;��H;H�H;��H;��H; �H;O�H;��H;��H;��H;5�H;��H;��H;�H;ɯH;��H;O�H;C�H;UpH;�YH;k?H;� H; �G;u�G;}G;G;�F;��E;�E;)D;�C;-�A;��@;�?;-�>;�Y>;      ��C;qD;�AD;2�D;	E;��E;� F;�vF;!�F;)<G;+�G;�G;��G;"H;�3H;�LH;*cH;5wH;�H;c�H;��H;ΰH;�H;��H;<�H;��H;��H;^�H;c�H;��H;��H;f�H;��H;?�H;��H;C�H;L�H;C�H;��H;?�H;��H;f�H;��H;��H;c�H;^�H;��H;��H;<�H;��H;�H;ΰH;��H;c�H;�H;5wH;*cH;�LH;�3H;"H;��G;�G;+�G;)<G;!�F;�vF;� F;��E;	E;2�D;�AD;qD;      �vF;�~F;ՕF;�F;:�F;�G;�MG;I�G;|�G;
�G;��G;iH;�0H;GH;�[H;�nH;�H;7�H;��H;v�H;��H;��H;U�H;��H;��H;W�H;$�H;�H;��H;��H;�H;S�H;6�H;��H;m�H;��H;��H;��H;m�H;��H;6�H;S�H;�H;��H;��H;�H;$�H;W�H;��H;��H;U�H;��H;��H;v�H;��H;7�H;�H;�nH;�[H;GH;�0H;iH;��G;
�G;|�G;I�G;�MG;�G;:�F;�F;ՕF;�~F;      �G;\�G;�G;�G;P�G;2�G;��G;��G;�H;�#H;@7H;wIH;�ZH;lkH;{H;o�H;m�H;�H;r�H;��H;��H;��H;L�H;5�H;��H;$�H;�H;h�H;J�H;��H;7�H;�H;��H;��H;��H;�H;�H;�H;��H;��H;��H;�H;7�H;��H;J�H;h�H;�H;$�H;��H;5�H;L�H;��H;��H;��H;r�H;�H;m�H;o�H;{H;lkH;�ZH;wIH;@7H;�#H;�H;��G;��G;2�G;P�G;�G;�G;\�G;      ��G;+H;�H;�H;�H;s H;9,H;�8H;�EH;jSH;aH;`nH;m{H;�H;��H;~�H;:�H;	�H;�H;�H;N�H;��H; �H;��H;^�H;�H;h�H;\�H;��H;�H;�H;��H;z�H;��H;�H;^�H;g�H;^�H;�H;��H;z�H;��H;�H;�H;��H;\�H;h�H;�H;^�H;��H; �H;��H;N�H;�H;�H;	�H;:�H;~�H;��H;�H;m{H;`nH;aH;jSH;�EH;�8H;9,H;s H;�H;�H;�H;+H;      >H;�>H;UAH;�EH;EKH;DRH;sZH;\cH;�lH;�vH;��H;��H;��H;��H;��H;��H;<�H;�H;)�H;t�H;�H;2�H;��H;��H;c�H;��H;J�H;��H;$�H;��H;��H;k�H;��H;5�H;p�H;��H;��H;��H;p�H;5�H;��H;k�H;��H;��H;$�H;��H;J�H;��H;c�H;��H;��H;2�H;�H;t�H;)�H;�H;<�H;��H;��H;��H;��H;��H;��H;�vH;�lH;\cH;sZH;DRH;EKH;�EH;UAH;�>H;      �gH;�hH;jH;�mH;�qH;�vH;�|H;x�H;��H;�H;Z�H;��H;֧H;��H;P�H;��H;>�H;H�H;��H;��H;��H;��H;��H;��H;��H;��H;��H;�H;��H;��H;t�H;��H;$�H;y�H;��H;��H;��H;��H;��H;y�H;$�H;��H;t�H;��H;��H;�H;��H;��H;��H;��H;��H;��H;��H;��H;��H;H�H;>�H;��H;P�H;��H;֧H;��H;Z�H;�H;��H;x�H;�|H;�vH;�qH;�mH;jH;�hH;      Z�H;�H;\�H;��H;��H;v�H;ǖH;��H;��H;�H;��H;�H;�H;ȻH;��H;Z�H;��H;^�H;��H;$�H;��H;^�H;u�H;O�H;��H;�H;7�H;�H;��H;t�H;��H;.�H;��H;��H;��H;��H;��H;��H;��H;��H;��H;.�H;��H;t�H;��H;�H;7�H;�H;��H;O�H;u�H;^�H;��H;$�H;��H;^�H;��H;Z�H;��H;ȻH;�H;�H;��H;�H;��H;��H;ǖH;v�H;��H;��H;\�H;�H;      v�H;�H;ߟH;}�H;ɣH;��H;©H;[�H;8�H;E�H;l�H;��H;��H;��H;5�H;��H;��H;�H;��H;�H;A�H;�H;��H; �H;f�H;S�H;�H;��H;k�H;��H;.�H;z�H;��H;��H;��H;�H;�H;�H;��H;��H;��H;z�H;.�H;��H;k�H;��H;�H;S�H;f�H; �H;��H;�H;A�H;�H;��H;�H;��H;��H;5�H;��H;��H;��H;l�H;E�H;8�H;[�H;©H;��H;ɣH;}�H;ߟH;�H;      8�H;q�H;(�H;j�H;�H;:�H;��H;e�H;d�H;t�H;��H;��H;��H;��H;��H;H�H;��H;�H;?�H;�H;��H;0�H;o�H;��H;��H;6�H;��H;z�H;��H;$�H;��H;��H;��H;��H;�H;�H;�H;�H;�H;��H;��H;��H;��H;$�H;��H;z�H;��H;6�H;��H;��H;o�H;0�H;��H;�H;?�H;�H;��H;H�H;��H;��H;��H;��H;��H;t�H;d�H;e�H;��H;:�H;�H;j�H;(�H;q�H;      �H;7�H;ԻH;ۼH;�H;��H;��H;��H;��H;4�H;��H;�H;|�H;��H;B�H;_�H;[�H;�H;��H;D�H;��H;��H;��H;��H;?�H;��H;��H;��H;5�H;y�H;��H;��H;��H; �H;-�H;8�H;�H;8�H;-�H; �H;��H;��H;��H;y�H;5�H;��H;��H;��H;?�H;��H;��H;��H;��H;D�H;��H;�H;[�H;_�H;B�H;��H;|�H;�H;��H;4�H;��H;��H;��H;��H;�H;ۼH;ԻH;7�H;      ��H;��H;k�H;4�H;.�H;r�H;��H;��H;��H;��H;{�H;��H;��H;g�H;A�H;��H;��H;*�H;��H;��H;��H;��H;��H;H�H;��H;m�H;��H;�H;p�H;��H;��H;��H;�H;-�H;�H;-�H;J�H;-�H;�H;-�H;�H;��H;��H;��H;p�H;�H;��H;m�H;��H;H�H;��H;��H;��H;��H;��H;*�H;��H;��H;A�H;g�H;��H;��H;{�H;��H;��H;��H;��H;r�H;.�H;4�H;k�H;��H;      (�H;S�H;��H;O�H;D�H;u�H;��H;K�H;��H;��H;A�H;�H;��H;^�H;��H;��H;��H;E�H;{�H;��H;��H;P�H;�H;��H;C�H;��H;�H;^�H;��H;��H;��H;�H;�H;8�H;-�H;$�H;6�H;$�H;-�H;8�H;�H;�H;��H;��H;��H;^�H;�H;��H;C�H;��H;�H;P�H;��H;��H;{�H;E�H;��H;��H;��H;^�H;��H;�H;A�H;��H;��H;K�H;��H;u�H;D�H;O�H;��H;S�H;      ��H;��H;B�H;��H;��H;��H;��H;f�H;��H;n�H;.�H;��H;d�H;�H;��H;�H;s�H;��H;��H;��H;��H;��H;\�H;��H;L�H;��H;�H;g�H;��H;��H;��H;�H;�H;�H;J�H;6�H;#�H;6�H;J�H;�H;�H;�H;��H;��H;��H;g�H;�H;��H;L�H;��H;\�H;��H;��H;��H;��H;��H;s�H;�H;��H;�H;d�H;��H;.�H;n�H;��H;f�H;��H;��H;��H;��H;B�H;��H;      (�H;S�H;��H;O�H;D�H;u�H;��H;K�H;��H;��H;A�H;�H;��H;^�H;��H;��H;��H;E�H;{�H;��H;��H;P�H;�H;��H;C�H;��H;�H;^�H;��H;��H;��H;�H;�H;8�H;-�H;$�H;6�H;$�H;-�H;8�H;�H;�H;��H;��H;��H;^�H;�H;��H;C�H;��H;�H;P�H;��H;��H;{�H;E�H;��H;��H;��H;^�H;��H;�H;A�H;��H;��H;K�H;��H;u�H;D�H;O�H;��H;S�H;      ��H;��H;k�H;4�H;.�H;r�H;��H;��H;��H;��H;{�H;��H;��H;g�H;A�H;��H;��H;*�H;��H;��H;��H;��H;��H;H�H;��H;m�H;��H;�H;p�H;��H;��H;��H;�H;-�H;�H;-�H;J�H;-�H;�H;-�H;�H;��H;��H;��H;p�H;�H;��H;m�H;��H;H�H;��H;��H;��H;��H;��H;*�H;��H;��H;A�H;g�H;��H;��H;{�H;��H;��H;��H;��H;r�H;.�H;4�H;k�H;��H;      �H;7�H;ԻH;ۼH;�H;��H;��H;��H;��H;4�H;��H;�H;|�H;��H;B�H;_�H;[�H;�H;��H;D�H;��H;��H;��H;��H;?�H;��H;��H;��H;5�H;y�H;��H;��H;��H; �H;-�H;8�H;�H;8�H;-�H; �H;��H;��H;��H;y�H;5�H;��H;��H;��H;?�H;��H;��H;��H;��H;D�H;��H;�H;[�H;_�H;B�H;��H;|�H;�H;��H;4�H;��H;��H;��H;��H;�H;ۼH;ԻH;7�H;      8�H;q�H;(�H;j�H;�H;:�H;��H;e�H;d�H;t�H;��H;��H;��H;��H;��H;H�H;��H;�H;?�H;�H;��H;0�H;o�H;��H;��H;6�H;��H;z�H;��H;$�H;��H;��H;��H;��H;�H;�H;�H;�H;�H;��H;��H;��H;��H;$�H;��H;z�H;��H;6�H;��H;��H;o�H;0�H;��H;�H;?�H;�H;��H;H�H;��H;��H;��H;��H;��H;t�H;d�H;e�H;��H;:�H;�H;j�H;(�H;q�H;      v�H;�H;ߟH;}�H;ɣH;��H;©H;[�H;8�H;E�H;l�H;��H;��H;��H;5�H;��H;��H;�H;��H;�H;A�H;�H;��H; �H;f�H;S�H;�H;��H;k�H;��H;.�H;z�H;��H;��H;��H;�H;�H;�H;��H;��H;��H;z�H;.�H;��H;k�H;��H;�H;S�H;f�H; �H;��H;�H;A�H;�H;��H;�H;��H;��H;5�H;��H;��H;��H;l�H;E�H;8�H;[�H;©H;��H;ɣH;}�H;ߟH;�H;      Z�H;�H;\�H;��H;��H;v�H;ǖH;��H;��H;�H;��H;�H;�H;ȻH;��H;Z�H;��H;^�H;��H;$�H;��H;^�H;u�H;O�H;��H;�H;7�H;�H;��H;t�H;��H;.�H;��H;��H;��H;��H;��H;��H;��H;��H;��H;.�H;��H;t�H;��H;�H;7�H;�H;��H;O�H;u�H;^�H;��H;$�H;��H;^�H;��H;Z�H;��H;ȻH;�H;�H;��H;�H;��H;��H;ǖH;v�H;��H;��H;\�H;�H;      �gH;�hH;jH;�mH;�qH;�vH;�|H;x�H;��H;�H;Z�H;��H;֧H;��H;P�H;��H;>�H;H�H;��H;��H;��H;��H;��H;��H;��H;��H;��H;�H;��H;��H;t�H;��H;$�H;y�H;��H;��H;��H;��H;��H;y�H;$�H;��H;t�H;��H;��H;�H;��H;��H;��H;��H;��H;��H;��H;��H;��H;H�H;>�H;��H;P�H;��H;֧H;��H;Z�H;�H;��H;x�H;�|H;�vH;�qH;�mH;jH;�hH;      >H;�>H;UAH;�EH;EKH;DRH;sZH;\cH;�lH;�vH;��H;��H;��H;��H;��H;��H;<�H;�H;)�H;t�H;�H;2�H;��H;��H;c�H;��H;J�H;��H;$�H;��H;��H;k�H;��H;5�H;p�H;��H;��H;��H;p�H;5�H;��H;k�H;��H;��H;$�H;��H;J�H;��H;c�H;��H;��H;2�H;�H;t�H;)�H;�H;<�H;��H;��H;��H;��H;��H;��H;�vH;�lH;\cH;sZH;DRH;EKH;�EH;UAH;�>H;      ��G;+H;�H;�H;�H;s H;9,H;�8H;�EH;jSH;aH;`nH;m{H;�H;��H;~�H;:�H;	�H;�H;�H;N�H;��H; �H;��H;^�H;�H;h�H;\�H;��H;�H;�H;��H;z�H;��H;�H;^�H;g�H;^�H;�H;��H;z�H;��H;�H;�H;��H;\�H;h�H;�H;^�H;��H; �H;��H;N�H;�H;�H;	�H;:�H;~�H;��H;�H;m{H;`nH;aH;jSH;�EH;�8H;9,H;s H;�H;�H;�H;+H;      �G;\�G;�G;�G;P�G;2�G;��G;��G;�H;�#H;@7H;wIH;�ZH;lkH;{H;o�H;m�H;�H;r�H;��H;��H;��H;L�H;5�H;��H;$�H;�H;h�H;J�H;��H;7�H;�H;��H;��H;��H;�H;�H;�H;��H;��H;��H;�H;7�H;��H;J�H;h�H;�H;$�H;��H;5�H;L�H;��H;��H;��H;r�H;�H;m�H;o�H;{H;lkH;�ZH;wIH;@7H;�#H;�H;��G;��G;2�G;P�G;�G;�G;\�G;      �vF;�~F;ՕF;�F;:�F;�G;�MG;I�G;|�G;
�G;��G;iH;�0H;GH;�[H;�nH;�H;7�H;��H;v�H;��H;��H;U�H;��H;��H;W�H;$�H;�H;��H;��H;�H;S�H;6�H;��H;m�H;��H;��H;��H;m�H;��H;6�H;S�H;�H;��H;��H;�H;$�H;W�H;��H;��H;U�H;��H;��H;v�H;��H;7�H;�H;�nH;�[H;GH;�0H;iH;��G;
�G;|�G;I�G;�MG;�G;:�F;�F;ՕF;�~F;      ��C;qD;�AD;2�D;	E;��E;� F;�vF;!�F;)<G;+�G;�G;��G;"H;�3H;�LH;*cH;5wH;�H;c�H;��H;ΰH;�H;��H;<�H;��H;��H;^�H;c�H;��H;��H;f�H;��H;?�H;��H;C�H;L�H;C�H;��H;?�H;��H;f�H;��H;��H;c�H;^�H;��H;��H;<�H;��H;�H;ΰH;��H;c�H;�H;5wH;*cH;�LH;�3H;"H;��G;�G;+�G;)<G;!�F;�vF;� F;��E;	E;2�D;�AD;qD;      n+>;�Y>;-�>;�?;��@;-�A;�C;)D;�E;��E;�F;G;}G;u�G; �G;� H;k?H;�YH;UpH;C�H;O�H;��H;ɯH;�H;��H;��H;5�H;��H;��H;��H;O�H; �H;��H;��H;H�H;��H;��H;��H;H�H;��H;��H; �H;O�H;��H;��H;��H;5�H;��H;��H;�H;ɯH;��H;O�H;C�H;UpH;�YH;k?H;� H; �G;u�G;}G;G;�F;��E;�E;)D;�C;-�A;��@;�?;-�>;�Y>;      ��1;�I2;�f3;�#5;�X7;5�9;�f<;s�>;1A;�C;S�D;N�E;��F;O)G;a�G;d�G;�H;�4H;RH;qkH;.�H;��H;�H;ɯH;�H;U�H;L�H; �H;��H;��H;u�H;��H;o�H;��H;��H;�H;\�H;�H;��H;��H;o�H;��H;u�H;��H;��H; �H;L�H;U�H;�H;ɯH;�H;��H;.�H;qkH;RH;�4H;�H;d�G;a�G;O)G;��F;N�E;S�D;�C;1A;s�>;�f<;5�9;�X7;�#5;�f3;�I2;      2;%�;n
;!z ; �$;��);�
/;o4;T�8;��<;G#@;��B;d�D;��E;J�F;�bG;��G;�H;�,H;�MH;�hH;B�H;��H;��H;ΰH;��H;��H;��H;2�H;��H;^�H;�H;0�H;��H;��H;P�H;��H;P�H;��H;��H;0�H;�H;^�H;��H;2�H;��H;��H;��H;ΰH;��H;��H;B�H;�hH;�MH;�,H;�H;��G;�bG;J�F;��E;d�D;��B;G#@;��<;T�8;o4;�
/;��); �$;!z ;n
;%�;      e�:���:��:_��:1;�X;';��;��(;�0;/Y7;��<;G�@;-`C;QBE;�vF;�7G;��G;q�G;�(H;�KH;�hH;.�H;O�H;��H;��H;��H;N�H;�H;��H;��H;A�H;��H;��H;��H;��H;��H;��H;��H;��H;��H;A�H;��H;��H;�H;N�H;��H;��H;��H;O�H;.�H;�hH;�KH;�(H;q�G;��G;�7G;�vF;QBE;-`C;G�@;��<;/Y7;�0;��(;��;';�X;1;_��:��:���:      Q�:Ο:�1<:1(i:�s�:��:u~�:�*�:	Y;��;�)';�1;}�8;�Y>;/B;?�D;�1F;>G;��G;%�G;�(H;�MH;qkH;C�H;c�H;v�H;��H;�H;t�H;��H;$�H;�H;�H;D�H;��H;��H;��H;��H;��H;D�H;�H;�H;$�H;��H;t�H;�H;��H;v�H;c�H;C�H;qkH;�MH;�(H;%�G;��G;>G;�1F;?�D;/B;�Y>;}�8;�1;�)';��;	Y;�*�:u~�:��:�s�:1(i:�1<:Ο:      a���tX��R!��q�=�ݷ�դ8<�:�O�:�O�:���:�_;�
;��*;<$5;�f<;9<A;4BD;/F;�G;��G;q�G;�,H;RH;UpH;�H;��H;r�H;�H;)�H;��H;��H;��H;?�H;��H;��H;{�H;��H;{�H;��H;��H;?�H;��H;��H;��H;)�H;�H;r�H;��H;�H;UpH;RH;�,H;q�G;��G;�G;/F;4BD;9<A;�f<;<$5;��*;�
;�_;���:�O�:�O�:<�:դ8ݷ�q�=�R!��tX��      �1��(Ȅ�Ѩu��PV��.�����W��y��U�9�)i:�:�*�:��;�s%;1J2;�;;�@;�D;/F;>G;��G;�H;�4H;�YH;5wH;7�H;�H;	�H;�H;H�H;^�H;�H;�H;�H;*�H;E�H;��H;E�H;*�H;�H;�H;�H;^�H;H�H;�H;	�H;�H;7�H;5wH;�YH;�4H;�H;��G;>G;/F;�D;�@;�;;1J2;�s%;��;�*�:�:�)i:�U�9y���W������.��PV�Ѩu�(Ȅ�      E��8�	����ǘ�Tʻ�R��3|�x.�jȺ����V�9^t�:��:;Y;��!;�0;-�:;�@;4BD;�1F;�7G;��G;�H;k?H;*cH;�H;m�H;:�H;<�H;>�H;��H;��H;��H;[�H;��H;��H;s�H;��H;��H;[�H;��H;��H;��H;>�H;<�H;:�H;m�H;�H;*cH;k?H;�H;��G;�7G;�1F;4BD;�@;-�:;�0;��!;;Y;��:^t�:�V�9���jȺx.�3|��R��Tʻǘ����8�	�      ��x��[t���g�-T�?�:������������1��b�(��W��?�t�xm`:v��:_\;pz ;�0;�;;9<A;?�D;�vF;�bG;d�G;� H;�LH;�nH;o�H;~�H;��H;��H;Z�H;��H;H�H;_�H;��H;��H;�H;��H;��H;_�H;H�H;��H;Z�H;��H;��H;~�H;o�H;�nH;�LH;� H;d�G;�bG;�vF;?�D;9<A;�;;�0;pz ;_\;v��:xm`:?�t��W��b�(��1������������?�:�-T���g��[t�      ,˼x�Ǽ�"��x뮼�v��G���[�Ey-�����.��͕b��0㺉ڷ��3<:L�:_\;��!;1J2;�f<;/B;QBE;J�F;a�G; �G;�3H;�[H;{H;��H;��H;P�H;��H;5�H;��H;B�H;A�H;��H;��H;��H;A�H;B�H;��H;5�H;��H;P�H;��H;��H;{H;�[H;�3H; �G;a�G;J�F;QBE;/B;�f<;1J2;��!;_\;L�:�3<:�ڷ��0�͕b��.�����Ey-��[�G���v��x뮼�"��x�Ǽ      ���k���1v�Rt��Ѽt뮼X��H�W������׻�Ǆ�1�����3<:v��:;Y;�s%;<$5;�Y>;-`C;��E;O)G;u�G;"H;GH;lkH;�H;��H;��H;ȻH;��H;��H;��H;g�H;^�H;�H;^�H;g�H;��H;��H;��H;ȻH;��H;��H;�H;lkH;GH;"H;u�G;O)G;��E;-`C;�Y>;<$5;�s%;;Y;v��:�3<:���1���Ǆ���׻���H�W�X��t뮼�ѼRt�1v����k�      m��Fi��&^�;�L�/�6������|ռPT��z�x���0��������1���ڷ�xm`:��:��;��*;}�8;G�@;d�D;��F;}G;��G;�0H;�ZH;m{H;��H;֧H;�H;��H;��H;|�H;��H;��H;d�H;��H;��H;|�H;��H;��H;�H;֧H;��H;m{H;�ZH;�0H;��G;}G;��F;d�D;G�@;}�8;��*;��;��:xm`:�ڷ�1��������껣�0�z�x�PT���|ռ����/�6�;�L��&^��Fi�      0��W;��&������n섽Q�e���?��k�Ot��跼G��ee7�����Ǆ��0�?�t�^t�:�*�:�
;�1;��<;��B;N�E;G;�G;iH;wIH;`nH;��H;��H;�H;��H;��H;�H;��H;�H;��H;�H;��H;�H;��H;��H;�H;��H;��H;`nH;wIH;iH;�G;G;N�E;��B;��<;�1;�
;�*�:^t�:?�t��0��Ǆ����ee7�G���跼Ot�k���?�Q�e�n섽���&���W;��      J��� ��s��ӽ~'��%�������Z�kQ+�����"��G����0���׻͕b��W���V�9�:�_;�)';/Y7;G#@;S�D;�F;+�G;��G;@7H;aH;��H;Z�H;��H;l�H;��H;��H;{�H;A�H;.�H;A�H;{�H;��H;��H;l�H;��H;Z�H;��H;aH;@7H;��G;+�G;�F;S�D;G#@;/Y7;�)';�_;�:�V�9�W��͕b���׻��0�G���"�����kQ+��Z����%���~'���ӽ�s� ��      �!,� )��K ����x��ͻ޽ ������Fi���0�����跼z�x�����.��b�(�����)i:���:��;�0;��<;�C;��E;)<G;
�G;�#H;jSH;�vH;�H;�H;E�H;t�H;4�H;��H;��H;n�H;��H;��H;4�H;t�H;E�H;�H;�H;�vH;jSH;�#H;
�G;)<G;��E;�C;��<;�0;��;���:�)i:���b�(��.�����z�x��跼�����0��Fi���� ��ͻ޽x������K � )�      	�j�ȟf��Z�]�F��>/��^�H�����Ž- ���Fi�kQ+�Ot�PT��H�W�����1��jȺ�U�9�O�:	Y;��(;T�8;1A;�E;!�F;|�G;�H;�EH;�lH;��H;��H;8�H;d�H;��H;��H;��H;��H;��H;��H;��H;d�H;8�H;��H;��H;�lH;�EH;�H;|�G;!�F;�E;1A;T�8;��(;	Y;�O�:�U�9jȺ�1�����H�W�PT��Ot�kQ+��Fi�- ����ŽH����^��>/�]�F��Z�ȟf�      ��b���f�6���ȟf�rSC��K �Gn����Ž����Z��k��|ռX��Ey-����x.�y���O�:�*�:��;o4;s�>;)D;�vF;I�G;��G;�8H;\cH;x�H;��H;[�H;e�H;��H;��H;K�H;f�H;K�H;��H;��H;e�H;[�H;��H;x�H;\cH;�8H;��G;I�G;�vF;)D;s�>;o4;��;�*�:�O�:y��x.����Ey-�X���|ռ�k��Z������ŽGn���K �rSC�ȟf�6���f�b���      {�˾��Ǿi���
���C͓�9�x�ؘJ��K �H��� �������?���t뮼�[�����3|��W��<�:u~�:';�
/;�f<;�C;� F;�MG;��G;9,H;sZH;�|H;ǖH;©H;��H;��H;��H;��H;��H;��H;��H;��H;��H;©H;ǖH;�|H;sZH;9,H;��G;�MG;� F;�C;�f<;�
/;';u~�:<�:�W��3|������[�t뮼����?���� ��H����K �ؘJ�9�x�C͓�
���i�����Ǿ      e� ������쾻{ԾS���b���9�x�rSC��^�ͻ޽%���Q�e����ѼG������R�����դ8��:�X;��);5�9;-�A;��E;�G;2�G;s H;DRH;�vH;v�H;��H;:�H;��H;r�H;u�H;��H;u�H;r�H;��H;:�H;��H;v�H;�vH;DRH;s H;2�G;�G;��E;-�A;5�9;��);�X;��:դ8����R�����G���Ѽ��Q�e�%���ͻ޽�^�rSC�9�x�b���S����{Ծ�쾃���      ����D��k�e� �<�ݾS���C͓�ȟf��>/�x��~'��n섽/�6�Rt��v��?�:�Tʻ�.�ݷ��s�:1; �$;�X7;��@;	E;:�F;P�G;�H;EKH;�qH;��H;ɣH;�H;�H;.�H;D�H;��H;D�H;.�H;�H;�H;ɣH;��H;�qH;EKH;�H;P�G;:�F;	E;��@;�X7; �$;1;�s�:ݷ��.�Tʻ?�:��v��Rt�/�6�n섽~'��x���>/�ȟf�C͓�S���<�ݾe� ��k��D�      ߛ7�v3��'����e� ��{Ծ
���6���]�F�����ӽ���;�L�1v�x뮼-T�ǘ��PV�q�=�1(i:_��:!z ;�#5;�?;2�D;�F;�G;�H;�EH;�mH;��H;}�H;j�H;ۼH;4�H;O�H;��H;O�H;4�H;ۼH;j�H;}�H;��H;�mH;�EH;�H;�G;�F;2�D;�?;�#5;!z ;_��:1(i:q�=��PV�ǘ�-T�x뮼1v�;�L�����ӽ���]�F�6���
����{Ծe� �����'�v3�      tN��TI���;��'��k���i���f󐾖Z��K ��s�&����&^����"����g����Ѩu�R!���1<:��:n
;�f3;-�>;�AD;ՕF;�G;�H;UAH;jH;\�H;ߟH;(�H;ԻH;k�H;��H;B�H;��H;k�H;ԻH;(�H;ߟH;\�H;jH;UAH;�H;�G;ՕF;�AD;-�>;�f3;n
;��:�1<:R!��Ѩu������g��"�����&^�&����s潎K ��Z�f�i������k��'���;��TI�      I]�N�W��TI�v3��D�������Ǿb���ȟf� )� ��W;���Fi��k�x�Ǽ�[t�8�	�(Ȅ�tX��Ο:���:%�;�I2;�Y>;qD;�~F;\�G;+H;�>H;�hH;�H;�H;q�H;7�H;��H;S�H;��H;S�H;��H;7�H;q�H;�H;�H;�hH;�>H;+H;\�G;�~F;qD;�Y>;�I2;%�;���:Ο:tX��(Ȅ�8�	��[t�x�Ǽ�k��Fi�W;�� �� )�ȟf�b�����Ǿ�����D�v3��TI�N�W�      �?��ph��1v��� ��$�X��O/�#y�-�;Ѱ��j+X�����ѽ����Gn;�>�＿����B(�暩����$�e9��:^;Y.;��<;�VC;?ZF;�G;4/H;tiH;X�H;s�H;��H;E�H;��H;~�H;��H;��H;��H;~�H;��H;E�H;��H;s�H;X�H;tiH;4/H;�G;?ZF;�VC;��<;Y.;^;��:$�e9���暩��B(�����>��Gn;�������ѽ��j+X�Ѱ��-�;#y��O/�$�X�� ��1v��ph��      ph��"���V�����y�EvS�aM+��v� 9ɾ�����T�]��[ν����`\8�����x���%�\��������9B,�:��;�.;M�<; nC;�cF;�G;�0H;!jH;ǋH;ѣH;��H;��H;��H;��H;��H;��H;��H;��H;��H;��H;��H;ѣH;ǋH;!jH;�0H;�G;�cF; nC;M�<;�.;��;B,�:��9���\����%��x�����`\8������[ν]��T����� 9ɾ�v�aM+�EvS���y�V���"���      1v��V���L ��M�h�%E�I��R���i㼾n���nH�È�a�ý�Ȅ��s/��o༼#�����4J���к��9#f�:Ml;�0;P\=; �C;5�F;��G;Q5H;^lH;H�H;ϤH;��H;�H;b�H;��H;#�H; �H;#�H;��H;b�H;�H;��H;ϤH;H�H;^lH;Q5H;��G;5�F; �C;P\=;�0;Ml;#f�:��9�к4J������#���o��s/��Ȅ�a�ýÈ��nH�n��i㼾R���I��%E�M�h�L ��V���      � ����y�M�h�ބN��O/����-�߾�A���*|�ؕ6�a}��㳽KSt�(�!�Wrμ(F{��_�Y��h����:���:VZ;2;�N>;�D;��F;��G;J<H;�oH;��H;t�H;��H;��H;��H;��H;��H;�H;��H;��H;��H;��H;��H;t�H;��H;�oH;J<H;��G;��F;�D;�N>;2;VZ;���:�:h���Y���_�(F{�Wrμ(�!�KSt��㳽a}�ؕ6��*|��A��-�߾����O/�ބN�M�h���y�      $�X�EvS�%E��O/��S�1W����������4S\�� �q�&�����Y�h��������]�}���T�b��Y���Y:~�:�_;��4;�?;|�D;�F;/�G;5EH;tH;�H;��H;��H;3�H;��H;D�H;7�H;�H;7�H;D�H;��H;3�H;��H;��H;�H;tH;5EH;/�G;�F;|�D;�?;��4;�_;~�:��Y:�Y�T�b�}�����]�����h����Y�&���q�� �4S\���������1W���S��O/�%E�EvS�      �O/�aM+�I�����1W�� 9ɾ0���Mw�� :�Y��_�ý�L��Dn;�>���bv���E<��˻)�-����x�:^;%;�7;��@;V4E;�!G;,�G;hOH;0zH;��H;��H;��H;��H;�H;2�H;�H;��H;�H;2�H;�H;��H;��H;��H;��H;0zH;hOH;,�G;�!G;V4E;��@;�7;%;^;�x�:��)�-��˻�E<�bv��>���Dn;��L��_�ýY��� :��Mw�0�� 9ɾ1W�����I��aM+�      #y��v�R���-�߾����0��1����nH���(Ὁu��r�d�O�Prμ="�����	��3���k89v:�:��;+;�{:;�6B;)�E;EaG;�H;ZH;��H;M�H;ĮH;�H;e�H;e�H;*�H;��H;��H;��H;*�H;e�H;e�H;�H;ĮH;M�H;��H;ZH;�H;EaG;)�E;�6B;�{:;+;��;v:�:�k893��	�����="��PrμO�r�d��u��(����nH�1���0������-�߾R����v�      -�; 9ɾi㼾�A�������Mw��nH�����Z��㳽����Z\8�P#�������]N�J��.�b�YJx�w5:��:��;8�0;v\=;u�C;�ZF;�G;)H;eH;��H;F�H;g�H;��H;7�H;��H;P�H;��H;��H;��H;P�H;��H;7�H;��H;g�H;F�H;��H;eH;)H;�G;�ZF;u�C;v\=;8�0;��;��:w5:YJx�.�b�J���]N�����P#��Z\8������㳽�Z񽞯��nH��Mw������A��i㼾 9ɾ      Ѱ������n���*|�4S\�� :����Z�U$������K�c���Oļ����������y&�-��O.�:0^;��#;G6;��?;-�D;��F;��G;)?H;�oH;�H;��H;9�H;q�H;J�H;��H;��H;��H;��H;��H;��H;��H;J�H;q�H;9�H;��H;�H;�oH;)?H;��G;��F;-�D;��?;G6;��#;0^;O.�:-��y&������������Oļc���K����U$���Z���� :�4S\��*|�n������      j+X��T��nH�ؕ6�� �Y��(��㳽����mR����ټ�����E<��?ݻbd\�c ��#:�c�:8�;y�,;��:;�6B;ͱE;�KG;iH;�RH;�zH;��H;
�H;9�H;`�H;n�H;+�H;��H;�H;��H;�H;��H;+�H;n�H;`�H;9�H;
�H;��H;�zH;�RH;iH;�KG;ͱE;�6B;��:;y�,;8�;�c�:#:c ��bd\��?ݻ�E<������ټ���mR�����㳽(�Y��� �ؕ6��nH��T�      ��]�È�a}�q�_�ý�u�������K����o�Wv���&R���f^����R@���:�A;�";��4;��>;�D;��F;,�G; )H;�cH;��H;5�H;��H;N�H;M�H;��H;��H;<�H;(�H;��H;(�H;<�H;��H;��H;M�H;N�H;��H;5�H;��H;�cH; )H;,�G;��F;�D;��>;��4;�";�A;��:R@���f^�����&R�Wv���o����K������u��_�ýq�a}�È�]�      ��ѽ�[νa�ý�㳽&����L��r�d�Z\8�c���ټWv����Y��_����z��]���Y:?��:�l;r-;Q�:;��A;qnE;�!G;��G;�FH;�rH;�H;��H;�H;J�H;5�H;��H;��H;��H;B�H;�H;B�H;��H;��H;��H;5�H;J�H;�H;��H;�H;�rH;�FH;��G;�!G;qnE;��A;Q�:;r-;�l;?��:��Y:]�z������_���Y�Wv���ټc��Z\8�r�d��L��&����㳽a�ý�[ν      ���������Ȅ�KSt���Y�Dn;�O�P#���Oļ�����&R��_������N3�/�Y�-2:�:9�;@?&;(G6;�W?;�D;fwF;�G;c H;�]H;��H;�H;�H;a�H;#�H;�H;��H;(�H;��H;i�H;$�H;i�H;��H;(�H;��H;�H;#�H;a�H;�H;�H;��H;�]H;c H;�G;fwF;�D;�W?;(G6;@?&;9�;�:-2:/�Y��N3������_��&R������OļP#��O�Dn;���Y�KSt��Ȅ�����      Gn;�`\8��s/�(�!�h��>���Prμ��������E<�������N3��Ix�a�9��:T^;� ;~2;��<;.�B;�E;e4G;1�G;^EH;�pH;��H;h�H;ϳH;k�H;��H;��H;�H;��H;1�H;��H;�H;��H;1�H;��H;�H;��H;��H;k�H;ϳH;h�H;��H;�pH;^EH;1�G;e4G;�E;.�B;��<;~2;� ;T^;��:a�9�Ix��N3�������E<��������Prμ>���h��(�!��s/�`\8�      >�Ｘ���o�Wrμ����bv��="���]N�����?ݻf^��z��/�Y�a�9��:���:B�;��.;�{:;2>A;��D;`�F;ߵG;
)H;D`H;5�H;��H;�H;R�H;6�H;R�H;t�H;�H;.�H;k�H;��H;��H;��H;k�H;.�H;�H;t�H;R�H;6�H;R�H;�H;��H;5�H;D`H;
)H;ߵG;`�F;��D;2>A;�{:;��.;B�;���:��:a�9/�Y�z��f^���?ݻ����]N�="��bv������Wrμ�o༸��      �����x���#��(F{���]��E<����J�뻲���bd\���]�-2:��:���:�Z;��,;/�8;` @;0D;�ZF;PzG;
H;iOH;=uH;�H;[�H;�H;B�H;z�H;��H;��H;��H;��H;��H;��H;��H;��H;��H;��H;��H;��H;��H;z�H;B�H;�H;[�H;�H;=uH;iOH;
H;PzG;�ZF;0D;` @;/�8;��,;�Z;���:��:-2:]���bd\�����J�뻛���E<���]�(F{��#���x��      �B(��%�����_�}����˻	��.�b�y&�c ��R@���Y:�:T^;B�;��,;Z_8;��?;��C;�F;FG;t�G;?H;FjH;#�H; �H;
�H;k�H;��H;~�H;��H;/�H;��H;��H;��H;��H;��H;��H;��H;��H;��H;/�H;��H;~�H;��H;k�H;
�H; �H;#�H;FjH;?H;t�G;FG;�F;��C;��?;Z_8;��,;B�;T^;�:��Y:R@�c ��y&�.�b�	���˻}����_�����%�      暩�\���4J��Y��T�b�)�-�3��YJx�-��#:��:?��:9�;� ;��.;/�8;��?;2�C;�E;e"G;�G;1H;aH;gH;��H;��H;��H;��H;s�H;(�H;I�H;J�H;��H;(�H;��H;G�H;��H;G�H;��H;(�H;��H;J�H;I�H;(�H;s�H;��H;��H;��H;��H;gH;aH;1H;�G;e"G;�E;2�C;��?;/�8;��.;� ;9�;?��:��:#:-��YJx�3��)�-�T�b�Y��4J��\���      �����뺸кh����Y����k89w5:O.�:�c�:�A;�l;@?&;~2;�{:;` @;��C;�E;�G;�G;}'H;ZH;�yH;W�H;��H;��H;{�H;��H;��H;l�H;��H;
�H;[�H;<�H;W�H;
�H;��H;
�H;W�H;<�H;[�H;
�H;��H;l�H;��H;��H;{�H;��H;��H;W�H;�yH;ZH;}'H;�G;�G;�E;��C;` @;�{:;~2;@?&;�l;�A;�c�:O.�:w5:�k89���Y�h����к���      $�e9��9��9�:��Y:�x�:v:�:��:0^;8�;�";r-;(G6;��<;2>A;0D;�F;e"G;�G;$H;VH;�uH;��H;X�H;b�H;��H;!�H;��H;��H;E�H;��H;��H;��H;6�H;�H;��H;�H;��H;�H;6�H;��H;��H;��H;E�H;��H;��H;!�H;��H;b�H;X�H;��H;�uH;VH;$H;�G;e"G;�F;0D;2>A;��<;(G6;r-;�";8�;0^;��:v:�:�x�:��Y:�:��9��9      ��:B,�:#f�:���:~�:^;��;��;��#;y�,;��4;Q�:;�W?;.�B;��D;�ZF;FG;�G;}'H;VH;�tH;��H;.�H;�H;<�H;	�H;��H;��H;��H;��H;��H;��H;��H;��H;��H;^�H;b�H;^�H;��H;��H;��H;��H;��H;��H;��H;��H;��H;	�H;<�H;�H;.�H;��H;�tH;VH;}'H;�G;FG;�ZF;��D;.�B;�W?;Q�:;��4;y�,;��#;��;��;^;~�:���:#f�:B,�:      ^;��;Ml;VZ;�_;%;+;8�0;G6;��:;��>;��A;�D;�E;`�F;PzG;t�G;1H;ZH;�uH;��H;g�H;ܫH;߷H;��H;e�H;��H;��H;��H;��H;H�H;G�H;��H;��H;p�H;��H;��H;��H;p�H;��H;��H;G�H;H�H;��H;��H;��H;��H;e�H;��H;߷H;ܫH;g�H;��H;�uH;ZH;1H;t�G;PzG;`�F;�E;�D;��A;��>;��:;G6;8�0;+;%;�_;VZ;Ml;��;      Y.;�.;�0;2;��4;�7;�{:;v\=;��?;�6B;�D;qnE;fwF;e4G;ߵG;
H;?H;aH;�yH;��H;.�H;ܫH;`�H;��H;�H;��H;��H;�H;)�H;��H;��H;h�H;c�H;O�H;��H;(�H;P�H;(�H;��H;O�H;c�H;h�H;��H;��H;)�H;�H;��H;��H;�H;��H;`�H;ܫH;.�H;��H;�yH;aH;?H;
H;ߵG;e4G;fwF;qnE;�D;�6B;��?;v\=;�{:;�7;��4;2;�0;�.;      ��<;M�<;P\=;�N>;�?;��@;�6B;u�C;-�D;ͱE;��F;�!G;�G;1�G;
)H;iOH;FjH;gH;W�H;X�H;�H;߷H;��H;H�H;I�H;E�H;W�H;��H;,�H;B�H;�H;�H;�H;��H;H�H;��H;��H;��H;H�H;��H;�H;�H;�H;B�H;,�H;��H;W�H;E�H;I�H;H�H;��H;߷H;�H;X�H;W�H;gH;FjH;iOH;
)H;1�G;�G;�!G;��F;ͱE;-�D;u�C;�6B;��@;�?;�N>;P\=;M�<;      �VC; nC; �C;�D;|�D;V4E;)�E;�ZF;��F;�KG;,�G;��G;c H;^EH;D`H;=uH;#�H;��H;��H;b�H;<�H;��H;�H;I�H;�H;�H;O�H;��H;��H;��H;��H;��H;��H;=�H;��H;��H;��H;��H;��H;=�H;��H;��H;��H;��H;��H;��H;O�H;�H;�H;I�H;�H;��H;<�H;b�H;��H;��H;#�H;=uH;D`H;^EH;c H;��G;,�G;�KG;��F;�ZF;)�E;V4E;|�D;�D; �C; nC;      ?ZF;�cF;5�F;��F;�F;�!G;EaG;�G;��G;iH; )H;�FH;�]H;�pH;5�H;�H; �H;��H;��H;��H;	�H;e�H;��H;E�H;�H;5�H;��H;��H;t�H;��H;��H;��H;,�H;~�H;��H;�H;�H;�H;��H;~�H;,�H;��H;��H;��H;t�H;��H;��H;5�H;�H;E�H;��H;e�H;	�H;��H;��H;��H; �H;�H;5�H;�pH;�]H;�FH; )H;iH;��G;�G;EaG;�!G;�F;��F;5�F;�cF;      �G;�G;��G;��G;/�G;,�G;�H;)H;)?H;�RH;�cH;�rH;��H;��H;��H;[�H;
�H;��H;{�H;!�H;��H;��H;��H;W�H;O�H;��H;��H;J�H;��H;��H;j�H; �H;}�H;��H;�H;;�H;Y�H;;�H;�H;��H;}�H; �H;j�H;��H;��H;J�H;��H;��H;O�H;W�H;��H;��H;��H;!�H;{�H;��H;
�H;[�H;��H;��H;��H;�rH;�cH;�RH;)?H;)H;�H;,�G;/�G;��G;��G;�G;      4/H;�0H;Q5H;J<H;5EH;hOH;ZH;eH;�oH;�zH;��H;�H;�H;h�H;�H;�H;k�H;��H;��H;��H;��H;��H;�H;��H;��H;��H;J�H;��H;e�H;S�H;�H;i�H;��H;�H;E�H;[�H;M�H;[�H;E�H;�H;��H;i�H;�H;S�H;e�H;��H;J�H;��H;��H;��H;�H;��H;��H;��H;��H;��H;k�H;�H;�H;h�H;�H;�H;��H;�zH;�oH;eH;ZH;hOH;5EH;J<H;Q5H;�0H;      tiH;!jH;^lH;�oH;tH;0zH;��H;��H;�H;��H;5�H;��H;�H;ϳH;R�H;B�H;��H;s�H;��H;��H;��H;��H;)�H;,�H;��H;t�H;��H;e�H;[�H;��H;Y�H;��H;��H;5�H;e�H;o�H;b�H;o�H;e�H;5�H;��H;��H;Y�H;��H;[�H;e�H;��H;t�H;��H;,�H;)�H;��H;��H;��H;��H;s�H;��H;B�H;R�H;ϳH;�H;��H;5�H;��H;�H;��H;��H;0zH;tH;�oH;^lH;!jH;      X�H;ǋH;H�H;��H;�H;��H;M�H;F�H;��H;
�H;��H;�H;a�H;k�H;6�H;z�H;~�H;(�H;l�H;E�H;��H;��H;��H;B�H;��H;��H;��H;S�H;��H;K�H;��H;��H;6�H;]�H;h�H;��H;��H;��H;h�H;]�H;6�H;��H;��H;K�H;��H;S�H;��H;��H;��H;B�H;��H;��H;��H;E�H;l�H;(�H;~�H;z�H;6�H;k�H;a�H;�H;��H;
�H;��H;F�H;M�H;��H;�H;��H;H�H;ǋH;      s�H;ѣH;ϤH;t�H;��H;��H;ĮH;g�H;9�H;9�H;N�H;J�H;#�H;��H;R�H;��H;��H;I�H;��H;��H;��H;H�H;��H;�H;��H;��H;j�H;�H;Y�H;��H;��H;)�H;a�H;o�H;��H;��H;��H;��H;��H;o�H;a�H;)�H;��H;��H;Y�H;�H;j�H;��H;��H;�H;��H;H�H;��H;��H;��H;I�H;��H;��H;R�H;��H;#�H;J�H;N�H;9�H;9�H;g�H;ĮH;��H;��H;t�H;ϤH;ѣH;      ��H;��H;��H;��H;��H;��H;�H;��H;q�H;`�H;M�H;5�H;�H;��H;t�H;��H;/�H;J�H;
�H;��H;��H;G�H;h�H;�H;��H;��H; �H;i�H;��H;��H;)�H;A�H;k�H;��H;��H;��H;��H;��H;��H;��H;k�H;A�H;)�H;��H;��H;i�H; �H;��H;��H;�H;h�H;G�H;��H;��H;
�H;J�H;/�H;��H;t�H;��H;�H;5�H;M�H;`�H;q�H;��H;�H;��H;��H;��H;��H;��H;      E�H;��H;�H;��H;3�H;��H;e�H;7�H;J�H;n�H;��H;��H;��H;�H;�H;��H;��H;��H;[�H;��H;��H;��H;c�H;�H;��H;,�H;}�H;��H;��H;6�H;a�H;k�H;{�H;��H;��H;��H;��H;��H;��H;��H;{�H;k�H;a�H;6�H;��H;��H;}�H;,�H;��H;�H;c�H;��H;��H;��H;[�H;��H;��H;��H;�H;�H;��H;��H;��H;n�H;J�H;7�H;e�H;��H;3�H;��H;�H;��H;      ��H;��H;b�H;��H;��H;�H;e�H;��H;��H;+�H;��H;��H;(�H;��H;.�H;��H;��H;(�H;<�H;6�H;��H;��H;O�H;��H;=�H;~�H;��H;�H;5�H;]�H;o�H;��H;��H;��H;��H;��H;��H;��H;��H;��H;��H;��H;o�H;]�H;5�H;�H;��H;~�H;=�H;��H;O�H;��H;��H;6�H;<�H;(�H;��H;��H;.�H;��H;(�H;��H;��H;+�H;��H;��H;e�H;�H;��H;��H;b�H;��H;      ~�H;��H;��H;��H;D�H;2�H;*�H;P�H;��H;��H;<�H;��H;��H;1�H;k�H;��H;��H;��H;W�H;�H;��H;p�H;��H;H�H;��H;��H;�H;E�H;e�H;h�H;��H;��H;��H;��H;��H;��H;��H;��H;��H;��H;��H;��H;��H;h�H;e�H;E�H;�H;��H;��H;H�H;��H;p�H;��H;�H;W�H;��H;��H;��H;k�H;1�H;��H;��H;<�H;��H;��H;P�H;*�H;2�H;D�H;��H;��H;��H;      ��H;��H;#�H;��H;7�H;�H;��H;��H;��H;�H;(�H;B�H;i�H;��H;��H;��H;��H;G�H;
�H;��H;^�H;��H;(�H;��H;��H;�H;;�H;[�H;o�H;��H;��H;��H;��H;��H;��H;��H;��H;��H;��H;��H;��H;��H;��H;��H;o�H;[�H;;�H;�H;��H;��H;(�H;��H;^�H;��H;
�H;G�H;��H;��H;��H;��H;i�H;B�H;(�H;�H;��H;��H;��H;�H;7�H;��H;#�H;��H;      ��H;��H; �H;�H;�H;��H;��H;��H;��H;��H;��H;�H;$�H;�H;��H;��H;��H;��H;��H;�H;b�H;��H;P�H;��H;��H;�H;Y�H;M�H;b�H;��H;��H;��H;��H;��H;��H;��H;��H;��H;��H;��H;��H;��H;��H;��H;b�H;M�H;Y�H;�H;��H;��H;P�H;��H;b�H;�H;��H;��H;��H;��H;��H;�H;$�H;�H;��H;��H;��H;��H;��H;��H;�H;�H; �H;��H;      ��H;��H;#�H;��H;7�H;�H;��H;��H;��H;�H;(�H;B�H;i�H;��H;��H;��H;��H;G�H;
�H;��H;^�H;��H;(�H;��H;��H;�H;;�H;[�H;o�H;��H;��H;��H;��H;��H;��H;��H;��H;��H;��H;��H;��H;��H;��H;��H;o�H;[�H;;�H;�H;��H;��H;(�H;��H;^�H;��H;
�H;G�H;��H;��H;��H;��H;i�H;B�H;(�H;�H;��H;��H;��H;�H;7�H;��H;#�H;��H;      ~�H;��H;��H;��H;D�H;2�H;*�H;P�H;��H;��H;<�H;��H;��H;1�H;k�H;��H;��H;��H;W�H;�H;��H;p�H;��H;H�H;��H;��H;�H;E�H;e�H;h�H;��H;��H;��H;��H;��H;��H;��H;��H;��H;��H;��H;��H;��H;h�H;e�H;E�H;�H;��H;��H;H�H;��H;p�H;��H;�H;W�H;��H;��H;��H;k�H;1�H;��H;��H;<�H;��H;��H;P�H;*�H;2�H;D�H;��H;��H;��H;      ��H;��H;b�H;��H;��H;�H;e�H;��H;��H;+�H;��H;��H;(�H;��H;.�H;��H;��H;(�H;<�H;6�H;��H;��H;O�H;��H;=�H;~�H;��H;�H;5�H;]�H;o�H;��H;��H;��H;��H;��H;��H;��H;��H;��H;��H;��H;o�H;]�H;5�H;�H;��H;~�H;=�H;��H;O�H;��H;��H;6�H;<�H;(�H;��H;��H;.�H;��H;(�H;��H;��H;+�H;��H;��H;e�H;�H;��H;��H;b�H;��H;      E�H;��H;�H;��H;3�H;��H;e�H;7�H;J�H;n�H;��H;��H;��H;�H;�H;��H;��H;��H;[�H;��H;��H;��H;c�H;�H;��H;,�H;}�H;��H;��H;6�H;a�H;k�H;{�H;��H;��H;��H;��H;��H;��H;��H;{�H;k�H;a�H;6�H;��H;��H;}�H;,�H;��H;�H;c�H;��H;��H;��H;[�H;��H;��H;��H;�H;�H;��H;��H;��H;n�H;J�H;7�H;e�H;��H;3�H;��H;�H;��H;      ��H;��H;��H;��H;��H;��H;�H;��H;q�H;`�H;M�H;5�H;�H;��H;t�H;��H;/�H;J�H;
�H;��H;��H;G�H;h�H;�H;��H;��H; �H;i�H;��H;��H;)�H;A�H;k�H;��H;��H;��H;��H;��H;��H;��H;k�H;A�H;)�H;��H;��H;i�H; �H;��H;��H;�H;h�H;G�H;��H;��H;
�H;J�H;/�H;��H;t�H;��H;�H;5�H;M�H;`�H;q�H;��H;�H;��H;��H;��H;��H;��H;      s�H;ѣH;ϤH;t�H;��H;��H;ĮH;g�H;9�H;9�H;N�H;J�H;#�H;��H;R�H;��H;��H;I�H;��H;��H;��H;H�H;��H;�H;��H;��H;j�H;�H;Y�H;��H;��H;)�H;a�H;o�H;��H;��H;��H;��H;��H;o�H;a�H;)�H;��H;��H;Y�H;�H;j�H;��H;��H;�H;��H;H�H;��H;��H;��H;I�H;��H;��H;R�H;��H;#�H;J�H;N�H;9�H;9�H;g�H;ĮH;��H;��H;t�H;ϤH;ѣH;      X�H;ǋH;H�H;��H;�H;��H;M�H;F�H;��H;
�H;��H;�H;a�H;k�H;6�H;z�H;~�H;(�H;l�H;E�H;��H;��H;��H;B�H;��H;��H;��H;S�H;��H;K�H;��H;��H;6�H;]�H;h�H;��H;��H;��H;h�H;]�H;6�H;��H;��H;K�H;��H;S�H;��H;��H;��H;B�H;��H;��H;��H;E�H;l�H;(�H;~�H;z�H;6�H;k�H;a�H;�H;��H;
�H;��H;F�H;M�H;��H;�H;��H;H�H;ǋH;      tiH;!jH;^lH;�oH;tH;0zH;��H;��H;�H;��H;5�H;��H;�H;ϳH;R�H;B�H;��H;s�H;��H;��H;��H;��H;)�H;,�H;��H;t�H;��H;e�H;[�H;��H;Y�H;��H;��H;5�H;e�H;o�H;b�H;o�H;e�H;5�H;��H;��H;Y�H;��H;[�H;e�H;��H;t�H;��H;,�H;)�H;��H;��H;��H;��H;s�H;��H;B�H;R�H;ϳH;�H;��H;5�H;��H;�H;��H;��H;0zH;tH;�oH;^lH;!jH;      4/H;�0H;Q5H;J<H;5EH;hOH;ZH;eH;�oH;�zH;��H;�H;�H;h�H;�H;�H;k�H;��H;��H;��H;��H;��H;�H;��H;��H;��H;J�H;��H;e�H;S�H;�H;i�H;��H;�H;E�H;[�H;M�H;[�H;E�H;�H;��H;i�H;�H;S�H;e�H;��H;J�H;��H;��H;��H;�H;��H;��H;��H;��H;��H;k�H;�H;�H;h�H;�H;�H;��H;�zH;�oH;eH;ZH;hOH;5EH;J<H;Q5H;�0H;      �G;�G;��G;��G;/�G;,�G;�H;)H;)?H;�RH;�cH;�rH;��H;��H;��H;[�H;
�H;��H;{�H;!�H;��H;��H;��H;W�H;O�H;��H;��H;J�H;��H;��H;j�H; �H;}�H;��H;�H;;�H;Y�H;;�H;�H;��H;}�H; �H;j�H;��H;��H;J�H;��H;��H;O�H;W�H;��H;��H;��H;!�H;{�H;��H;
�H;[�H;��H;��H;��H;�rH;�cH;�RH;)?H;)H;�H;,�G;/�G;��G;��G;�G;      ?ZF;�cF;5�F;��F;�F;�!G;EaG;�G;��G;iH; )H;�FH;�]H;�pH;5�H;�H; �H;��H;��H;��H;	�H;e�H;��H;E�H;�H;5�H;��H;��H;t�H;��H;��H;��H;,�H;~�H;��H;�H;�H;�H;��H;~�H;,�H;��H;��H;��H;t�H;��H;��H;5�H;�H;E�H;��H;e�H;	�H;��H;��H;��H; �H;�H;5�H;�pH;�]H;�FH; )H;iH;��G;�G;EaG;�!G;�F;��F;5�F;�cF;      �VC; nC; �C;�D;|�D;V4E;)�E;�ZF;��F;�KG;,�G;��G;c H;^EH;D`H;=uH;#�H;��H;��H;b�H;<�H;��H;�H;I�H;�H;�H;O�H;��H;��H;��H;��H;��H;��H;=�H;��H;��H;��H;��H;��H;=�H;��H;��H;��H;��H;��H;��H;O�H;�H;�H;I�H;�H;��H;<�H;b�H;��H;��H;#�H;=uH;D`H;^EH;c H;��G;,�G;�KG;��F;�ZF;)�E;V4E;|�D;�D; �C; nC;      ��<;M�<;P\=;�N>;�?;��@;�6B;u�C;-�D;ͱE;��F;�!G;�G;1�G;
)H;iOH;FjH;gH;W�H;X�H;�H;߷H;��H;H�H;I�H;E�H;W�H;��H;,�H;B�H;�H;�H;�H;��H;H�H;��H;��H;��H;H�H;��H;�H;�H;�H;B�H;,�H;��H;W�H;E�H;I�H;H�H;��H;߷H;�H;X�H;W�H;gH;FjH;iOH;
)H;1�G;�G;�!G;��F;ͱE;-�D;u�C;�6B;��@;�?;�N>;P\=;M�<;      Y.;�.;�0;2;��4;�7;�{:;v\=;��?;�6B;�D;qnE;fwF;e4G;ߵG;
H;?H;aH;�yH;��H;.�H;ܫH;`�H;��H;�H;��H;��H;�H;)�H;��H;��H;h�H;c�H;O�H;��H;(�H;P�H;(�H;��H;O�H;c�H;h�H;��H;��H;)�H;�H;��H;��H;�H;��H;`�H;ܫH;.�H;��H;�yH;aH;?H;
H;ߵG;e4G;fwF;qnE;�D;�6B;��?;v\=;�{:;�7;��4;2;�0;�.;      ^;��;Ml;VZ;�_;%;+;8�0;G6;��:;��>;��A;�D;�E;`�F;PzG;t�G;1H;ZH;�uH;��H;g�H;ܫH;߷H;��H;e�H;��H;��H;��H;��H;H�H;G�H;��H;��H;p�H;��H;��H;��H;p�H;��H;��H;G�H;H�H;��H;��H;��H;��H;e�H;��H;߷H;ܫH;g�H;��H;�uH;ZH;1H;t�G;PzG;`�F;�E;�D;��A;��>;��:;G6;8�0;+;%;�_;VZ;Ml;��;      ��:B,�:#f�:���:~�:^;��;��;��#;y�,;��4;Q�:;�W?;.�B;��D;�ZF;FG;�G;}'H;VH;�tH;��H;.�H;�H;<�H;	�H;��H;��H;��H;��H;��H;��H;��H;��H;��H;^�H;b�H;^�H;��H;��H;��H;��H;��H;��H;��H;��H;��H;	�H;<�H;�H;.�H;��H;�tH;VH;}'H;�G;FG;�ZF;��D;.�B;�W?;Q�:;��4;y�,;��#;��;��;^;~�:���:#f�:B,�:      $�e9��9��9�:��Y:�x�:v:�:��:0^;8�;�";r-;(G6;��<;2>A;0D;�F;e"G;�G;$H;VH;�uH;��H;X�H;b�H;��H;!�H;��H;��H;E�H;��H;��H;��H;6�H;�H;��H;�H;��H;�H;6�H;��H;��H;��H;E�H;��H;��H;!�H;��H;b�H;X�H;��H;�uH;VH;$H;�G;e"G;�F;0D;2>A;��<;(G6;r-;�";8�;0^;��:v:�:�x�:��Y:�:��9��9      �����뺸кh����Y����k89w5:O.�:�c�:�A;�l;@?&;~2;�{:;` @;��C;�E;�G;�G;}'H;ZH;�yH;W�H;��H;��H;{�H;��H;��H;l�H;��H;
�H;[�H;<�H;W�H;
�H;��H;
�H;W�H;<�H;[�H;
�H;��H;l�H;��H;��H;{�H;��H;��H;W�H;�yH;ZH;}'H;�G;�G;�E;��C;` @;�{:;~2;@?&;�l;�A;�c�:O.�:w5:�k89���Y�h����к���      暩�\���4J��Y��T�b�)�-�3��YJx�-��#:��:?��:9�;� ;��.;/�8;��?;2�C;�E;e"G;�G;1H;aH;gH;��H;��H;��H;��H;s�H;(�H;I�H;J�H;��H;(�H;��H;G�H;��H;G�H;��H;(�H;��H;J�H;I�H;(�H;s�H;��H;��H;��H;��H;gH;aH;1H;�G;e"G;�E;2�C;��?;/�8;��.;� ;9�;?��:��:#:-��YJx�3��)�-�T�b�Y��4J��\���      �B(��%�����_�}����˻	��.�b�y&�c ��R@���Y:�:T^;B�;��,;Z_8;��?;��C;�F;FG;t�G;?H;FjH;#�H; �H;
�H;k�H;��H;~�H;��H;/�H;��H;��H;��H;��H;��H;��H;��H;��H;��H;/�H;��H;~�H;��H;k�H;
�H; �H;#�H;FjH;?H;t�G;FG;�F;��C;��?;Z_8;��,;B�;T^;�:��Y:R@�c ��y&�.�b�	���˻}����_�����%�      �����x���#��(F{���]��E<����J�뻲���bd\���]�-2:��:���:�Z;��,;/�8;` @;0D;�ZF;PzG;
H;iOH;=uH;�H;[�H;�H;B�H;z�H;��H;��H;��H;��H;��H;��H;��H;��H;��H;��H;��H;��H;��H;z�H;B�H;�H;[�H;�H;=uH;iOH;
H;PzG;�ZF;0D;` @;/�8;��,;�Z;���:��:-2:]���bd\�����J�뻛���E<���]�(F{��#���x��      >�Ｘ���o�Wrμ����bv��="���]N�����?ݻf^��z��/�Y�a�9��:���:B�;��.;�{:;2>A;��D;`�F;ߵG;
)H;D`H;5�H;��H;�H;R�H;6�H;R�H;t�H;�H;.�H;k�H;��H;��H;��H;k�H;.�H;�H;t�H;R�H;6�H;R�H;�H;��H;5�H;D`H;
)H;ߵG;`�F;��D;2>A;�{:;��.;B�;���:��:a�9/�Y�z��f^���?ݻ����]N�="��bv������Wrμ�o༸��      Gn;�`\8��s/�(�!�h��>���Prμ��������E<�������N3��Ix�a�9��:T^;� ;~2;��<;.�B;�E;e4G;1�G;^EH;�pH;��H;h�H;ϳH;k�H;��H;��H;�H;��H;1�H;��H;�H;��H;1�H;��H;�H;��H;��H;k�H;ϳH;h�H;��H;�pH;^EH;1�G;e4G;�E;.�B;��<;~2;� ;T^;��:a�9�Ix��N3�������E<��������Prμ>���h��(�!��s/�`\8�      ���������Ȅ�KSt���Y�Dn;�O�P#���Oļ�����&R��_������N3�/�Y�-2:�:9�;@?&;(G6;�W?;�D;fwF;�G;c H;�]H;��H;�H;�H;a�H;#�H;�H;��H;(�H;��H;i�H;$�H;i�H;��H;(�H;��H;�H;#�H;a�H;�H;�H;��H;�]H;c H;�G;fwF;�D;�W?;(G6;@?&;9�;�:-2:/�Y��N3������_��&R������OļP#��O�Dn;���Y�KSt��Ȅ�����      ��ѽ�[νa�ý�㳽&����L��r�d�Z\8�c���ټWv����Y��_����z��]���Y:?��:�l;r-;Q�:;��A;qnE;�!G;��G;�FH;�rH;�H;��H;�H;J�H;5�H;��H;��H;��H;B�H;�H;B�H;��H;��H;��H;5�H;J�H;�H;��H;�H;�rH;�FH;��G;�!G;qnE;��A;Q�:;r-;�l;?��:��Y:]�z������_���Y�Wv���ټc��Z\8�r�d��L��&����㳽a�ý�[ν      ��]�È�a}�q�_�ý�u�������K����o�Wv���&R���f^����R@���:�A;�";��4;��>;�D;��F;,�G; )H;�cH;��H;5�H;��H;N�H;M�H;��H;��H;<�H;(�H;��H;(�H;<�H;��H;��H;M�H;N�H;��H;5�H;��H;�cH; )H;,�G;��F;�D;��>;��4;�";�A;��:R@���f^�����&R�Wv���o����K������u��_�ýq�a}�È�]�      j+X��T��nH�ؕ6�� �Y��(��㳽����mR����ټ�����E<��?ݻbd\�c ��#:�c�:8�;y�,;��:;�6B;ͱE;�KG;iH;�RH;�zH;��H;
�H;9�H;`�H;n�H;+�H;��H;�H;��H;�H;��H;+�H;n�H;`�H;9�H;
�H;��H;�zH;�RH;iH;�KG;ͱE;�6B;��:;y�,;8�;�c�:#:c ��bd\��?ݻ�E<������ټ���mR�����㳽(�Y��� �ؕ6��nH��T�      Ѱ������n���*|�4S\�� :����Z�U$������K�c���Oļ����������y&�-��O.�:0^;��#;G6;��?;-�D;��F;��G;)?H;�oH;�H;��H;9�H;q�H;J�H;��H;��H;��H;��H;��H;��H;��H;J�H;q�H;9�H;��H;�H;�oH;)?H;��G;��F;-�D;��?;G6;��#;0^;O.�:-��y&������������Oļc���K����U$���Z���� :�4S\��*|�n������      -�; 9ɾi㼾�A�������Mw��nH�����Z��㳽����Z\8�P#�������]N�J��.�b�YJx�w5:��:��;8�0;v\=;u�C;�ZF;�G;)H;eH;��H;F�H;g�H;��H;7�H;��H;P�H;��H;��H;��H;P�H;��H;7�H;��H;g�H;F�H;��H;eH;)H;�G;�ZF;u�C;v\=;8�0;��;��:w5:YJx�.�b�J���]N�����P#��Z\8������㳽�Z񽞯��nH��Mw������A��i㼾 9ɾ      #y��v�R���-�߾����0��1����nH���(Ὁu��r�d�O�Prμ="�����	��3���k89v:�:��;+;�{:;�6B;)�E;EaG;�H;ZH;��H;M�H;ĮH;�H;e�H;e�H;*�H;��H;��H;��H;*�H;e�H;e�H;�H;ĮH;M�H;��H;ZH;�H;EaG;)�E;�6B;�{:;+;��;v:�:�k893��	�����="��PrμO�r�d��u��(����nH�1���0������-�߾R����v�      �O/�aM+�I�����1W�� 9ɾ0���Mw�� :�Y��_�ý�L��Dn;�>���bv���E<��˻)�-����x�:^;%;�7;��@;V4E;�!G;,�G;hOH;0zH;��H;��H;��H;��H;�H;2�H;�H;��H;�H;2�H;�H;��H;��H;��H;��H;0zH;hOH;,�G;�!G;V4E;��@;�7;%;^;�x�:��)�-��˻�E<�bv��>���Dn;��L��_�ýY��� :��Mw�0�� 9ɾ1W�����I��aM+�      $�X�EvS�%E��O/��S�1W����������4S\�� �q�&�����Y�h��������]�}���T�b��Y���Y:~�:�_;��4;�?;|�D;�F;/�G;5EH;tH;�H;��H;��H;3�H;��H;D�H;7�H;�H;7�H;D�H;��H;3�H;��H;��H;�H;tH;5EH;/�G;�F;|�D;�?;��4;�_;~�:��Y:�Y�T�b�}�����]�����h����Y�&���q�� �4S\���������1W���S��O/�%E�EvS�      � ����y�M�h�ބN��O/����-�߾�A���*|�ؕ6�a}��㳽KSt�(�!�Wrμ(F{��_�Y��h����:���:VZ;2;�N>;�D;��F;��G;J<H;�oH;��H;t�H;��H;��H;��H;��H;��H;�H;��H;��H;��H;��H;��H;t�H;��H;�oH;J<H;��G;��F;�D;�N>;2;VZ;���:�:h���Y���_�(F{�Wrμ(�!�KSt��㳽a}�ؕ6��*|��A��-�߾����O/�ބN�M�h���y�      1v��V���L ��M�h�%E�I��R���i㼾n���nH�È�a�ý�Ȅ��s/��o༼#�����4J���к��9#f�:Ml;�0;P\=; �C;5�F;��G;Q5H;^lH;H�H;ϤH;��H;�H;b�H;��H;#�H; �H;#�H;��H;b�H;�H;��H;ϤH;H�H;^lH;Q5H;��G;5�F; �C;P\=;�0;Ml;#f�:��9�к4J������#���o��s/��Ȅ�a�ýÈ��nH�n��i㼾R���I��%E�M�h�L ��V���      ph��"���V�����y�EvS�aM+��v� 9ɾ�����T�]��[ν����`\8�����x���%�\��������9B,�:��;�.;M�<; nC;�cF;�G;�0H;!jH;ǋH;ѣH;��H;��H;��H;��H;��H;��H;��H;��H;��H;��H;��H;ѣH;ǋH;!jH;�0H;�G;�cF; nC;M�<;�.;��;B,�:��9���\����%��x�����`\8������[ν]��T����� 9ɾ�v�aM+�EvS���y�V���"���      Vܿ%�ֿ�aǿ2^��&���Io���7����iþ�(���-=��` ��@����_�&]�&p����I�r�ѻ��)��R�[�:��
;*;C�:;�B;UHF;=�G;�kH;3�H;��H;h�H;��H;��H;o�H;��H;(�H;��H;(�H;��H;o�H;��H;��H;h�H;��H;3�H;�kH;=�G;UHF;�B;C�:;*;��
;[�:�R���)�r�ѻ��I�&p��&]���_��@���` ��-=��(���iþ����7�Io�&���2^���aǿ%�ֿ      %�ֿ5pѿ֊¿������PXi�Õ3��
�GD��;l��1�9�j.���R��\� �\x��1�E��ͻ��$�� ����:��;��*;[�:;.�B;3TF;��G;ZmH;ϠH;ܶH;��H;��H;��H;�H;��H;<�H;��H;<�H;��H;�H;��H;��H;��H;ܶH;ϠH;ZmH;��G;3TF;.�B;[�:;��*;��;���:� ���$��ͻ1�E�\x�� �\��R��j.��1�9�;l��GD���
�Õ3�PXi�������֊¿5pѿ      �aǿ֊¿���������s"Y��f'�����)o���.}��k/�m��ڟ�<Q�%#�ע��(;�P������#�7���:I�;�,;��;;�C;RvF;/�G;�qH;[�H;��H;=�H;�H;�H;��H;��H;j�H;��H;j�H;��H;��H;�H;�H;=�H;��H;[�H;�qH;/�G;RvF;�C;��;;�,;I�;��:#�7����P����(;�ע�%#�<Q�ڟ�m���k/��.}�)o�������f'�s"Y����������֊¿      2^������b���Io���@���޾����&ce�"����ڽ绒��f@������R���O*�mG�����v<^9Ѳ�:[;�c.;'�<;ՏC;F�F;��G;�xH;äH;7�H;I�H;��H;��H;��H;�H;��H;6�H;��H;�H;��H;��H;��H;I�H;7�H;äH;�xH;��G;F�F;ՏC;'�<;�c.;[;Ѳ�:v<^9���mG���O*��R�������f@�绒���ڽ"��&ce������޾���@�Io�b�������      &����������Io��!J�@�#��\��HD������jPH�����b��C��t +�u�ټ%��������������:���:��;�X1;3>;�/D;��F;�H;r�H;��H;)�H;��H;��H;)�H;��H;p�H;��H;~�H;��H;p�H;��H;)�H;��H;��H;)�H;��H;r�H;�H;��F;�/D;3>;�X1;��;���:��:����������%��u�ټt +�C���b�����jPH�����HD���\��@�#��!J�Io��������      Io�PXi�s"Y���@�@�#��
��о�A�� �i���(�i��gr����_��5��ɺ�o�`��<����d�@�\�M�X:OO�:6`;#�4;�?;��D;�7G;�/H;ȊH;��H;��H;.�H;��H;��H;�H;��H;-�H;��H;-�H;��H;�H;��H;��H;.�H;��H;��H;ȊH;�/H;�7G;��D;�?;#�4;6`;OO�:M�X:@�\���d��<��o�`��ɺ��5���_�gr��i����(� �i��A���о�
�@�#���@�s"Y�PXi�      ��7�Õ3��f'���\���о�����.}��-=�o
�y�ĽO��:����������7�@GĻ+�$�S�����:�z;�C&;E+8;EIA;0�E;��G;�KH;�H;��H;R�H;�H;(�H;��H;��H;@�H;��H;5�H;��H;@�H;��H;��H;(�H;�H;R�H;��H;�H;�KH;��G;0�E;EIA;E+8;�C&;�z;���:S��+�$�@GĻ�7���������:�O��y�Ľo
��-=��.}������о�\����f'�Õ3�      ���
������޾HD���A���.}��D�[t���ڽ�!��\����P�ļ�
v�F�����Jɺ�N�9���:h';�-;ӊ;;��B;�HF;��G;?eH;ʜH;�H;N�H;��H;��H;��H;{�H;��H;�H;��H;�H;��H;{�H;��H;��H;��H;N�H;�H;ʜH;?eH;��G;�HF;��B;ӊ;;�-;h';���:�N�9�Jɺ��F���
v�P�ļ���\��!����ڽ[t��D��.}��A��HD���޾�����
�      �iþGD��)o���������� �i��-=�[t����R��Tys�m +����s񗼗(;�H�ѻt@�χ!��1j:�O�:4�;�C3;}�>;CED;��F;�H;_{H;��H;��H;V�H;�H;�H;��H;9�H;R�H;��H;�H;��H;R�H;9�H;��H;�H;�H;V�H;��H;��H;_{H;�H;��F;CED;}�>;�C3;4�;�O�:�1j:χ!�t@�H�ѻ�(;�s����m +�Tys��R����[t��-=� �i���������)o��GD��      �(��;l���.}�&ce�jPH���(�o
���ڽ�R����{�4�6�� �$p��\�`�ר�-��JҺ�C^9`��:=�;�}(;t�8;IA;5{E;FiG;�<H;i�H; �H;H�H;�H;N�H;��H;��H;��H;��H;�H;i�H;�H;��H;��H;��H;��H;N�H;�H;H�H; �H;i�H;�<H;FiG;5{E;IA;t�8;�}(;=�;`��:�C^9JҺ-��ר�\�`�$p��� �4�6���{��R����ڽo
���(�jPH�&ce��.}�;l��      �-=�1�9��k/�"�����i��y�Ľ�!��Tys�4�6�#��ɺ��vz����c^��̃$������r:���:7�;�X1;>H=;jwC;WvF;R�G;/eH;m�H;��H;��H;��H;u�H;�H;��H;��H;��H;��H;��H;��H;��H;��H;��H;�H;u�H;��H;��H;��H;m�H;/eH;R�G;WvF;jwC;>H=;�X1;7�;���:��r:���̃$�c^������vz��ɺ�#�4�6�Tys��!��y�Ľi���"���k/�1�9�      �` �j.��m��ڽ�b��gr��O��\�m +�� ��ɺ�<��O*�bͻQ6R��ǅ���:���:ڃ;�);6t8;��@;�)E;�7G;t#H;p�H;c�H;�H;I�H;��H;��H;��H;�H;m�H;�H; �H;>�H; �H;�H;m�H;�H;��H;��H;��H;I�H;�H;c�H;p�H;t#H;�7G;�)E;��@;6t8;�);ڃ;���:��:�ǅ�Q6R�bͻ�O*�<��ɺ�� �m +�\�O��gr���b����ڽm��j.��      �@���R��ڟ�绒�C����_�:�������$p���vz��O*�5ֻfk������09�:_0;�� ;�C3;��=;�C;kF;��G;�[H;H;o�H;%�H;b�H;��H;��H;��H;�H;'�H;��H;n�H;��H;n�H;��H;'�H;�H;��H;��H;��H;b�H;%�H;o�H;H;�[H;��G;kF;�C;��=;�C3;�� ;_0;�:��09���fk�5ֻ�O*��vz�$p����輙��:���_�C��绒�ڟ��R��      ��_�\�<Q��f@�t +��5�����P�ļs�\�`����bͻfk��Iɺ6
7��:�O�:x�;%d.;��:;Z�A;c{E;�MG;q&H;/�H;�H;��H;��H;I�H;n�H;|�H;R�H;�H;��H;*�H;��H;�H;��H;*�H;��H;�H;R�H;|�H;n�H;I�H;��H;��H;�H;/�H;q&H;�MG;c{E;Z�A;��:;%d.;x�;�O�:�:6
7��Iɺfk�bͻ���\�`�s�P�ļ�����5�t +��f@�<Q�\�      &]� �%#�����u�ټ�ɺ������
v��(;�ר�c^��Q6R����6
7����:���:N�;k�*;+8;� @;��D;��F;'�G; eH;��H;��H;ľH;��H;�H;��H;A�H;��H;��H;��H;��H;B�H;u�H;B�H;��H;��H;��H;��H;A�H;��H;�H;��H;ľH;��H;��H; eH;'�G;��F;��D;� @;+8;k�*;N�;���:���:6
7����Q6R�c^��ר��(;��
v������ɺ�u�ټ����%#� �      &p��\x��ע��R��%��o�`��7�F��H�ѻ-��̃$��ǅ���09�:���:�; ~(;�Y6;��>;�C;&HF;�G;DH;s�H;�H;θH;2�H;K�H;2�H;�H;��H;��H;��H;,�H;�H;��H;��H;��H;�H;,�H;��H;��H;��H;�H;2�H;K�H;2�H;θH;�H;s�H;DH;�G;&HF;�C;��>;�Y6; ~(;�;���:�:��09�ǅ�̃$�-��H�ѻF���7�o�`�%���R��ע�\x��      ��I�1�E��(;��O*�����<��@GĻ��t@�JҺ���:�:�O�:N�; ~(;R�5;>;pC;k�E;�bG;k#H;"{H;^�H;I�H;��H;��H;Y�H;��H;:�H;w�H;��H;h�H;��H;Y�H;��H;�H;��H;Y�H;��H;h�H;��H;w�H;:�H;��H;Y�H;��H;��H;I�H;^�H;"{H;k#H;�bG;k�E;pC;>;R�5; ~(;N�;�O�:�:��:���JҺt@���@GĻ�<������O*��(;�1�E�      r�ѻ�ͻP���mG�������d�+�$��Jɺχ!��C^9��r:���:_0;x�;k�*;�Y6;>;n�B;��E;8G;�H;,mH;A�H;m�H;μH;��H;��H;��H;g�H;�H;��H;��H;�H;�H;��H;�H;<�H;�H;��H;�H;�H;��H;��H;�H;g�H;��H;��H;��H;μH;m�H;A�H;,mH;�H;8G;��E;n�B;>;�Y6;k�*;x�;_0;���:��r:�C^9χ!��Jɺ+�$���d����mG��P����ͻ      ��)���$�����������@�\�S���N�9�1j:`��:���:ڃ;�� ;%d.;+8;��>;pC;��E;�(G;��G;>cH;��H;��H;��H;��H;T�H;��H;��H;��H;��H;��H;a�H;��H;w�H;�H;I�H;b�H;I�H;�H;w�H;��H;a�H;��H;��H;��H;��H;��H;T�H;��H;��H;��H;��H;>cH;��G;�(G;��E;pC;��>;+8;%d.;�� ;ڃ;���:`��:�1j:�N�9S��@�\�������������$�      �R�� �#�7�v<^9��:M�X:���:���:�O�:=�;7�;�);�C3;��:;� @;�C;k�E;8G;��G;�_H;��H;?�H;?�H;��H;d�H;Q�H;h�H;w�H;��H;��H;��H;$�H;��H;��H;@�H;{�H;{�H;{�H;@�H;��H;��H;$�H;��H;��H;��H;w�H;h�H;Q�H;d�H;��H;?�H;?�H;��H;�_H;��G;8G;k�E;�C;� @;��:;�C3;�);7�;=�;�O�:���:���:M�X:��:v<^9#�7�� �      [�:���:��:Ѳ�:���:OO�:�z;h';4�;�}(;�X1;6t8;��=;Z�A;��D;&HF;�bG;�H;>cH;��H;m�H;��H;R�H;�H;��H;Y�H;d�H;��H;<�H;��H;��H;��H;l�H;��H;X�H;��H;��H;��H;X�H;��H;l�H;��H;��H;��H;<�H;��H;d�H;Y�H;��H;�H;R�H;��H;m�H;��H;>cH;�H;�bG;&HF;��D;Z�A;��=;6t8;�X1;�}(;4�;h';�z;OO�:���:Ѳ�:��:���:      ��
;��;I�;[;��;6`;�C&;�-;�C3;t�8;>H=;��@;�C;c{E;��F;�G;k#H;,mH;��H;?�H;��H;��H;Y�H;:�H;��H;��H;��H;��H;~�H;�H;4�H;�H;��H;1�H;r�H;��H;��H;��H;r�H;1�H;��H;�H;4�H;�H;~�H;��H;��H;��H;��H;:�H;Y�H;��H;��H;?�H;��H;,mH;k#H;�G;��F;c{E;�C;��@;>H=;t�8;�C3;�-;�C&;6`;��;[;I�;��;      *;��*;�,;�c.;�X1;#�4;E+8;ӊ;;}�>;IA;jwC;�)E;kF;�MG;'�G;DH;"{H;A�H;��H;?�H;R�H;Y�H;��H;�H;�H;w�H;"�H;�H;��H;��H;��H;��H;��H;L�H;��H;��H;��H;��H;��H;L�H;��H;��H;��H;��H;��H;�H;"�H;w�H;�H;�H;��H;Y�H;R�H;?�H;��H;A�H;"{H;DH;'�G;�MG;kF;�)E;jwC;IA;}�>;ӊ;;E+8;#�4;�X1;�c.;�,;��*;      C�:;[�:;��;;'�<;3>;�?;EIA;��B;CED;5{E;WvF;�7G;��G;q&H; eH;s�H;^�H;m�H;��H;��H;�H;:�H;�H;��H;5�H;��H;��H;G�H;��H;~�H;(�H;��H;,�H;l�H;��H;��H;��H;��H;��H;l�H;,�H;��H;(�H;~�H;��H;G�H;��H;��H;5�H;��H;�H;:�H;�H;��H;��H;m�H;^�H;s�H; eH;q&H;��G;�7G;WvF;5{E;CED;��B;EIA;�?;3>;'�<;��;;[�:;      �B;.�B;�C;ՏC;�/D;��D;0�E;�HF;��F;FiG;R�G;t#H;�[H;/�H;��H;�H;I�H;μH;��H;d�H;��H;��H;�H;5�H;��H;��H;�H;T�H;8�H;�H;��H;��H;=�H;��H;��H;��H;��H;��H;��H;��H;=�H;��H;��H;�H;8�H;T�H;�H;��H;��H;5�H;�H;��H;��H;d�H;��H;μH;I�H;�H;��H;/�H;�[H;t#H;R�G;FiG;��F;�HF;0�E;��D;�/D;ՏC;�C;.�B;      UHF;3TF;RvF;F�F;��F;�7G;��G;��G;�H;�<H;/eH;p�H;H;�H;��H;θH;��H;��H;T�H;Q�H;Y�H;��H;w�H;��H;��H;	�H;9�H;�H;��H;R�H;��H;.�H;C�H;}�H;��H;��H;��H;��H;��H;}�H;C�H;.�H;��H;R�H;��H;�H;9�H;	�H;��H;��H;w�H;��H;Y�H;Q�H;T�H;��H;��H;θH;��H;�H;H;p�H;/eH;�<H;�H;��G;��G;�7G;��F;F�F;RvF;3TF;      =�G;��G;/�G;��G;�H;�/H;�KH;?eH;_{H;i�H;m�H;c�H;o�H;��H;ľH;2�H;��H;��H;��H;h�H;d�H;��H;"�H;��H;�H;9�H;�H;��H;[�H;��H;��H;<�H;\�H;�H;��H;��H;��H;��H;��H;�H;\�H;<�H;��H;��H;[�H;��H;�H;9�H;�H;��H;"�H;��H;d�H;h�H;��H;��H;��H;2�H;ľH;��H;o�H;c�H;m�H;i�H;_{H;?eH;�KH;�/H;�H;��G;/�G;��G;      �kH;ZmH;�qH;�xH;r�H;ȊH;�H;ʜH;��H; �H;��H;�H;%�H;��H;��H;K�H;Y�H;��H;��H;w�H;��H;��H;�H;G�H;T�H;�H;��H;B�H;��H;��H;�H;B�H;k�H;l�H;��H;��H;��H;��H;��H;l�H;k�H;B�H;�H;��H;��H;B�H;��H;�H;T�H;G�H;�H;��H;��H;w�H;��H;��H;Y�H;K�H;��H;��H;%�H;�H;��H; �H;��H;ʜH;�H;ȊH;r�H;�xH;�qH;ZmH;      3�H;ϠH;[�H;äH;��H;��H;��H;�H;��H;H�H;��H;I�H;b�H;I�H;�H;2�H;��H;g�H;��H;��H;<�H;~�H;��H;��H;8�H;��H;[�H;��H;��H;�H;6�H;S�H;j�H;k�H;j�H;u�H;u�H;u�H;j�H;k�H;j�H;S�H;6�H;�H;��H;��H;[�H;��H;8�H;��H;��H;~�H;<�H;��H;��H;g�H;��H;2�H;�H;I�H;b�H;I�H;��H;H�H;��H;�H;��H;��H;��H;äH;[�H;ϠH;      ��H;ܶH;��H;7�H;)�H;��H;R�H;N�H;V�H;�H;��H;��H;��H;n�H;��H;�H;:�H;�H;��H;��H;��H;�H;��H;~�H;�H;R�H;��H;��H;�H;+�H;J�H;I�H;X�H;h�H;P�H;b�H;{�H;b�H;P�H;h�H;X�H;I�H;J�H;+�H;�H;��H;��H;R�H;�H;~�H;��H;�H;��H;��H;��H;�H;:�H;�H;��H;n�H;��H;��H;��H;�H;V�H;N�H;R�H;��H;)�H;7�H;��H;ܶH;      h�H;��H;=�H;I�H;��H;.�H;�H;��H;�H;N�H;u�H;��H;��H;|�H;A�H;��H;w�H;��H;��H;��H;��H;4�H;��H;(�H;��H;��H;��H;�H;6�H;J�H;a�H;T�H;E�H;E�H;c�H;U�H;6�H;U�H;c�H;E�H;E�H;T�H;a�H;J�H;6�H;�H;��H;��H;��H;(�H;��H;4�H;��H;��H;��H;��H;w�H;��H;A�H;|�H;��H;��H;u�H;N�H;�H;��H;�H;.�H;��H;I�H;=�H;��H;      ��H;��H;�H;��H;��H;��H;(�H;��H;�H;��H;�H;��H;��H;R�H;��H;��H;��H;��H;a�H;$�H;��H;�H;��H;��H;��H;.�H;<�H;B�H;S�H;I�H;T�H;Z�H;C�H;=�H;O�H;4�H;+�H;4�H;O�H;=�H;C�H;Z�H;T�H;I�H;S�H;B�H;<�H;.�H;��H;��H;��H;�H;��H;$�H;a�H;��H;��H;��H;��H;R�H;��H;��H;�H;��H;�H;��H;(�H;��H;��H;��H;�H;��H;      ��H;��H;�H;��H;)�H;��H;��H;��H;��H;��H;��H;�H;�H;�H;��H;��H;h�H;�H;��H;��H;l�H;��H;��H;,�H;=�H;C�H;\�H;k�H;j�H;X�H;E�H;C�H;G�H;C�H;"�H;#�H;S�H;#�H;"�H;C�H;G�H;C�H;E�H;X�H;j�H;k�H;\�H;C�H;=�H;,�H;��H;��H;l�H;��H;��H;�H;h�H;��H;��H;�H;�H;�H;��H;��H;��H;��H;��H;��H;)�H;��H;�H;��H;      o�H;�H;��H;��H;��H;�H;��H;{�H;9�H;��H;��H;m�H;'�H;��H;��H;,�H;��H;�H;w�H;��H;��H;1�H;L�H;l�H;��H;}�H;�H;l�H;k�H;h�H;E�H;=�H;C�H;-�H;�H;$�H;)�H;$�H;�H;-�H;C�H;=�H;E�H;h�H;k�H;l�H;�H;}�H;��H;l�H;L�H;1�H;��H;��H;w�H;�H;��H;,�H;��H;��H;'�H;m�H;��H;��H;9�H;{�H;��H;�H;��H;��H;��H;�H;      ��H;��H;��H;�H;p�H;��H;@�H;��H;R�H;��H;��H;�H;��H;*�H;��H;�H;Y�H;��H;�H;@�H;X�H;r�H;��H;��H;��H;��H;��H;��H;j�H;P�H;c�H;O�H;"�H;�H;'�H;�H;�H;�H;'�H;�H;"�H;O�H;c�H;P�H;j�H;��H;��H;��H;��H;��H;��H;r�H;X�H;@�H;�H;��H;Y�H;�H;��H;*�H;��H;�H;��H;��H;R�H;��H;@�H;��H;p�H;�H;��H;��H;      (�H;<�H;j�H;��H;��H;-�H;��H;�H;��H;�H;��H; �H;n�H;��H;B�H;��H;��H;�H;I�H;{�H;��H;��H;��H;��H;��H;��H;��H;��H;u�H;b�H;U�H;4�H;#�H;$�H;�H;�H;�H;�H;�H;$�H;#�H;4�H;U�H;b�H;u�H;��H;��H;��H;��H;��H;��H;��H;��H;{�H;I�H;�H;��H;��H;B�H;��H;n�H; �H;��H;�H;��H;�H;��H;-�H;��H;��H;j�H;<�H;      ��H;��H;��H;6�H;~�H;��H;5�H;��H;�H;i�H;��H;>�H;��H;�H;u�H;��H;�H;<�H;b�H;{�H;��H;��H;��H;��H;��H;��H;��H;��H;u�H;{�H;6�H;+�H;S�H;)�H;�H;�H;�H;�H;�H;)�H;S�H;+�H;6�H;{�H;u�H;��H;��H;��H;��H;��H;��H;��H;��H;{�H;b�H;<�H;�H;��H;u�H;�H;��H;>�H;��H;i�H;�H;��H;5�H;��H;~�H;6�H;��H;��H;      (�H;<�H;j�H;��H;��H;-�H;��H;�H;��H;�H;��H; �H;n�H;��H;B�H;��H;��H;�H;I�H;{�H;��H;��H;��H;��H;��H;��H;��H;��H;u�H;b�H;U�H;4�H;#�H;$�H;�H;�H;�H;�H;�H;$�H;#�H;4�H;U�H;b�H;u�H;��H;��H;��H;��H;��H;��H;��H;��H;{�H;I�H;�H;��H;��H;B�H;��H;n�H; �H;��H;�H;��H;�H;��H;-�H;��H;��H;j�H;<�H;      ��H;��H;��H;�H;p�H;��H;@�H;��H;R�H;��H;��H;�H;��H;*�H;��H;�H;Y�H;��H;�H;@�H;X�H;r�H;��H;��H;��H;��H;��H;��H;j�H;P�H;c�H;O�H;"�H;�H;'�H;�H;�H;�H;'�H;�H;"�H;O�H;c�H;P�H;j�H;��H;��H;��H;��H;��H;��H;r�H;X�H;@�H;�H;��H;Y�H;�H;��H;*�H;��H;�H;��H;��H;R�H;��H;@�H;��H;p�H;�H;��H;��H;      o�H;�H;��H;��H;��H;�H;��H;{�H;9�H;��H;��H;m�H;'�H;��H;��H;,�H;��H;�H;w�H;��H;��H;1�H;L�H;l�H;��H;}�H;�H;l�H;k�H;h�H;E�H;=�H;C�H;-�H;�H;$�H;)�H;$�H;�H;-�H;C�H;=�H;E�H;h�H;k�H;l�H;�H;}�H;��H;l�H;L�H;1�H;��H;��H;w�H;�H;��H;,�H;��H;��H;'�H;m�H;��H;��H;9�H;{�H;��H;�H;��H;��H;��H;�H;      ��H;��H;�H;��H;)�H;��H;��H;��H;��H;��H;��H;�H;�H;�H;��H;��H;h�H;�H;��H;��H;l�H;��H;��H;,�H;=�H;C�H;\�H;k�H;j�H;X�H;E�H;C�H;G�H;C�H;"�H;#�H;S�H;#�H;"�H;C�H;G�H;C�H;E�H;X�H;j�H;k�H;\�H;C�H;=�H;,�H;��H;��H;l�H;��H;��H;�H;h�H;��H;��H;�H;�H;�H;��H;��H;��H;��H;��H;��H;)�H;��H;�H;��H;      ��H;��H;�H;��H;��H;��H;(�H;��H;�H;��H;�H;��H;��H;R�H;��H;��H;��H;��H;a�H;$�H;��H;�H;��H;��H;��H;.�H;<�H;B�H;S�H;I�H;T�H;Z�H;C�H;=�H;O�H;4�H;+�H;4�H;O�H;=�H;C�H;Z�H;T�H;I�H;S�H;B�H;<�H;.�H;��H;��H;��H;�H;��H;$�H;a�H;��H;��H;��H;��H;R�H;��H;��H;�H;��H;�H;��H;(�H;��H;��H;��H;�H;��H;      h�H;��H;=�H;I�H;��H;.�H;�H;��H;�H;N�H;u�H;��H;��H;|�H;A�H;��H;w�H;��H;��H;��H;��H;4�H;��H;(�H;��H;��H;��H;�H;6�H;J�H;a�H;T�H;E�H;E�H;c�H;U�H;6�H;U�H;c�H;E�H;E�H;T�H;a�H;J�H;6�H;�H;��H;��H;��H;(�H;��H;4�H;��H;��H;��H;��H;w�H;��H;A�H;|�H;��H;��H;u�H;N�H;�H;��H;�H;.�H;��H;I�H;=�H;��H;      ��H;ܶH;��H;7�H;)�H;��H;R�H;N�H;V�H;�H;��H;��H;��H;n�H;��H;�H;:�H;�H;��H;��H;��H;�H;��H;~�H;�H;R�H;��H;��H;�H;+�H;J�H;I�H;X�H;h�H;P�H;b�H;{�H;b�H;P�H;h�H;X�H;I�H;J�H;+�H;�H;��H;��H;R�H;�H;~�H;��H;�H;��H;��H;��H;�H;:�H;�H;��H;n�H;��H;��H;��H;�H;V�H;N�H;R�H;��H;)�H;7�H;��H;ܶH;      3�H;ϠH;[�H;äH;��H;��H;��H;�H;��H;H�H;��H;I�H;b�H;I�H;�H;2�H;��H;g�H;��H;��H;<�H;~�H;��H;��H;8�H;��H;[�H;��H;��H;�H;6�H;S�H;j�H;k�H;j�H;u�H;u�H;u�H;j�H;k�H;j�H;S�H;6�H;�H;��H;��H;[�H;��H;8�H;��H;��H;~�H;<�H;��H;��H;g�H;��H;2�H;�H;I�H;b�H;I�H;��H;H�H;��H;�H;��H;��H;��H;äH;[�H;ϠH;      �kH;ZmH;�qH;�xH;r�H;ȊH;�H;ʜH;��H; �H;��H;�H;%�H;��H;��H;K�H;Y�H;��H;��H;w�H;��H;��H;�H;G�H;T�H;�H;��H;B�H;��H;��H;�H;B�H;k�H;l�H;��H;��H;��H;��H;��H;l�H;k�H;B�H;�H;��H;��H;B�H;��H;�H;T�H;G�H;�H;��H;��H;w�H;��H;��H;Y�H;K�H;��H;��H;%�H;�H;��H; �H;��H;ʜH;�H;ȊH;r�H;�xH;�qH;ZmH;      =�G;��G;/�G;��G;�H;�/H;�KH;?eH;_{H;i�H;m�H;c�H;o�H;��H;ľH;2�H;��H;��H;��H;h�H;d�H;��H;"�H;��H;�H;9�H;�H;��H;[�H;��H;��H;<�H;\�H;�H;��H;��H;��H;��H;��H;�H;\�H;<�H;��H;��H;[�H;��H;�H;9�H;�H;��H;"�H;��H;d�H;h�H;��H;��H;��H;2�H;ľH;��H;o�H;c�H;m�H;i�H;_{H;?eH;�KH;�/H;�H;��G;/�G;��G;      UHF;3TF;RvF;F�F;��F;�7G;��G;��G;�H;�<H;/eH;p�H;H;�H;��H;θH;��H;��H;T�H;Q�H;Y�H;��H;w�H;��H;��H;	�H;9�H;�H;��H;R�H;��H;.�H;C�H;}�H;��H;��H;��H;��H;��H;}�H;C�H;.�H;��H;R�H;��H;�H;9�H;	�H;��H;��H;w�H;��H;Y�H;Q�H;T�H;��H;��H;θH;��H;�H;H;p�H;/eH;�<H;�H;��G;��G;�7G;��F;F�F;RvF;3TF;      �B;.�B;�C;ՏC;�/D;��D;0�E;�HF;��F;FiG;R�G;t#H;�[H;/�H;��H;�H;I�H;μH;��H;d�H;��H;��H;�H;5�H;��H;��H;�H;T�H;8�H;�H;��H;��H;=�H;��H;��H;��H;��H;��H;��H;��H;=�H;��H;��H;�H;8�H;T�H;�H;��H;��H;5�H;�H;��H;��H;d�H;��H;μH;I�H;�H;��H;/�H;�[H;t#H;R�G;FiG;��F;�HF;0�E;��D;�/D;ՏC;�C;.�B;      C�:;[�:;��;;'�<;3>;�?;EIA;��B;CED;5{E;WvF;�7G;��G;q&H; eH;s�H;^�H;m�H;��H;��H;�H;:�H;�H;��H;5�H;��H;��H;G�H;��H;~�H;(�H;��H;,�H;l�H;��H;��H;��H;��H;��H;l�H;,�H;��H;(�H;~�H;��H;G�H;��H;��H;5�H;��H;�H;:�H;�H;��H;��H;m�H;^�H;s�H; eH;q&H;��G;�7G;WvF;5{E;CED;��B;EIA;�?;3>;'�<;��;;[�:;      *;��*;�,;�c.;�X1;#�4;E+8;ӊ;;}�>;IA;jwC;�)E;kF;�MG;'�G;DH;"{H;A�H;��H;?�H;R�H;Y�H;��H;�H;�H;w�H;"�H;�H;��H;��H;��H;��H;��H;L�H;��H;��H;��H;��H;��H;L�H;��H;��H;��H;��H;��H;�H;"�H;w�H;�H;�H;��H;Y�H;R�H;?�H;��H;A�H;"{H;DH;'�G;�MG;kF;�)E;jwC;IA;}�>;ӊ;;E+8;#�4;�X1;�c.;�,;��*;      ��
;��;I�;[;��;6`;�C&;�-;�C3;t�8;>H=;��@;�C;c{E;��F;�G;k#H;,mH;��H;?�H;��H;��H;Y�H;:�H;��H;��H;��H;��H;~�H;�H;4�H;�H;��H;1�H;r�H;��H;��H;��H;r�H;1�H;��H;�H;4�H;�H;~�H;��H;��H;��H;��H;:�H;Y�H;��H;��H;?�H;��H;,mH;k#H;�G;��F;c{E;�C;��@;>H=;t�8;�C3;�-;�C&;6`;��;[;I�;��;      [�:���:��:Ѳ�:���:OO�:�z;h';4�;�}(;�X1;6t8;��=;Z�A;��D;&HF;�bG;�H;>cH;��H;m�H;��H;R�H;�H;��H;Y�H;d�H;��H;<�H;��H;��H;��H;l�H;��H;X�H;��H;��H;��H;X�H;��H;l�H;��H;��H;��H;<�H;��H;d�H;Y�H;��H;�H;R�H;��H;m�H;��H;>cH;�H;�bG;&HF;��D;Z�A;��=;6t8;�X1;�}(;4�;h';�z;OO�:���:Ѳ�:��:���:      �R�� �#�7�v<^9��:M�X:���:���:�O�:=�;7�;�);�C3;��:;� @;�C;k�E;8G;��G;�_H;��H;?�H;?�H;��H;d�H;Q�H;h�H;w�H;��H;��H;��H;$�H;��H;��H;@�H;{�H;{�H;{�H;@�H;��H;��H;$�H;��H;��H;��H;w�H;h�H;Q�H;d�H;��H;?�H;?�H;��H;�_H;��G;8G;k�E;�C;� @;��:;�C3;�);7�;=�;�O�:���:���:M�X:��:v<^9#�7�� �      ��)���$�����������@�\�S���N�9�1j:`��:���:ڃ;�� ;%d.;+8;��>;pC;��E;�(G;��G;>cH;��H;��H;��H;��H;T�H;��H;��H;��H;��H;��H;a�H;��H;w�H;�H;I�H;b�H;I�H;�H;w�H;��H;a�H;��H;��H;��H;��H;��H;T�H;��H;��H;��H;��H;>cH;��G;�(G;��E;pC;��>;+8;%d.;�� ;ڃ;���:`��:�1j:�N�9S��@�\�������������$�      r�ѻ�ͻP���mG�������d�+�$��Jɺχ!��C^9��r:���:_0;x�;k�*;�Y6;>;n�B;��E;8G;�H;,mH;A�H;m�H;μH;��H;��H;��H;g�H;�H;��H;��H;�H;�H;��H;�H;<�H;�H;��H;�H;�H;��H;��H;�H;g�H;��H;��H;��H;μH;m�H;A�H;,mH;�H;8G;��E;n�B;>;�Y6;k�*;x�;_0;���:��r:�C^9χ!��Jɺ+�$���d����mG��P����ͻ      ��I�1�E��(;��O*�����<��@GĻ��t@�JҺ���:�:�O�:N�; ~(;R�5;>;pC;k�E;�bG;k#H;"{H;^�H;I�H;��H;��H;Y�H;��H;:�H;w�H;��H;h�H;��H;Y�H;��H;�H;��H;Y�H;��H;h�H;��H;w�H;:�H;��H;Y�H;��H;��H;I�H;^�H;"{H;k#H;�bG;k�E;pC;>;R�5; ~(;N�;�O�:�:��:���JҺt@���@GĻ�<������O*��(;�1�E�      &p��\x��ע��R��%��o�`��7�F��H�ѻ-��̃$��ǅ���09�:���:�; ~(;�Y6;��>;�C;&HF;�G;DH;s�H;�H;θH;2�H;K�H;2�H;�H;��H;��H;��H;,�H;�H;��H;��H;��H;�H;,�H;��H;��H;��H;�H;2�H;K�H;2�H;θH;�H;s�H;DH;�G;&HF;�C;��>;�Y6; ~(;�;���:�:��09�ǅ�̃$�-��H�ѻF���7�o�`�%���R��ע�\x��      &]� �%#�����u�ټ�ɺ������
v��(;�ר�c^��Q6R����6
7����:���:N�;k�*;+8;� @;��D;��F;'�G; eH;��H;��H;ľH;��H;�H;��H;A�H;��H;��H;��H;��H;B�H;u�H;B�H;��H;��H;��H;��H;A�H;��H;�H;��H;ľH;��H;��H; eH;'�G;��F;��D;� @;+8;k�*;N�;���:���:6
7����Q6R�c^��ר��(;��
v������ɺ�u�ټ����%#� �      ��_�\�<Q��f@�t +��5�����P�ļs�\�`����bͻfk��Iɺ6
7��:�O�:x�;%d.;��:;Z�A;c{E;�MG;q&H;/�H;�H;��H;��H;I�H;n�H;|�H;R�H;�H;��H;*�H;��H;�H;��H;*�H;��H;�H;R�H;|�H;n�H;I�H;��H;��H;�H;/�H;q&H;�MG;c{E;Z�A;��:;%d.;x�;�O�:�:6
7��Iɺfk�bͻ���\�`�s�P�ļ�����5�t +��f@�<Q�\�      �@���R��ڟ�绒�C����_�:�������$p���vz��O*�5ֻfk������09�:_0;�� ;�C3;��=;�C;kF;��G;�[H;H;o�H;%�H;b�H;��H;��H;��H;�H;'�H;��H;n�H;��H;n�H;��H;'�H;�H;��H;��H;��H;b�H;%�H;o�H;H;�[H;��G;kF;�C;��=;�C3;�� ;_0;�:��09���fk�5ֻ�O*��vz�$p����輙��:���_�C��绒�ڟ��R��      �` �j.��m��ڽ�b��gr��O��\�m +�� ��ɺ�<��O*�bͻQ6R��ǅ���:���:ڃ;�);6t8;��@;�)E;�7G;t#H;p�H;c�H;�H;I�H;��H;��H;��H;�H;m�H;�H; �H;>�H; �H;�H;m�H;�H;��H;��H;��H;I�H;�H;c�H;p�H;t#H;�7G;�)E;��@;6t8;�);ڃ;���:��:�ǅ�Q6R�bͻ�O*�<��ɺ�� �m +�\�O��gr���b����ڽm��j.��      �-=�1�9��k/�"�����i��y�Ľ�!��Tys�4�6�#��ɺ��vz����c^��̃$������r:���:7�;�X1;>H=;jwC;WvF;R�G;/eH;m�H;��H;��H;��H;u�H;�H;��H;��H;��H;��H;��H;��H;��H;��H;��H;�H;u�H;��H;��H;��H;m�H;/eH;R�G;WvF;jwC;>H=;�X1;7�;���:��r:���̃$�c^������vz��ɺ�#�4�6�Tys��!��y�Ľi���"���k/�1�9�      �(��;l���.}�&ce�jPH���(�o
���ڽ�R����{�4�6�� �$p��\�`�ר�-��JҺ�C^9`��:=�;�}(;t�8;IA;5{E;FiG;�<H;i�H; �H;H�H;�H;N�H;��H;��H;��H;��H;�H;i�H;�H;��H;��H;��H;��H;N�H;�H;H�H; �H;i�H;�<H;FiG;5{E;IA;t�8;�}(;=�;`��:�C^9JҺ-��ר�\�`�$p��� �4�6���{��R����ڽo
���(�jPH�&ce��.}�;l��      �iþGD��)o���������� �i��-=�[t����R��Tys�m +����s񗼗(;�H�ѻt@�χ!��1j:�O�:4�;�C3;}�>;CED;��F;�H;_{H;��H;��H;V�H;�H;�H;��H;9�H;R�H;��H;�H;��H;R�H;9�H;��H;�H;�H;V�H;��H;��H;_{H;�H;��F;CED;}�>;�C3;4�;�O�:�1j:χ!�t@�H�ѻ�(;�s����m +�Tys��R����[t��-=� �i���������)o��GD��      ���
������޾HD���A���.}��D�[t���ڽ�!��\����P�ļ�
v�F�����Jɺ�N�9���:h';�-;ӊ;;��B;�HF;��G;?eH;ʜH;�H;N�H;��H;��H;��H;{�H;��H;�H;��H;�H;��H;{�H;��H;��H;��H;N�H;�H;ʜH;?eH;��G;�HF;��B;ӊ;;�-;h';���:�N�9�Jɺ��F���
v�P�ļ���\��!����ڽ[t��D��.}��A��HD���޾�����
�      ��7�Õ3��f'���\���о�����.}��-=�o
�y�ĽO��:����������7�@GĻ+�$�S�����:�z;�C&;E+8;EIA;0�E;��G;�KH;�H;��H;R�H;�H;(�H;��H;��H;@�H;��H;5�H;��H;@�H;��H;��H;(�H;�H;R�H;��H;�H;�KH;��G;0�E;EIA;E+8;�C&;�z;���:S��+�$�@GĻ�7���������:�O��y�Ľo
��-=��.}������о�\����f'�Õ3�      Io�PXi�s"Y���@�@�#��
��о�A�� �i���(�i��gr����_��5��ɺ�o�`��<����d�@�\�M�X:OO�:6`;#�4;�?;��D;�7G;�/H;ȊH;��H;��H;.�H;��H;��H;�H;��H;-�H;��H;-�H;��H;�H;��H;��H;.�H;��H;��H;ȊH;�/H;�7G;��D;�?;#�4;6`;OO�:M�X:@�\���d��<��o�`��ɺ��5���_�gr��i����(� �i��A���о�
�@�#���@�s"Y�PXi�      &����������Io��!J�@�#��\��HD������jPH�����b��C��t +�u�ټ%��������������:���:��;�X1;3>;�/D;��F;�H;r�H;��H;)�H;��H;��H;)�H;��H;p�H;��H;~�H;��H;p�H;��H;)�H;��H;��H;)�H;��H;r�H;�H;��F;�/D;3>;�X1;��;���:��:����������%��u�ټt +�C���b�����jPH�����HD���\��@�#��!J�Io��������      2^������b���Io���@���޾����&ce�"����ڽ绒��f@������R���O*�mG�����v<^9Ѳ�:[;�c.;'�<;ՏC;F�F;��G;�xH;äH;7�H;I�H;��H;��H;��H;�H;��H;6�H;��H;�H;��H;��H;��H;I�H;7�H;äH;�xH;��G;F�F;ՏC;'�<;�c.;[;Ѳ�:v<^9���mG���O*��R�������f@�绒���ڽ"��&ce������޾���@�Io�b�������      �aǿ֊¿���������s"Y��f'�����)o���.}��k/�m��ڟ�<Q�%#�ע��(;�P������#�7���:I�;�,;��;;�C;RvF;/�G;�qH;[�H;��H;=�H;�H;�H;��H;��H;j�H;��H;j�H;��H;��H;�H;�H;=�H;��H;[�H;�qH;/�G;RvF;�C;��;;�,;I�;��:#�7����P����(;�ע�%#�<Q�ڟ�m���k/��.}�)o�������f'�s"Y����������֊¿      %�ֿ5pѿ֊¿������PXi�Õ3��
�GD��;l��1�9�j.���R��\� �\x��1�E��ͻ��$�� ����:��;��*;[�:;.�B;3TF;��G;ZmH;ϠH;ܶH;��H;��H;��H;�H;��H;<�H;��H;<�H;��H;�H;��H;��H;��H;ܶH;ϠH;ZmH;��G;3TF;.�B;[�:;��*;��;���:� ���$��ͻ1�E�\x�� �\��R��j.��1�9�;l��GD���
�Õ3�PXi�������֊¿5pѿ      ���$������꿥�ſ�ޞ�3s��2�/����� j���nHͽ������'�B<ͼ��n������Q^�0.��:�V;�R%;~n8;��A;mCF;�H;��H;��H;��H;L�H;>�H;C�H;��H;��H;��H;+�H;��H;��H;��H;C�H;>�H;L�H;��H;��H;��H;�H;mCF;��A;~n8;�R%;�V;�:0.��Q^�������n�B<ͼ��'�����nHͽ�� j���/����2�3s��ޞ���ſ������$�      $��������~�����cm�L�-�����Fh��Ide�-�̪ɽ�v��#�$���ɼ�mj�o����X�7��mĆ:�w;i�%;M�8;B;{QF;H;5�H;U�H;�H;p�H;B�H;5�H;��H;��H;��H;$�H;��H;��H;��H;5�H;B�H;p�H;�H;U�H;5�H;H;{QF;B;M�8;i�%;�w;mĆ:7���X�o����mj���ɼ#�$��v��̪ɽ-�Ide�Fh������L�-�cm����~���忖����      ������{���ԿBw�����/�\��"����b��M0X�}���;����w����������]�X��VF�0��nȒ:0�;^�';׎9;1oB;�yF;� H;��H;7�H;�H;��H;F�H;:�H;��H;��H;��H;�H;��H;��H;��H;:�H;F�H;��H;�H;7�H;��H;� H;�yF;1oB;׎9;^�';0�;nȒ:0��VF�X�黼�]����������w��;��}��M0X�b������"�/�\����Bw���Կ{�𿖏�      ������Կp���ޞ�RF�]�C�$E��;�I��sD�|�"��]�c�y��֯���J�P�ѻ]�)���K����:Q�
;M*;��:;�C;�F;�7H;Z�H;��H;w�H;��H;>�H;9�H;��H;��H;��H;��H;��H;��H;��H;9�H;>�H;��H;w�H;��H;Z�H;�7H;�F;�C;��:;M*;Q�
;���:��K�]�)�P�ѻ��J��֯�y�]�c�"��|�sD��I���;$E�]�C�RF��ޞ�p���Կ��      ��ſ~��Bw���ޞ�|���3�W�,�%�����^ɰ��|x�\{+�ű����J��  �Ҷ��n�1�f����+�
9q�:�;4�-;��<;��C;�G;�SH;Q�H;��H;��H;��H;V�H;2�H;��H;��H;��H;��H;��H;��H;��H;2�H;V�H;��H;��H;��H;Q�H;�SH;�G;��C;��<;4�-;�;q�:
9�+�f���n�1�Ҷ���  ��J���ű�\{+��|x�^ɰ�����,�%�3�W�|����ޞ�Bw��~��      �ޞ�������RF�3�W�M�-���4Kɾ�G����O�z��ƽ����Ȅ-���ۼㄼL4�[ǐ�-ж��Z:n��:�;ʕ1;
c>;{�D;�[G;KrH;��H;i�H;e�H;'�H;u�H;)�H;h�H;��H;|�H;��H;|�H;��H;h�H;)�H;u�H;'�H;e�H;i�H;��H;KrH;�[G;{�D;
c>;ʕ1;�;n��:�Z:-ж�[ǐ�L4�ㄼ��ۼȄ-�����ƽz����O��G��4Kɾ��M�-�3�W�RF�������      3s�cm�/�\�]�C�,�%����TҾa����i��C(����UP����[�x������Y�l���X���<���k:���:)� ;�5;ZQ@;otE;�G;9�H;L�H;��H;�H;I�H;l�H;$�H;c�H;s�H;W�H;��H;W�H;s�H;c�H;$�H;l�H;I�H;�H;��H;L�H;9�H;�G;otE;ZQ@;�5;)� ;���:��k:��<��X�l����Y����x���[�UP����콡C(���i�a���TҾ��,�%�]�C�/�\�cm�      �2�L�-��"�$E�����4Kɾa��w�s�.�5�y�k㻽�v��z0��;��+��-�*�S����6�CjS� L�:��	;��(;5�9;�.B;�CF;YH;ԪH;��H;��H;��H;w�H;��H;�H;0�H;C�H;<�H;Y�H;<�H;C�H;0�H;�H;��H;w�H;��H;��H;��H;ԪH;YH;�CF;�.B;5�9;��(;��	; L�:CjS��6�S���-�*��+���;�z0��v��k㻽y�.�5�w�s�a��4Kɾ����$E��"�L�-�      /�����������;^ɰ��G����i�.�5��	�ĪɽR����J�p���沼��]�J���V
x��
��k:5��:v;��/;�,=;��C;N�F;#HH;��H;(�H;��H;#�H;��H;��H;��H;�H;�H;�H;$�H;�H;�H;�H;��H;��H;��H;#�H;��H;(�H;��H;#HH;N�F;��C;�,=;��/;v;5��:k:�
��V
x�J�����]��沼p���J�R���Īɽ�	�.�5���i��G��^ɰ��;��徨���      ��Fh��b���I���|x���O��C(�y�Īɽ����JDX�D��'<ͼㄼ�X!�t��hX��K����:�x;7�#;$H6;IQ@;�OE;��G;��H;��H;1�H;��H;��H;��H;v�H;��H;��H;��H;��H;��H;��H;��H;��H;��H;v�H;��H;��H;��H;1�H;��H;��H;��G;�OE;IQ@;$H6;7�#;�x;���:�K�hX�t���X!�ㄼ'<ͼD��JDX�����Īɽy��C(���O��|x��I��b��Fh��       j�Ide�M0X�sD�\{+�z�����k㻽R���JDX������ۼо����;�>ۻ�X���y�<<":I��:��;��-;��;;�B;�yF;�H;��H;|�H;&�H;��H;��H;��H;m�H;��H;��H;��H;��H;z�H;��H;��H;��H;��H;m�H;��H;��H;��H;&�H;|�H;��H;�H;�yF;�B;��;;��-;��;I��:<<":��y��X�>ۻ��;�о����ۼ���JDX�R���k㻽���z��\{+�sD�M0X�Ide�      ��-�}��|�ű�ƽUP���v���J�D����ۼ��v�J������+���sѺ&
9fL�:�;�$;#�5;�?;��D;j[G;eH;��H;��H;��H;��H;!�H;��H;T�H;n�H;Y�H;T�H;a�H;7�H;a�H;T�H;Y�H;n�H;T�H;��H;!�H;��H;��H;��H;��H;eH;j[G;��D;�?;#�5;�$;�;fL�:&
9�sѺ�+������v�J�����ۼD���J��v��UP��ƽű�|�}��-�      nHͽ̪ɽ�;��"����������[�z0�p��'<ͼо��v�J���k��+��(����:�`�:|�;�/;�K<; C;9lF;��G;�H;
�H;�H;�H;A�H;T�H;��H;%�H;/�H;�H;�H;�H;��H;�H;�H;�H;/�H;%�H;��H;T�H;A�H;�H;�H;
�H;�H;��G;9lF; C;�K<;�/;|�;�`�:���:�(�+�k����v�J�о��'<ͼp��z0���[�������"���;��̪ɽ      �����v����w�]�c��J�Ȅ-�x��;缈沼ㄼ��;�����k��66�h��K<Q:֣�:�h;M*;��8;��@;�OE;�tG;DhH;��H;��H;�H;#�H;��H;y�H;��H;��H;��H;��H;��H;��H;��H;��H;��H;��H;��H;��H;��H;y�H;��H;#�H;�H;��H;��H;DhH;�tG;�OE;��@;��8;M*;�h;֣�:K<Q:h��66�k��������;�ㄼ�沼�;�x�Ȅ-��J�]�c���w��v��      ��'�#�$����y��  ���ۼ����+����]��X!�>ۻ�+��+�h���>:\��:@�;Z�%;	�5;��>;�'D;�F;� H;8�H;[�H;��H;��H;��H;��H;k�H;��H;��H;��H;��H;g�H;K�H;m�H;K�H;g�H;��H;��H;��H;��H;k�H;��H;��H;��H;��H;[�H;8�H;� H;�F;�'D;��>;	�5;Z�%;@�;\��:�>:h��+��+��>ۻ�X!���]��+�������ۼ�  �y����#�$�      B<ͼ��ɼ�����֯�Ҷ��ㄼ��Y�-�*�J���t���X��sѺ�(�K<Q:\��:��
;u�#;��3;�b=;#C;3CF;�G;�H;��H;�H;8�H;��H;W�H;!�H;d�H;��H;b�H;5�H;O�H;	�H;��H;�H;��H;	�H;O�H;5�H;b�H;��H;d�H;!�H;W�H;��H;8�H;�H;��H;�H;�G;3CF;#C;�b=;��3;u�#;��
;\��:K<Q:�(��sѺ�X�t��J���-�*���Y�ㄼҶ���֯�������ɼ      ��n��mj���]���J�n�1�L4�l��S���V
x�hX���y�&
9���:֣�:@�;u�#;v�2;�<;�oB;7�E;��G;�dH;��H;8�H;��H;��H;��H;��H;9�H;F�H;7�H;�H;��H;��H;��H;��H;��H;��H;��H;��H;��H;�H;7�H;F�H;9�H;��H;��H;��H;��H;8�H;��H;�dH;��G;7�E;�oB;�<;v�2;u�#;@�;֣�:���:&
9��y�hX�V
x�S���l��L4�n�1���J���]��mj�      ����o���X��P�ѻf���[ǐ��X��6��
���K�<<":fL�:�`�:�h;Z�%;��3;�<;Y/B;��E;�[G;�GH;N�H;��H;a�H;�H;7�H;=�H;��H;�H;�H;��H;��H;��H;]�H;O�H;K�H;'�H;K�H;O�H;]�H;��H;��H;��H;�H;�H;��H;=�H;7�H;�H;a�H;��H;N�H;�GH;�[G;��E;Y/B;�<;��3;Z�%;�h;�`�:fL�:<<":�K��
���6��X�[ǐ�f���P�ѻX��o���      �Q^��X�VF�]�)��+�-ж���<�CjS�k:���:I��:�;|�;M*;	�5;�b=;�oB;��E;�IG;\7H;s�H;��H;�H;-�H;��H;��H;��H;��H;��H;��H;��H;t�H;P�H;��H;��H;��H;��H;��H;��H;��H;P�H;t�H;��H;��H;��H;��H;��H;��H;��H;-�H;�H;��H;s�H;\7H;�IG;��E;�oB;�b=;	�5;M*;|�;�;I��:���:k:CjS���<�-ж��+�]�)�VF��X�      0.�7��0�깤�K�
9�Z:��k: L�:5��:�x;��;�$;�/;��8;��>;#C;7�E;�[G;\7H;̤H;�H;&�H;��H;5�H;��H;P�H;��H;��H;��H;z�H;5�H;�H;��H;��H;��H;��H;u�H;��H;��H;��H;��H;�H;5�H;z�H;��H;��H;��H;P�H;��H;5�H;��H;&�H;�H;̤H;\7H;�[G;7�E;#C;��>;��8;�/;�$;��;�x;5��: L�:��k:�Z:
9��K�0��7��      �:mĆ:nȒ:���:q�:n��:���:��	;v;7�#;��-;#�5;�K<;��@;�'D;3CF;��G;�GH;s�H;�H;��H;O�H;��H;\�H;"�H;��H;��H;��H;[�H;�H;��H;��H;m�H;[�H;)�H;�H;�H;�H;)�H;[�H;m�H;��H;��H;�H;[�H;��H;��H;��H;"�H;\�H;��H;O�H;��H;�H;s�H;�GH;��G;3CF;�'D;��@;�K<;#�5;��-;7�#;v;��	;���:n��:q�:���:nȒ:mĆ:      �V;�w;0�;Q�
;�;�;)� ;��(;��/;$H6;��;;�?; C;�OE;�F;�G;�dH;N�H;��H;&�H;O�H;��H;0�H;��H;e�H;�H;��H;a�H;��H;��H;��H;A�H;�H;�H;��H;��H;��H;��H;��H;�H;�H;A�H;��H;��H;��H;a�H;��H;�H;e�H;��H;0�H;��H;O�H;&�H;��H;N�H;�dH;�G;�F;�OE; C;�?;��;;$H6;��/;��(;)� ;�;�;Q�
;0�;�w;      �R%;i�%;^�';M*;4�-;ʕ1;�5;5�9;�,=;IQ@;�B;��D;9lF;�tG;� H;�H;��H;��H;�H;��H;��H;0�H;�H;a�H;��H;r�H;5�H;��H;��H;��H;�H;��H;��H;��H;|�H;e�H;L�H;e�H;|�H;��H;��H;��H;�H;��H;��H;��H;5�H;r�H;��H;a�H;�H;0�H;��H;��H;�H;��H;��H;�H;� H;�tG;9lF;��D;�B;IQ@;�,=;5�9;�5;ʕ1;4�-;M*;^�';i�%;      ~n8;M�8;׎9;��:;��<;
c>;ZQ@;�.B;��C;�OE;�yF;j[G;��G;DhH;8�H;��H;8�H;a�H;-�H;5�H;\�H;��H;a�H;k�H;i�H;D�H;��H;��H;e�H;	�H;��H;��H;Y�H;(�H;"�H;�H;��H;�H;"�H;(�H;Y�H;��H;��H;	�H;e�H;��H;��H;D�H;i�H;k�H;a�H;��H;\�H;5�H;-�H;a�H;8�H;��H;8�H;DhH;��G;j[G;�yF;�OE;��C;�.B;ZQ@;
c>;��<;��:;׎9;M�8;      ��A;B;1oB;�C;��C;{�D;otE;�CF;N�F;��G;�H;eH;�H;��H;[�H;�H;��H;�H;��H;��H;"�H;e�H;��H;i�H;-�H;��H;��H;i�H; �H;��H;r�H;@�H;
�H;��H;��H;��H;��H;��H;��H;��H;
�H;@�H;r�H;��H; �H;i�H;��H;��H;-�H;i�H;��H;e�H;"�H;��H;��H;�H;��H;�H;[�H;��H;�H;eH;�H;��G;N�F;�CF;otE;{�D;��C;�C;1oB;B;      mCF;{QF;�yF;�F;�G;�[G;�G;YH;#HH;��H;��H;��H;
�H;��H;��H;8�H;��H;7�H;��H;P�H;��H;�H;r�H;D�H;��H;��H;_�H;��H;��H;`�H;�H;��H;��H;��H;o�H;\�H;n�H;\�H;o�H;��H;��H;��H;�H;`�H;��H;��H;_�H;��H;��H;D�H;r�H;�H;��H;P�H;��H;7�H;��H;8�H;��H;��H;
�H;��H;��H;��H;#HH;YH;�G;�[G;�G;�F;�yF;{QF;      �H;H;� H;�7H;�SH;KrH;9�H;ԪH;��H;��H;|�H;��H;�H;�H;��H;��H;��H;=�H;��H;��H;��H;��H;5�H;��H;��H;_�H;��H;��H;H�H;�H;��H;��H;b�H;C�H;(�H;�H;�H;�H;(�H;C�H;b�H;��H;��H;�H;H�H;��H;��H;_�H;��H;��H;5�H;��H;��H;��H;��H;=�H;��H;��H;��H;�H;�H;��H;|�H;��H;��H;ԪH;9�H;KrH;�SH;�7H;� H;H;      ��H;5�H;��H;Z�H;Q�H;��H;L�H;��H;(�H;1�H;&�H;��H;�H;#�H;��H;W�H;��H;��H;��H;��H;��H;a�H;��H;��H;i�H;��H;��H;W�H;�H;��H;u�H;F�H; �H;��H;��H;��H;��H;��H;��H;��H; �H;F�H;u�H;��H;�H;W�H;��H;��H;i�H;��H;��H;a�H;��H;��H;��H;��H;��H;W�H;��H;#�H;�H;��H;&�H;1�H;(�H;��H;L�H;��H;Q�H;Z�H;��H;5�H;      ��H;U�H;7�H;��H;��H;i�H;��H;��H;��H;��H;��H;��H;A�H;��H;��H;!�H;9�H;�H;��H;��H;[�H;��H;��H;e�H; �H;��H;H�H;�H;��H;k�H;7�H;��H;��H;��H;��H;��H;�H;��H;��H;��H;��H;��H;7�H;k�H;��H;�H;H�H;��H; �H;e�H;��H;��H;[�H;��H;��H;�H;9�H;!�H;��H;��H;A�H;��H;��H;��H;��H;��H;��H;i�H;��H;��H;7�H;U�H;      ��H;�H;�H;w�H;��H;e�H;�H;��H;#�H;��H;��H;!�H;T�H;y�H;k�H;d�H;F�H;�H;��H;z�H;�H;��H;��H;	�H;��H;`�H;�H;��H;k�H;-�H;��H;��H;��H;��H;c�H;K�H;A�H;K�H;c�H;��H;��H;��H;��H;-�H;k�H;��H;�H;`�H;��H;	�H;��H;��H;�H;z�H;��H;�H;F�H;d�H;k�H;y�H;T�H;!�H;��H;��H;#�H;��H;�H;e�H;��H;w�H;�H;�H;      L�H;p�H;��H;��H;��H;'�H;I�H;w�H;��H;��H;��H;��H;��H;��H;��H;��H;7�H;��H;��H;5�H;��H;��H;�H;��H;r�H;�H;��H;u�H;7�H;��H;��H;��H;w�H;?�H;�H;'�H;(�H;'�H;�H;?�H;w�H;��H;��H;��H;7�H;u�H;��H;�H;r�H;��H;�H;��H;��H;5�H;��H;��H;7�H;��H;��H;��H;��H;��H;��H;��H;��H;w�H;I�H;'�H;��H;��H;��H;p�H;      >�H;B�H;F�H;>�H;V�H;u�H;l�H;��H;��H;v�H;m�H;T�H;%�H;��H;��H;b�H;�H;��H;t�H;�H;��H;A�H;��H;��H;@�H;��H;��H;F�H;��H;��H;��H;_�H;A�H;�H;��H;��H;��H;��H;��H;�H;A�H;_�H;��H;��H;��H;F�H;��H;��H;@�H;��H;��H;A�H;��H;�H;t�H;��H;�H;b�H;��H;��H;%�H;T�H;m�H;v�H;��H;��H;l�H;u�H;V�H;>�H;F�H;B�H;      C�H;5�H;:�H;9�H;2�H;)�H;$�H;�H;��H;��H;��H;n�H;/�H;��H;��H;5�H;��H;��H;P�H;��H;m�H;�H;��H;Y�H;
�H;��H;b�H; �H;��H;��H;w�H;A�H;��H;��H;��H;��H;��H;��H;��H;��H;��H;A�H;w�H;��H;��H; �H;b�H;��H;
�H;Y�H;��H;�H;m�H;��H;P�H;��H;��H;5�H;��H;��H;/�H;n�H;��H;��H;��H;�H;$�H;)�H;2�H;9�H;:�H;5�H;      ��H;��H;��H;��H;��H;h�H;c�H;0�H;�H;��H;��H;Y�H;�H;��H;��H;O�H;��H;]�H;��H;��H;[�H;�H;��H;(�H;��H;��H;C�H;��H;��H;��H;?�H;�H;��H;��H;��H;��H;��H;��H;��H;��H;��H;�H;?�H;��H;��H;��H;C�H;��H;��H;(�H;��H;�H;[�H;��H;��H;]�H;��H;O�H;��H;��H;�H;Y�H;��H;��H;�H;0�H;c�H;h�H;��H;��H;��H;��H;      ��H;��H;��H;��H;��H;��H;s�H;C�H;�H;��H;��H;T�H;�H;��H;g�H;	�H;��H;O�H;��H;��H;)�H;��H;|�H;"�H;��H;o�H;(�H;��H;��H;c�H;�H;��H;��H;��H;��H;��H;��H;��H;��H;��H;��H;��H;�H;c�H;��H;��H;(�H;o�H;��H;"�H;|�H;��H;)�H;��H;��H;O�H;��H;	�H;g�H;��H;�H;T�H;��H;��H;�H;C�H;s�H;��H;��H;��H;��H;��H;      ��H;��H;��H;��H;��H;|�H;W�H;<�H;�H;��H;��H;a�H;�H;��H;K�H;��H;��H;K�H;��H;��H;�H;��H;e�H;�H;��H;\�H;�H;��H;��H;K�H;'�H;��H;��H;��H;��H;��H;��H;��H;��H;��H;��H;��H;'�H;K�H;��H;��H;�H;\�H;��H;�H;e�H;��H;�H;��H;��H;K�H;��H;��H;K�H;��H;�H;a�H;��H;��H;�H;<�H;W�H;|�H;��H;��H;��H;��H;      +�H;$�H;�H;��H;��H;��H;��H;Y�H;$�H;��H;z�H;7�H;��H;��H;m�H;�H;��H;'�H;��H;u�H;�H;��H;L�H;��H;��H;n�H;�H;��H;�H;A�H;(�H;��H;��H;��H;��H;��H;~�H;��H;��H;��H;��H;��H;(�H;A�H;�H;��H;�H;n�H;��H;��H;L�H;��H;�H;u�H;��H;'�H;��H;�H;m�H;��H;��H;7�H;z�H;��H;$�H;Y�H;��H;��H;��H;��H;�H;$�H;      ��H;��H;��H;��H;��H;|�H;W�H;<�H;�H;��H;��H;a�H;�H;��H;K�H;��H;��H;K�H;��H;��H;�H;��H;e�H;�H;��H;\�H;�H;��H;��H;K�H;'�H;��H;��H;��H;��H;��H;��H;��H;��H;��H;��H;��H;'�H;K�H;��H;��H;�H;\�H;��H;�H;e�H;��H;�H;��H;��H;K�H;��H;��H;K�H;��H;�H;a�H;��H;��H;�H;<�H;W�H;|�H;��H;��H;��H;��H;      ��H;��H;��H;��H;��H;��H;s�H;C�H;�H;��H;��H;T�H;�H;��H;g�H;	�H;��H;O�H;��H;��H;)�H;��H;|�H;"�H;��H;o�H;(�H;��H;��H;c�H;�H;��H;��H;��H;��H;��H;��H;��H;��H;��H;��H;��H;�H;c�H;��H;��H;(�H;o�H;��H;"�H;|�H;��H;)�H;��H;��H;O�H;��H;	�H;g�H;��H;�H;T�H;��H;��H;�H;C�H;s�H;��H;��H;��H;��H;��H;      ��H;��H;��H;��H;��H;h�H;c�H;0�H;�H;��H;��H;Y�H;�H;��H;��H;O�H;��H;]�H;��H;��H;[�H;�H;��H;(�H;��H;��H;C�H;��H;��H;��H;?�H;�H;��H;��H;��H;��H;��H;��H;��H;��H;��H;�H;?�H;��H;��H;��H;C�H;��H;��H;(�H;��H;�H;[�H;��H;��H;]�H;��H;O�H;��H;��H;�H;Y�H;��H;��H;�H;0�H;c�H;h�H;��H;��H;��H;��H;      C�H;5�H;:�H;9�H;2�H;)�H;$�H;�H;��H;��H;��H;n�H;/�H;��H;��H;5�H;��H;��H;P�H;��H;m�H;�H;��H;Y�H;
�H;��H;b�H; �H;��H;��H;w�H;A�H;��H;��H;��H;��H;��H;��H;��H;��H;��H;A�H;w�H;��H;��H; �H;b�H;��H;
�H;Y�H;��H;�H;m�H;��H;P�H;��H;��H;5�H;��H;��H;/�H;n�H;��H;��H;��H;�H;$�H;)�H;2�H;9�H;:�H;5�H;      >�H;B�H;F�H;>�H;V�H;u�H;l�H;��H;��H;v�H;m�H;T�H;%�H;��H;��H;b�H;�H;��H;t�H;�H;��H;A�H;��H;��H;@�H;��H;��H;F�H;��H;��H;��H;_�H;A�H;�H;��H;��H;��H;��H;��H;�H;A�H;_�H;��H;��H;��H;F�H;��H;��H;@�H;��H;��H;A�H;��H;�H;t�H;��H;�H;b�H;��H;��H;%�H;T�H;m�H;v�H;��H;��H;l�H;u�H;V�H;>�H;F�H;B�H;      L�H;p�H;��H;��H;��H;'�H;I�H;w�H;��H;��H;��H;��H;��H;��H;��H;��H;7�H;��H;��H;5�H;��H;��H;�H;��H;r�H;�H;��H;u�H;7�H;��H;��H;��H;w�H;?�H;�H;'�H;(�H;'�H;�H;?�H;w�H;��H;��H;��H;7�H;u�H;��H;�H;r�H;��H;�H;��H;��H;5�H;��H;��H;7�H;��H;��H;��H;��H;��H;��H;��H;��H;w�H;I�H;'�H;��H;��H;��H;p�H;      ��H;�H;�H;w�H;��H;e�H;�H;��H;#�H;��H;��H;!�H;T�H;y�H;k�H;d�H;F�H;�H;��H;z�H;�H;��H;��H;	�H;��H;`�H;�H;��H;k�H;-�H;��H;��H;��H;��H;c�H;K�H;A�H;K�H;c�H;��H;��H;��H;��H;-�H;k�H;��H;�H;`�H;��H;	�H;��H;��H;�H;z�H;��H;�H;F�H;d�H;k�H;y�H;T�H;!�H;��H;��H;#�H;��H;�H;e�H;��H;w�H;�H;�H;      ��H;U�H;7�H;��H;��H;i�H;��H;��H;��H;��H;��H;��H;A�H;��H;��H;!�H;9�H;�H;��H;��H;[�H;��H;��H;e�H; �H;��H;H�H;�H;��H;k�H;7�H;��H;��H;��H;��H;��H;�H;��H;��H;��H;��H;��H;7�H;k�H;��H;�H;H�H;��H; �H;e�H;��H;��H;[�H;��H;��H;�H;9�H;!�H;��H;��H;A�H;��H;��H;��H;��H;��H;��H;i�H;��H;��H;7�H;U�H;      ��H;5�H;��H;Z�H;Q�H;��H;L�H;��H;(�H;1�H;&�H;��H;�H;#�H;��H;W�H;��H;��H;��H;��H;��H;a�H;��H;��H;i�H;��H;��H;W�H;�H;��H;u�H;F�H; �H;��H;��H;��H;��H;��H;��H;��H; �H;F�H;u�H;��H;�H;W�H;��H;��H;i�H;��H;��H;a�H;��H;��H;��H;��H;��H;W�H;��H;#�H;�H;��H;&�H;1�H;(�H;��H;L�H;��H;Q�H;Z�H;��H;5�H;      �H;H;� H;�7H;�SH;KrH;9�H;ԪH;��H;��H;|�H;��H;�H;�H;��H;��H;��H;=�H;��H;��H;��H;��H;5�H;��H;��H;_�H;��H;��H;H�H;�H;��H;��H;b�H;C�H;(�H;�H;�H;�H;(�H;C�H;b�H;��H;��H;�H;H�H;��H;��H;_�H;��H;��H;5�H;��H;��H;��H;��H;=�H;��H;��H;��H;�H;�H;��H;|�H;��H;��H;ԪH;9�H;KrH;�SH;�7H;� H;H;      mCF;{QF;�yF;�F;�G;�[G;�G;YH;#HH;��H;��H;��H;
�H;��H;��H;8�H;��H;7�H;��H;P�H;��H;�H;r�H;D�H;��H;��H;_�H;��H;��H;`�H;�H;��H;��H;��H;o�H;\�H;n�H;\�H;o�H;��H;��H;��H;�H;`�H;��H;��H;_�H;��H;��H;D�H;r�H;�H;��H;P�H;��H;7�H;��H;8�H;��H;��H;
�H;��H;��H;��H;#HH;YH;�G;�[G;�G;�F;�yF;{QF;      ��A;B;1oB;�C;��C;{�D;otE;�CF;N�F;��G;�H;eH;�H;��H;[�H;�H;��H;�H;��H;��H;"�H;e�H;��H;i�H;-�H;��H;��H;i�H; �H;��H;r�H;@�H;
�H;��H;��H;��H;��H;��H;��H;��H;
�H;@�H;r�H;��H; �H;i�H;��H;��H;-�H;i�H;��H;e�H;"�H;��H;��H;�H;��H;�H;[�H;��H;�H;eH;�H;��G;N�F;�CF;otE;{�D;��C;�C;1oB;B;      ~n8;M�8;׎9;��:;��<;
c>;ZQ@;�.B;��C;�OE;�yF;j[G;��G;DhH;8�H;��H;8�H;a�H;-�H;5�H;\�H;��H;a�H;k�H;i�H;D�H;��H;��H;e�H;	�H;��H;��H;Y�H;(�H;"�H;�H;��H;�H;"�H;(�H;Y�H;��H;��H;	�H;e�H;��H;��H;D�H;i�H;k�H;a�H;��H;\�H;5�H;-�H;a�H;8�H;��H;8�H;DhH;��G;j[G;�yF;�OE;��C;�.B;ZQ@;
c>;��<;��:;׎9;M�8;      �R%;i�%;^�';M*;4�-;ʕ1;�5;5�9;�,=;IQ@;�B;��D;9lF;�tG;� H;�H;��H;��H;�H;��H;��H;0�H;�H;a�H;��H;r�H;5�H;��H;��H;��H;�H;��H;��H;��H;|�H;e�H;L�H;e�H;|�H;��H;��H;��H;�H;��H;��H;��H;5�H;r�H;��H;a�H;�H;0�H;��H;��H;�H;��H;��H;�H;� H;�tG;9lF;��D;�B;IQ@;�,=;5�9;�5;ʕ1;4�-;M*;^�';i�%;      �V;�w;0�;Q�
;�;�;)� ;��(;��/;$H6;��;;�?; C;�OE;�F;�G;�dH;N�H;��H;&�H;O�H;��H;0�H;��H;e�H;�H;��H;a�H;��H;��H;��H;A�H;�H;�H;��H;��H;��H;��H;��H;�H;�H;A�H;��H;��H;��H;a�H;��H;�H;e�H;��H;0�H;��H;O�H;&�H;��H;N�H;�dH;�G;�F;�OE; C;�?;��;;$H6;��/;��(;)� ;�;�;Q�
;0�;�w;      �:mĆ:nȒ:���:q�:n��:���:��	;v;7�#;��-;#�5;�K<;��@;�'D;3CF;��G;�GH;s�H;�H;��H;O�H;��H;\�H;"�H;��H;��H;��H;[�H;�H;��H;��H;m�H;[�H;)�H;�H;�H;�H;)�H;[�H;m�H;��H;��H;�H;[�H;��H;��H;��H;"�H;\�H;��H;O�H;��H;�H;s�H;�GH;��G;3CF;�'D;��@;�K<;#�5;��-;7�#;v;��	;���:n��:q�:���:nȒ:mĆ:      0.�7��0�깤�K�
9�Z:��k: L�:5��:�x;��;�$;�/;��8;��>;#C;7�E;�[G;\7H;̤H;�H;&�H;��H;5�H;��H;P�H;��H;��H;��H;z�H;5�H;�H;��H;��H;��H;��H;u�H;��H;��H;��H;��H;�H;5�H;z�H;��H;��H;��H;P�H;��H;5�H;��H;&�H;�H;̤H;\7H;�[G;7�E;#C;��>;��8;�/;�$;��;�x;5��: L�:��k:�Z:
9��K�0��7��      �Q^��X�VF�]�)��+�-ж���<�CjS�k:���:I��:�;|�;M*;	�5;�b=;�oB;��E;�IG;\7H;s�H;��H;�H;-�H;��H;��H;��H;��H;��H;��H;��H;t�H;P�H;��H;��H;��H;��H;��H;��H;��H;P�H;t�H;��H;��H;��H;��H;��H;��H;��H;-�H;�H;��H;s�H;\7H;�IG;��E;�oB;�b=;	�5;M*;|�;�;I��:���:k:CjS���<�-ж��+�]�)�VF��X�      ����o���X��P�ѻf���[ǐ��X��6��
���K�<<":fL�:�`�:�h;Z�%;��3;�<;Y/B;��E;�[G;�GH;N�H;��H;a�H;�H;7�H;=�H;��H;�H;�H;��H;��H;��H;]�H;O�H;K�H;'�H;K�H;O�H;]�H;��H;��H;��H;�H;�H;��H;=�H;7�H;�H;a�H;��H;N�H;�GH;�[G;��E;Y/B;�<;��3;Z�%;�h;�`�:fL�:<<":�K��
���6��X�[ǐ�f���P�ѻX��o���      ��n��mj���]���J�n�1�L4�l��S���V
x�hX���y�&
9���:֣�:@�;u�#;v�2;�<;�oB;7�E;��G;�dH;��H;8�H;��H;��H;��H;��H;9�H;F�H;7�H;�H;��H;��H;��H;��H;��H;��H;��H;��H;��H;�H;7�H;F�H;9�H;��H;��H;��H;��H;8�H;��H;�dH;��G;7�E;�oB;�<;v�2;u�#;@�;֣�:���:&
9��y�hX�V
x�S���l��L4�n�1���J���]��mj�      B<ͼ��ɼ�����֯�Ҷ��ㄼ��Y�-�*�J���t���X��sѺ�(�K<Q:\��:��
;u�#;��3;�b=;#C;3CF;�G;�H;��H;�H;8�H;��H;W�H;!�H;d�H;��H;b�H;5�H;O�H;	�H;��H;�H;��H;	�H;O�H;5�H;b�H;��H;d�H;!�H;W�H;��H;8�H;�H;��H;�H;�G;3CF;#C;�b=;��3;u�#;��
;\��:K<Q:�(��sѺ�X�t��J���-�*���Y�ㄼҶ���֯�������ɼ      ��'�#�$����y��  ���ۼ����+����]��X!�>ۻ�+��+�h���>:\��:@�;Z�%;	�5;��>;�'D;�F;� H;8�H;[�H;��H;��H;��H;��H;k�H;��H;��H;��H;��H;g�H;K�H;m�H;K�H;g�H;��H;��H;��H;��H;k�H;��H;��H;��H;��H;[�H;8�H;� H;�F;�'D;��>;	�5;Z�%;@�;\��:�>:h��+��+��>ۻ�X!���]��+�������ۼ�  �y����#�$�      �����v����w�]�c��J�Ȅ-�x��;缈沼ㄼ��;�����k��66�h��K<Q:֣�:�h;M*;��8;��@;�OE;�tG;DhH;��H;��H;�H;#�H;��H;y�H;��H;��H;��H;��H;��H;��H;��H;��H;��H;��H;��H;��H;��H;y�H;��H;#�H;�H;��H;��H;DhH;�tG;�OE;��@;��8;M*;�h;֣�:K<Q:h��66�k��������;�ㄼ�沼�;�x�Ȅ-��J�]�c���w��v��      nHͽ̪ɽ�;��"����������[�z0�p��'<ͼо��v�J���k��+��(����:�`�:|�;�/;�K<; C;9lF;��G;�H;
�H;�H;�H;A�H;T�H;��H;%�H;/�H;�H;�H;�H;��H;�H;�H;�H;/�H;%�H;��H;T�H;A�H;�H;�H;
�H;�H;��G;9lF; C;�K<;�/;|�;�`�:���:�(�+�k����v�J�о��'<ͼp��z0���[�������"���;��̪ɽ      ��-�}��|�ű�ƽUP���v���J�D����ۼ��v�J������+���sѺ&
9fL�:�;�$;#�5;�?;��D;j[G;eH;��H;��H;��H;��H;!�H;��H;T�H;n�H;Y�H;T�H;a�H;7�H;a�H;T�H;Y�H;n�H;T�H;��H;!�H;��H;��H;��H;��H;eH;j[G;��D;�?;#�5;�$;�;fL�:&
9�sѺ�+������v�J�����ۼD���J��v��UP��ƽű�|�}��-�       j�Ide�M0X�sD�\{+�z�����k㻽R���JDX������ۼо����;�>ۻ�X���y�<<":I��:��;��-;��;;�B;�yF;�H;��H;|�H;&�H;��H;��H;��H;m�H;��H;��H;��H;��H;z�H;��H;��H;��H;��H;m�H;��H;��H;��H;&�H;|�H;��H;�H;�yF;�B;��;;��-;��;I��:<<":��y��X�>ۻ��;�о����ۼ���JDX�R���k㻽���z��\{+�sD�M0X�Ide�      ��Fh��b���I���|x���O��C(�y�Īɽ����JDX�D��'<ͼㄼ�X!�t��hX��K����:�x;7�#;$H6;IQ@;�OE;��G;��H;��H;1�H;��H;��H;��H;v�H;��H;��H;��H;��H;��H;��H;��H;��H;��H;v�H;��H;��H;��H;1�H;��H;��H;��G;�OE;IQ@;$H6;7�#;�x;���:�K�hX�t���X!�ㄼ'<ͼD��JDX�����Īɽy��C(���O��|x��I��b��Fh��      /�����������;^ɰ��G����i�.�5��	�ĪɽR����J�p���沼��]�J���V
x��
��k:5��:v;��/;�,=;��C;N�F;#HH;��H;(�H;��H;#�H;��H;��H;��H;�H;�H;�H;$�H;�H;�H;�H;��H;��H;��H;#�H;��H;(�H;��H;#HH;N�F;��C;�,=;��/;v;5��:k:�
��V
x�J�����]��沼p���J�R���Īɽ�	�.�5���i��G��^ɰ��;��徨���      �2�L�-��"�$E�����4Kɾa��w�s�.�5�y�k㻽�v��z0��;��+��-�*�S����6�CjS� L�:��	;��(;5�9;�.B;�CF;YH;ԪH;��H;��H;��H;w�H;��H;�H;0�H;C�H;<�H;Y�H;<�H;C�H;0�H;�H;��H;w�H;��H;��H;��H;ԪH;YH;�CF;�.B;5�9;��(;��	; L�:CjS��6�S���-�*��+���;�z0��v��k㻽y�.�5�w�s�a��4Kɾ����$E��"�L�-�      3s�cm�/�\�]�C�,�%����TҾa����i��C(����UP����[�x������Y�l���X���<���k:���:)� ;�5;ZQ@;otE;�G;9�H;L�H;��H;�H;I�H;l�H;$�H;c�H;s�H;W�H;��H;W�H;s�H;c�H;$�H;l�H;I�H;�H;��H;L�H;9�H;�G;otE;ZQ@;�5;)� ;���:��k:��<��X�l����Y����x���[�UP����콡C(���i�a���TҾ��,�%�]�C�/�\�cm�      �ޞ�������RF�3�W�M�-���4Kɾ�G����O�z��ƽ����Ȅ-���ۼㄼL4�[ǐ�-ж��Z:n��:�;ʕ1;
c>;{�D;�[G;KrH;��H;i�H;e�H;'�H;u�H;)�H;h�H;��H;|�H;��H;|�H;��H;h�H;)�H;u�H;'�H;e�H;i�H;��H;KrH;�[G;{�D;
c>;ʕ1;�;n��:�Z:-ж�[ǐ�L4�ㄼ��ۼȄ-�����ƽz����O��G��4Kɾ��M�-�3�W�RF�������      ��ſ~��Bw���ޞ�|���3�W�,�%�����^ɰ��|x�\{+�ű����J��  �Ҷ��n�1�f����+�
9q�:�;4�-;��<;��C;�G;�SH;Q�H;��H;��H;��H;V�H;2�H;��H;��H;��H;��H;��H;��H;��H;2�H;V�H;��H;��H;��H;Q�H;�SH;�G;��C;��<;4�-;�;q�:
9�+�f���n�1�Ҷ���  ��J���ű�\{+��|x�^ɰ�����,�%�3�W�|����ޞ�Bw��~��      ������Կp���ޞ�RF�]�C�$E��;�I��sD�|�"��]�c�y��֯���J�P�ѻ]�)���K����:Q�
;M*;��:;�C;�F;�7H;Z�H;��H;w�H;��H;>�H;9�H;��H;��H;��H;��H;��H;��H;��H;9�H;>�H;��H;w�H;��H;Z�H;�7H;�F;�C;��:;M*;Q�
;���:��K�]�)�P�ѻ��J��֯�y�]�c�"��|�sD��I���;$E�]�C�RF��ޞ�p���Կ��      ������{���ԿBw�����/�\��"����b��M0X�}���;����w����������]�X��VF�0��nȒ:0�;^�';׎9;1oB;�yF;� H;��H;7�H;�H;��H;F�H;:�H;��H;��H;��H;�H;��H;��H;��H;:�H;F�H;��H;�H;7�H;��H;� H;�yF;1oB;׎9;^�';0�;nȒ:0��VF�X�黼�]����������w��;��}��M0X�b������"�/�\����Bw���Կ{�𿖏�      $��������~�����cm�L�-�����Fh��Ide�-�̪ɽ�v��#�$���ɼ�mj�o����X�7��mĆ:�w;i�%;M�8;B;{QF;H;5�H;U�H;�H;p�H;B�H;5�H;��H;��H;��H;$�H;��H;��H;��H;5�H;B�H;p�H;�H;U�H;5�H;H;{QF;B;M�8;i�%;�w;mĆ:7���X�o����mj���ɼ#�$��v��̪ɽ-�Ide�Fh������L�-�cm����~���忖����      �>���8���*�O������˿�o��<�b�=\�+m־^��K�:��J�&��F�B�F���������/��������>:�r�:do ;�I6;DA;�HF;�MH;�H;!I;�I;I;�I;mI;I;q�H;��H;*�H;��H;q�H;I;mI;�I;I;�I;!I;�H;�MH;�HF;DA;�I6;do ;�r�:��>:�����/���������F��F�B�&���J�K�:�^��+m־=\�<�b��o���˿����O���*���8�      ��8��4��g&�0��2����<ƿ벗��>]����G�Ѿ�p���*7����"W��MR?�	}鼀8����s������8�G:���: !;&�6;(kA;�XF;�SH;s�H;!I;�I;�I;�I;FI;�I;e�H;��H;�H;��H;e�H;�I;FI;�I;�I;�I;!I;s�H;�SH;�XF;(kA;&�6; !;���:8�G:���s������8��	}�MR?�"W�����*7��p��G�Ѿ����>]�벗��<ƿ2���0���g&��4�      ��*��g&��#�o�K[�jL�������M�l5��>ľ
����,��D�撐��5�;�ݼ���q
���x��wk�~�b:�j�:#;ږ7;��A;�F;�cH;�I;\!I;I;oI;AI;�I;�I; �H;x�H;��H;x�H; �H;�I;�I;AI;oI;I;\!I;�I;�cH;�F;��A;ږ7;#;�j�:~�b:�wk���x��q
���;�ݼ�5�撐��Dὤ�,�
���>ľl5���M����jL��K[�o��#��g&�      O�0��o����˿:1��-�y���6��z �����)�l�+��ͽ!�����&���˼_�k�q���k�X��� �г�:o�;)&;�9;��B;�F;�|H;�I;e!I;5I;�I;�
I;qI;FI;��H;"�H;��H;"�H;��H;FI;qI;�
I;�I;5I;e!I;�I;�|H;�F;��B;�9;)&;o�;г�:�� �k�X�q���_�k���˼��&�!����ͽ+�)�l������z ���6�-�y�:1���˿���o�0��      ����2���K[忭˿�T��蟉�s�R�����E۾̗����M�~�	������j��3�"d��ɆO���׻c�/��
�����:��	;%*;l;;�iC;�&G;�H;�I;
!I;�I;�I;�	I;�I;� I;I�H;��H; �H;��H;I�H;� I;�I;�	I;�I;�I;
!I;�I;�H;�&G;�iC;l;;%*;��	;���:�
��c�/���׻ɆO�"d���3���j����~�	���M�̗���E۾���s�R�蟉��T���˿K[�2���      �˿�<ƿjL��:1��蟉��>]���)��$���ճ���{���,�j��$��Q`I��J��-��4/�S,��˻ ��!69	3�:�;o.;0-=;o`D;�G;o�H;�I;? I;aI;SI;�I;�I;��H;��H;�H;d�H;�H;��H;��H;�I;�I;SI;aI;? I;�I;o�H;�G;o`D;0-=;o.;�;	3�:�!69˻ �S,��4/�-���J��Q`I�$��j�齞�,���{��ճ��$����)��>]�蟉�:1��jL���<ƿ      �o��벗����-�y�s�R���)�iv��>ľ�]����I�Tl�~��������&�߮Ҽ	�}�VB�"���������!:>)�:Vy;�3;li?;�[E;��G;��H;tI;�I;�I;�I;|I;�I;�H;��H;c�H;��H;c�H;��H;�H;�I;|I;�I;�I;�I;tI;��H;��G;�[E;li?;�3;Vy;>)�:��!:����"���VB�	�}�߮Ҽ��&����~���Tl���I��]���>ľiv���)�s�R�-�y����벗�      <�b��>]���M���6�����$���>ľq��q�Z�+�K9ݽW����L����0F��&�G�\�׻�;�u�Ǌ:�h;5O$;�7;y�A;IF;9BH;��H;�I;mI;xI;I;-I;�I;�H;��H;��H;�H;��H;��H;�H;�I;-I;I;xI;mI;�I;��H;9BH;IF;y�A;�7;5O$;�h;Ǌ:u칹;�\�׻&�G�0F�������L�W��K9ݽ+�q�Z�q���>ľ�$�������6���M��>]�      =\����l5��z ��E۾�ճ��]��q�Z�F?#����A����j�(��Oϼ��������Snۺl3�9�2�:o�;y�,;��;;C�C;�G;Q�H;�
I;� I;�I;FI;.
I;�I;> I;�H;�H;��H;!�H;��H;�H;�H;> I;�I;.
I;FI;�I;� I;�
I;Q�H;�G;C�C;��;;y�,;o�;�2�:l3�9Snۺ��������Oϼ(����j��A�����F?#�q�Z��]���ճ��E۾�z �l5����      +m־G�Ѿ�>ľ����̗����{���I�+����V���{�?�/�.���,��c=���һ�@�<� ���k:B�:#a;��3;Ai?;v1E;��G;p�H;7I;wI;�I;�I;%I;�I;��H;��H;��H;��H;V�H;��H;��H;��H;��H;�I;%I;�I;�I;wI;7I;p�H;��G;v1E;Ai?;��3;#a;B�:��k:<� ��@���һc=��,��.��?�/��{��V�����+���I���{�̗�������>ľG�Ѿ      ^���p��
��)�l���M���,�Tl�K9ݽ�A���{���5��J��;���T[�I?������Q���I�9�:��;:*;4�9;jjB;چF;�MH;��H; I;�I;�I;"I;I;@I;^�H;��H;��H;��H;j�H;��H;��H;��H;^�H;@I;I;"I;�I;�I; I;��H;�MH;چF;jjB;4�9;:*;��;�:�I�9�Q������I?��T[�;���J����5��{��A��K9ݽTl���,���M�)�l�
���p��      K�:��*7���,�+�~�	�j��~���W����j�?�/��J���I��%�k���c.������;Ǌ:�m�:';mq3;1�>;8�D;t�G;R�H;I;/ I;�I;�I;�	I;�I;`�H;��H;��H;��H;��H;^�H;��H;��H;��H;��H;`�H;�I;�	I;�I;�I;/ I;I;R�H;t�G;8�D;1�>;mq3;';�m�:;Ǌ:����c.����%�k��I���J��?�/���j�W��~���j��~�	�+���,��*7�      �J���D��ͽ���$�������L�(��.��;��%�k����I����/��"/�)�>:���:�A;v�,;��:;>�B;�wF;�;H;��H;	I;�I;�I;AI;�I;�I;��H;s�H;4�H;n�H;��H;l�H;��H;n�H;4�H;s�H;��H;�I;�I;AI;�I;�I;	I;��H;�;H;�wF;>�B;��:;v�,;�A;���:)�>:�"/���/��I����%�k�;��.��(����L����$������ͽ�Dὼ��      &��"W��撐�!�����j�Q`I���&����Oϼ�,���T[����I��;��qk�k:h3�:� ;!&;�6;� @;C1E;�G;��H;�I;�I;OI;I;�	I;:I;u�H;��H;�H;��H;^�H;��H;D�H;��H;^�H;��H;�H;��H;u�H;:I;�	I;I;OI;�I;�I;��H;�G;C1E;� @;�6;!&;� ;h3�:k:�qk�;��I�����T[��,��Oϼ�����&�Q`I���j�!���撐�"W��      F�B�MR?��5���&��3��J��߮Ҽ0F����c=�I?�c.����/��qk����9�ճ:�;J!;l3;��=;��C;*�F;cH;��H;�I;I;�I;$I;�I;�I;C�H;��H;��H;|�H;?�H;|�H;3�H;|�H;?�H;|�H;��H;��H;C�H;�I;�I;$I;�I;I;�I;��H;cH;*�F;��C;��=;l3;J!;�;�ճ:���9�qk���/�c.��I?�c=���0F��߮Ҽ�J���3���&��5�MR?�      F��	}�;�ݼ��˼"d��-��	�}�&�G������һ�������"/�k:�ճ:#�;�a;Ģ0;�<;��B;�HF;uH;,�H;�I;yI;I;8I;Y	I;�I;�H;/�H;T�H;�H;#�H;�H;r�H;5�H;r�H;�H;#�H;�H;T�H;/�H;�H;�I;Y	I;8I;I;yI;�I;,�H;uH;�HF;��B;�<;Ģ0;�a;#�;�ճ:k:�"/���������һ���&�G�	�}�-��"d����˼;�ݼ	}�      �����8����_�k�ɆO�4/�VB�\�׻����@��Q����)�>:h3�:�;�a;��/;=;;J�A;��E;ɾG;��H;�	I;gI;I;�I;�I;�I;� I;��H;;�H;��H;��H;��H;�H;c�H;)�H;c�H;�H;��H;��H;��H;;�H;��H;� I;�I;�I;�I;I;gI;�	I;��H;ɾG;��E;J�A;=;;��/;�a;�;h3�:)�>:���Q���@����\�׻VB�4/�ɆO�_�k����8��      ������q
�q�����׻S,��"����;�Snۺ<� ��I�9;Ǌ:���:� ;J!;Ģ0;=;;̒A;�oE;|�G;ӍH;��H;�I;9I;ZI; I;�I;oI;��H;=�H;x�H;�H;�H;��H;��H;[�H;1�H;[�H;��H;��H;�H;�H;x�H;=�H;��H;oI;�I; I;ZI;9I;�I;��H;ӍH;|�G;�oE;̒A;=;;Ģ0;J!;� ;���:;Ǌ:�I�9<� �Snۺ�;�"���S,����׻q����q
���      �/��s�����x�k�X�c�/�˻ �����u�l3�9��k:�:�m�:�A;!&;l3;�<;J�A;�oE;hsG;�{H;.�H;,I;rI;CI;�I;i	I;�I;L�H;I�H;�H;��H;x�H;��H;��H;��H;l�H;\�H;l�H;��H;��H;��H;x�H;��H;�H;I�H;L�H;�I;i	I;�I;CI;rI;,I;.�H;�{H;hsG;�oE;J�A;�<;l3;!&;�A;�m�:�:��k:l3�9u칋���˻ �c�/�k�X���x�s���      ��������wk��� ��
���!69��!:Ǌ:�2�:B�:��;';v�,;�6;��=;��B;��E;|�G;�{H;��H;zI;I;�I;WI;�
I;"I;� I;A�H;��H;4�H;��H;�H;��H;��H;��H;}�H;k�H;}�H;��H;��H;��H;�H;��H;4�H;��H;A�H;� I;"I;�
I;WI;�I;I;zI;��H;�{H;|�G;��E;��B;��=;�6;v�,;';��;B�:�2�:Ǌ:��!:�!69�
���� ��wk����      ��>:8�G:~�b:г�:���:	3�:>)�:�h;o�;#a;:*;mq3;��:;� @;��C;�HF;ɾG;ӍH;.�H;zI;I;BI;9I;�I;I;VI;�H;��H;��H;o�H;B�H;��H;��H;��H;	�H;��H;y�H;��H;	�H;��H;��H;��H;B�H;o�H;��H;��H;�H;VI;I;�I;9I;BI;I;zI;.�H;ӍH;ɾG;�HF;��C;� @;��:;mq3;:*;#a;o�;�h;>)�:	3�:���:г�:~�b:8�G:      �r�:���:�j�:o�;��	;�;Vy;5O$;y�,;��3;4�9;1�>;>�B;C1E;*�F;uH;��H;��H;,I;I;BI;�I;6I;�I;�I;��H;�H;F�H;��H;��H;��H;��H;��H;��H;)�H;��H;��H;��H;)�H;��H;��H;��H;��H;��H;��H;F�H;�H;��H;�I;�I;6I;�I;BI;I;,I;��H;��H;uH;*�F;C1E;>�B;1�>;4�9;��3;y�,;5O$;Vy;�;��	;o�;�j�:���:      do ; !;#;)&;%*;o.;�3;�7;��;;Ai?;jjB;8�D;�wF;�G;cH;,�H;�	I;�I;rI;�I;9I;6I;�I;RI;4�H;��H;��H; �H;��H;�H;��H;x�H;��H;��H;E�H;�H;��H;�H;E�H;��H;��H;x�H;��H;�H;��H; �H;��H;��H;4�H;RI;�I;6I;9I;�I;rI;�I;�	I;,�H;cH;�G;�wF;8�D;jjB;Ai?;��;;�7;�3;o.;%*;)&;#; !;      �I6;&�6;ږ7;�9;l;;0-=;li?;y�A;C�C;v1E;چF;t�G;�;H;��H;��H;�I;gI;9I;CI;WI;�I;�I;RI;E�H;��H;��H;Y�H;$�H;0�H;��H;~�H;e�H;��H;�H;��H;]�H;:�H;]�H;��H;�H;��H;e�H;~�H;��H;0�H;$�H;Y�H;��H;��H;E�H;RI;�I;�I;WI;CI;9I;gI;�I;��H;��H;�;H;t�G;چF;v1E;C�C;y�A;li?;0-=;l;;�9;ږ7;&�6;      DA;(kA;��A;��B;�iC;o`D;�[E;IF;�G;��G;�MH;R�H;��H;�I;�I;yI;I;ZI;�I;�
I;I;�I;4�H;��H;��H;w�H;-�H;@�H;��H;��H;`�H;u�H;��H;O�H;��H;��H;��H;��H;��H;O�H;��H;u�H;`�H;��H;��H;@�H;-�H;w�H;��H;��H;4�H;�I;I;�
I;�I;ZI;I;yI;�I;�I;��H;R�H;�MH;��G;�G;IF;�[E;o`D;�iC;��B;��A;(kA;      �HF;�XF;�F;�F;�&G;�G;��G;9BH;Q�H;p�H;��H;I;	I;�I;I;I;�I; I;i	I;"I;VI;��H;��H;��H;w�H;S�H;Z�H;��H;��H;i�H;X�H;��H;&�H;��H;@�H;"�H;�H;"�H;@�H;��H;&�H;��H;X�H;i�H;��H;��H;Z�H;S�H;w�H;��H;��H;��H;VI;"I;i	I; I;�I;I;I;�I;	I;I;��H;p�H;Q�H;9BH;��G;�G;�&G;�F;�F;�XF;      �MH;�SH;�cH;�|H;�H;o�H;��H;��H;�
I;7I; I;/ I;�I;OI;�I;8I;�I;�I;�I;� I;�H;�H;��H;Y�H;-�H;Z�H;��H;��H;X�H;Z�H;��H;��H;d�H;��H;��H;��H;��H;��H;��H;��H;d�H;��H;��H;Z�H;X�H;��H;��H;Z�H;-�H;Y�H;��H;�H;�H;� I;�I;�I;�I;8I;�I;OI;�I;/ I; I;7I;�
I;��H;��H;o�H;�H;�|H;�cH;�SH;      �H;s�H;�I;�I;�I;�I;tI;�I;� I;wI;�I;�I;�I;I;$I;Y	I;�I;oI;L�H;A�H;��H;F�H; �H;$�H;@�H;��H;��H;k�H;O�H;��H;��H;;�H;��H;|�H;9�H;
�H;�H;
�H;9�H;|�H;��H;;�H;��H;��H;O�H;k�H;��H;��H;@�H;$�H; �H;F�H;��H;A�H;L�H;oI;�I;Y	I;$I;I;�I;�I;�I;wI;� I;�I;tI;�I;�I;�I;�I;s�H;      !I;!I;\!I;e!I;
!I;? I;�I;mI;�I;�I;�I;�I;AI;�	I;�I;�I;� I;��H;I�H;��H;��H;��H;��H;0�H;��H;��H;X�H;O�H;��H;��H;/�H;��H;M�H;��H;��H;��H;��H;��H;��H;��H;M�H;��H;/�H;��H;��H;O�H;X�H;��H;��H;0�H;��H;��H;��H;��H;I�H;��H;� I;�I;�I;�	I;AI;�I;�I;�I;�I;mI;�I;? I;
!I;e!I;\!I;!I;      �I;�I;I;5I;�I;aI;�I;xI;FI;�I;"I;�	I;�I;:I;�I;�H;��H;=�H;�H;4�H;o�H;��H;�H;��H;��H;i�H;Z�H;��H;��H;�H;��H;C�H;��H;��H;g�H;J�H;9�H;J�H;g�H;��H;��H;C�H;��H;�H;��H;��H;Z�H;i�H;��H;��H;�H;��H;o�H;4�H;�H;=�H;��H;�H;�I;:I;�I;�	I;"I;�I;FI;xI;�I;aI;�I;5I;I;�I;      I;�I;oI;�I;�I;SI;�I;I;.
I;%I;I;�I;�I;u�H;C�H;/�H;;�H;x�H;��H;��H;B�H;��H;��H;~�H;`�H;X�H;��H;��H;/�H;��H;'�H;��H;v�H;<�H;	�H;��H;��H;��H;	�H;<�H;v�H;��H;'�H;��H;/�H;��H;��H;X�H;`�H;~�H;��H;��H;B�H;��H;��H;x�H;;�H;/�H;C�H;u�H;�I;�I;I;%I;.
I;I;�I;SI;�I;�I;oI;�I;      �I;�I;AI;�
I;�	I;�I;|I;-I;�I;�I;@I;`�H;��H;��H;��H;T�H;��H;�H;x�H;�H;��H;��H;x�H;e�H;u�H;��H;��H;;�H;��H;C�H;��H;R�H;!�H;��H;��H;��H;��H;��H;��H;��H;!�H;R�H;��H;C�H;��H;;�H;��H;��H;u�H;e�H;x�H;��H;��H;�H;x�H;�H;��H;T�H;��H;��H;��H;`�H;@I;�I;�I;-I;|I;�I;�	I;�
I;AI;�I;      mI;FI;�I;qI;�I;�I;�I;�I;> I;��H;^�H;��H;s�H;�H;��H;�H;��H;�H;��H;��H;��H;��H;��H;��H;��H;&�H;d�H;��H;M�H;��H;v�H;!�H;��H;��H;��H;m�H;f�H;m�H;��H;��H;��H;!�H;v�H;��H;M�H;��H;d�H;&�H;��H;��H;��H;��H;��H;��H;��H;�H;��H;�H;��H;�H;s�H;��H;^�H;��H;> I;�I;�I;�I;�I;qI;�I;FI;      I;�I;�I;FI;� I;��H;�H;�H;�H;��H;��H;��H;4�H;��H;|�H;#�H;��H;��H;��H;��H;��H;��H;��H;�H;O�H;��H;��H;|�H;��H;��H;<�H;��H;��H;n�H;V�H;J�H;9�H;J�H;V�H;n�H;��H;��H;<�H;��H;��H;|�H;��H;��H;O�H;�H;��H;��H;��H;��H;��H;��H;��H;#�H;|�H;��H;4�H;��H;��H;��H;�H;�H;�H;��H;� I;FI;�I;�I;      q�H;e�H; �H;��H;I�H;��H;��H;��H;�H;��H;��H;��H;n�H;^�H;?�H;�H;�H;��H;��H;��H;	�H;)�H;E�H;��H;��H;@�H;��H;9�H;��H;g�H;	�H;��H;��H;V�H;1�H;&�H;(�H;&�H;1�H;V�H;��H;��H;	�H;g�H;��H;9�H;��H;@�H;��H;��H;E�H;)�H;	�H;��H;��H;��H;�H;�H;?�H;^�H;n�H;��H;��H;��H;�H;��H;��H;��H;I�H;��H; �H;e�H;      ��H;��H;x�H;"�H;��H;�H;c�H;��H;��H;��H;��H;��H;��H;��H;|�H;r�H;c�H;[�H;l�H;}�H;��H;��H;�H;]�H;��H;"�H;��H;
�H;��H;J�H;��H;��H;m�H;J�H;&�H;
�H;�H;
�H;&�H;J�H;m�H;��H;��H;J�H;��H;
�H;��H;"�H;��H;]�H;�H;��H;��H;}�H;l�H;[�H;c�H;r�H;|�H;��H;��H;��H;��H;��H;��H;��H;c�H;�H;��H;"�H;x�H;��H;      *�H;�H;��H;��H; �H;d�H;��H;�H;!�H;V�H;j�H;^�H;l�H;D�H;3�H;5�H;)�H;1�H;\�H;k�H;y�H;��H;��H;:�H;��H;�H;��H;�H;��H;9�H;��H;��H;f�H;9�H;(�H;�H;	�H;�H;(�H;9�H;f�H;��H;��H;9�H;��H;�H;��H;�H;��H;:�H;��H;��H;y�H;k�H;\�H;1�H;)�H;5�H;3�H;D�H;l�H;^�H;j�H;V�H;!�H;�H;��H;d�H; �H;��H;��H;�H;      ��H;��H;x�H;"�H;��H;�H;c�H;��H;��H;��H;��H;��H;��H;��H;|�H;r�H;c�H;[�H;l�H;}�H;��H;��H;�H;]�H;��H;"�H;��H;
�H;��H;J�H;��H;��H;m�H;J�H;&�H;
�H;�H;
�H;&�H;J�H;m�H;��H;��H;J�H;��H;
�H;��H;"�H;��H;]�H;�H;��H;��H;}�H;l�H;[�H;c�H;r�H;|�H;��H;��H;��H;��H;��H;��H;��H;c�H;�H;��H;"�H;x�H;��H;      q�H;e�H; �H;��H;I�H;��H;��H;��H;�H;��H;��H;��H;n�H;^�H;?�H;�H;�H;��H;��H;��H;	�H;)�H;E�H;��H;��H;@�H;��H;9�H;��H;g�H;	�H;��H;��H;V�H;1�H;&�H;(�H;&�H;1�H;V�H;��H;��H;	�H;g�H;��H;9�H;��H;@�H;��H;��H;E�H;)�H;	�H;��H;��H;��H;�H;�H;?�H;^�H;n�H;��H;��H;��H;�H;��H;��H;��H;I�H;��H; �H;e�H;      I;�I;�I;FI;� I;��H;�H;�H;�H;��H;��H;��H;4�H;��H;|�H;#�H;��H;��H;��H;��H;��H;��H;��H;�H;O�H;��H;��H;|�H;��H;��H;<�H;��H;��H;n�H;V�H;J�H;9�H;J�H;V�H;n�H;��H;��H;<�H;��H;��H;|�H;��H;��H;O�H;�H;��H;��H;��H;��H;��H;��H;��H;#�H;|�H;��H;4�H;��H;��H;��H;�H;�H;�H;��H;� I;FI;�I;�I;      mI;FI;�I;qI;�I;�I;�I;�I;> I;��H;^�H;��H;s�H;�H;��H;�H;��H;�H;��H;��H;��H;��H;��H;��H;��H;&�H;d�H;��H;M�H;��H;v�H;!�H;��H;��H;��H;m�H;f�H;m�H;��H;��H;��H;!�H;v�H;��H;M�H;��H;d�H;&�H;��H;��H;��H;��H;��H;��H;��H;�H;��H;�H;��H;�H;s�H;��H;^�H;��H;> I;�I;�I;�I;�I;qI;�I;FI;      �I;�I;AI;�
I;�	I;�I;|I;-I;�I;�I;@I;`�H;��H;��H;��H;T�H;��H;�H;x�H;�H;��H;��H;x�H;e�H;u�H;��H;��H;;�H;��H;C�H;��H;R�H;!�H;��H;��H;��H;��H;��H;��H;��H;!�H;R�H;��H;C�H;��H;;�H;��H;��H;u�H;e�H;x�H;��H;��H;�H;x�H;�H;��H;T�H;��H;��H;��H;`�H;@I;�I;�I;-I;|I;�I;�	I;�
I;AI;�I;      I;�I;oI;�I;�I;SI;�I;I;.
I;%I;I;�I;�I;u�H;C�H;/�H;;�H;x�H;��H;��H;B�H;��H;��H;~�H;`�H;X�H;��H;��H;/�H;��H;'�H;��H;v�H;<�H;	�H;��H;��H;��H;	�H;<�H;v�H;��H;'�H;��H;/�H;��H;��H;X�H;`�H;~�H;��H;��H;B�H;��H;��H;x�H;;�H;/�H;C�H;u�H;�I;�I;I;%I;.
I;I;�I;SI;�I;�I;oI;�I;      �I;�I;I;5I;�I;aI;�I;xI;FI;�I;"I;�	I;�I;:I;�I;�H;��H;=�H;�H;4�H;o�H;��H;�H;��H;��H;i�H;Z�H;��H;��H;�H;��H;C�H;��H;��H;g�H;J�H;9�H;J�H;g�H;��H;��H;C�H;��H;�H;��H;��H;Z�H;i�H;��H;��H;�H;��H;o�H;4�H;�H;=�H;��H;�H;�I;:I;�I;�	I;"I;�I;FI;xI;�I;aI;�I;5I;I;�I;      !I;!I;\!I;e!I;
!I;? I;�I;mI;�I;�I;�I;�I;AI;�	I;�I;�I;� I;��H;I�H;��H;��H;��H;��H;0�H;��H;��H;X�H;O�H;��H;��H;/�H;��H;M�H;��H;��H;��H;��H;��H;��H;��H;M�H;��H;/�H;��H;��H;O�H;X�H;��H;��H;0�H;��H;��H;��H;��H;I�H;��H;� I;�I;�I;�	I;AI;�I;�I;�I;�I;mI;�I;? I;
!I;e!I;\!I;!I;      �H;s�H;�I;�I;�I;�I;tI;�I;� I;wI;�I;�I;�I;I;$I;Y	I;�I;oI;L�H;A�H;��H;F�H; �H;$�H;@�H;��H;��H;k�H;O�H;��H;��H;;�H;��H;|�H;9�H;
�H;�H;
�H;9�H;|�H;��H;;�H;��H;��H;O�H;k�H;��H;��H;@�H;$�H; �H;F�H;��H;A�H;L�H;oI;�I;Y	I;$I;I;�I;�I;�I;wI;� I;�I;tI;�I;�I;�I;�I;s�H;      �MH;�SH;�cH;�|H;�H;o�H;��H;��H;�
I;7I; I;/ I;�I;OI;�I;8I;�I;�I;�I;� I;�H;�H;��H;Y�H;-�H;Z�H;��H;��H;X�H;Z�H;��H;��H;d�H;��H;��H;��H;��H;��H;��H;��H;d�H;��H;��H;Z�H;X�H;��H;��H;Z�H;-�H;Y�H;��H;�H;�H;� I;�I;�I;�I;8I;�I;OI;�I;/ I; I;7I;�
I;��H;��H;o�H;�H;�|H;�cH;�SH;      �HF;�XF;�F;�F;�&G;�G;��G;9BH;Q�H;p�H;��H;I;	I;�I;I;I;�I; I;i	I;"I;VI;��H;��H;��H;w�H;S�H;Z�H;��H;��H;i�H;X�H;��H;&�H;��H;@�H;"�H;�H;"�H;@�H;��H;&�H;��H;X�H;i�H;��H;��H;Z�H;S�H;w�H;��H;��H;��H;VI;"I;i	I; I;�I;I;I;�I;	I;I;��H;p�H;Q�H;9BH;��G;�G;�&G;�F;�F;�XF;      DA;(kA;��A;��B;�iC;o`D;�[E;IF;�G;��G;�MH;R�H;��H;�I;�I;yI;I;ZI;�I;�
I;I;�I;4�H;��H;��H;w�H;-�H;@�H;��H;��H;`�H;u�H;��H;O�H;��H;��H;��H;��H;��H;O�H;��H;u�H;`�H;��H;��H;@�H;-�H;w�H;��H;��H;4�H;�I;I;�
I;�I;ZI;I;yI;�I;�I;��H;R�H;�MH;��G;�G;IF;�[E;o`D;�iC;��B;��A;(kA;      �I6;&�6;ږ7;�9;l;;0-=;li?;y�A;C�C;v1E;چF;t�G;�;H;��H;��H;�I;gI;9I;CI;WI;�I;�I;RI;E�H;��H;��H;Y�H;$�H;0�H;��H;~�H;e�H;��H;�H;��H;]�H;:�H;]�H;��H;�H;��H;e�H;~�H;��H;0�H;$�H;Y�H;��H;��H;E�H;RI;�I;�I;WI;CI;9I;gI;�I;��H;��H;�;H;t�G;چF;v1E;C�C;y�A;li?;0-=;l;;�9;ږ7;&�6;      do ; !;#;)&;%*;o.;�3;�7;��;;Ai?;jjB;8�D;�wF;�G;cH;,�H;�	I;�I;rI;�I;9I;6I;�I;RI;4�H;��H;��H; �H;��H;�H;��H;x�H;��H;��H;E�H;�H;��H;�H;E�H;��H;��H;x�H;��H;�H;��H; �H;��H;��H;4�H;RI;�I;6I;9I;�I;rI;�I;�	I;,�H;cH;�G;�wF;8�D;jjB;Ai?;��;;�7;�3;o.;%*;)&;#; !;      �r�:���:�j�:o�;��	;�;Vy;5O$;y�,;��3;4�9;1�>;>�B;C1E;*�F;uH;��H;��H;,I;I;BI;�I;6I;�I;�I;��H;�H;F�H;��H;��H;��H;��H;��H;��H;)�H;��H;��H;��H;)�H;��H;��H;��H;��H;��H;��H;F�H;�H;��H;�I;�I;6I;�I;BI;I;,I;��H;��H;uH;*�F;C1E;>�B;1�>;4�9;��3;y�,;5O$;Vy;�;��	;o�;�j�:���:      ��>:8�G:~�b:г�:���:	3�:>)�:�h;o�;#a;:*;mq3;��:;� @;��C;�HF;ɾG;ӍH;.�H;zI;I;BI;9I;�I;I;VI;�H;��H;��H;o�H;B�H;��H;��H;��H;	�H;��H;y�H;��H;	�H;��H;��H;��H;B�H;o�H;��H;��H;�H;VI;I;�I;9I;BI;I;zI;.�H;ӍH;ɾG;�HF;��C;� @;��:;mq3;:*;#a;o�;�h;>)�:	3�:���:г�:~�b:8�G:      ��������wk��� ��
���!69��!:Ǌ:�2�:B�:��;';v�,;�6;��=;��B;��E;|�G;�{H;��H;zI;I;�I;WI;�
I;"I;� I;A�H;��H;4�H;��H;�H;��H;��H;��H;}�H;k�H;}�H;��H;��H;��H;�H;��H;4�H;��H;A�H;� I;"I;�
I;WI;�I;I;zI;��H;�{H;|�G;��E;��B;��=;�6;v�,;';��;B�:�2�:Ǌ:��!:�!69�
���� ��wk����      �/��s�����x�k�X�c�/�˻ �����u�l3�9��k:�:�m�:�A;!&;l3;�<;J�A;�oE;hsG;�{H;.�H;,I;rI;CI;�I;i	I;�I;L�H;I�H;�H;��H;x�H;��H;��H;��H;l�H;\�H;l�H;��H;��H;��H;x�H;��H;�H;I�H;L�H;�I;i	I;�I;CI;rI;,I;.�H;�{H;hsG;�oE;J�A;�<;l3;!&;�A;�m�:�:��k:l3�9u칋���˻ �c�/�k�X���x�s���      ������q
�q�����׻S,��"����;�Snۺ<� ��I�9;Ǌ:���:� ;J!;Ģ0;=;;̒A;�oE;|�G;ӍH;��H;�I;9I;ZI; I;�I;oI;��H;=�H;x�H;�H;�H;��H;��H;[�H;1�H;[�H;��H;��H;�H;�H;x�H;=�H;��H;oI;�I; I;ZI;9I;�I;��H;ӍH;|�G;�oE;̒A;=;;Ģ0;J!;� ;���:;Ǌ:�I�9<� �Snۺ�;�"���S,����׻q����q
���      �����8����_�k�ɆO�4/�VB�\�׻����@��Q����)�>:h3�:�;�a;��/;=;;J�A;��E;ɾG;��H;�	I;gI;I;�I;�I;�I;� I;��H;;�H;��H;��H;��H;�H;c�H;)�H;c�H;�H;��H;��H;��H;;�H;��H;� I;�I;�I;�I;I;gI;�	I;��H;ɾG;��E;J�A;=;;��/;�a;�;h3�:)�>:���Q���@����\�׻VB�4/�ɆO�_�k����8��      F��	}�;�ݼ��˼"d��-��	�}�&�G������һ�������"/�k:�ճ:#�;�a;Ģ0;�<;��B;�HF;uH;,�H;�I;yI;I;8I;Y	I;�I;�H;/�H;T�H;�H;#�H;�H;r�H;5�H;r�H;�H;#�H;�H;T�H;/�H;�H;�I;Y	I;8I;I;yI;�I;,�H;uH;�HF;��B;�<;Ģ0;�a;#�;�ճ:k:�"/���������һ���&�G�	�}�-��"d����˼;�ݼ	}�      F�B�MR?��5���&��3��J��߮Ҽ0F����c=�I?�c.����/��qk����9�ճ:�;J!;l3;��=;��C;*�F;cH;��H;�I;I;�I;$I;�I;�I;C�H;��H;��H;|�H;?�H;|�H;3�H;|�H;?�H;|�H;��H;��H;C�H;�I;�I;$I;�I;I;�I;��H;cH;*�F;��C;��=;l3;J!;�;�ճ:���9�qk���/�c.��I?�c=���0F��߮Ҽ�J���3���&��5�MR?�      &��"W��撐�!�����j�Q`I���&����Oϼ�,���T[����I��;��qk�k:h3�:� ;!&;�6;� @;C1E;�G;��H;�I;�I;OI;I;�	I;:I;u�H;��H;�H;��H;^�H;��H;D�H;��H;^�H;��H;�H;��H;u�H;:I;�	I;I;OI;�I;�I;��H;�G;C1E;� @;�6;!&;� ;h3�:k:�qk�;��I�����T[��,��Oϼ�����&�Q`I���j�!���撐�"W��      �J���D��ͽ���$�������L�(��.��;��%�k����I����/��"/�)�>:���:�A;v�,;��:;>�B;�wF;�;H;��H;	I;�I;�I;AI;�I;�I;��H;s�H;4�H;n�H;��H;l�H;��H;n�H;4�H;s�H;��H;�I;�I;AI;�I;�I;	I;��H;�;H;�wF;>�B;��:;v�,;�A;���:)�>:�"/���/��I����%�k�;��.��(����L����$������ͽ�Dὼ��      K�:��*7���,�+�~�	�j��~���W����j�?�/��J���I��%�k���c.������;Ǌ:�m�:';mq3;1�>;8�D;t�G;R�H;I;/ I;�I;�I;�	I;�I;`�H;��H;��H;��H;��H;^�H;��H;��H;��H;��H;`�H;�I;�	I;�I;�I;/ I;I;R�H;t�G;8�D;1�>;mq3;';�m�:;Ǌ:����c.����%�k��I���J��?�/���j�W��~���j��~�	�+���,��*7�      ^���p��
��)�l���M���,�Tl�K9ݽ�A���{���5��J��;���T[�I?������Q���I�9�:��;:*;4�9;jjB;چF;�MH;��H; I;�I;�I;"I;I;@I;^�H;��H;��H;��H;j�H;��H;��H;��H;^�H;@I;I;"I;�I;�I; I;��H;�MH;چF;jjB;4�9;:*;��;�:�I�9�Q������I?��T[�;���J����5��{��A��K9ݽTl���,���M�)�l�
���p��      +m־G�Ѿ�>ľ����̗����{���I�+����V���{�?�/�.���,��c=���һ�@�<� ���k:B�:#a;��3;Ai?;v1E;��G;p�H;7I;wI;�I;�I;%I;�I;��H;��H;��H;��H;V�H;��H;��H;��H;��H;�I;%I;�I;�I;wI;7I;p�H;��G;v1E;Ai?;��3;#a;B�:��k:<� ��@���һc=��,��.��?�/��{��V�����+���I���{�̗�������>ľG�Ѿ      =\����l5��z ��E۾�ճ��]��q�Z�F?#����A����j�(��Oϼ��������Snۺl3�9�2�:o�;y�,;��;;C�C;�G;Q�H;�
I;� I;�I;FI;.
I;�I;> I;�H;�H;��H;!�H;��H;�H;�H;> I;�I;.
I;FI;�I;� I;�
I;Q�H;�G;C�C;��;;y�,;o�;�2�:l3�9Snۺ��������Oϼ(����j��A�����F?#�q�Z��]���ճ��E۾�z �l5����      <�b��>]���M���6�����$���>ľq��q�Z�+�K9ݽW����L����0F��&�G�\�׻�;�u�Ǌ:�h;5O$;�7;y�A;IF;9BH;��H;�I;mI;xI;I;-I;�I;�H;��H;��H;�H;��H;��H;�H;�I;-I;I;xI;mI;�I;��H;9BH;IF;y�A;�7;5O$;�h;Ǌ:u칹;�\�׻&�G�0F�������L�W��K9ݽ+�q�Z�q���>ľ�$�������6���M��>]�      �o��벗����-�y�s�R���)�iv��>ľ�]����I�Tl�~��������&�߮Ҽ	�}�VB�"���������!:>)�:Vy;�3;li?;�[E;��G;��H;tI;�I;�I;�I;|I;�I;�H;��H;c�H;��H;c�H;��H;�H;�I;|I;�I;�I;�I;tI;��H;��G;�[E;li?;�3;Vy;>)�:��!:����"���VB�	�}�߮Ҽ��&����~���Tl���I��]���>ľiv���)�s�R�-�y����벗�      �˿�<ƿjL��:1��蟉��>]���)��$���ճ���{���,�j��$��Q`I��J��-��4/�S,��˻ ��!69	3�:�;o.;0-=;o`D;�G;o�H;�I;? I;aI;SI;�I;�I;��H;��H;�H;d�H;�H;��H;��H;�I;�I;SI;aI;? I;�I;o�H;�G;o`D;0-=;o.;�;	3�:�!69˻ �S,��4/�-���J��Q`I�$��j�齞�,���{��ճ��$����)��>]�蟉�:1��jL���<ƿ      ����2���K[忭˿�T��蟉�s�R�����E۾̗����M�~�	������j��3�"d��ɆO���׻c�/��
�����:��	;%*;l;;�iC;�&G;�H;�I;
!I;�I;�I;�	I;�I;� I;I�H;��H; �H;��H;I�H;� I;�I;�	I;�I;�I;
!I;�I;�H;�&G;�iC;l;;%*;��	;���:�
��c�/���׻ɆO�"d���3���j����~�	���M�̗���E۾���s�R�蟉��T���˿K[�2���      O�0��o����˿:1��-�y���6��z �����)�l�+��ͽ!�����&���˼_�k�q���k�X��� �г�:o�;)&;�9;��B;�F;�|H;�I;e!I;5I;�I;�
I;qI;FI;��H;"�H;��H;"�H;��H;FI;qI;�
I;�I;5I;e!I;�I;�|H;�F;��B;�9;)&;o�;г�:�� �k�X�q���_�k���˼��&�!����ͽ+�)�l������z ���6�-�y�:1���˿���o�0��      ��*��g&��#�o�K[�jL�������M�l5��>ľ
����,��D�撐��5�;�ݼ���q
���x��wk�~�b:�j�:#;ږ7;��A;�F;�cH;�I;\!I;I;oI;AI;�I;�I; �H;x�H;��H;x�H; �H;�I;�I;AI;oI;I;\!I;�I;�cH;�F;��A;ږ7;#;�j�:~�b:�wk���x��q
���;�ݼ�5�撐��Dὤ�,�
���>ľl5���M����jL��K[�o��#��g&�      ��8��4��g&�0��2����<ƿ벗��>]����G�Ѿ�p���*7����"W��MR?�	}鼀8����s������8�G:���: !;&�6;(kA;�XF;�SH;s�H;!I;�I;�I;�I;FI;�I;e�H;��H;�H;��H;e�H;�I;FI;�I;�I;�I;!I;s�H;�SH;�XF;(kA;&�6; !;���:8�G:���s������8��	}�MR?�"W�����*7��p��G�Ѿ����>]�벗��<ƿ2���0���g&��4�      �Aq���i���U�A:�@�����6���q���uA�a5�� ��y^Z�����A���]�����d��|",�6��:�Ѻ���9'��:d�;dX4;p�@;�UF;��H;�FI;�aI;2NI;A9I;�(I;=I;�I;�I;�I;�
I;�I;�I;�I;=I;�(I;A9I;2NI;�aI;�FI;��H;�UF;p�@;dX4;d�;'��:���9:�Ѻ6��|",��d������]��A�����y^Z�� ��a5�uA�q���6�������@�A:���U���i�      ��i���b�T�O�.5�-i������������q<�����e��[
V�FE	�!���IY�s9�Z����(� S����Ⱥ��:���:'�;L�4;h�@;kgF;��H;4HI;�aI;�MI;�8I;�(I;I;~I;�I;{I;x
I;{I;�I;~I;I;�(I;�8I;�MI;�aI;4HI;��H;kgF;h�@;L�4;'�;���:��:��Ⱥ S���(�Z���s9��IY�!��FE	�[
V��e������q<������������-i�.5�T�O���b�      ��U�T�O�B-?�(�'���F�`欿Y�{�aa/���뾙���I����e���ZN�o5��Ǩ��nH�� ������ݧ":��:��;��5;�_A;ٚF;Z�H;<LI;aI;�LI;�7I;(I;aI;I;_I;&I;&
I;&I;_I;I;aI;(I;�7I;�LI;aI;<LI;Z�H;ٚF;�_A;��5;��;��:ݧ":����� ��nH�Ǩ��o5���ZN�e������I�������aa/�Y�{��欿F����(�'�B-?�T�O�      A:�.5�(�'��������dȿ���e$_���Q�Ҿؕ��
�6�����*���`=�P���)��{G��6��B����Q:�:/";�7;�%B;�F;��H;RI;�_I;�JI;C6I;�&I;ZI;7I;�I;�
I;�	I;�
I;�I;7I;ZI;�&I;C6I;�JI;�_I;RI;��H;�F;�%B;�7;/";�:��Q:B���6��{G��)��P���`=��*�����
�6�ؕ��Q�Ҿ��e$_����dȿ�������(�'�.5�      @�-i�������B�ѿf�������q<��:��a����q����Wн齅���'�ib̼�zl�/���X�z�� �:��;
�&;٪9;KC;wLG;�H;]XI;�]I;�GI;4I;�$I;I;'I;�I;�	I;�I;�	I;�I;'I;I;�$I;4I;�GI;�]I;]XI;�H;wLG;KC;٪9;
�&;��; �:z���X�/���zl�ib̼��'�齅��Wн����q��a���:��q<����f���B�ѿ������-i�      �������F��dȿf���������O���u]׾w���	�I�����A��C�d�v��֮�<RH�Kkλ �$�s5����:mM;˅+;�<;"3D;�G;�I;�]I;�ZI;	DI;H1I;�"I;`I;�I;�I;�I;�I;�I;�I;�I;`I;�"I;H1I;	DI;�ZI;�]I;�I;�G;"3D;�<;˅+;mM;���:s5� �$�Kkλ<RH��֮�v�C�d��A�����	�I�w���u]׾����O�����f���dȿF�ῢ��      6��������欿��������O�}x����� ���l���"��ܽ���`=�Ý��l"��R���ۺO��9�=�:�K;��0;͞>;�LE;|"H;�$I;�`I;(VI;�?I;.I;` I;[I;"I;/
I;lI;�I;lI;/
I;"I;[I;` I;.I;�?I;(VI;�`I;�$I;|"H;�LE;͞>;��0;�K;�=�:O��9�ۺ�R��l"����Ý��`=����ܽ��"��l�� �����}x���O��������欿����      q�������Y�{�e$_��q<�������}��w���6�����!��!�h��������� d��.��g_e�TL[���Z:���:�+ ;��5;�A;�UF;˃H;@I;�aI;�PI;;I;e*I;�I;+I;WI;�I;I;LI;I;�I;WI;+I;�I;e*I;;I;�PI;�aI;@I;˃H;�UF;�A;��5;�+ ;���:��Z:TL[�g_e��.��� d��������!�h�!�������6�w���}��������q<�e$_�Y�{�����      uA��q<�aa/����:�u]׾� ��w��>�BE	�����ܽ����3�r�꼰���>",�X��3��LAQ�خ�:�L
;�e);ބ:;D?C;?G;|�H;fSI;�^I;KJI;6I;t&I;�I;�I;ZI;�I;�I;�I;�I;�I;ZI;�I;�I;t&I;6I;KJI;�^I;fSI;|�H;?G;D?C;ބ:;�e);�L
;خ�:LAQ�3��X��>",�����r�꼠�3�ܽ������BE	�>�w��� ��u]׾�:���aa/��q<�      a5�������Q�Ҿ�a��w����l��6�BE	���Ƚk���aG����z֮�C�W����:�k����U`,:���:�;��1;m�>;^E;L�G;BI;G^I;hYI;ZCI;�0I;V"I;cI;I;#	I;,I;�I;=I;�I;,I;#	I;I;cI;V"I;�0I;ZCI;hYI;G^I;BI;L�G;^E;m�>;��1;�;���:U`,:���:�k����C�W�z֮�����aG�k����ȽBE	��6��l�w����a��Q�Ҿ������      � ���e�����ؕ����q�	�I���"���������k���ZN�c�6¼~�y��$�PR��]� ���[��:G/;J�&;
w8;��A;��F;��H;?I;aI;�QI;:<I;7+I;�I;I;uI;�I;WI;9I;� I;9I;WI;�I;uI;I;�I;7+I;:<I;�QI;aI;?I;��H;��F;��A;
w8;J�&;G/;�:��[�]� �PR���$�~�y�6¼c��ZN�k������������"�	�I���q�ؕ������e��      y^Z�[
V��I�
�6�������ܽ!��ܽ���aG�c��ȼ�)����(����H5���.�Z:k�:7R;/&1;��=;ПD;P�G;�H;�WI;9]I;�HI;5I;�%I;�I;�I;�	I;�I;mI;|�H;��H;|�H;mI;�I;�	I;�I;�I;�%I;5I;�HI;9]I;�WI;�H;P�G;ПD;��=;/&1;7R;k�:.�Z:��H5������(��)���ȼc��aG�ܽ��!���ܽ�����
�6��I�[
V�      ���FE	��������Wн�A����!�h���3����6¼�)��ax/�v�һC�X� %����9���:�=;[e);�_9;�%B;ډF;�|H;�5I;u`I;�TI;�?I;�-I; I;jI;DI;�I;jI;q�H;��H;�H;��H;q�H;jI;�I;DI;jI; I;�-I;�?I;�TI;u`I;�5I;�|H;ډF;�%B;�_9;[e);�=;���:��9 %��C�X�v�һax/��)��6¼�����3�!�h��󑽢A���Wн��콹��FE	�      �A��!��e���*��齅�C�d��`=����r��z֮�~�y���(�v�һj^e����� �f9���:X�;m0";A�4;�l?;E;��G;��H;�VI;�]I;(JI;�6I;'I;�I;FI;�	I;>I;7 I;��H;��H;V�H;��H;��H;7 I;>I;�	I;FI;�I;'I;�6I;(JI;�]I;�VI;��H;��G;E;�l?;A�4;m0";X�;���: �f9����j^e�v�һ��(�~�y�z֮�r�꼠���`=�C�d�齅��*��e��!��      �]��IY��ZN��`=���'�v�Ý���������C�W��$����C�X������9�ޚ:���:��;˷0;�<;v�C;GG;�H;�>I;P`I;�SI;^?I;1.I;z I;�I;.I;�I;�I;��H;��H;&�H;��H;&�H;��H;��H;�I;�I;.I;�I;z I;1.I;^?I;�SI;P`I;�>I;�H;GG;v�C;�<;˷0;��;���:�ޚ:�9����C�X�����$�C�W���������Ý�v���'��`=��ZN��IY�      ���s9�o5��P��ib̼�֮����� d�>",����PR��H5� %�� �f9�ޚ:��:6�;��-;��:;KB;_UF;:JH; I;�[I;G[I;�GI;%5I;<&I;7I;�I;9	I;^I;�H;��H;��H;n�H;�H;n�H;��H;��H;�H;^I;9	I;�I;7I;<&I;%5I;�GI;G[I;�[I; I;:JH;_UF;KB;��:;��-;6�;��:�ޚ: �f9 %��H5�PR�����>",�� d�����֮�ib̼P��o5��s9�      �d��Z���Ǩ���)���zl�<RH�l"��.��X��:�k�]� �����9���:���:6�;�-;�9;j`A;۹E;J�G;��H;#RI;4_I;OI;�;I;�+I;�I;MI;)I;�I;p I;��H;��H;��H;��H;|�H;��H;��H;��H;��H;p I;�I;)I;MI;�I;�+I;�;I;OI;4_I;#RI;��H;J�G;۹E;j`A;�9;�-;6�;���:���:��9��]� �:�k�X���.��l"�<RH��zl��)��Ǩ��Z���      |",��(�nH�{G�/��Kkλ�R��g_e�3�������[�.�Z:���:X�;��;��-;�9;�A;�bE;D�G;��H;tFI;`I;�TI;bAI;�0I;#I;�I;I;�I;I;��H;b�H;��H;!�H;,�H;��H;,�H;!�H;��H;b�H;��H;I;�I;I;�I;#I;�0I;bAI;�TI;`I;tFI;��H;D�G;�bE;�A;�9;��-;��;X�;���:.�Z:��[����3��g_e��R��Kkλ/��{G�nH��(�      6�� S��� ���6���X� �$��ۺTL[�LAQ�U`,:�:k�:�=;m0";˷0;��:;j`A;�bE;�G;��H;�<I;N_I;�XI;FI;5I;�&I;I;�I;
I;�I;��H;�H;6�H;�H;��H;��H;S�H;��H;��H;�H;6�H;�H;��H;�I;
I;�I;I;�&I;5I;FI;�XI;N_I;�<I;��H;�G;�bE;j`A;��:;˷0;m0";�=;k�:�:U`,:LAQ�TL[��ۺ �$��X��6��� �� S��      :�Ѻ��Ⱥ����B��z��s5�O��9��Z:خ�:���:G/;7R;[e);A�4;�<;KB;۹E;D�G;��H;�9I;q^I;�ZI;?II;8I;�)I;�I;I;I;vI;$ I;��H;��H;%�H;C�H;�H;F�H;��H;F�H;�H;C�H;%�H;��H;��H;$ I;vI;I;I;�I;�)I;8I;?II;�ZI;q^I;�9I;��H;D�G;۹E;KB;�<;A�4;[e);7R;G/;���:خ�:��Z:O��9s5�z��B��������Ⱥ      ���9��:ݧ":��Q: �:���:�=�:���:�L
;�;J�&;/&1;�_9;�l?;v�C;_UF;J�G;��H;�<I;q^I;1[I;�JI;1:I;�+I;�I;I;�I;�I;`I;��H;K�H;��H;J�H;��H;��H;��H;��H;��H;��H;��H;J�H;��H;K�H;��H;`I;�I;�I;I;�I;�+I;1:I;�JI;1[I;q^I;�<I;��H;J�G;_UF;v�C;�l?;�_9;/&1;J�&;�;�L
;���:�=�:���: �:��Q:ݧ":��:      '��:���:��:�:��;mM;�K;�+ ;�e);��1;
w8;��=;�%B;E;GG;:JH;��H;tFI;N_I;�ZI;�JI;�:I;-I;H!I;QI;*I;0I;xI;��H;��H;��H;}�H;��H;-�H;R�H;��H;y�H;��H;R�H;-�H;��H;}�H;��H;��H;��H;xI;0I;*I;QI;H!I;-I;�:I;�JI;�ZI;N_I;tFI;��H;:JH;GG;E;�%B;��=;
w8;��1;�e);�+ ;�K;mM;��;�:��:���:      d�;'�;��;/";
�&;˅+;��0;��5;ބ:;m�>;��A;ПD;ډF;��G;�H; I;#RI;`I;�XI;?II;1:I;-I;�!I;I;�I;	I;BI;]�H;��H;j�H;��H;��H;�H;��H; �H;��H;p�H;��H; �H;��H;�H;��H;��H;j�H;��H;]�H;BI;	I;�I;I;�!I;-I;1:I;?II;�XI;`I;#RI; I;�H;��G;ډF;ПD;��A;m�>;ބ:;��5;��0;˅+;
�&;/";��;'�;      dX4;L�4;��5;�7;٪9;�<;͞>;�A;D?C;^E;��F;P�G;�|H;��H;�>I;�[I;4_I;�TI;FI;8I;�+I;H!I;I;9I;v	I;�I; �H;��H;��H;��H;��H;�H;��H;��H;��H;��H;u�H;��H;��H;��H;��H;�H;��H;��H;��H;��H; �H;�I;v	I;9I;I;H!I;�+I;8I;FI;�TI;4_I;�[I;�>I;��H;�|H;P�G;��F;^E;D?C;�A;͞>;�<;٪9;�7;��5;L�4;      p�@;h�@;�_A;�%B;KC;"3D;�LE;�UF;?G;L�G;��H;�H;�5I;�VI;P`I;G[I;OI;bAI;5I;�)I;�I;QI;�I;v	I;I;.�H;D�H;��H;0�H;��H;�H;��H;[�H;��H;��H;��H;r�H;��H;��H;��H;[�H;��H;�H;��H;0�H;��H;D�H;.�H;I;v	I;�I;QI;�I;�)I;5I;bAI;OI;G[I;P`I;�VI;�5I;�H;��H;L�G;?G;�UF;�LE;"3D;KC;�%B;�_A;h�@;      �UF;kgF;ٚF;�F;wLG;�G;|"H;˃H;|�H;BI;?I;�WI;u`I;�]I;�SI;�GI;�;I;�0I;�&I;�I;I;*I;	I;�I;.�H;V�H;'�H;i�H;��H;�H;��H;V�H;L�H;��H;�H;��H;��H;��H;�H;��H;L�H;V�H;��H;�H;��H;i�H;'�H;V�H;.�H;�I;	I;*I;I;�I;�&I;�0I;�;I;�GI;�SI;�]I;u`I;�WI;?I;BI;|�H;˃H;|"H;�G;wLG;�F;ٚF;kgF;      ��H;��H;Z�H;��H;�H;�I;�$I;@I;fSI;G^I;aI;9]I;�TI;(JI;^?I;%5I;�+I;#I;I;I;�I;0I;BI; �H;D�H;'�H;\�H;�H;7�H;|�H;7�H;�H;F�H;��H;@�H;��H;��H;��H;@�H;��H;F�H;�H;7�H;|�H;7�H;�H;\�H;'�H;D�H; �H;BI;0I;�I;I;I;#I;�+I;%5I;^?I;(JI;�TI;9]I;aI;G^I;fSI;@I;�$I;�I;�H;��H;Z�H;��H;      �FI;4HI;<LI;RI;]XI;�]I;�`I;�aI;�^I;hYI;�QI;�HI;�?I;�6I;1.I;<&I;�I;�I;�I;I;�I;xI;]�H;��H;��H;i�H;�H;�H;��H;2�H;�H;�H;p�H;��H;|�H;F�H;@�H;F�H;|�H;��H;p�H;�H;�H;2�H;��H;�H;�H;i�H;��H;��H;]�H;xI;�I;I;�I;�I;�I;<&I;1.I;�6I;�?I;�HI;�QI;hYI;�^I;�aI;�`I;�]I;]XI;RI;<LI;4HI;      �aI;�aI;aI;�_I;�]I;�ZI;(VI;�PI;KJI;ZCI;:<I;5I;�-I;'I;z I;7I;MI;I;
I;vI;`I;��H;��H;��H;0�H;��H;7�H;��H;)�H;�H; �H;B�H;��H;2�H;��H;��H;��H;��H;��H;2�H;��H;B�H; �H;�H;)�H;��H;7�H;��H;0�H;��H;��H;��H;`I;vI;
I;I;MI;7I;z I;'I;�-I;5I;:<I;ZCI;KJI;�PI;(VI;�ZI;�]I;�_I;aI;�aI;      2NI;�MI;�LI;�JI;�GI;	DI;�?I;;I;6I;�0I;7+I;�%I; I;�I;�I;�I;)I;�I;�I;$ I;��H;��H;j�H;��H;��H;�H;|�H;2�H;�H;�H;1�H;��H;��H;��H;H�H;(�H;%�H;(�H;H�H;��H;��H;��H;1�H;�H;�H;2�H;|�H;�H;��H;��H;j�H;��H;��H;$ I;�I;�I;)I;�I;�I;�I; I;�%I;7+I;�0I;6I;;I;�?I;	DI;�GI;�JI;�LI;�MI;      A9I;�8I;�7I;C6I;4I;H1I;.I;e*I;t&I;V"I;�I;�I;jI;FI;.I;9	I;�I;I;��H;��H;K�H;��H;��H;��H;�H;��H;7�H;�H; �H;1�H;��H;��H;d�H;�H;��H;��H;��H;��H;��H;�H;d�H;��H;��H;1�H; �H;�H;7�H;��H;�H;��H;��H;��H;K�H;��H;��H;I;�I;9	I;.I;FI;jI;�I;�I;V"I;t&I;e*I;.I;H1I;4I;C6I;�7I;�8I;      �(I;�(I;(I;�&I;�$I;�"I;` I;�I;�I;cI;I;�I;DI;�	I;�I;^I;p I;��H;�H;��H;��H;}�H;��H;�H;��H;V�H;�H;�H;B�H;��H;��H;{�H;��H;��H;z�H;T�H;>�H;T�H;z�H;��H;��H;{�H;��H;��H;B�H;�H;�H;V�H;��H;�H;��H;}�H;��H;��H;�H;��H;p I;^I;�I;�	I;DI;�I;I;cI;�I;�I;` I;�"I;�$I;�&I;(I;�(I;      =I;I;aI;ZI;I;`I;[I;+I;�I;I;uI;�	I;�I;>I;�I;�H;��H;b�H;6�H;%�H;J�H;��H;�H;��H;[�H;L�H;F�H;p�H;��H;��H;d�H;��H;��H;\�H;�H;�H;�H;�H;�H;\�H;��H;��H;d�H;��H;��H;p�H;F�H;L�H;[�H;��H;�H;��H;J�H;%�H;6�H;b�H;��H;�H;�I;>I;�I;�	I;uI;I;�I;+I;[I;`I;I;ZI;aI;I;      �I;~I;I;7I;'I;�I;"I;WI;ZI;#	I;�I;�I;jI;7 I;��H;��H;��H;��H;�H;C�H;��H;-�H;��H;��H;��H;��H;��H;��H;2�H;��H;�H;��H;\�H; �H;��H;��H;��H;��H;��H; �H;\�H;��H;�H;��H;2�H;��H;��H;��H;��H;��H;��H;-�H;��H;C�H;�H;��H;��H;��H;��H;7 I;jI;�I;�I;#	I;ZI;WI;"I;�I;'I;7I;I;~I;      �I;�I;_I;�I;�I;�I;/
I;�I;�I;,I;WI;mI;q�H;��H;��H;��H;��H;!�H;��H;�H;��H;R�H; �H;��H;��H;�H;@�H;|�H;��H;H�H;��H;z�H;�H;��H;��H;��H;��H;��H;��H;��H;�H;z�H;��H;H�H;��H;|�H;@�H;�H;��H;��H; �H;R�H;��H;�H;��H;!�H;��H;��H;��H;��H;q�H;mI;WI;,I;�I;�I;/
I;�I;�I;�I;_I;�I;      �I;{I;&I;�
I;�	I;�I;lI;I;�I;�I;9I;|�H;��H;��H;&�H;n�H;��H;,�H;��H;F�H;��H;��H;��H;��H;��H;��H;��H;F�H;��H;(�H;��H;T�H;�H;��H;��H;��H;}�H;��H;��H;��H;�H;T�H;��H;(�H;��H;F�H;��H;��H;��H;��H;��H;��H;��H;F�H;��H;,�H;��H;n�H;&�H;��H;��H;|�H;9I;�I;�I;I;lI;�I;�	I;�
I;&I;{I;      �
I;x
I;&
I;�	I;�I;�I;�I;LI;�I;=I;� I;��H;�H;V�H;��H;�H;|�H;��H;S�H;��H;��H;y�H;p�H;u�H;r�H;��H;��H;@�H;��H;%�H;��H;>�H;�H;��H;��H;}�H;��H;}�H;��H;��H;�H;>�H;��H;%�H;��H;@�H;��H;��H;r�H;u�H;p�H;y�H;��H;��H;S�H;��H;|�H;�H;��H;V�H;�H;��H;� I;=I;�I;LI;�I;�I;�I;�	I;&
I;x
I;      �I;{I;&I;�
I;�	I;�I;lI;I;�I;�I;9I;|�H;��H;��H;&�H;n�H;��H;,�H;��H;F�H;��H;��H;��H;��H;��H;��H;��H;F�H;��H;(�H;��H;T�H;�H;��H;��H;��H;}�H;��H;��H;��H;�H;T�H;��H;(�H;��H;F�H;��H;��H;��H;��H;��H;��H;��H;F�H;��H;,�H;��H;n�H;&�H;��H;��H;|�H;9I;�I;�I;I;lI;�I;�	I;�
I;&I;{I;      �I;�I;_I;�I;�I;�I;/
I;�I;�I;,I;WI;mI;q�H;��H;��H;��H;��H;!�H;��H;�H;��H;R�H; �H;��H;��H;�H;@�H;|�H;��H;H�H;��H;z�H;�H;��H;��H;��H;��H;��H;��H;��H;�H;z�H;��H;H�H;��H;|�H;@�H;�H;��H;��H; �H;R�H;��H;�H;��H;!�H;��H;��H;��H;��H;q�H;mI;WI;,I;�I;�I;/
I;�I;�I;�I;_I;�I;      �I;~I;I;7I;'I;�I;"I;WI;ZI;#	I;�I;�I;jI;7 I;��H;��H;��H;��H;�H;C�H;��H;-�H;��H;��H;��H;��H;��H;��H;2�H;��H;�H;��H;\�H; �H;��H;��H;��H;��H;��H; �H;\�H;��H;�H;��H;2�H;��H;��H;��H;��H;��H;��H;-�H;��H;C�H;�H;��H;��H;��H;��H;7 I;jI;�I;�I;#	I;ZI;WI;"I;�I;'I;7I;I;~I;      =I;I;aI;ZI;I;`I;[I;+I;�I;I;uI;�	I;�I;>I;�I;�H;��H;b�H;6�H;%�H;J�H;��H;�H;��H;[�H;L�H;F�H;p�H;��H;��H;d�H;��H;��H;\�H;�H;�H;�H;�H;�H;\�H;��H;��H;d�H;��H;��H;p�H;F�H;L�H;[�H;��H;�H;��H;J�H;%�H;6�H;b�H;��H;�H;�I;>I;�I;�	I;uI;I;�I;+I;[I;`I;I;ZI;aI;I;      �(I;�(I;(I;�&I;�$I;�"I;` I;�I;�I;cI;I;�I;DI;�	I;�I;^I;p I;��H;�H;��H;��H;}�H;��H;�H;��H;V�H;�H;�H;B�H;��H;��H;{�H;��H;��H;z�H;T�H;>�H;T�H;z�H;��H;��H;{�H;��H;��H;B�H;�H;�H;V�H;��H;�H;��H;}�H;��H;��H;�H;��H;p I;^I;�I;�	I;DI;�I;I;cI;�I;�I;` I;�"I;�$I;�&I;(I;�(I;      A9I;�8I;�7I;C6I;4I;H1I;.I;e*I;t&I;V"I;�I;�I;jI;FI;.I;9	I;�I;I;��H;��H;K�H;��H;��H;��H;�H;��H;7�H;�H; �H;1�H;��H;��H;d�H;�H;��H;��H;��H;��H;��H;�H;d�H;��H;��H;1�H; �H;�H;7�H;��H;�H;��H;��H;��H;K�H;��H;��H;I;�I;9	I;.I;FI;jI;�I;�I;V"I;t&I;e*I;.I;H1I;4I;C6I;�7I;�8I;      2NI;�MI;�LI;�JI;�GI;	DI;�?I;;I;6I;�0I;7+I;�%I; I;�I;�I;�I;)I;�I;�I;$ I;��H;��H;j�H;��H;��H;�H;|�H;2�H;�H;�H;1�H;��H;��H;��H;H�H;(�H;%�H;(�H;H�H;��H;��H;��H;1�H;�H;�H;2�H;|�H;�H;��H;��H;j�H;��H;��H;$ I;�I;�I;)I;�I;�I;�I; I;�%I;7+I;�0I;6I;;I;�?I;	DI;�GI;�JI;�LI;�MI;      �aI;�aI;aI;�_I;�]I;�ZI;(VI;�PI;KJI;ZCI;:<I;5I;�-I;'I;z I;7I;MI;I;
I;vI;`I;��H;��H;��H;0�H;��H;7�H;��H;)�H;�H; �H;B�H;��H;2�H;��H;��H;��H;��H;��H;2�H;��H;B�H; �H;�H;)�H;��H;7�H;��H;0�H;��H;��H;��H;`I;vI;
I;I;MI;7I;z I;'I;�-I;5I;:<I;ZCI;KJI;�PI;(VI;�ZI;�]I;�_I;aI;�aI;      �FI;4HI;<LI;RI;]XI;�]I;�`I;�aI;�^I;hYI;�QI;�HI;�?I;�6I;1.I;<&I;�I;�I;�I;I;�I;xI;]�H;��H;��H;i�H;�H;�H;��H;2�H;�H;�H;p�H;��H;|�H;F�H;@�H;F�H;|�H;��H;p�H;�H;�H;2�H;��H;�H;�H;i�H;��H;��H;]�H;xI;�I;I;�I;�I;�I;<&I;1.I;�6I;�?I;�HI;�QI;hYI;�^I;�aI;�`I;�]I;]XI;RI;<LI;4HI;      ��H;��H;Z�H;��H;�H;�I;�$I;@I;fSI;G^I;aI;9]I;�TI;(JI;^?I;%5I;�+I;#I;I;I;�I;0I;BI; �H;D�H;'�H;\�H;�H;7�H;|�H;7�H;�H;F�H;��H;@�H;��H;��H;��H;@�H;��H;F�H;�H;7�H;|�H;7�H;�H;\�H;'�H;D�H; �H;BI;0I;�I;I;I;#I;�+I;%5I;^?I;(JI;�TI;9]I;aI;G^I;fSI;@I;�$I;�I;�H;��H;Z�H;��H;      �UF;kgF;ٚF;�F;wLG;�G;|"H;˃H;|�H;BI;?I;�WI;u`I;�]I;�SI;�GI;�;I;�0I;�&I;�I;I;*I;	I;�I;.�H;V�H;'�H;i�H;��H;�H;��H;V�H;L�H;��H;�H;��H;��H;��H;�H;��H;L�H;V�H;��H;�H;��H;i�H;'�H;V�H;.�H;�I;	I;*I;I;�I;�&I;�0I;�;I;�GI;�SI;�]I;u`I;�WI;?I;BI;|�H;˃H;|"H;�G;wLG;�F;ٚF;kgF;      p�@;h�@;�_A;�%B;KC;"3D;�LE;�UF;?G;L�G;��H;�H;�5I;�VI;P`I;G[I;OI;bAI;5I;�)I;�I;QI;�I;v	I;I;.�H;D�H;��H;0�H;��H;�H;��H;[�H;��H;��H;��H;r�H;��H;��H;��H;[�H;��H;�H;��H;0�H;��H;D�H;.�H;I;v	I;�I;QI;�I;�)I;5I;bAI;OI;G[I;P`I;�VI;�5I;�H;��H;L�G;?G;�UF;�LE;"3D;KC;�%B;�_A;h�@;      dX4;L�4;��5;�7;٪9;�<;͞>;�A;D?C;^E;��F;P�G;�|H;��H;�>I;�[I;4_I;�TI;FI;8I;�+I;H!I;I;9I;v	I;�I; �H;��H;��H;��H;��H;�H;��H;��H;��H;��H;u�H;��H;��H;��H;��H;�H;��H;��H;��H;��H; �H;�I;v	I;9I;I;H!I;�+I;8I;FI;�TI;4_I;�[I;�>I;��H;�|H;P�G;��F;^E;D?C;�A;͞>;�<;٪9;�7;��5;L�4;      d�;'�;��;/";
�&;˅+;��0;��5;ބ:;m�>;��A;ПD;ډF;��G;�H; I;#RI;`I;�XI;?II;1:I;-I;�!I;I;�I;	I;BI;]�H;��H;j�H;��H;��H;�H;��H; �H;��H;p�H;��H; �H;��H;�H;��H;��H;j�H;��H;]�H;BI;	I;�I;I;�!I;-I;1:I;?II;�XI;`I;#RI; I;�H;��G;ډF;ПD;��A;m�>;ބ:;��5;��0;˅+;
�&;/";��;'�;      '��:���:��:�:��;mM;�K;�+ ;�e);��1;
w8;��=;�%B;E;GG;:JH;��H;tFI;N_I;�ZI;�JI;�:I;-I;H!I;QI;*I;0I;xI;��H;��H;��H;}�H;��H;-�H;R�H;��H;y�H;��H;R�H;-�H;��H;}�H;��H;��H;��H;xI;0I;*I;QI;H!I;-I;�:I;�JI;�ZI;N_I;tFI;��H;:JH;GG;E;�%B;��=;
w8;��1;�e);�+ ;�K;mM;��;�:��:���:      ���9��:ݧ":��Q: �:���:�=�:���:�L
;�;J�&;/&1;�_9;�l?;v�C;_UF;J�G;��H;�<I;q^I;1[I;�JI;1:I;�+I;�I;I;�I;�I;`I;��H;K�H;��H;J�H;��H;��H;��H;��H;��H;��H;��H;J�H;��H;K�H;��H;`I;�I;�I;I;�I;�+I;1:I;�JI;1[I;q^I;�<I;��H;J�G;_UF;v�C;�l?;�_9;/&1;J�&;�;�L
;���:�=�:���: �:��Q:ݧ":��:      :�Ѻ��Ⱥ����B��z��s5�O��9��Z:خ�:���:G/;7R;[e);A�4;�<;KB;۹E;D�G;��H;�9I;q^I;�ZI;?II;8I;�)I;�I;I;I;vI;$ I;��H;��H;%�H;C�H;�H;F�H;��H;F�H;�H;C�H;%�H;��H;��H;$ I;vI;I;I;�I;�)I;8I;?II;�ZI;q^I;�9I;��H;D�G;۹E;KB;�<;A�4;[e);7R;G/;���:خ�:��Z:O��9s5�z��B��������Ⱥ      6�� S��� ���6���X� �$��ۺTL[�LAQ�U`,:�:k�:�=;m0";˷0;��:;j`A;�bE;�G;��H;�<I;N_I;�XI;FI;5I;�&I;I;�I;
I;�I;��H;�H;6�H;�H;��H;��H;S�H;��H;��H;�H;6�H;�H;��H;�I;
I;�I;I;�&I;5I;FI;�XI;N_I;�<I;��H;�G;�bE;j`A;��:;˷0;m0";�=;k�:�:U`,:LAQ�TL[��ۺ �$��X��6��� �� S��      |",��(�nH�{G�/��Kkλ�R��g_e�3�������[�.�Z:���:X�;��;��-;�9;�A;�bE;D�G;��H;tFI;`I;�TI;bAI;�0I;#I;�I;I;�I;I;��H;b�H;��H;!�H;,�H;��H;,�H;!�H;��H;b�H;��H;I;�I;I;�I;#I;�0I;bAI;�TI;`I;tFI;��H;D�G;�bE;�A;�9;��-;��;X�;���:.�Z:��[����3��g_e��R��Kkλ/��{G�nH��(�      �d��Z���Ǩ���)���zl�<RH�l"��.��X��:�k�]� �����9���:���:6�;�-;�9;j`A;۹E;J�G;��H;#RI;4_I;OI;�;I;�+I;�I;MI;)I;�I;p I;��H;��H;��H;��H;|�H;��H;��H;��H;��H;p I;�I;)I;MI;�I;�+I;�;I;OI;4_I;#RI;��H;J�G;۹E;j`A;�9;�-;6�;���:���:��9��]� �:�k�X���.��l"�<RH��zl��)��Ǩ��Z���      ���s9�o5��P��ib̼�֮����� d�>",����PR��H5� %�� �f9�ޚ:��:6�;��-;��:;KB;_UF;:JH; I;�[I;G[I;�GI;%5I;<&I;7I;�I;9	I;^I;�H;��H;��H;n�H;�H;n�H;��H;��H;�H;^I;9	I;�I;7I;<&I;%5I;�GI;G[I;�[I; I;:JH;_UF;KB;��:;��-;6�;��:�ޚ: �f9 %��H5�PR�����>",�� d�����֮�ib̼P��o5��s9�      �]��IY��ZN��`=���'�v�Ý���������C�W��$����C�X������9�ޚ:���:��;˷0;�<;v�C;GG;�H;�>I;P`I;�SI;^?I;1.I;z I;�I;.I;�I;�I;��H;��H;&�H;��H;&�H;��H;��H;�I;�I;.I;�I;z I;1.I;^?I;�SI;P`I;�>I;�H;GG;v�C;�<;˷0;��;���:�ޚ:�9����C�X�����$�C�W���������Ý�v���'��`=��ZN��IY�      �A��!��e���*��齅�C�d��`=����r��z֮�~�y���(�v�һj^e����� �f9���:X�;m0";A�4;�l?;E;��G;��H;�VI;�]I;(JI;�6I;'I;�I;FI;�	I;>I;7 I;��H;��H;V�H;��H;��H;7 I;>I;�	I;FI;�I;'I;�6I;(JI;�]I;�VI;��H;��G;E;�l?;A�4;m0";X�;���: �f9����j^e�v�һ��(�~�y�z֮�r�꼠���`=�C�d�齅��*��e��!��      ���FE	��������Wн�A����!�h���3����6¼�)��ax/�v�һC�X� %����9���:�=;[e);�_9;�%B;ډF;�|H;�5I;u`I;�TI;�?I;�-I; I;jI;DI;�I;jI;q�H;��H;�H;��H;q�H;jI;�I;DI;jI; I;�-I;�?I;�TI;u`I;�5I;�|H;ډF;�%B;�_9;[e);�=;���:��9 %��C�X�v�һax/��)��6¼�����3�!�h��󑽢A���Wн��콹��FE	�      y^Z�[
V��I�
�6�������ܽ!��ܽ���aG�c��ȼ�)����(����H5���.�Z:k�:7R;/&1;��=;ПD;P�G;�H;�WI;9]I;�HI;5I;�%I;�I;�I;�	I;�I;mI;|�H;��H;|�H;mI;�I;�	I;�I;�I;�%I;5I;�HI;9]I;�WI;�H;P�G;ПD;��=;/&1;7R;k�:.�Z:��H5������(��)���ȼc��aG�ܽ��!���ܽ�����
�6��I�[
V�      � ���e�����ؕ����q�	�I���"���������k���ZN�c�6¼~�y��$�PR��]� ���[��:G/;J�&;
w8;��A;��F;��H;?I;aI;�QI;:<I;7+I;�I;I;uI;�I;WI;9I;� I;9I;WI;�I;uI;I;�I;7+I;:<I;�QI;aI;?I;��H;��F;��A;
w8;J�&;G/;�:��[�]� �PR���$�~�y�6¼c��ZN�k������������"�	�I���q�ؕ������e��      a5�������Q�Ҿ�a��w����l��6�BE	���Ƚk���aG����z֮�C�W����:�k����U`,:���:�;��1;m�>;^E;L�G;BI;G^I;hYI;ZCI;�0I;V"I;cI;I;#	I;,I;�I;=I;�I;,I;#	I;I;cI;V"I;�0I;ZCI;hYI;G^I;BI;L�G;^E;m�>;��1;�;���:U`,:���:�k����C�W�z֮�����aG�k����ȽBE	��6��l�w����a��Q�Ҿ������      uA��q<�aa/����:�u]׾� ��w��>�BE	�����ܽ����3�r�꼰���>",�X��3��LAQ�خ�:�L
;�e);ބ:;D?C;?G;|�H;fSI;�^I;KJI;6I;t&I;�I;�I;ZI;�I;�I;�I;�I;�I;ZI;�I;�I;t&I;6I;KJI;�^I;fSI;|�H;?G;D?C;ބ:;�e);�L
;خ�:LAQ�3��X��>",�����r�꼠�3�ܽ������BE	�>�w��� ��u]׾�:���aa/��q<�      q�������Y�{�e$_��q<�������}��w���6�����!��!�h��������� d��.��g_e�TL[���Z:���:�+ ;��5;�A;�UF;˃H;@I;�aI;�PI;;I;e*I;�I;+I;WI;�I;I;LI;I;�I;WI;+I;�I;e*I;;I;�PI;�aI;@I;˃H;�UF;�A;��5;�+ ;���:��Z:TL[�g_e��.��� d��������!�h�!�������6�w���}��������q<�e$_�Y�{�����      6��������欿��������O�}x����� ���l���"��ܽ���`=�Ý��l"��R���ۺO��9�=�:�K;��0;͞>;�LE;|"H;�$I;�`I;(VI;�?I;.I;` I;[I;"I;/
I;lI;�I;lI;/
I;"I;[I;` I;.I;�?I;(VI;�`I;�$I;|"H;�LE;͞>;��0;�K;�=�:O��9�ۺ�R��l"����Ý��`=����ܽ��"��l�� �����}x���O��������欿����      �������F��dȿf���������O���u]׾w���	�I�����A��C�d�v��֮�<RH�Kkλ �$�s5����:mM;˅+;�<;"3D;�G;�I;�]I;�ZI;	DI;H1I;�"I;`I;�I;�I;�I;�I;�I;�I;�I;`I;�"I;H1I;	DI;�ZI;�]I;�I;�G;"3D;�<;˅+;mM;���:s5� �$�Kkλ<RH��֮�v�C�d��A�����	�I�w���u]׾����O�����f���dȿF�ῢ��      @�-i�������B�ѿf�������q<��:��a����q����Wн齅���'�ib̼�zl�/���X�z�� �:��;
�&;٪9;KC;wLG;�H;]XI;�]I;�GI;4I;�$I;I;'I;�I;�	I;�I;�	I;�I;'I;I;�$I;4I;�GI;�]I;]XI;�H;wLG;KC;٪9;
�&;��; �:z���X�/���zl�ib̼��'�齅��Wн����q��a���:��q<����f���B�ѿ������-i�      A:�.5�(�'��������dȿ���e$_���Q�Ҿؕ��
�6�����*���`=�P���)��{G��6��B����Q:�:/";�7;�%B;�F;��H;RI;�_I;�JI;C6I;�&I;ZI;7I;�I;�
I;�	I;�
I;�I;7I;ZI;�&I;C6I;�JI;�_I;RI;��H;�F;�%B;�7;/";�:��Q:B���6��{G��)��P���`=��*�����
�6�ؕ��Q�Ҿ��e$_����dȿ�������(�'�.5�      ��U�T�O�B-?�(�'���F�`欿Y�{�aa/���뾙���I����e���ZN�o5��Ǩ��nH�� ������ݧ":��:��;��5;�_A;ٚF;Z�H;<LI;aI;�LI;�7I;(I;aI;I;_I;&I;&
I;&I;_I;I;aI;(I;�7I;�LI;aI;<LI;Z�H;ٚF;�_A;��5;��;��:ݧ":����� ��nH�Ǩ��o5���ZN�e������I�������aa/�Y�{��欿F����(�'�B-?�T�O�      ��i���b�T�O�.5�-i������������q<�����e��[
V�FE	�!���IY�s9�Z����(� S����Ⱥ��:���:'�;L�4;h�@;kgF;��H;4HI;�aI;�MI;�8I;�(I;I;~I;�I;{I;x
I;{I;�I;~I;I;�(I;�8I;�MI;�aI;4HI;��H;kgF;h�@;L�4;'�;���:��:��Ⱥ S���(�Z���s9��IY�!��FE	�[
V��e������q<������������-i�.5�T�O���b�      ݶ��O���ά��(�_���7�w�}߿���~,b��V�*l¾Fx�c.���Ž��t�6�����*�?��N�����sx9���:��;��2;T?@;�eF;C�H;��I;��I;9{I;�ZI;�BI;#1I;�$I;�I;�I;NI;�I;�I;�$I;#1I;�BI;�ZI;9{I;��I;��I;C�H;�eF;T?@;��2;��;���:�sx9���N��*�?����6����t���Žc.�Fx�*l¾�V�~,b����}߿w���7�(�_�ά��O���      O���A���}��+Y��3�����$ڿ"����\����(���s��3�9�����p�p�p���<<����e������9{��:�;V$3;ho@;yF;��H;�I;�I;�zI;sZI;yBI;�0I;t$I;EI;tI; I;tI;EI;t$I;�0I;yBI;sZI;�zI;�I;�I;��H;yF;ho@;V$3;�;{��:���9e�������<<�p��p���p�9����3��s�(�������\�"���$ڿ����3��+Y�}�A���      ά��}�8tf��lG�Ң%��p�*�ʿV����>M����S����d�ɤ�̷�9�d��
��I��@�1���������9���:N;�T4;��@;�F;@�H;�I;ܙI;�xI;�XI;bAI;�/I;�#I;�I;�I;�I;�I;�I;�#I;�/I;bAI;�XI;�xI;ܙI;�I;@�H;�F;��@;�T4;N;���:��9������@�1��I���
�9�d�̷�ɤ��d�S�������>M�V���*�ʿ�p�Ң%��lG�8tf�}�      (�_��+Y��lG�f.�w���꿭���J䂿��5���󾋰��M�N�W��V��-�Q�*�������;i!��g��,󳺏:��:�;e06;��A;tG;I;Z�I;��I;�uI;qVI;�?I;�.I;�"I;�I;'I;�I;'I;�I;�"I;�.I;�?I;qVI;�uI;��I;Z�I;I;tG;��A;e06;�;��:�:,��g��;i!�����*���-�Q�V��W��M�N���������5�J䂿�������w�f.��lG��+Y�      ��7��3�Ң%�w��<����ſ�����\�9����Ͼ����`�3����z����9�z�ἷ���z��8}�ht�H�^:�)�:΢#;��8;��B;ArG;�$I;јI;�I;$qI;6SI;=I;�,I;0!I;nI;I;�I;I;nI;0!I;�,I;=I;6SI;$qI;�I;јI;�$I;ArG;��B;��8;΢#;�)�:H�^:ht��8}��z����z�Ἁ�9��z����`�3�������Ͼ9����\������ſ�<��w�Ң%��3�      w�����p������ſ!��{Ps���1�-r���d���d�}I�҈Ž��}�l*�fC��W�^�RC�f�D�(N๪��:��;�);.6;;KD;e�G;kGI;ΜI;ȎI;�kI;OI;�9I;3*I;8I;�I;�I;KI;�I;�I;8I;3*I;�9I;OI;�kI;ȎI;ΜI;kGI;e�G;KD;.6;;�);��;���:(N�f�D�RC�W�^�fC��l*���}�҈Ž}I��d��d��-r����1�{Ps�!����ſ��꿀p����      }߿�$ڿ*�ʿ�������{Ps�MX:����#l¾�ǆ���7����<5��$�Q�����t��85�������"��8 ȼ:��;��.;��=;�DE;�XH;�gI;G�I;ڇI;GeI;@JI;E6I;a'I;�I;I;�I;�I;�I;I;�I;a'I;E6I;@JI;GeI;ڇI;G�I;�gI;�XH;�DE;��=;��.;��; ȼ:"��8������85��t�����$�Q�<5�������7��ǆ�#l¾���MX:�{Ps��������*�ʿ�$ڿ      ���"��V���J䂿��\���1�����J˾睒�C�N�y��L������c�'���Ҽ �|��z�ko��z��'�&:�N�:˧;�V4;�@;HfF;��H;.�I;A�I;UI;=^I;�DI;&2I;<$I;bI;�I;I;�I;I;�I;bI;<$I;&2I;�DI;=^I;UI;A�I;.�I;��H;HfF;�@;�V4;˧;�N�:'�&:z��ko���z� �|���Ҽc�'����L���y��C�N�睒��J˾�����1���\�J䂿V���"��      ~,b���\��>M���5�9��-r��#l¾睒�"&W��3�<Sؽ�z��fG�����I���?��̻{�-����K��:��;Ͽ&;B{9;�C;�cG;sI;]�I;r�I;ruI;�VI;O?I;�-I;� I;�I;yI;�I;�I;�I;yI;�I;� I;�-I;O?I;�VI;ruI;r�I;]�I;sI;�cG;�C;B{9;Ͽ&;��;K��:���{�-��̻�?��I�����fG��z��<Sؽ�3�"&W�睒�#l¾-r��9����5��>M���\�      �V������������Ͼ�d���ǆ�C�N��3��c�[����\�@��EC��N�o�Ъ	�t숻0�L��9J��:�g;o�/;\�=;bE;2H;�VI;؜I;�I;�jI;�NI;G9I;)I;=I;�I;I;�I;�
I;�I;I;�I;=I;)I;G9I;�NI;�jI;�I;؜I;�VI;2H;bE;\�=;o�/;�g;J��:L��90�t숻Ъ	�N�o�EC��@����\�[���cཱ3�C�N��ǆ��d����Ͼ���������      *l¾(��S������������d���7�y��<Sؽ[�� �d�P*�kּI\����'�����S������
�:�Y;�#;Y<7;M�A;2�F;{�H;��I;	�I;րI;	`I;�FI;3I;B$I;�I;�I;vI;i	I;iI;i	I;vI;�I;�I;B$I;3I;�FI;	`I;րI;	�I;��I;{�H;2�F;M�A;Y<7;�#;�Y;�
�:�����S������'�I\��kּP*� �d�[��<Sؽy����7��d���������S���(��      Fx��s��d�M�N�`�3�}I����L����z����\�P*�'�ݼe���j<<���ڻ��V��gt�r�&:���:[B;�;/;nC=;��D;��G;8I;�I;ÓI;3sI;IUI;}>I;�,I;�I;�I;xI;�	I;I;.I;I;�	I;xI;�I;�I;�,I;}>I;IUI;3sI;ÓI;�I;8I;��G;��D;nC=;�;/;[B;���:r�&:�gt���V���ڻj<<�e���'�ݼP*���\��z��L������}I�`�3�M�N��d��s�      c.��3�ɤ�W����҈Ž<5�����fG�@��kּe���:yC�?�W7}�𮼺K�x9���:&	;O�&;�:8;��A;F;ϸH;WxI;��I;�I;PeI;�JI;m6I;�&I;�I;�I;uI;/I;�I;�I;�I;/I;uI;�I;�I;�&I;m6I;�JI;PeI;�I;��I;WxI;ϸH;F;��A;�:8;O�&;&	;���:K�x9𮼺W7}�?�:yC�e���kּ@��fG����<5��҈Ž��W��ɤ��3�      ��Ž9���̷�V���z����}�$�Q�c�'����EC��I\��j<<�?��n����YU�b��:Z��:,�;�&3;��>;�E;�H;};I;�I;ÔI;�uI;�WI;�@I;�.I;� I;�I;I;oI;�I;<I;�I;<I;�I;oI;I;�I;� I;�.I;�@I;�WI;�uI;ÔI;�I;};I;�H;�E;��>;�&3;,�;Z��:b��:YU����n��?�j<<�I\��EC�����c�'�$�Q���}��z��V��̷�9���      ��t���p�9�d�-�Q���9�l*������Ҽ�I��N�o���'���ڻW7}���pH��߄:�k�:��;�.;5<;�nC;^6G;��H;�I;��I;�I;;eI;^KI;7I;�&I;�I;�I;h
I;cI;�I;��H;l�H;��H;�I;cI;h
I;�I;�I;�&I;7I;^KI;;eI;�I;��I;�I;��H;^6G;�nC;5<;�.;��;�k�:�߄:pH���W7}���ڻ��'�N�o��I����Ҽ���l*���9�-�Q�9�d���p�      6��p��
�*���z��fC���t�� �|��?�Ъ	������V�𮼺YU��߄:��:�g;6�+;�9;��A;�eF;w�H;�^I;��I;��I; rI;�UI;�?I;�-I; I;uI;(I;�I;�I;i�H;��H;�H;��H;i�H;�I;�I;(I;uI; I;�-I;�?I;�UI; rI;��I;��I;�^I;w�H;�eF;��A;�9;6�+;�g;��:�߄:YU�𮼺��V����Ъ	��?� �|��t��fC��z��*����
�p�      ���p���I���������W�^�85��z��̻t숻�S��gt�K�x9b��:�k�:�g;y�*;�8;�@; �E;W'H;�7I;ߒI;2�I;o}I;�_I;�GI;�4I;y%I;�I;RI;	I;�I;��H;�H;i�H;��H;i�H;�H;��H;�I;	I;RI;�I;y%I;�4I;�GI;�_I;o}I;2�I;ߒI;�7I;W'H; �E;�@;�8;y�*;�g;�k�:b��:K�x9�gt��S�t숻�̻�z�85�W�^���������I��p��      *�?��<<�@�1�;i!��z�RC����ko��{�-�0򳺱���r�&:���:Z��:��;6�+;�8;W�@;]E;��G;eI;	�I;l�I;P�I;�hI;UOI;";I;�*I;�I;�I;nI;EI;� I;��H;��H;d�H;��H;d�H;��H;��H;� I;EI;nI;�I;�I;�*I;";I;UOI;�hI;P�I;l�I;	�I;eI;��G;]E;W�@;�8;6�+;��;Z��:���:r�&:����0�{�-�ko�����RC��z�;i!�@�1��<<�      �N����������g���8}�f�D����z�����L��9�
�:���:&	;,�;�.;�9;�@;]E;��G;]I;�~I;#�I;g�I;�oI;�UI;�@I;�/I;�!I;�I;I;I;�I;��H;s�H;��H;r�H;��H;r�H;��H;s�H;��H;�I;I;I;�I;�!I;�/I;�@I;�UI;�oI;g�I;#�I;�~I;]I;��G;]E;�@;�9;�.;,�;&	;���:�
�:L��9���z�����f�D��8}��g���������      ��e�����,�ht�(N�"��8'�&:K��:J��:�Y;[B;O�&;�&3;5<;��A; �E;��G;]I;w{I;��I;��I;�tI;�ZI;*EI;�3I;E%I;�I;bI;�I;I;O�H;��H;I�H;��H;��H;1�H;��H;��H;I�H;��H;O�H;I;�I;bI;�I;E%I;�3I;*EI;�ZI;�tI;��I;��I;w{I;]I;��G; �E;��A;5<;�&3;O�&;[B;�Y;J��:K��:'�&:"��8(N�ht�,���e���      �sx9���9��9�:H�^:���: ȼ:�N�:��;�g;�#;�;/;�:8;��>;�nC;�eF;W'H;eI;�~I;��I;ːI;wI;�]I;QHI;�6I;(I;#I;�I;�
I;\I;b�H;]�H;h�H;L�H;��H;��H;��H;��H;��H;L�H;h�H;]�H;b�H;\I;�
I;�I;#I;(I;�6I;QHI;�]I;wI;ːI;��I;�~I;eI;W'H;�eF;�nC;��>;�:8;�;/;�#;�g;��;�N�: ȼ:���:H�^:�:��9���9      ���:{��:���:��:�)�:��;��;˧;Ͽ&;o�/;Y<7;nC=;��A;�E;^6G;w�H;�7I;	�I;#�I;��I;wI;�^I;�II;�8I;*I;I;LI;QI;�I;L I;�H;��H;*�H;M�H;��H;�H;��H;�H;��H;M�H;*�H;��H;�H;L I;�I;QI;LI;I;*I;�8I;�II;�^I;wI;��I;#�I;	�I;�7I;w�H;^6G;�E;��A;nC=;Y<7;o�/;Ͽ&;˧;��;��;�)�:��:���:{��:      ��;�;N;�;΢#;�);��.;�V4;B{9;\�=;M�A;��D;F;�H;��H;�^I;ߒI;l�I;g�I;�tI;�]I;�II;=9I;6+I;VI;�I;gI;�I;4I;��H;�H;F�H;�H;{�H;p�H;��H;b�H;��H;p�H;{�H;�H;F�H;�H;��H;4I;�I;gI;�I;VI;6+I;=9I;�II;�]I;�tI;g�I;l�I;ߒI;�^I;��H;�H;F;��D;M�A;\�=;B{9;�V4;��.;�);΢#;�;N;�;      ��2;V$3;�T4;e06;��8;.6;;��=;�@;�C;bE;2�F;��G;ϸH;};I;�I;��I;2�I;P�I;�oI;�ZI;QHI;�8I;6+I;�I;5I;2I;iI;�I;Y�H;t�H;q�H;:�H;L�H;��H;��H;i�H;�H;i�H;��H;��H;L�H;:�H;q�H;t�H;Y�H;�I;iI;2I;5I;�I;6+I;�8I;QHI;�ZI;�oI;P�I;2�I;��I;�I;};I;ϸH;��G;2�F;bE;�C;�@;��=;.6;;��8;e06;�T4;V$3;      T?@;ho@;��@;��A;��B;KD;�DE;HfF;�cG;2H;{�H;8I;WxI;�I;��I;��I;o}I;�hI;�UI;*EI;�6I;*I;VI;5I;tI;�I;QI;��H;��H;��H;.�H;0�H;��H;}�H;��H;,�H;	�H;,�H;��H;}�H;��H;0�H;.�H;��H;��H;��H;QI;�I;tI;5I;VI;*I;�6I;*EI;�UI;�hI;o}I;��I;��I;�I;WxI;8I;{�H;2H;�cG;HfF;�DE;KD;��B;��A;��@;ho@;      �eF;yF;�F;tG;ArG;e�G;�XH;��H;sI;�VI;��I;�I;��I;ÔI;�I; rI;�_I;UOI;�@I;�3I;(I;I;�I;2I;�I;jI;��H;�H;��H;b�H;?�H;q�H;#�H;9�H;|�H;�H;�H;�H;|�H;9�H;#�H;q�H;?�H;b�H;��H;�H;��H;jI;�I;2I;�I;I;(I;�3I;�@I;UOI;�_I; rI;�I;ÔI;��I;�I;��I;�VI;sI;��H;�XH;e�G;ArG;tG;�F;yF;      C�H;��H;@�H;I;�$I;kGI;�gI;.�I;]�I;؜I;	�I;ÓI;�I;�uI;;eI;�UI;�GI;";I;�/I;E%I;#I;LI;gI;iI;QI;��H;�H;��H;s�H;@�H;{�H; �H;��H;�H;q�H;�H;�H;�H;q�H;�H;��H; �H;{�H;@�H;s�H;��H;�H;��H;QI;iI;gI;LI;#I;E%I;�/I;";I;�GI;�UI;;eI;�uI;�I;ÓI;	�I;؜I;]�I;.�I;�gI;kGI;�$I;I;@�H;��H;      ��I;�I;�I;Z�I;јI;ΜI;G�I;A�I;r�I;�I;րI;3sI;PeI;�WI;^KI;�?I;�4I;�*I;�!I;�I;�I;QI;�I;�I;��H;�H;��H;k�H;Q�H;j�H;��H;��H;��H;�H;��H;H�H;1�H;H�H;��H;�H;��H;��H;��H;j�H;Q�H;k�H;��H;�H;��H;�I;�I;QI;�I;�I;�!I;�*I;�4I;�?I;^KI;�WI;PeI;3sI;րI;�I;r�I;A�I;G�I;ΜI;јI;Z�I;�I;�I;      ��I;�I;ܙI;��I;�I;ȎI;ڇI;UI;ruI;�jI;	`I;IUI;�JI;�@I;7I;�-I;y%I;�I;�I;bI;�
I;�I;4I;Y�H;��H;��H;s�H;Q�H;j�H;��H;��H;��H;��H;-�H;��H;��H;Y�H;��H;��H;-�H;��H;��H;��H;��H;j�H;Q�H;s�H;��H;��H;Y�H;4I;�I;�
I;bI;�I;�I;y%I;�-I;7I;�@I;�JI;IUI;	`I;�jI;ruI;UI;ڇI;ȎI;�I;��I;ܙI;�I;      9{I;�zI;�xI;�uI;$qI;�kI;GeI;=^I;�VI;�NI;�FI;}>I;m6I;�.I;�&I; I;�I;�I;I;�I;\I;L I;��H;t�H;��H;b�H;@�H;j�H;��H;��H;��H;��H;�H;��H;�H;��H;��H;��H;�H;��H;�H;��H;��H;��H;��H;j�H;@�H;b�H;��H;t�H;��H;L I;\I;�I;I;�I;�I; I;�&I;�.I;m6I;}>I;�FI;�NI;�VI;=^I;GeI;�kI;$qI;�uI;�xI;�zI;      �ZI;sZI;�XI;qVI;6SI;OI;@JI;�DI;O?I;G9I;3I;�,I;�&I;� I;�I;uI;RI;nI;I;I;b�H;�H;�H;q�H;.�H;?�H;{�H;��H;��H;��H;��H;��H;_�H;��H;|�H;c�H;Z�H;c�H;|�H;��H;_�H;��H;��H;��H;��H;��H;{�H;?�H;.�H;q�H;�H;�H;b�H;I;I;nI;RI;uI;�I;� I;�&I;�,I;3I;G9I;O?I;�DI;@JI;OI;6SI;qVI;�XI;sZI;      �BI;yBI;bAI;�?I;=I;�9I;E6I;&2I;�-I;)I;B$I;�I;�I;�I;�I;(I;	I;EI;�I;O�H;]�H;��H;F�H;:�H;0�H;q�H; �H;��H;��H;��H;��H;I�H;��H;U�H;�H;��H;��H;��H;�H;U�H;��H;I�H;��H;��H;��H;��H; �H;q�H;0�H;:�H;F�H;��H;]�H;O�H;�I;EI;	I;(I;�I;�I;�I;�I;B$I;)I;�-I;&2I;E6I;�9I;=I;�?I;bAI;yBI;      #1I;�0I;�/I;�.I;�,I;3*I;a'I;<$I;� I;=I;�I;�I;�I;I;h
I;�I;�I;� I;��H;��H;h�H;*�H;�H;L�H;��H;#�H;��H;��H;��H;�H;_�H;��H;9�H;��H;��H;��H;t�H;��H;��H;��H;9�H;��H;_�H;�H;��H;��H;��H;#�H;��H;L�H;�H;*�H;h�H;��H;��H;� I;�I;�I;h
I;I;�I;�I;�I;=I;� I;<$I;a'I;3*I;�,I;�.I;�/I;�0I;      �$I;t$I;�#I;�"I;0!I;8I;�I;bI;�I;�I;�I;xI;uI;oI;cI;�I;��H;��H;s�H;I�H;L�H;M�H;{�H;��H;}�H;9�H;�H;�H;-�H;��H;��H;U�H;��H;��H;b�H;@�H;)�H;@�H;b�H;��H;��H;U�H;��H;��H;-�H;�H;�H;9�H;}�H;��H;{�H;M�H;L�H;I�H;s�H;��H;��H;�I;cI;oI;uI;xI;�I;�I;�I;bI;�I;8I;0!I;�"I;�#I;t$I;      �I;EI;�I;�I;nI;�I;I;�I;yI;I;vI;�	I;/I;�I;�I;i�H;�H;��H;��H;��H;��H;��H;p�H;��H;��H;|�H;q�H;��H;��H;�H;|�H;�H;��H;b�H;�H;�H;�H;�H;�H;b�H;��H;�H;|�H;�H;��H;��H;q�H;|�H;��H;��H;p�H;��H;��H;��H;��H;��H;�H;i�H;�I;�I;/I;�	I;vI;I;yI;�I;I;�I;nI;�I;�I;EI;      �I;tI;�I;'I;I;�I;�I;I;�I;�I;i	I;I;�I;<I;��H;��H;i�H;d�H;r�H;��H;��H;�H;��H;i�H;,�H;�H;�H;H�H;��H;��H;c�H;��H;��H;@�H;�H;��H;��H;��H;�H;@�H;��H;��H;c�H;��H;��H;H�H;�H;�H;,�H;i�H;��H;�H;��H;��H;r�H;d�H;i�H;��H;��H;<I;�I;I;i	I;�I;�I;I;�I;�I;I;'I;�I;tI;      NI; I;�I;�I;�I;KI;�I;�I;�I;�
I;iI;.I;�I;�I;l�H;�H;��H;��H;��H;1�H;��H;��H;b�H;�H;	�H;�H;�H;1�H;Y�H;��H;Z�H;��H;t�H;)�H;�H;��H;��H;��H;�H;)�H;t�H;��H;Z�H;��H;Y�H;1�H;�H;�H;	�H;�H;b�H;��H;��H;1�H;��H;��H;��H;�H;l�H;�I;�I;.I;iI;�
I;�I;�I;�I;KI;�I;�I;�I; I;      �I;tI;�I;'I;I;�I;�I;I;�I;�I;i	I;I;�I;<I;��H;��H;i�H;d�H;r�H;��H;��H;�H;��H;i�H;,�H;�H;�H;H�H;��H;��H;c�H;��H;��H;@�H;�H;��H;��H;��H;�H;@�H;��H;��H;c�H;��H;��H;H�H;�H;�H;,�H;i�H;��H;�H;��H;��H;r�H;d�H;i�H;��H;��H;<I;�I;I;i	I;�I;�I;I;�I;�I;I;'I;�I;tI;      �I;EI;�I;�I;nI;�I;I;�I;yI;I;vI;�	I;/I;�I;�I;i�H;�H;��H;��H;��H;��H;��H;p�H;��H;��H;|�H;q�H;��H;��H;�H;|�H;�H;��H;b�H;�H;�H;�H;�H;�H;b�H;��H;�H;|�H;�H;��H;��H;q�H;|�H;��H;��H;p�H;��H;��H;��H;��H;��H;�H;i�H;�I;�I;/I;�	I;vI;I;yI;�I;I;�I;nI;�I;�I;EI;      �$I;t$I;�#I;�"I;0!I;8I;�I;bI;�I;�I;�I;xI;uI;oI;cI;�I;��H;��H;s�H;I�H;L�H;M�H;{�H;��H;}�H;9�H;�H;�H;-�H;��H;��H;U�H;��H;��H;b�H;@�H;)�H;@�H;b�H;��H;��H;U�H;��H;��H;-�H;�H;�H;9�H;}�H;��H;{�H;M�H;L�H;I�H;s�H;��H;��H;�I;cI;oI;uI;xI;�I;�I;�I;bI;�I;8I;0!I;�"I;�#I;t$I;      #1I;�0I;�/I;�.I;�,I;3*I;a'I;<$I;� I;=I;�I;�I;�I;I;h
I;�I;�I;� I;��H;��H;h�H;*�H;�H;L�H;��H;#�H;��H;��H;��H;�H;_�H;��H;9�H;��H;��H;��H;t�H;��H;��H;��H;9�H;��H;_�H;�H;��H;��H;��H;#�H;��H;L�H;�H;*�H;h�H;��H;��H;� I;�I;�I;h
I;I;�I;�I;�I;=I;� I;<$I;a'I;3*I;�,I;�.I;�/I;�0I;      �BI;yBI;bAI;�?I;=I;�9I;E6I;&2I;�-I;)I;B$I;�I;�I;�I;�I;(I;	I;EI;�I;O�H;]�H;��H;F�H;:�H;0�H;q�H; �H;��H;��H;��H;��H;I�H;��H;U�H;�H;��H;��H;��H;�H;U�H;��H;I�H;��H;��H;��H;��H; �H;q�H;0�H;:�H;F�H;��H;]�H;O�H;�I;EI;	I;(I;�I;�I;�I;�I;B$I;)I;�-I;&2I;E6I;�9I;=I;�?I;bAI;yBI;      �ZI;sZI;�XI;qVI;6SI;OI;@JI;�DI;O?I;G9I;3I;�,I;�&I;� I;�I;uI;RI;nI;I;I;b�H;�H;�H;q�H;.�H;?�H;{�H;��H;��H;��H;��H;��H;_�H;��H;|�H;c�H;Z�H;c�H;|�H;��H;_�H;��H;��H;��H;��H;��H;{�H;?�H;.�H;q�H;�H;�H;b�H;I;I;nI;RI;uI;�I;� I;�&I;�,I;3I;G9I;O?I;�DI;@JI;OI;6SI;qVI;�XI;sZI;      9{I;�zI;�xI;�uI;$qI;�kI;GeI;=^I;�VI;�NI;�FI;}>I;m6I;�.I;�&I; I;�I;�I;I;�I;\I;L I;��H;t�H;��H;b�H;@�H;j�H;��H;��H;��H;��H;�H;��H;�H;��H;��H;��H;�H;��H;�H;��H;��H;��H;��H;j�H;@�H;b�H;��H;t�H;��H;L I;\I;�I;I;�I;�I; I;�&I;�.I;m6I;}>I;�FI;�NI;�VI;=^I;GeI;�kI;$qI;�uI;�xI;�zI;      ��I;�I;ܙI;��I;�I;ȎI;ڇI;UI;ruI;�jI;	`I;IUI;�JI;�@I;7I;�-I;y%I;�I;�I;bI;�
I;�I;4I;Y�H;��H;��H;s�H;Q�H;j�H;��H;��H;��H;��H;-�H;��H;��H;Y�H;��H;��H;-�H;��H;��H;��H;��H;j�H;Q�H;s�H;��H;��H;Y�H;4I;�I;�
I;bI;�I;�I;y%I;�-I;7I;�@I;�JI;IUI;	`I;�jI;ruI;UI;ڇI;ȎI;�I;��I;ܙI;�I;      ��I;�I;�I;Z�I;јI;ΜI;G�I;A�I;r�I;�I;րI;3sI;PeI;�WI;^KI;�?I;�4I;�*I;�!I;�I;�I;QI;�I;�I;��H;�H;��H;k�H;Q�H;j�H;��H;��H;��H;�H;��H;H�H;1�H;H�H;��H;�H;��H;��H;��H;j�H;Q�H;k�H;��H;�H;��H;�I;�I;QI;�I;�I;�!I;�*I;�4I;�?I;^KI;�WI;PeI;3sI;րI;�I;r�I;A�I;G�I;ΜI;јI;Z�I;�I;�I;      C�H;��H;@�H;I;�$I;kGI;�gI;.�I;]�I;؜I;	�I;ÓI;�I;�uI;;eI;�UI;�GI;";I;�/I;E%I;#I;LI;gI;iI;QI;��H;�H;��H;s�H;@�H;{�H; �H;��H;�H;q�H;�H;�H;�H;q�H;�H;��H; �H;{�H;@�H;s�H;��H;�H;��H;QI;iI;gI;LI;#I;E%I;�/I;";I;�GI;�UI;;eI;�uI;�I;ÓI;	�I;؜I;]�I;.�I;�gI;kGI;�$I;I;@�H;��H;      �eF;yF;�F;tG;ArG;e�G;�XH;��H;sI;�VI;��I;�I;��I;ÔI;�I; rI;�_I;UOI;�@I;�3I;(I;I;�I;2I;�I;jI;��H;�H;��H;b�H;?�H;q�H;#�H;9�H;|�H;�H;�H;�H;|�H;9�H;#�H;q�H;?�H;b�H;��H;�H;��H;jI;�I;2I;�I;I;(I;�3I;�@I;UOI;�_I; rI;�I;ÔI;��I;�I;��I;�VI;sI;��H;�XH;e�G;ArG;tG;�F;yF;      T?@;ho@;��@;��A;��B;KD;�DE;HfF;�cG;2H;{�H;8I;WxI;�I;��I;��I;o}I;�hI;�UI;*EI;�6I;*I;VI;5I;tI;�I;QI;��H;��H;��H;.�H;0�H;��H;}�H;��H;,�H;	�H;,�H;��H;}�H;��H;0�H;.�H;��H;��H;��H;QI;�I;tI;5I;VI;*I;�6I;*EI;�UI;�hI;o}I;��I;��I;�I;WxI;8I;{�H;2H;�cG;HfF;�DE;KD;��B;��A;��@;ho@;      ��2;V$3;�T4;e06;��8;.6;;��=;�@;�C;bE;2�F;��G;ϸH;};I;�I;��I;2�I;P�I;�oI;�ZI;QHI;�8I;6+I;�I;5I;2I;iI;�I;Y�H;t�H;q�H;:�H;L�H;��H;��H;i�H;�H;i�H;��H;��H;L�H;:�H;q�H;t�H;Y�H;�I;iI;2I;5I;�I;6+I;�8I;QHI;�ZI;�oI;P�I;2�I;��I;�I;};I;ϸH;��G;2�F;bE;�C;�@;��=;.6;;��8;e06;�T4;V$3;      ��;�;N;�;΢#;�);��.;�V4;B{9;\�=;M�A;��D;F;�H;��H;�^I;ߒI;l�I;g�I;�tI;�]I;�II;=9I;6+I;VI;�I;gI;�I;4I;��H;�H;F�H;�H;{�H;p�H;��H;b�H;��H;p�H;{�H;�H;F�H;�H;��H;4I;�I;gI;�I;VI;6+I;=9I;�II;�]I;�tI;g�I;l�I;ߒI;�^I;��H;�H;F;��D;M�A;\�=;B{9;�V4;��.;�);΢#;�;N;�;      ���:{��:���:��:�)�:��;��;˧;Ͽ&;o�/;Y<7;nC=;��A;�E;^6G;w�H;�7I;	�I;#�I;��I;wI;�^I;�II;�8I;*I;I;LI;QI;�I;L I;�H;��H;*�H;M�H;��H;�H;��H;�H;��H;M�H;*�H;��H;�H;L I;�I;QI;LI;I;*I;�8I;�II;�^I;wI;��I;#�I;	�I;�7I;w�H;^6G;�E;��A;nC=;Y<7;o�/;Ͽ&;˧;��;��;�)�:��:���:{��:      �sx9���9��9�:H�^:���: ȼ:�N�:��;�g;�#;�;/;�:8;��>;�nC;�eF;W'H;eI;�~I;��I;ːI;wI;�]I;QHI;�6I;(I;#I;�I;�
I;\I;b�H;]�H;h�H;L�H;��H;��H;��H;��H;��H;L�H;h�H;]�H;b�H;\I;�
I;�I;#I;(I;�6I;QHI;�]I;wI;ːI;��I;�~I;eI;W'H;�eF;�nC;��>;�:8;�;/;�#;�g;��;�N�: ȼ:���:H�^:�:��9���9      ��e�����,�ht�(N�"��8'�&:K��:J��:�Y;[B;O�&;�&3;5<;��A; �E;��G;]I;w{I;��I;��I;�tI;�ZI;*EI;�3I;E%I;�I;bI;�I;I;O�H;��H;I�H;��H;��H;1�H;��H;��H;I�H;��H;O�H;I;�I;bI;�I;E%I;�3I;*EI;�ZI;�tI;��I;��I;w{I;]I;��G; �E;��A;5<;�&3;O�&;[B;�Y;J��:K��:'�&:"��8(N�ht�,���e���      �N����������g���8}�f�D����z�����L��9�
�:���:&	;,�;�.;�9;�@;]E;��G;]I;�~I;#�I;g�I;�oI;�UI;�@I;�/I;�!I;�I;I;I;�I;��H;s�H;��H;r�H;��H;r�H;��H;s�H;��H;�I;I;I;�I;�!I;�/I;�@I;�UI;�oI;g�I;#�I;�~I;]I;��G;]E;�@;�9;�.;,�;&	;���:�
�:L��9���z�����f�D��8}��g���������      *�?��<<�@�1�;i!��z�RC����ko��{�-�0򳺱���r�&:���:Z��:��;6�+;�8;W�@;]E;��G;eI;	�I;l�I;P�I;�hI;UOI;";I;�*I;�I;�I;nI;EI;� I;��H;��H;d�H;��H;d�H;��H;��H;� I;EI;nI;�I;�I;�*I;";I;UOI;�hI;P�I;l�I;	�I;eI;��G;]E;W�@;�8;6�+;��;Z��:���:r�&:����0�{�-�ko�����RC��z�;i!�@�1��<<�      ���p���I���������W�^�85��z��̻t숻�S��gt�K�x9b��:�k�:�g;y�*;�8;�@; �E;W'H;�7I;ߒI;2�I;o}I;�_I;�GI;�4I;y%I;�I;RI;	I;�I;��H;�H;i�H;��H;i�H;�H;��H;�I;	I;RI;�I;y%I;�4I;�GI;�_I;o}I;2�I;ߒI;�7I;W'H; �E;�@;�8;y�*;�g;�k�:b��:K�x9�gt��S�t숻�̻�z�85�W�^���������I��p��      6��p��
�*���z��fC���t�� �|��?�Ъ	������V�𮼺YU��߄:��:�g;6�+;�9;��A;�eF;w�H;�^I;��I;��I; rI;�UI;�?I;�-I; I;uI;(I;�I;�I;i�H;��H;�H;��H;i�H;�I;�I;(I;uI; I;�-I;�?I;�UI; rI;��I;��I;�^I;w�H;�eF;��A;�9;6�+;�g;��:�߄:YU�𮼺��V����Ъ	��?� �|��t��fC��z��*����
�p�      ��t���p�9�d�-�Q���9�l*������Ҽ�I��N�o���'���ڻW7}���pH��߄:�k�:��;�.;5<;�nC;^6G;��H;�I;��I;�I;;eI;^KI;7I;�&I;�I;�I;h
I;cI;�I;��H;l�H;��H;�I;cI;h
I;�I;�I;�&I;7I;^KI;;eI;�I;��I;�I;��H;^6G;�nC;5<;�.;��;�k�:�߄:pH���W7}���ڻ��'�N�o��I����Ҽ���l*���9�-�Q�9�d���p�      ��Ž9���̷�V���z����}�$�Q�c�'����EC��I\��j<<�?��n����YU�b��:Z��:,�;�&3;��>;�E;�H;};I;�I;ÔI;�uI;�WI;�@I;�.I;� I;�I;I;oI;�I;<I;�I;<I;�I;oI;I;�I;� I;�.I;�@I;�WI;�uI;ÔI;�I;};I;�H;�E;��>;�&3;,�;Z��:b��:YU����n��?�j<<�I\��EC�����c�'�$�Q���}��z��V��̷�9���      c.��3�ɤ�W����҈Ž<5�����fG�@��kּe���:yC�?�W7}�𮼺K�x9���:&	;O�&;�:8;��A;F;ϸH;WxI;��I;�I;PeI;�JI;m6I;�&I;�I;�I;uI;/I;�I;�I;�I;/I;uI;�I;�I;�&I;m6I;�JI;PeI;�I;��I;WxI;ϸH;F;��A;�:8;O�&;&	;���:K�x9𮼺W7}�?�:yC�e���kּ@��fG����<5��҈Ž��W��ɤ��3�      Fx��s��d�M�N�`�3�}I����L����z����\�P*�'�ݼe���j<<���ڻ��V��gt�r�&:���:[B;�;/;nC=;��D;��G;8I;�I;ÓI;3sI;IUI;}>I;�,I;�I;�I;xI;�	I;I;.I;I;�	I;xI;�I;�I;�,I;}>I;IUI;3sI;ÓI;�I;8I;��G;��D;nC=;�;/;[B;���:r�&:�gt���V���ڻj<<�e���'�ݼP*���\��z��L������}I�`�3�M�N��d��s�      *l¾(��S������������d���7�y��<Sؽ[�� �d�P*�kּI\����'�����S������
�:�Y;�#;Y<7;M�A;2�F;{�H;��I;	�I;րI;	`I;�FI;3I;B$I;�I;�I;vI;i	I;iI;i	I;vI;�I;�I;B$I;3I;�FI;	`I;րI;	�I;��I;{�H;2�F;M�A;Y<7;�#;�Y;�
�:�����S������'�I\��kּP*� �d�[��<Sؽy����7��d���������S���(��      �V������������Ͼ�d���ǆ�C�N��3��c�[����\�@��EC��N�o�Ъ	�t숻0�L��9J��:�g;o�/;\�=;bE;2H;�VI;؜I;�I;�jI;�NI;G9I;)I;=I;�I;I;�I;�
I;�I;I;�I;=I;)I;G9I;�NI;�jI;�I;؜I;�VI;2H;bE;\�=;o�/;�g;J��:L��90�t숻Ъ	�N�o�EC��@����\�[���cཱ3�C�N��ǆ��d����Ͼ���������      ~,b���\��>M���5�9��-r��#l¾睒�"&W��3�<Sؽ�z��fG�����I���?��̻{�-����K��:��;Ͽ&;B{9;�C;�cG;sI;]�I;r�I;ruI;�VI;O?I;�-I;� I;�I;yI;�I;�I;�I;yI;�I;� I;�-I;O?I;�VI;ruI;r�I;]�I;sI;�cG;�C;B{9;Ͽ&;��;K��:���{�-��̻�?��I�����fG��z��<Sؽ�3�"&W�睒�#l¾-r��9����5��>M���\�      ���"��V���J䂿��\���1�����J˾睒�C�N�y��L������c�'���Ҽ �|��z�ko��z��'�&:�N�:˧;�V4;�@;HfF;��H;.�I;A�I;UI;=^I;�DI;&2I;<$I;bI;�I;I;�I;I;�I;bI;<$I;&2I;�DI;=^I;UI;A�I;.�I;��H;HfF;�@;�V4;˧;�N�:'�&:z��ko���z� �|���Ҽc�'����L���y��C�N�睒��J˾�����1���\�J䂿V���"��      }߿�$ڿ*�ʿ�������{Ps�MX:����#l¾�ǆ���7����<5��$�Q�����t��85�������"��8 ȼ:��;��.;��=;�DE;�XH;�gI;G�I;ڇI;GeI;@JI;E6I;a'I;�I;I;�I;�I;�I;I;�I;a'I;E6I;@JI;GeI;ڇI;G�I;�gI;�XH;�DE;��=;��.;��; ȼ:"��8������85��t�����$�Q�<5�������7��ǆ�#l¾���MX:�{Ps��������*�ʿ�$ڿ      w�����p������ſ!��{Ps���1�-r���d���d�}I�҈Ž��}�l*�fC��W�^�RC�f�D�(N๪��:��;�);.6;;KD;e�G;kGI;ΜI;ȎI;�kI;OI;�9I;3*I;8I;�I;�I;KI;�I;�I;8I;3*I;�9I;OI;�kI;ȎI;ΜI;kGI;e�G;KD;.6;;�);��;���:(N�f�D�RC�W�^�fC��l*���}�҈Ž}I��d��d��-r����1�{Ps�!����ſ��꿀p����      ��7��3�Ң%�w��<����ſ�����\�9����Ͼ����`�3����z����9�z�ἷ���z��8}�ht�H�^:�)�:΢#;��8;��B;ArG;�$I;јI;�I;$qI;6SI;=I;�,I;0!I;nI;I;�I;I;nI;0!I;�,I;=I;6SI;$qI;�I;јI;�$I;ArG;��B;��8;΢#;�)�:H�^:ht��8}��z����z�Ἁ�9��z����`�3�������Ͼ9����\������ſ�<��w�Ң%��3�      (�_��+Y��lG�f.�w���꿭���J䂿��5���󾋰��M�N�W��V��-�Q�*�������;i!��g��,󳺏:��:�;e06;��A;tG;I;Z�I;��I;�uI;qVI;�?I;�.I;�"I;�I;'I;�I;'I;�I;�"I;�.I;�?I;qVI;�uI;��I;Z�I;I;tG;��A;e06;�;��:�:,��g��;i!�����*���-�Q�V��W��M�N���������5�J䂿�������w�f.��lG��+Y�      ά��}�8tf��lG�Ң%��p�*�ʿV����>M����S����d�ɤ�̷�9�d��
��I��@�1���������9���:N;�T4;��@;�F;@�H;�I;ܙI;�xI;�XI;bAI;�/I;�#I;�I;�I;�I;�I;�I;�#I;�/I;bAI;�XI;�xI;ܙI;�I;@�H;�F;��@;�T4;N;���:��9������@�1��I���
�9�d�̷�ɤ��d�S�������>M�V���*�ʿ�p�Ң%��lG�8tf�}�      O���A���}��+Y��3�����$ڿ"����\����(���s��3�9�����p�p�p���<<����e������9{��:�;V$3;ho@;yF;��H;�I;�I;�zI;sZI;yBI;�0I;t$I;EI;tI; I;tI;EI;t$I;�0I;yBI;sZI;�zI;�I;�I;��H;yF;ho@;V$3;�;{��:���9e�������<<�p��p���p�9����3��s�(�������\�"���$ڿ����3��+Y�}�A���      ����,������Q���F�Q�Ù$�.���~�7�}�E(�>�׾�T���L+���սr����@L��jO�9�ͻ�����l8�m�:��;T�1;��?;uF;s�H;��I;��I;��I;�uI;�VI;�@I;1I;�&I;� I;I;� I;�&I;1I;�@I;�VI;�uI;��I;��I;��I;s�H;uF;��?;T�1;��;�m�:��l8���9�ͻjO�@L����r����ս�L+��T��>�׾E(�7�}�~�.���Ù$�F�Q�Q��������,��      �,��^�� P���{��K��x �����n�����w��$���Ҿf��� (���ѽٷ��7����$�K��ɻ����8���:��;��1;@;��F;.I;�I;4�I;ĝI;�tI;NVI;�@I;�0I;�&I;� I;�I;� I;�&I;�0I;�@I;NVI;�tI;ĝI;4�I;�I;.I;��F;@;��1;��;���:��8���ɻ$�K����7�ٷ����ѽ (�f�����Ҿ�$���w�n��������x ��K��{� P��^��      ���� P�������d���;� ����㿰���#f�b��ž��z���C�ƽ40v�e5�R����o@����pj��Pu9]I�:=\;�63;@�@;�F;WI;��I;{�I;o�I;�rI;�TI;^?I;0I;&I;, I;MI;, I;&I;0I;^?I;�TI;�rI;o�I;{�I;��I;WI;�F;@�@;�63;=\;]I�:�Pu9pj�����o@�R���e5�40v�C�ƽ����z�žb��#f�������� ����;���d���� P��      Q����{���d��F�Ù$�7����ɿ,蒿��K�O���j�� Zb�H�8�����a����`���%�.� e��W�غƨ�9�W�:VW;�15;?�A;� G;Z6I;��I;k�I;m�I;�oI;�RI;�=I;�.I;�$I;AI;OI;AI;�$I;�.I;�=I;�RI;�oI;m�I;k�I;��I;Z6I;� G;?�A;�15;VW;�W�:ƨ�9W�غ e��%�.�`��������a�8���H� Zb��j��O����K�,蒿��ɿ7��Ù$��F���d��{�      F�Q��K���;�Ù$��;
��޿�����w�o,���澝���(�D������I��3�G�����N��Ǩ�2��:�����9:���:�m!;��7;۸B;}�G;
YI;L�I;��I;ؑI;�kI;�OI;4;I;�,I;3#I;�I;�I;�I;3#I;�,I;4;I;�OI;�kI;ؑI;��I;L�I;
YI;}�G;۸B;��7;�m!;���:��9::���2��Ǩ��N�����3�G��I������(�D��������o,���w�����޿�;
�Ù$���;��K�      Ù$��x � ��7���޿m���ǅ����F�{�
��~����z��$���ս$���P2+���ϼXPp����K�]��*�"��:,�;�7';��:;�C;+H;�|I;?�I;��I;��I;�fI;�KI;98I;V*I;D!I;I;GI;I;D!I;V*I;98I;�KI;�fI;��I;��I;?�I;�|I;+H;�C;��:;�7';,�;"��:�*�K�]����XPp���ϼP2+�$�����ս�$���z��~��{�
���F�ǅ��m����޿7�� ���x �      .���������㿆�ɿ���ǅ����P�b��:�׾�`��U�H����@��a�a�"����!D�Hɻ�!������U�:�~;�H-;H{=;ABE;ȄH;)�I; �I;��I;ւI;�`I;BGI;�4I;�'I;�I; I;pI; I;�I;�'I;�4I;BGI;�`I;ւI;��I; �I;)�I;ȄH;ABE;H{=;�H-;�~;�U�:�����!�Hɻ!D���"��a�a��@����U�H��`��:�׾b����P�ǅ�������ɿ��㿯���      ~�n�������,蒿��w���F�b��Ȱ�����Yb�+����ѽ�%��'D4����@X��ʨ��H���轺K��9bp�:�; 93;;P@;�uF;9�H;%�I;��I;��I;�yI;�YI;2BI;�0I;�$I;dI;�I;@I;�I;dI;�$I;�0I;2BI;�YI;�yI;��I;��I;%�I;9�H;�uF;;P@; 93;�;bp�:K��9�轺�H��ʨ�@X�����'D4��%����ѽ+���Yb����Ȱ�b����F���w�,蒿����n���      7�}���w�#f���K�o,�{�
�:�׾�����k���'�lz꽥I���;V�LM�*����iO��G�npE����b�:S� ;��$;˳8;q�B;�G;VJI;1�I;9�I;a�I;*pI;�RI;�<I;�,I;%!I;�I;9I;�I;9I;�I;%!I;�,I;�<I;�RI;*pI;a�I;9�I;1�I;VJI;�G;q�B;˳8;��$;S� ;b�:���npE��G��iO�*���LM��;V��I��lz���'���k����:�׾{�
�o,���K�#f���w�      E(��$�b��O������~���`���Yb���'��U�N$��S�m�5����ϼ0�����_�����غ�0�9c��: F;�F.;3{=;aE;�[H;B�I;��I;��I;�I;%fI;%KI;7I;&(I;�I;�I;�I;DI;�I;�I;�I;&(I;7I;%KI;%fI;�I;��I;��I;B�I;�[H;aE;3{=;�F.; F;c��:�0�9��غ_������0����ϼ5��S�m�N$���U���'��Yb��`���~�����O��b���$�      >�׾��Ҿž�j��������z�U�H�+��lz�N$��0v�!2+����9���5�-ɻ44�0�����:���:Nn!;*O6;(kA;��F;��H;��I;��I;�I;k|I;�[I;~CI;%1I;�#I;�I;jI;�I;�I;�I;jI;�I;�#I;%1I;~CI;�[I;k|I;�I;��I;��I;��H;��F;(kA;*O6;Nn!;���:���:0��44�-ɻ�5�9�����!2+�0v�N$��lz�+��U�H���z������j��ž��Ҿ      �T��f�����z� Zb�(�D��$�����ѽ�I��S�m�!2+��������K��ﻙ�p�;������9LR�:�.;��-;��<;iyD;uH;�lI;�I;��I;��I;�nI;�QI;�;I;!+I;�I;*I;NI;�I;�I;�I;NI;*I;�I;!+I;�;I;�QI;�nI;��I;��I;�I;�lI;uH;iyD;��<;��-;�.;LR�:���9;�����p��ﻍ�K������!2+�S�m��I����ѽ���$�(�D� Zb���z�f���      �L+� (���H�������ս�@���%���;V�5���������MS�������zF���n8o�:�;��$;^7;K�A;��F;�H;��I;��I;��I;��I;uaI;�GI;-4I;A%I;II;ZI;I;�	I; 	I;�	I;I;ZI;II;A%I;-4I;�GI;uaI;��I;��I;��I;��I;�H;��F;K�A;^7;��$;�;o�:��n8zF⺧������MS�������5���;V��%���@����ս����H��� (�      ��ս��ѽC�ƽ8����I��$���a�a�'D4�LM���ϼ9����K�����G��]g�p�o���:�@�:�X;��1;jk>;�
E;
/H;;pI;"�I;	�I;��I;!rI;�TI;>I;�,I;~I;�I;�I;�	I;/I;MI;/I;�	I;�I;�I;~I;�,I;>I;�TI;!rI;��I;	�I;"�I;;pI;
/H;�
E;jk>;��1;�X;�@�:��:p�o�]g��G�������K�9����ϼLM�'D4�a�a�$����I��8���C�ƽ��ѽ      r��ٷ��40v���a�3�G�P2+�"�����*���0���5��ﻧ��]g��ହ�g:^�:�;1H-;3f;;NC;)RG;�I;�I;@�I;�I;%�I;+bI;�HI;�4I;�%I;�I;PI;�
I;�I;eI;sI;eI;�I;�
I;PI;�I;�%I;�4I;�HI;+bI;%�I;�I;@�I;�I;�I;)RG;NC;3f;;1H-;�;^�:�g:�ହ]g�������5�0��*������"��P2+�3�G���a�40v�ٷ��      ��7�e5���������ϼ��@X���iO����-ɻ��p�zF�p�o��g:^�:YF;�*;�9;��A;�tF;;�H;�I;��I;ɺI;e�I;�oI;SSI;n=I;9,I;�I;�I;I;pI;�I;�I;� I;�I;�I;pI;I;�I;�I;9,I;n=I;SSI;�oI;e�I;ɺI;��I;�I;;�H;�tF;��A;�9;�*;YF;^�:�g:p�o�zF⺙�p�-ɻ����iO�@X������ϼ������e5�7�      @L�����R���`����N��XPp�!D�ʨ��G�_���44�;�����n8��:^�:YF;�(;��7;v�@;��E;mPH;5lI;��I;�I;��I;C|I;�]I;�EI;�2I;�#I;zI;�I;		I;(I;� I; �H;h�H; �H;� I;(I;		I;�I;zI;�#I;�2I;�EI;�]I;C|I;��I;�I;��I;5lI;mPH;��E;v�@;��7;�(;YF;^�:��:��n8;���44�_����G�ʨ�!D�XPp��N��`���R������      jO�$�K��o@�%�.�Ǩ����Hɻ�H��npE���غ0�����9o�:�@�:�;�*;��7;�O@;�[E;H;�HI;��I;��I;)�I;|�I;ZgI;�MI;z9I;W)I;�I;�I;�
I;,I;'I;G�H;s�H;��H;s�H;G�H;'I;,I;�
I;�I;�I;W)I;z9I;�MI;ZgI;|�I;)�I;��I;��I;�HI;H;�[E;�O@;��7;�*;�;�@�:o�:���90����غnpE��H��Hɻ���Ǩ�%�.��o@�$�K�      9�ͻ�ɻ��� e��2��K�]��!��轺����0�9���:LR�:�;�X;1H-;�9;v�@;�[E;��G;Q4I;ճI;d�I;��I;m�I;�oI;�TI;q?I;M.I;� I;�I;YI;�I;�I;6�H;��H;,�H;��H;,�H;��H;6�H;�I;�I;YI;�I;� I;M.I;q?I;�TI;�oI;m�I;��I;d�I;ճI;Q4I;��G;�[E;v�@;�9;1H-;�X;�;LR�:���:�0�9����轺�!�K�]�2�� e������ɻ      �����pj�W�غ:����*�����K��9b�:c��:���:�.;��$;��1;3f;;��A;��E;H;Q4I;W�I;��I;m�I;��I;�uI;tZI;xDI;�2I;K$I;�I;�I;hI;�I;��H;s�H;7�H;��H;��H;��H;7�H;s�H;��H;�I;hI;�I;�I;K$I;�2I;xDI;tZI;�uI;��I;m�I;��I;W�I;Q4I;H;��E;��A;3f;;��1;��$;�.;���:c��:b�:K��9�����*�:���W�غpj���      ��l8��8�Pu9ƨ�9��9:"��:�U�:bp�:S� ; F;Nn!;��-;^7;jk>;NC;�tF;mPH;�HI;ճI;��I;ϺI;әI;�yI;�^I;aHI;d6I;}'I;vI;�I;1
I;�I;>�H;��H;��H;�H;��H;��H;��H;�H;��H;��H;>�H;�I;1
I;�I;vI;}'I;d6I;aHI;�^I;�yI;әI;ϺI;��I;ճI;�HI;mPH;�tF;NC;jk>;^7;��-;Nn!; F;S� ;bp�:�U�:"��:��9:ƨ�9�Pu9��8      �m�:���:]I�:�W�:���:,�;�~;�;��$;�F.;*O6;��<;K�A;�
E;)RG;;�H;5lI;��I;d�I;m�I;әI;�zI;�`I;�JI;�8I;�)I;�I;�I;�I;9I; I;�H;��H;{�H; �H;�H;��H;�H; �H;{�H;��H;�H; I;9I;�I;�I;�I;�)I;�8I;�JI;�`I;�zI;әI;m�I;d�I;��I;5lI;;�H;)RG;�
E;K�A;��<;*O6;�F.;��$;�;�~;,�;���:�W�:]I�:���:      ��;��;=\;VW;�m!;�7';�H-; 93;˳8;3{=;(kA;iyD;��F;
/H;�I;�I;��I;��I;��I;��I;�yI;�`I;�KI;4:I;+I;EI;8I;I;MI;� I;��H;�H;w�H;~�H;�H;a�H;2�H;a�H;�H;~�H;w�H;�H;��H;� I;MI;I;8I;EI;+I;4:I;�KI;�`I;�yI;��I;��I;��I;��I;�I;�I;
/H;��F;iyD;(kA;3{=;˳8; 93;�H-;�7';�m!;VW;=\;��;      T�1;��1;�63;�15;��7;��:;H{=;;P@;q�B;aE;��F;uH;�H;;pI;�I;��I;�I;)�I;m�I;�uI;�^I;�JI;4:I;�+I; I;+I;�I;*I;�I;�H;��H;~�H;4�H;��H;z�H;��H;��H;��H;z�H;��H;4�H;~�H;��H;�H;�I;*I;�I;+I; I;�+I;4:I;�JI;�^I;�uI;m�I;)�I;�I;��I;�I;;pI;�H;uH;��F;aE;q�B;;P@;H{=;��:;��7;�15;�63;��1;      ��?;@;@�@;?�A;۸B;�C;ABE;�uF;�G;�[H;��H;�lI;��I;"�I;@�I;ɺI;��I;|�I;�oI;tZI;aHI;�8I;+I; I;�I;sI;�I;I;s�H;��H;��H;;�H;d�H;��H;��H;f�H;=�H;f�H;��H;��H;d�H;;�H;��H;��H;s�H;I;�I;sI;�I; I;+I;�8I;aHI;tZI;�oI;|�I;��I;ɺI;@�I;"�I;��I;�lI;��H;�[H;�G;�uF;ABE;�C;۸B;?�A;@�@;@;      uF;��F;�F;� G;}�G;+H;ȄH;9�H;VJI;B�I;��I;�I;��I;	�I;�I;e�I;C|I;ZgI;�TI;xDI;d6I;�)I;EI;+I;sI;�I;ZI;��H;��H;��H;6�H;I�H;��H;j�H;��H;$�H;��H;$�H;��H;j�H;��H;I�H;6�H;��H;��H;��H;ZI;�I;sI;+I;EI;�)I;d6I;xDI;�TI;ZgI;C|I;e�I;�I;	�I;��I;�I;��I;B�I;VJI;9�H;ȄH;+H;}�G;� G;�F;��F;      s�H;.I;WI;Z6I;
YI;�|I;)�I;%�I;1�I;��I;��I;��I;��I;��I;%�I;�oI;�]I;�MI;q?I;�2I;}'I;�I;8I;�I;�I;ZI;��H;2�H;��H;@�H;1�H;s�H;%�H;#�H;��H;�H;��H;�H;��H;#�H;%�H;s�H;1�H;@�H;��H;2�H;��H;ZI;�I;�I;8I;�I;}'I;�2I;q?I;�MI;�]I;�oI;%�I;��I;��I;��I;��I;��I;1�I;%�I;)�I;�|I;
YI;Z6I;WI;.I;      ��I;�I;��I;��I;L�I;?�I; �I;��I;9�I;��I;�I;��I;��I;!rI;+bI;SSI;�EI;z9I;M.I;K$I;vI;�I;I;*I;I;��H;2�H;�H;L�H;-�H;d�H;��H;��H;
�H;b�H;�H;��H;�H;b�H;
�H;��H;��H;d�H;-�H;L�H;�H;2�H;��H;I;*I;I;�I;vI;K$I;M.I;z9I;�EI;SSI;+bI;!rI;��I;��I;�I;��I;9�I;��I; �I;?�I;L�I;��I;��I;�I;      ��I;4�I;{�I;k�I;��I;��I;��I;��I;a�I;�I;k|I;�nI;uaI;�TI;�HI;n=I;�2I;W)I;� I;�I;�I;�I;MI;�I;s�H;��H;��H;L�H;8�H;a�H;��H;��H;��H;�H;��H;<�H;4�H;<�H;��H;�H;��H;��H;��H;a�H;8�H;L�H;��H;��H;s�H;�I;MI;�I;�I;�I;� I;W)I;�2I;n=I;�HI;�TI;uaI;�nI;k|I;�I;a�I;��I;��I;��I;��I;k�I;{�I;4�I;      ��I;ĝI;o�I;m�I;ؑI;��I;ւI;�yI;*pI;%fI;�[I;�QI;�GI;>I;�4I;9,I;�#I;�I;�I;�I;1
I;9I;� I;�H;��H;��H;@�H;-�H;a�H;��H;��H;��H;��H;"�H;��H;��H;c�H;��H;��H;"�H;��H;��H;��H;��H;a�H;-�H;@�H;��H;��H;�H;� I;9I;1
I;�I;�I;�I;�#I;9,I;�4I;>I;�GI;�QI;�[I;%fI;*pI;�yI;ւI;��I;ؑI;m�I;o�I;ĝI;      �uI;�tI;�rI;�oI;�kI;�fI;�`I;�YI;�RI;%KI;~CI;�;I;-4I;�,I;�%I;�I;zI;�I;YI;hI;�I; I;��H;��H;��H;6�H;1�H;d�H;��H;��H;��H;��H;��H;c�H;�H;��H;��H;��H;�H;c�H;��H;��H;��H;��H;��H;d�H;1�H;6�H;��H;��H;��H; I;�I;hI;YI;�I;zI;�I;�%I;�,I;-4I;�;I;~CI;%KI;�RI;�YI;�`I;�fI;�kI;�oI;�rI;�tI;      �VI;NVI;�TI;�RI;�OI;�KI;BGI;2BI;�<I;7I;%1I;!+I;A%I;~I;�I;�I;�I;�
I;�I;�I;>�H;�H;�H;~�H;;�H;I�H;s�H;��H;��H;��H;��H;��H;K�H;��H;��H;J�H;P�H;J�H;��H;��H;K�H;��H;��H;��H;��H;��H;s�H;I�H;;�H;~�H;�H;�H;>�H;�I;�I;�
I;�I;�I;�I;~I;A%I;!+I;%1I;7I;�<I;2BI;BGI;�KI;�OI;�RI;�TI;NVI;      �@I;�@I;^?I;�=I;4;I;98I;�4I;�0I;�,I;&(I;�#I;�I;II;�I;PI;I;		I;,I;�I;��H;��H;��H;w�H;4�H;d�H;��H;%�H;��H;��H;��H;��H;K�H;��H;d�H;�H;��H;��H;��H;�H;d�H;��H;K�H;��H;��H;��H;��H;%�H;��H;d�H;4�H;w�H;��H;��H;��H;�I;,I;		I;I;PI;�I;II;�I;�#I;&(I;�,I;�0I;�4I;98I;4;I;�=I;^?I;�@I;      1I;�0I;0I;�.I;�,I;V*I;�'I;�$I;%!I;�I;�I;*I;ZI;�I;�
I;pI;(I;'I;6�H;s�H;��H;{�H;~�H;��H;��H;j�H;#�H;
�H;�H;"�H;c�H;��H;d�H;��H;��H;��H;��H;��H;��H;��H;d�H;��H;c�H;"�H;�H;
�H;#�H;j�H;��H;��H;~�H;{�H;��H;s�H;6�H;'I;(I;pI;�
I;�I;ZI;*I;�I;�I;%!I;�$I;�'I;V*I;�,I;�.I;0I;�0I;      �&I;�&I;&I;�$I;3#I;D!I;�I;dI;�I;�I;jI;NI;I;�	I;�I;�I;� I;G�H;��H;7�H;�H; �H;�H;z�H;��H;��H;��H;b�H;��H;��H;�H;��H;�H;��H;��H;d�H;[�H;d�H;��H;��H;�H;��H;�H;��H;��H;b�H;��H;��H;��H;z�H;�H; �H;�H;7�H;��H;G�H;� I;�I;�I;�	I;I;NI;jI;�I;�I;dI;�I;D!I;3#I;�$I;&I;�&I;      � I;� I;, I;AI;�I;I; I;�I;9I;�I;�I;�I;�	I;/I;eI;�I; �H;s�H;,�H;��H;��H;�H;a�H;��H;f�H;$�H;�H;�H;<�H;��H;��H;J�H;��H;��H;d�H;2�H;/�H;2�H;d�H;��H;��H;J�H;��H;��H;<�H;�H;�H;$�H;f�H;��H;a�H;�H;��H;��H;,�H;s�H; �H;�I;eI;/I;�	I;�I;�I;�I;9I;�I; I;I;�I;AI;, I;� I;      I;�I;MI;OI;�I;GI;pI;@I;�I;DI;�I;�I; 	I;MI;sI;� I;h�H;��H;��H;��H;��H;��H;2�H;��H;=�H;��H;��H;��H;4�H;c�H;��H;P�H;��H;��H;[�H;/�H;�H;/�H;[�H;��H;��H;P�H;��H;c�H;4�H;��H;��H;��H;=�H;��H;2�H;��H;��H;��H;��H;��H;h�H;� I;sI;MI; 	I;�I;�I;DI;�I;@I;pI;GI;�I;OI;MI;�I;      � I;� I;, I;AI;�I;I; I;�I;9I;�I;�I;�I;�	I;/I;eI;�I; �H;s�H;,�H;��H;��H;�H;a�H;��H;f�H;$�H;�H;�H;<�H;��H;��H;J�H;��H;��H;d�H;2�H;/�H;2�H;d�H;��H;��H;J�H;��H;��H;<�H;�H;�H;$�H;f�H;��H;a�H;�H;��H;��H;,�H;s�H; �H;�I;eI;/I;�	I;�I;�I;�I;9I;�I; I;I;�I;AI;, I;� I;      �&I;�&I;&I;�$I;3#I;D!I;�I;dI;�I;�I;jI;NI;I;�	I;�I;�I;� I;G�H;��H;7�H;�H; �H;�H;z�H;��H;��H;��H;b�H;��H;��H;�H;��H;�H;��H;��H;d�H;[�H;d�H;��H;��H;�H;��H;�H;��H;��H;b�H;��H;��H;��H;z�H;�H; �H;�H;7�H;��H;G�H;� I;�I;�I;�	I;I;NI;jI;�I;�I;dI;�I;D!I;3#I;�$I;&I;�&I;      1I;�0I;0I;�.I;�,I;V*I;�'I;�$I;%!I;�I;�I;*I;ZI;�I;�
I;pI;(I;'I;6�H;s�H;��H;{�H;~�H;��H;��H;j�H;#�H;
�H;�H;"�H;c�H;��H;d�H;��H;��H;��H;��H;��H;��H;��H;d�H;��H;c�H;"�H;�H;
�H;#�H;j�H;��H;��H;~�H;{�H;��H;s�H;6�H;'I;(I;pI;�
I;�I;ZI;*I;�I;�I;%!I;�$I;�'I;V*I;�,I;�.I;0I;�0I;      �@I;�@I;^?I;�=I;4;I;98I;�4I;�0I;�,I;&(I;�#I;�I;II;�I;PI;I;		I;,I;�I;��H;��H;��H;w�H;4�H;d�H;��H;%�H;��H;��H;��H;��H;K�H;��H;d�H;�H;��H;��H;��H;�H;d�H;��H;K�H;��H;��H;��H;��H;%�H;��H;d�H;4�H;w�H;��H;��H;��H;�I;,I;		I;I;PI;�I;II;�I;�#I;&(I;�,I;�0I;�4I;98I;4;I;�=I;^?I;�@I;      �VI;NVI;�TI;�RI;�OI;�KI;BGI;2BI;�<I;7I;%1I;!+I;A%I;~I;�I;�I;�I;�
I;�I;�I;>�H;�H;�H;~�H;;�H;I�H;s�H;��H;��H;��H;��H;��H;K�H;��H;��H;J�H;P�H;J�H;��H;��H;K�H;��H;��H;��H;��H;��H;s�H;I�H;;�H;~�H;�H;�H;>�H;�I;�I;�
I;�I;�I;�I;~I;A%I;!+I;%1I;7I;�<I;2BI;BGI;�KI;�OI;�RI;�TI;NVI;      �uI;�tI;�rI;�oI;�kI;�fI;�`I;�YI;�RI;%KI;~CI;�;I;-4I;�,I;�%I;�I;zI;�I;YI;hI;�I; I;��H;��H;��H;6�H;1�H;d�H;��H;��H;��H;��H;��H;c�H;�H;��H;��H;��H;�H;c�H;��H;��H;��H;��H;��H;d�H;1�H;6�H;��H;��H;��H; I;�I;hI;YI;�I;zI;�I;�%I;�,I;-4I;�;I;~CI;%KI;�RI;�YI;�`I;�fI;�kI;�oI;�rI;�tI;      ��I;ĝI;o�I;m�I;ؑI;��I;ւI;�yI;*pI;%fI;�[I;�QI;�GI;>I;�4I;9,I;�#I;�I;�I;�I;1
I;9I;� I;�H;��H;��H;@�H;-�H;a�H;��H;��H;��H;��H;"�H;��H;��H;c�H;��H;��H;"�H;��H;��H;��H;��H;a�H;-�H;@�H;��H;��H;�H;� I;9I;1
I;�I;�I;�I;�#I;9,I;�4I;>I;�GI;�QI;�[I;%fI;*pI;�yI;ւI;��I;ؑI;m�I;o�I;ĝI;      ��I;4�I;{�I;k�I;��I;��I;��I;��I;a�I;�I;k|I;�nI;uaI;�TI;�HI;n=I;�2I;W)I;� I;�I;�I;�I;MI;�I;s�H;��H;��H;L�H;8�H;a�H;��H;��H;��H;�H;��H;<�H;4�H;<�H;��H;�H;��H;��H;��H;a�H;8�H;L�H;��H;��H;s�H;�I;MI;�I;�I;�I;� I;W)I;�2I;n=I;�HI;�TI;uaI;�nI;k|I;�I;a�I;��I;��I;��I;��I;k�I;{�I;4�I;      ��I;�I;��I;��I;L�I;?�I; �I;��I;9�I;��I;�I;��I;��I;!rI;+bI;SSI;�EI;z9I;M.I;K$I;vI;�I;I;*I;I;��H;2�H;�H;L�H;-�H;d�H;��H;��H;
�H;b�H;�H;��H;�H;b�H;
�H;��H;��H;d�H;-�H;L�H;�H;2�H;��H;I;*I;I;�I;vI;K$I;M.I;z9I;�EI;SSI;+bI;!rI;��I;��I;�I;��I;9�I;��I; �I;?�I;L�I;��I;��I;�I;      s�H;.I;WI;Z6I;
YI;�|I;)�I;%�I;1�I;��I;��I;��I;��I;��I;%�I;�oI;�]I;�MI;q?I;�2I;}'I;�I;8I;�I;�I;ZI;��H;2�H;��H;@�H;1�H;s�H;%�H;#�H;��H;�H;��H;�H;��H;#�H;%�H;s�H;1�H;@�H;��H;2�H;��H;ZI;�I;�I;8I;�I;}'I;�2I;q?I;�MI;�]I;�oI;%�I;��I;��I;��I;��I;��I;1�I;%�I;)�I;�|I;
YI;Z6I;WI;.I;      uF;��F;�F;� G;}�G;+H;ȄH;9�H;VJI;B�I;��I;�I;��I;	�I;�I;e�I;C|I;ZgI;�TI;xDI;d6I;�)I;EI;+I;sI;�I;ZI;��H;��H;��H;6�H;I�H;��H;j�H;��H;$�H;��H;$�H;��H;j�H;��H;I�H;6�H;��H;��H;��H;ZI;�I;sI;+I;EI;�)I;d6I;xDI;�TI;ZgI;C|I;e�I;�I;	�I;��I;�I;��I;B�I;VJI;9�H;ȄH;+H;}�G;� G;�F;��F;      ��?;@;@�@;?�A;۸B;�C;ABE;�uF;�G;�[H;��H;�lI;��I;"�I;@�I;ɺI;��I;|�I;�oI;tZI;aHI;�8I;+I; I;�I;sI;�I;I;s�H;��H;��H;;�H;d�H;��H;��H;f�H;=�H;f�H;��H;��H;d�H;;�H;��H;��H;s�H;I;�I;sI;�I; I;+I;�8I;aHI;tZI;�oI;|�I;��I;ɺI;@�I;"�I;��I;�lI;��H;�[H;�G;�uF;ABE;�C;۸B;?�A;@�@;@;      T�1;��1;�63;�15;��7;��:;H{=;;P@;q�B;aE;��F;uH;�H;;pI;�I;��I;�I;)�I;m�I;�uI;�^I;�JI;4:I;�+I; I;+I;�I;*I;�I;�H;��H;~�H;4�H;��H;z�H;��H;��H;��H;z�H;��H;4�H;~�H;��H;�H;�I;*I;�I;+I; I;�+I;4:I;�JI;�^I;�uI;m�I;)�I;�I;��I;�I;;pI;�H;uH;��F;aE;q�B;;P@;H{=;��:;��7;�15;�63;��1;      ��;��;=\;VW;�m!;�7';�H-; 93;˳8;3{=;(kA;iyD;��F;
/H;�I;�I;��I;��I;��I;��I;�yI;�`I;�KI;4:I;+I;EI;8I;I;MI;� I;��H;�H;w�H;~�H;�H;a�H;2�H;a�H;�H;~�H;w�H;�H;��H;� I;MI;I;8I;EI;+I;4:I;�KI;�`I;�yI;��I;��I;��I;��I;�I;�I;
/H;��F;iyD;(kA;3{=;˳8; 93;�H-;�7';�m!;VW;=\;��;      �m�:���:]I�:�W�:���:,�;�~;�;��$;�F.;*O6;��<;K�A;�
E;)RG;;�H;5lI;��I;d�I;m�I;әI;�zI;�`I;�JI;�8I;�)I;�I;�I;�I;9I; I;�H;��H;{�H; �H;�H;��H;�H; �H;{�H;��H;�H; I;9I;�I;�I;�I;�)I;�8I;�JI;�`I;�zI;әI;m�I;d�I;��I;5lI;;�H;)RG;�
E;K�A;��<;*O6;�F.;��$;�;�~;,�;���:�W�:]I�:���:      ��l8��8�Pu9ƨ�9��9:"��:�U�:bp�:S� ; F;Nn!;��-;^7;jk>;NC;�tF;mPH;�HI;ճI;��I;ϺI;әI;�yI;�^I;aHI;d6I;}'I;vI;�I;1
I;�I;>�H;��H;��H;�H;��H;��H;��H;�H;��H;��H;>�H;�I;1
I;�I;vI;}'I;d6I;aHI;�^I;�yI;әI;ϺI;��I;ճI;�HI;mPH;�tF;NC;jk>;^7;��-;Nn!; F;S� ;bp�:�U�:"��:��9:ƨ�9�Pu9��8      �����pj�W�غ:����*�����K��9b�:c��:���:�.;��$;��1;3f;;��A;��E;H;Q4I;W�I;��I;m�I;��I;�uI;tZI;xDI;�2I;K$I;�I;�I;hI;�I;��H;s�H;7�H;��H;��H;��H;7�H;s�H;��H;�I;hI;�I;�I;K$I;�2I;xDI;tZI;�uI;��I;m�I;��I;W�I;Q4I;H;��E;��A;3f;;��1;��$;�.;���:c��:b�:K��9�����*�:���W�غpj���      9�ͻ�ɻ��� e��2��K�]��!��轺����0�9���:LR�:�;�X;1H-;�9;v�@;�[E;��G;Q4I;ճI;d�I;��I;m�I;�oI;�TI;q?I;M.I;� I;�I;YI;�I;�I;6�H;��H;,�H;��H;,�H;��H;6�H;�I;�I;YI;�I;� I;M.I;q?I;�TI;�oI;m�I;��I;d�I;ճI;Q4I;��G;�[E;v�@;�9;1H-;�X;�;LR�:���:�0�9����轺�!�K�]�2�� e������ɻ      jO�$�K��o@�%�.�Ǩ����Hɻ�H��npE���غ0�����9o�:�@�:�;�*;��7;�O@;�[E;H;�HI;��I;��I;)�I;|�I;ZgI;�MI;z9I;W)I;�I;�I;�
I;,I;'I;G�H;s�H;��H;s�H;G�H;'I;,I;�
I;�I;�I;W)I;z9I;�MI;ZgI;|�I;)�I;��I;��I;�HI;H;�[E;�O@;��7;�*;�;�@�:o�:���90����غnpE��H��Hɻ���Ǩ�%�.��o@�$�K�      @L�����R���`����N��XPp�!D�ʨ��G�_���44�;�����n8��:^�:YF;�(;��7;v�@;��E;mPH;5lI;��I;�I;��I;C|I;�]I;�EI;�2I;�#I;zI;�I;		I;(I;� I; �H;h�H; �H;� I;(I;		I;�I;zI;�#I;�2I;�EI;�]I;C|I;��I;�I;��I;5lI;mPH;��E;v�@;��7;�(;YF;^�:��:��n8;���44�_����G�ʨ�!D�XPp��N��`���R������      ��7�e5���������ϼ��@X���iO����-ɻ��p�zF�p�o��g:^�:YF;�*;�9;��A;�tF;;�H;�I;��I;ɺI;e�I;�oI;SSI;n=I;9,I;�I;�I;I;pI;�I;�I;� I;�I;�I;pI;I;�I;�I;9,I;n=I;SSI;�oI;e�I;ɺI;��I;�I;;�H;�tF;��A;�9;�*;YF;^�:�g:p�o�zF⺙�p�-ɻ����iO�@X������ϼ������e5�7�      r��ٷ��40v���a�3�G�P2+�"�����*���0���5��ﻧ��]g��ହ�g:^�:�;1H-;3f;;NC;)RG;�I;�I;@�I;�I;%�I;+bI;�HI;�4I;�%I;�I;PI;�
I;�I;eI;sI;eI;�I;�
I;PI;�I;�%I;�4I;�HI;+bI;%�I;�I;@�I;�I;�I;)RG;NC;3f;;1H-;�;^�:�g:�ହ]g�������5�0��*������"��P2+�3�G���a�40v�ٷ��      ��ս��ѽC�ƽ8����I��$���a�a�'D4�LM���ϼ9����K�����G��]g�p�o���:�@�:�X;��1;jk>;�
E;
/H;;pI;"�I;	�I;��I;!rI;�TI;>I;�,I;~I;�I;�I;�	I;/I;MI;/I;�	I;�I;�I;~I;�,I;>I;�TI;!rI;��I;	�I;"�I;;pI;
/H;�
E;jk>;��1;�X;�@�:��:p�o�]g��G�������K�9����ϼLM�'D4�a�a�$����I��8���C�ƽ��ѽ      �L+� (���H�������ս�@���%���;V�5���������MS�������zF���n8o�:�;��$;^7;K�A;��F;�H;��I;��I;��I;��I;uaI;�GI;-4I;A%I;II;ZI;I;�	I; 	I;�	I;I;ZI;II;A%I;-4I;�GI;uaI;��I;��I;��I;��I;�H;��F;K�A;^7;��$;�;o�:��n8zF⺧������MS�������5���;V��%���@����ս����H��� (�      �T��f�����z� Zb�(�D��$�����ѽ�I��S�m�!2+��������K��ﻙ�p�;������9LR�:�.;��-;��<;iyD;uH;�lI;�I;��I;��I;�nI;�QI;�;I;!+I;�I;*I;NI;�I;�I;�I;NI;*I;�I;!+I;�;I;�QI;�nI;��I;��I;�I;�lI;uH;iyD;��<;��-;�.;LR�:���9;�����p��ﻍ�K������!2+�S�m��I����ѽ���$�(�D� Zb���z�f���      >�׾��Ҿž�j��������z�U�H�+��lz�N$��0v�!2+����9���5�-ɻ44�0�����:���:Nn!;*O6;(kA;��F;��H;��I;��I;�I;k|I;�[I;~CI;%1I;�#I;�I;jI;�I;�I;�I;jI;�I;�#I;%1I;~CI;�[I;k|I;�I;��I;��I;��H;��F;(kA;*O6;Nn!;���:���:0��44�-ɻ�5�9�����!2+�0v�N$��lz�+��U�H���z������j��ž��Ҿ      E(��$�b��O������~���`���Yb���'��U�N$��S�m�5����ϼ0�����_�����غ�0�9c��: F;�F.;3{=;aE;�[H;B�I;��I;��I;�I;%fI;%KI;7I;&(I;�I;�I;�I;DI;�I;�I;�I;&(I;7I;%KI;%fI;�I;��I;��I;B�I;�[H;aE;3{=;�F.; F;c��:�0�9��غ_������0����ϼ5��S�m�N$���U���'��Yb��`���~�����O��b���$�      7�}���w�#f���K�o,�{�
�:�׾�����k���'�lz꽥I���;V�LM�*����iO��G�npE����b�:S� ;��$;˳8;q�B;�G;VJI;1�I;9�I;a�I;*pI;�RI;�<I;�,I;%!I;�I;9I;�I;9I;�I;%!I;�,I;�<I;�RI;*pI;a�I;9�I;1�I;VJI;�G;q�B;˳8;��$;S� ;b�:���npE��G��iO�*���LM��;V��I��lz���'���k����:�׾{�
�o,���K�#f���w�      ~�n�������,蒿��w���F�b��Ȱ�����Yb�+����ѽ�%��'D4����@X��ʨ��H���轺K��9bp�:�; 93;;P@;�uF;9�H;%�I;��I;��I;�yI;�YI;2BI;�0I;�$I;dI;�I;@I;�I;dI;�$I;�0I;2BI;�YI;�yI;��I;��I;%�I;9�H;�uF;;P@; 93;�;bp�:K��9�轺�H��ʨ�@X�����'D4��%����ѽ+���Yb����Ȱ�b����F���w�,蒿����n���      .���������㿆�ɿ���ǅ����P�b��:�׾�`��U�H����@��a�a�"����!D�Hɻ�!������U�:�~;�H-;H{=;ABE;ȄH;)�I; �I;��I;ւI;�`I;BGI;�4I;�'I;�I; I;pI; I;�I;�'I;�4I;BGI;�`I;ւI;��I; �I;)�I;ȄH;ABE;H{=;�H-;�~;�U�:�����!�Hɻ!D���"��a�a��@����U�H��`��:�׾b����P�ǅ�������ɿ��㿯���      Ù$��x � ��7���޿m���ǅ����F�{�
��~����z��$���ս$���P2+���ϼXPp����K�]��*�"��:,�;�7';��:;�C;+H;�|I;?�I;��I;��I;�fI;�KI;98I;V*I;D!I;I;GI;I;D!I;V*I;98I;�KI;�fI;��I;��I;?�I;�|I;+H;�C;��:;�7';,�;"��:�*�K�]����XPp���ϼP2+�$�����ս�$���z��~��{�
���F�ǅ��m����޿7�� ���x �      F�Q��K���;�Ù$��;
��޿�����w�o,���澝���(�D������I��3�G�����N��Ǩ�2��:�����9:���:�m!;��7;۸B;}�G;
YI;L�I;��I;ؑI;�kI;�OI;4;I;�,I;3#I;�I;�I;�I;3#I;�,I;4;I;�OI;�kI;ؑI;��I;L�I;
YI;}�G;۸B;��7;�m!;���:��9::���2��Ǩ��N�����3�G��I������(�D��������o,���w�����޿�;
�Ù$���;��K�      Q����{���d��F�Ù$�7����ɿ,蒿��K�O���j�� Zb�H�8�����a����`���%�.� e��W�غƨ�9�W�:VW;�15;?�A;� G;Z6I;��I;k�I;m�I;�oI;�RI;�=I;�.I;�$I;AI;OI;AI;�$I;�.I;�=I;�RI;�oI;m�I;k�I;��I;Z6I;� G;?�A;�15;VW;�W�:ƨ�9W�غ e��%�.�`��������a�8���H� Zb��j��O����K�,蒿��ɿ7��Ù$��F���d��{�      ���� P�������d���;� ����㿰���#f�b��ž��z���C�ƽ40v�e5�R����o@����pj��Pu9]I�:=\;�63;@�@;�F;WI;��I;{�I;o�I;�rI;�TI;^?I;0I;&I;, I;MI;, I;&I;0I;^?I;�TI;�rI;o�I;{�I;��I;WI;�F;@�@;�63;=\;]I�:�Pu9pj�����o@�R���e5�40v�C�ƽ����z�žb��#f�������� ����;���d���� P��      �,��^�� P���{��K��x �����n�����w��$���Ҿf��� (���ѽٷ��7����$�K��ɻ����8���:��;��1;@;��F;.I;�I;4�I;ĝI;�tI;NVI;�@I;�0I;�&I;� I;�I;� I;�&I;�0I;�@I;NVI;�tI;ĝI;4�I;�I;.I;��F;@;��1;��;���:��8���ɻ$�K����7�ٷ����ѽ (�f�����Ҿ�$���w�n��������x ��K��{� P��^��      A(��o'���o��L�d��X1�|x�Ŀ����3�v���x����4�s��b+���'�"�ü�yY�llٻq&�e�p�X��:_;��0;��?;�F;tI;�I;��I;H�I;��I;ucI;�JI;�8I;�-I;�&I;�$I;�&I;�-I;�8I;�JI;ucI;��I;H�I;��I;�I;tI;�F;��?;��0;_;X��:e�p�q&�llٻ�yY�"�ü�'�b+��s����4��x��v���3����Ŀ|x��X1�d�L��o��o'��      o'���X��c^�������]]���,�N9�3g��S�����/����o��j1��hܽ���-$��l��,}U��Ի~!� �-���:;�41;��?;m�F;N&I;��I;7�I;Y�I;ąI;�bI;\JI;�8I;E-I;�&I;�$I;�&I;E-I;�8I;\JI;�bI;ąI;Y�I;7�I;��I;N&I;m�F;��?;�41;;��: �-�~!��Ի,}U��l���-$����hܽj1��o���྘�/�S���3g��N9���,��]]�����c^���X��      �o��c^���ē��4z�1K�e��M��$ﱿQ�v��X#���Ѿń�	�&�w�нk̀�r��������I� ǻ�5��9�
�:W�;!�2;��@;�F;:I;�I;�I;��I;��I;qaI;II;�7I;~,I;�%I;�#I;�%I;~,I;�7I;II;qaI;��I;��I;�I;�I;:I;�F;��@;!�2;W�;�
�:�9�5� ǻ��I�����r��k̀�w�н	�&�ń���Ѿ�X#�Q�v�$ﱿM��e��1K��4z��ē�c^��      L������4z���V��X1��<�pؿ����RZ��	�(���KUo����fy��?l�l�S����7������𺢽�9��:��;\�4;�sA;�1G;�WI;��I;r�I;)�I;�I;�^I;GI;A6I;+I;�$I;�"I;�$I;+I;A6I;GI;�^I;�I;)�I;r�I;��I;�WI;�1G;�sA;\�4;��;��:���9�𺙼����7�S��l�?l�fy�����KUo�(����	��RZ����pؿ�<��X1���V��4z�����      d��]]�1K��X1�Xf���kQ��R���Z58��A���נ���O���h什�Q�,���cߓ��� �W��}谺�":��:# ;�/7;�B;`�G;{I;�I;��I;ԦI;]{I;Z[I;hDI;;4I;X)I;Q#I;G!I;Q#I;X)I;;4I;hDI;Z[I;]{I;ԦI;��I;�I;{I;`�G;�B;�/7;# ;��:�":}谺W���� �cߓ�,����Q�h什����O��נ��A��Z58�R���kQ����Xf��X1�1K��]]�      �X1���,�e���<���2g��c_���U�˂�ՌȾ	ń�-�-�q��Y ��8�2�.?ټ��{�G"��n��O���u:�O ;�&;5":;[�C;!%H;0�I;C�I;��I;�I;�uI;�VI;AI;�1I;3'I;c!I;}I;c!I;3'I;�1I;AI;�VI;�uI;�I;��I;C�I;0�I;!%H;[�C;5":;�&;�O ;��u:�O��n�G"���{�.?ټ8�2�Y ��q��-�-�	ń�ՌȾ˂��U�c_��2g���<�e����,�      |x�N9�M��pؿkQ��c_��4�_��X#�p���f��<�S�{�����-l�T�-w��f�M�#�Ի �+��LT���:�d;�[,;/=;�AE;|�H;��I;��I;��I;֕I;�nI;�QI;/=I;|.I;�$I;I;cI;I;�$I;|.I;/=I;�QI;�nI;֕I;��I;��I;��I;|�H;�AE;/=;�[,;�d;��:�LT� �+�#�Իf�M�-w��T�-l�����{�<�S��f��p���X#�4�_�c_��kQ��pؿM��N9�      Ŀ3g��$ﱿ���R����U��X#�r��d���JUo�
�#��hܽ����n<����`���҉ �;❻J�Ժ�l�9q��:�U;�2;�@;t�F;�I;�I;b�I;K�I;��I;%gI;.LI;�8I;+I;�!I;�I;�I;�I;�!I;+I;�8I;.LI;%gI;��I;K�I;b�I;�I;�I;t�F;�@;�2;�U;q��:�l�9J�Ժ;❻҉ �`�������n<�����hܽ
�#�JUo�d���r���X#��U�R������$ﱿ3g��      ���S���Q�v��RZ�Z58�˂�p��d���hoy�`1�gO��d什�`�`��7����yY���컟�T��1���u:��:\~#;.88;�B;��G;lI;-�I;!�I;L�I;��I;�^I;!FI;4I;C'I;�I;�I;)I;�I;�I;C'I;4I;!FI;�^I;��I;L�I;!�I;-�I;lI;��G;�B;.88;\~#;��:��u:�1���T���컷yY�7���`���`�d什gO��`1�hoy�d���p��˂�Z58��RZ�Q�v�S���      �3���/��X#��	��A��ՌȾ�f��JUo�`1�Ӱ���n���x��'��>ټ�@��-l�S���%���39�!�:;Q; d-;�.=;�E;~wH;��I;,�I;��I; �I;6uI;�VI;�?I;/I;B#I;_I;�I;TI;�I;_I;B#I;/I;�?I;�VI;6uI; �I;��I;,�I;��I;~wH;�E;�.=; d-;;Q;�!�:�39%��S���-l��@���>ټ�'��x��n��Ӱ��`1�JUo��f��ՌȾ�A���	��X#���/�      v���ྃ�Ѿ(����נ�	ń�<�S�
�#�gO���n��R̀��2�-������>���Ի��B��#�Ym:�E�:o ;��5;�EA;��F;�I;r�I;p�I;ŽI;��I;�iI;�MI;.9I;�)I;I;�I;�I;iI;�I;�I;I;�)I;.9I;�MI;�iI;��I;ŽI;p�I;r�I;�I;��F;�EA;��5;o ;�E�:Ym:�#���B���Ի��>���-���2�R̀��n��gO��
�#�<�S�	ń��נ�(�����Ѿ��      �x���o��ń�KUo���O�-�-�{��hܽd什�x��2��b��yR���|U��2�����$찺�m�9��:C;��,;�g<;�qD;g$H;�I;��I;��I;&�I;&I;�]I;(EI;r2I;�$I;�I;}I;�I;PI;�I;}I;�I;�$I;r2I;(EI;�]I;&I;&�I;��I;��I;�I;g$H;�qD;�g<;��,;C;��:�m�9$찺����2���|U�yR���b���2��x�d什�hܽ{�-�-���O�KUo�ń��o��      ��4�j1�	�&������q�ཌྷ�������`��'�-��yR����]�����V��	[����o����:{�;=~#;/�6;nsA;r�F;�I;��I;��I;��I;6�I;�oI;�RI;�<I;�+I;�I;�I;�I;`I;VI;`I;�I;�I;�I;�+I;�<I;�RI;�oI;6�I;��I;��I;��I;�I;r�F;nsA;/�6;=~#;{�;���:��o�	[���V�������]�yR��-��'��`��������q�������	�&�j1�      s�ཾhܽw�нfy��h什Y ��-l��n<�`���>ټ�𛼞|U����H᝻�2�������u:ij�:�;}61;j(>;rE;+IH;p�I;��I;��I;�I;��I;zaI;�GI;G4I;~%I;�I;�I;XI;<
I;6	I;<
I;XI;�I;�I;~%I;G4I;�GI;zaI;��I;�I;��I;��I;p�I;+IH;rE;j(>;}61;�;ij�:��u:�����2�H᝻����|U����>ټ`���n<�-l�Y ��h什fy��w�н�hܽ      b+����k̀�?l��Q�8�2�T����7����@����>��2���V���2���� R:���:�;�[,;P;;;C;�dG;w8I;��I;U�I;��I;^�I;�pI;�SI;=I;W,I;KI;�I;�I;�	I;+I;'I;+I;�	I;�I;�I;KI;W,I;=I;�SI;�pI;^�I;��I;U�I;��I;w8I;�dG;;C;P;;�[,;�;���: R:���2��V���2����>��@��7������T�8�2��Q�?l�k̀���      �'��-$�r��l�,���.?ټ-w��`����yY�-l���Ի���	[������ R:���:�Q;�);��8;��A;�F;R�H;I�I;��I;��I;ȨI;$�I;�_I;GI;�3I;�$I;cI;�I;�
I;�I;*I;]I;*I;�I;�
I;�I;cI;�$I;�3I;GI;�_I;$�I;ȨI;��I;��I;I�I;R�H;�F;��A;��8;�);�Q;���: R:����	[�������Ի-l��yY�`���-w��.?ټ,���l�r���-$�      "�ü�l������S��cߓ���{�f�M�҉ ����S�����B�$찺��o���u:���:�Q;D�';)07;ք@;�E;�kH;N�I;��I;��I;+�I;��I;�kI;�PI;D;I;�*I;�I;�I;|I;�I;[I;CI;� I;CI;[I;�I;|I;�I;�I;�*I;D;I;�PI;�kI;��I;+�I;��I;��I;N�I;�kH;�E;ք@;)07;D�';�Q;���:��u:��o�$찺��B�S������҉ �f�M���{�cߓ�S�������l��      �yY�,}U���I���7��� �G"�#�Ի;❻��T�%���#��m�9���:ij�:�;�);)07;D@;V\E;�#H;�jI;(�I;s�I;�I;L�I;�vI;�YI;�BI;�0I;g"I;CI;�I;EI;�I;N I;�H;�H;�H;N I;�I;EI;�I;CI;g"I;�0I;�BI;�YI;�vI;L�I;�I;s�I;(�I;�jI;�#H;V\E;D@;)07;�);�;ij�:���:�m�9�#�%���T�;❻#�ԻG"��� ���7���I�,}U�      llٻ�Ի ǻ����W���n� �+�J�Ժ�1��39Ym:��:{�;�;�[,;��8;ք@;V\E;�	H;jUI;��I;	�I;�I;}�I;#�I;�aI;}II;>6I;�&I;�I;GI;�	I;NI;O I;{�H;��H;��H;��H;{�H;O I;NI;�	I;GI;�I;�&I;>6I;}II;�aI;#�I;}�I;�I;	�I;��I;jUI;�	H;V\E;ք@;��8;�[,;�;{�;��:Ym:�39�1�J�Ժ �+��n�W������ ǻ�Ի      q&�~!��5���}谺�O��LT��l�9��u:�!�:�E�:C;=~#;}61;P;;��A;�E;�#H;jUI;,�I;��I;0�I;��I;�I;-hI;BOI;6;I;+I;3I;�I;�I;�I;� I;F�H;��H;��H;�H;��H;��H;F�H;� I;�I;�I;�I;3I;+I;6;I;BOI;-hI;�I;��I;0�I;��I;,�I;jUI;�#H;�E;��A;P;;}61;=~#;C;�E�:�!�:��u:�l�9�LT��O�}谺���5�~!�      e�p� �-��9���9�":��u:��:q��:��:;Q;o ;��,;/�6;j(>;;C;�F;�kH;�jI;��I;��I;��I;4�I;��I;�lI;�SI;??I;�.I;8!I;nI;�I;�I;�I;��H;��H;��H;c�H;��H;c�H;��H;��H;��H;�I;�I;�I;nI;8!I;�.I;??I;�SI;�lI;��I;4�I;��I;��I;��I;�jI;�kH;�F;;C;j(>;/�6;��,;o ;;Q;��:q��:��:��u:�":���9�9 �-�      X��:��:�
�:��:��:�O ;�d;�U;\~#; d-;��5;�g<;nsA;rE;�dG;R�H;N�I;(�I;	�I;0�I;4�I;�I;!oI;aVI;BI;X1I;�#I;�I;�I;VI;�I;�H;��H;�H;f�H;>�H;��H;>�H;f�H;�H;��H;�H;�I;VI;�I;�I;�#I;X1I;BI;aVI;!oI;�I;4�I;0�I;	�I;(�I;N�I;R�H;�dG;rE;nsA;�g<;��5; d-;\~#;�U;�d;�O ;��:��:�
�:��:      _;;W�;��;# ;�&;�[,;�2;.88;�.=;�EA;�qD;r�F;+IH;w8I;I�I;��I;s�I;�I;��I;��I;!oI;bWI;�CI;3I;r%I;7I;�I;�	I;�I;��H;��H;��H;��H;H�H;V�H;�H;V�H;H�H;��H;��H;��H;��H;�I;�	I;�I;7I;r%I;3I;�CI;bWI;!oI;��I;��I;�I;s�I;��I;I�I;w8I;+IH;r�F;�qD;�EA;�.=;.88;�2;�[,;�&;# ;��;W�;;      ��0;�41;!�2;\�4;�/7;5":;/=;�@;�B;�E;��F;g$H;�I;p�I;��I;��I;��I;�I;}�I;�I;�lI;aVI;�CI;�3I;Y&I;DI;I;�
I;II;>�H;A�H;��H;��H;��H;o�H;��H;w�H;��H;o�H;��H;��H;��H;A�H;>�H;II;�
I;I;DI;Y&I;�3I;�CI;aVI;�lI;�I;}�I;�I;��I;��I;��I;p�I;�I;g$H;��F;�E;�B;�@;/=;5":;�/7;\�4;!�2;�41;      ��?;��?;��@;�sA;�B;[�C;�AE;t�F;��G;~wH;�I;�I;��I;��I;U�I;��I;+�I;L�I;#�I;-hI;�SI;BI;3I;Y&I;�I;�I;)I;�I;��H;��H;&�H;z�H;p�H;��H;��H;5�H;�H;5�H;��H;��H;p�H;z�H;&�H;��H;��H;�I;)I;�I;�I;Y&I;3I;BI;�SI;-hI;#�I;L�I;+�I;��I;U�I;��I;��I;�I;�I;~wH;��G;t�F;�AE;[�C;�B;�sA;��@;��?;      �F;m�F;�F;�1G;`�G;!%H;|�H;�I;lI;��I;r�I;��I;��I;��I;��I;ȨI;��I;�vI;�aI;BOI;??I;X1I;r%I;DI;�I;OI;1I; I;��H;U�H;��H;c�H;��H;4�H;e�H;��H;��H;��H;e�H;4�H;��H;c�H;��H;U�H;��H; I;1I;OI;�I;DI;r%I;X1I;??I;BOI;�aI;�vI;��I;ȨI;��I;��I;��I;��I;r�I;��I;lI;�I;|�H;!%H;`�G;�1G;�F;m�F;      tI;N&I;:I;�WI;{I;0�I;��I;�I;-�I;,�I;p�I;��I;��I;�I;^�I;$�I;�kI;�YI;}II;6;I;�.I;�#I;7I;I;)I;1I; I;��H;}�H;��H;\�H;`�H;��H;��H;�H;��H;w�H;��H;�H;��H;��H;`�H;\�H;��H;}�H;��H; I;1I;)I;I;7I;�#I;�.I;6;I;}II;�YI;�kI;$�I;^�I;�I;��I;��I;p�I;,�I;-�I;�I;��I;0�I;{I;�WI;:I;N&I;      �I;��I;�I;��I;�I;C�I;��I;b�I;!�I;��I;ŽI;&�I;6�I;��I;�pI;�_I;�PI;�BI;>6I;+I;8!I;�I;�I;�
I;�I; I;��H;y�H;��H;c�H;a�H;��H;��H;��H;��H;��H;y�H;��H;��H;��H;��H;��H;a�H;c�H;��H;y�H;��H; I;�I;�
I;�I;�I;8!I;+I;>6I;�BI;�PI;�_I;�pI;��I;6�I;&�I;ŽI;��I;!�I;b�I;��I;C�I;�I;��I;�I;��I;      ��I;7�I;�I;r�I;��I;��I;��I;K�I;L�I; �I;��I;&I;�oI;zaI;�SI;GI;D;I;�0I;�&I;3I;nI;�I;�	I;II;��H;��H;}�H;��H;X�H;[�H;��H;Z�H;K�H;��H;��H;��H;��H;��H;��H;��H;K�H;Z�H;��H;[�H;X�H;��H;}�H;��H;��H;II;�	I;�I;nI;3I;�&I;�0I;D;I;GI;�SI;zaI;�oI;&I;��I; �I;L�I;K�I;��I;��I;��I;r�I;�I;7�I;      H�I;Y�I;��I;)�I;ԦI;�I;֕I;��I;��I;6uI;�iI;�]I;�RI;�GI;=I;�3I;�*I;g"I;�I;�I;�I;VI;�I;>�H;��H;U�H;��H;c�H;[�H;��H;6�H;�H;B�H;��H;�H;��H;��H;��H;�H;��H;B�H;�H;6�H;��H;[�H;c�H;��H;U�H;��H;>�H;�I;VI;�I;�I;�I;g"I;�*I;�3I;=I;�GI;�RI;�]I;�iI;6uI;��I;��I;֕I;�I;ԦI;)�I;��I;Y�I;      ��I;ąI;��I;�I;]{I;�uI;�nI;%gI;�^I;�VI;�MI;(EI;�<I;G4I;W,I;�$I;�I;CI;GI;�I;�I;�I;��H;A�H;&�H;��H;\�H;a�H;��H;6�H;�H;�H;\�H;��H;z�H;7�H;��H;7�H;z�H;��H;\�H;�H;�H;6�H;��H;a�H;\�H;��H;&�H;A�H;��H;�I;�I;�I;GI;CI;�I;�$I;W,I;G4I;�<I;(EI;�MI;�VI;�^I;%gI;�nI;�uI;]{I;�I;��I;ąI;      ucI;�bI;qaI;�^I;Z[I;�VI;�QI;.LI;!FI;�?I;.9I;r2I;�+I;~%I;KI;cI;�I;�I;�	I;�I;�I;�H;��H;��H;z�H;c�H;`�H;��H;Z�H;�H;�H;U�H;��H;,�H;��H;��H;��H;��H;��H;,�H;��H;U�H;�H;�H;Z�H;��H;`�H;c�H;z�H;��H;��H;�H;�I;�I;�	I;�I;�I;cI;KI;~%I;�+I;r2I;.9I;�?I;!FI;.LI;�QI;�VI;Z[I;�^I;qaI;�bI;      �JI;\JI;II;GI;hDI;AI;/=I;�8I;4I;/I;�)I;�$I;�I;�I;�I;�I;|I;EI;NI;� I;��H;��H;��H;��H;p�H;��H;��H;��H;K�H;B�H;\�H;��H;�H;��H;M�H;!�H;3�H;!�H;M�H;��H;�H;��H;\�H;B�H;K�H;��H;��H;��H;p�H;��H;��H;��H;��H;� I;NI;EI;|I;�I;�I;�I;�I;�$I;�)I;/I;4I;�8I;/=I;AI;hDI;GI;II;\JI;      �8I;�8I;�7I;A6I;;4I;�1I;|.I;+I;C'I;B#I;I;�I;�I;�I;�I;�
I;�I;�I;O I;F�H;��H;�H;��H;��H;��H;4�H;��H;��H;��H;��H;��H;,�H;��H;<�H;��H;��H;��H;��H;��H;<�H;��H;,�H;��H;��H;��H;��H;��H;4�H;��H;��H;��H;�H;��H;F�H;O I;�I;�I;�
I;�I;�I;�I;�I;I;B#I;C'I;+I;|.I;�1I;;4I;A6I;�7I;�8I;      �-I;E-I;~,I;+I;X)I;3'I;�$I;�!I;�I;_I;�I;}I;�I;XI;�	I;�I;[I;N I;{�H;��H;��H;f�H;H�H;o�H;��H;e�H;�H;��H;��H;�H;z�H;��H;M�H;��H;��H;��H;�H;��H;��H;��H;M�H;��H;z�H;�H;��H;��H;�H;e�H;��H;o�H;H�H;f�H;��H;��H;{�H;N I;[I;�I;�	I;XI;�I;}I;�I;_I;�I;�!I;�$I;3'I;X)I;+I;~,I;E-I;      �&I;�&I;�%I;�$I;Q#I;c!I;I;�I;�I;�I;�I;�I;`I;<
I;+I;*I;CI;�H;��H;��H;c�H;>�H;V�H;��H;5�H;��H;��H;��H;��H;��H;7�H;��H;!�H;��H;��H;k�H;q�H;k�H;��H;��H;!�H;��H;7�H;��H;��H;��H;��H;��H;5�H;��H;V�H;>�H;c�H;��H;��H;�H;CI;*I;+I;<
I;`I;�I;�I;�I;�I;�I;I;c!I;Q#I;�$I;�%I;�&I;      �$I;�$I;�#I;�"I;G!I;}I;cI;�I;)I;TI;iI;PI;VI;6	I;'I;]I;� I;�H;��H;�H;��H;��H;�H;w�H;�H;��H;w�H;y�H;��H;��H;��H;��H;3�H;��H;�H;q�H;w�H;q�H;�H;��H;3�H;��H;��H;��H;��H;y�H;w�H;��H;�H;w�H;�H;��H;��H;�H;��H;�H;� I;]I;'I;6	I;VI;PI;iI;TI;)I;�I;cI;}I;G!I;�"I;�#I;�$I;      �&I;�&I;�%I;�$I;Q#I;c!I;I;�I;�I;�I;�I;�I;`I;<
I;+I;*I;CI;�H;��H;��H;c�H;>�H;V�H;��H;5�H;��H;��H;��H;��H;��H;7�H;��H;!�H;��H;��H;k�H;q�H;k�H;��H;��H;!�H;��H;7�H;��H;��H;��H;��H;��H;5�H;��H;V�H;>�H;c�H;��H;��H;�H;CI;*I;+I;<
I;`I;�I;�I;�I;�I;�I;I;c!I;Q#I;�$I;�%I;�&I;      �-I;E-I;~,I;+I;X)I;3'I;�$I;�!I;�I;_I;�I;}I;�I;XI;�	I;�I;[I;N I;{�H;��H;��H;f�H;H�H;o�H;��H;e�H;�H;��H;��H;�H;z�H;��H;M�H;��H;��H;��H;�H;��H;��H;��H;M�H;��H;z�H;�H;��H;��H;�H;e�H;��H;o�H;H�H;f�H;��H;��H;{�H;N I;[I;�I;�	I;XI;�I;}I;�I;_I;�I;�!I;�$I;3'I;X)I;+I;~,I;E-I;      �8I;�8I;�7I;A6I;;4I;�1I;|.I;+I;C'I;B#I;I;�I;�I;�I;�I;�
I;�I;�I;O I;F�H;��H;�H;��H;��H;��H;4�H;��H;��H;��H;��H;��H;,�H;��H;<�H;��H;��H;��H;��H;��H;<�H;��H;,�H;��H;��H;��H;��H;��H;4�H;��H;��H;��H;�H;��H;F�H;O I;�I;�I;�
I;�I;�I;�I;�I;I;B#I;C'I;+I;|.I;�1I;;4I;A6I;�7I;�8I;      �JI;\JI;II;GI;hDI;AI;/=I;�8I;4I;/I;�)I;�$I;�I;�I;�I;�I;|I;EI;NI;� I;��H;��H;��H;��H;p�H;��H;��H;��H;K�H;B�H;\�H;��H;�H;��H;M�H;!�H;3�H;!�H;M�H;��H;�H;��H;\�H;B�H;K�H;��H;��H;��H;p�H;��H;��H;��H;��H;� I;NI;EI;|I;�I;�I;�I;�I;�$I;�)I;/I;4I;�8I;/=I;AI;hDI;GI;II;\JI;      ucI;�bI;qaI;�^I;Z[I;�VI;�QI;.LI;!FI;�?I;.9I;r2I;�+I;~%I;KI;cI;�I;�I;�	I;�I;�I;�H;��H;��H;z�H;c�H;`�H;��H;Z�H;�H;�H;U�H;��H;,�H;��H;��H;��H;��H;��H;,�H;��H;U�H;�H;�H;Z�H;��H;`�H;c�H;z�H;��H;��H;�H;�I;�I;�	I;�I;�I;cI;KI;~%I;�+I;r2I;.9I;�?I;!FI;.LI;�QI;�VI;Z[I;�^I;qaI;�bI;      ��I;ąI;��I;�I;]{I;�uI;�nI;%gI;�^I;�VI;�MI;(EI;�<I;G4I;W,I;�$I;�I;CI;GI;�I;�I;�I;��H;A�H;&�H;��H;\�H;a�H;��H;6�H;�H;�H;\�H;��H;z�H;7�H;��H;7�H;z�H;��H;\�H;�H;�H;6�H;��H;a�H;\�H;��H;&�H;A�H;��H;�I;�I;�I;GI;CI;�I;�$I;W,I;G4I;�<I;(EI;�MI;�VI;�^I;%gI;�nI;�uI;]{I;�I;��I;ąI;      H�I;Y�I;��I;)�I;ԦI;�I;֕I;��I;��I;6uI;�iI;�]I;�RI;�GI;=I;�3I;�*I;g"I;�I;�I;�I;VI;�I;>�H;��H;U�H;��H;c�H;[�H;��H;6�H;�H;B�H;��H;�H;��H;��H;��H;�H;��H;B�H;�H;6�H;��H;[�H;c�H;��H;U�H;��H;>�H;�I;VI;�I;�I;�I;g"I;�*I;�3I;=I;�GI;�RI;�]I;�iI;6uI;��I;��I;֕I;�I;ԦI;)�I;��I;Y�I;      ��I;7�I;�I;r�I;��I;��I;��I;K�I;L�I; �I;��I;&I;�oI;zaI;�SI;GI;D;I;�0I;�&I;3I;nI;�I;�	I;II;��H;��H;}�H;��H;X�H;[�H;��H;Z�H;K�H;��H;��H;��H;��H;��H;��H;��H;K�H;Z�H;��H;[�H;X�H;��H;}�H;��H;��H;II;�	I;�I;nI;3I;�&I;�0I;D;I;GI;�SI;zaI;�oI;&I;��I; �I;L�I;K�I;��I;��I;��I;r�I;�I;7�I;      �I;��I;�I;��I;�I;C�I;��I;b�I;!�I;��I;ŽI;&�I;6�I;��I;�pI;�_I;�PI;�BI;>6I;+I;8!I;�I;�I;�
I;�I; I;��H;y�H;��H;c�H;a�H;��H;��H;��H;��H;��H;y�H;��H;��H;��H;��H;��H;a�H;c�H;��H;y�H;��H; I;�I;�
I;�I;�I;8!I;+I;>6I;�BI;�PI;�_I;�pI;��I;6�I;&�I;ŽI;��I;!�I;b�I;��I;C�I;�I;��I;�I;��I;      tI;N&I;:I;�WI;{I;0�I;��I;�I;-�I;,�I;p�I;��I;��I;�I;^�I;$�I;�kI;�YI;}II;6;I;�.I;�#I;7I;I;)I;1I; I;��H;}�H;��H;\�H;`�H;��H;��H;�H;��H;w�H;��H;�H;��H;��H;`�H;\�H;��H;}�H;��H; I;1I;)I;I;7I;�#I;�.I;6;I;}II;�YI;�kI;$�I;^�I;�I;��I;��I;p�I;,�I;-�I;�I;��I;0�I;{I;�WI;:I;N&I;      �F;m�F;�F;�1G;`�G;!%H;|�H;�I;lI;��I;r�I;��I;��I;��I;��I;ȨI;��I;�vI;�aI;BOI;??I;X1I;r%I;DI;�I;OI;1I; I;��H;U�H;��H;c�H;��H;4�H;e�H;��H;��H;��H;e�H;4�H;��H;c�H;��H;U�H;��H; I;1I;OI;�I;DI;r%I;X1I;??I;BOI;�aI;�vI;��I;ȨI;��I;��I;��I;��I;r�I;��I;lI;�I;|�H;!%H;`�G;�1G;�F;m�F;      ��?;��?;��@;�sA;�B;[�C;�AE;t�F;��G;~wH;�I;�I;��I;��I;U�I;��I;+�I;L�I;#�I;-hI;�SI;BI;3I;Y&I;�I;�I;)I;�I;��H;��H;&�H;z�H;p�H;��H;��H;5�H;�H;5�H;��H;��H;p�H;z�H;&�H;��H;��H;�I;)I;�I;�I;Y&I;3I;BI;�SI;-hI;#�I;L�I;+�I;��I;U�I;��I;��I;�I;�I;~wH;��G;t�F;�AE;[�C;�B;�sA;��@;��?;      ��0;�41;!�2;\�4;�/7;5":;/=;�@;�B;�E;��F;g$H;�I;p�I;��I;��I;��I;�I;}�I;�I;�lI;aVI;�CI;�3I;Y&I;DI;I;�
I;II;>�H;A�H;��H;��H;��H;o�H;��H;w�H;��H;o�H;��H;��H;��H;A�H;>�H;II;�
I;I;DI;Y&I;�3I;�CI;aVI;�lI;�I;}�I;�I;��I;��I;��I;p�I;�I;g$H;��F;�E;�B;�@;/=;5":;�/7;\�4;!�2;�41;      _;;W�;��;# ;�&;�[,;�2;.88;�.=;�EA;�qD;r�F;+IH;w8I;I�I;��I;s�I;�I;��I;��I;!oI;bWI;�CI;3I;r%I;7I;�I;�	I;�I;��H;��H;��H;��H;H�H;V�H;�H;V�H;H�H;��H;��H;��H;��H;�I;�	I;�I;7I;r%I;3I;�CI;bWI;!oI;��I;��I;�I;s�I;��I;I�I;w8I;+IH;r�F;�qD;�EA;�.=;.88;�2;�[,;�&;# ;��;W�;;      X��:��:�
�:��:��:�O ;�d;�U;\~#; d-;��5;�g<;nsA;rE;�dG;R�H;N�I;(�I;	�I;0�I;4�I;�I;!oI;aVI;BI;X1I;�#I;�I;�I;VI;�I;�H;��H;�H;f�H;>�H;��H;>�H;f�H;�H;��H;�H;�I;VI;�I;�I;�#I;X1I;BI;aVI;!oI;�I;4�I;0�I;	�I;(�I;N�I;R�H;�dG;rE;nsA;�g<;��5; d-;\~#;�U;�d;�O ;��:��:�
�:��:      e�p� �-��9���9�":��u:��:q��:��:;Q;o ;��,;/�6;j(>;;C;�F;�kH;�jI;��I;��I;��I;4�I;��I;�lI;�SI;??I;�.I;8!I;nI;�I;�I;�I;��H;��H;��H;c�H;��H;c�H;��H;��H;��H;�I;�I;�I;nI;8!I;�.I;??I;�SI;�lI;��I;4�I;��I;��I;��I;�jI;�kH;�F;;C;j(>;/�6;��,;o ;;Q;��:q��:��:��u:�":���9�9 �-�      q&�~!��5���}谺�O��LT��l�9��u:�!�:�E�:C;=~#;}61;P;;��A;�E;�#H;jUI;,�I;��I;0�I;��I;�I;-hI;BOI;6;I;+I;3I;�I;�I;�I;� I;F�H;��H;��H;�H;��H;��H;F�H;� I;�I;�I;�I;3I;+I;6;I;BOI;-hI;�I;��I;0�I;��I;,�I;jUI;�#H;�E;��A;P;;}61;=~#;C;�E�:�!�:��u:�l�9�LT��O�}谺���5�~!�      llٻ�Ի ǻ����W���n� �+�J�Ժ�1��39Ym:��:{�;�;�[,;��8;ք@;V\E;�	H;jUI;��I;	�I;�I;}�I;#�I;�aI;}II;>6I;�&I;�I;GI;�	I;NI;O I;{�H;��H;��H;��H;{�H;O I;NI;�	I;GI;�I;�&I;>6I;}II;�aI;#�I;}�I;�I;	�I;��I;jUI;�	H;V\E;ք@;��8;�[,;�;{�;��:Ym:�39�1�J�Ժ �+��n�W������ ǻ�Ի      �yY�,}U���I���7��� �G"�#�Ի;❻��T�%���#��m�9���:ij�:�;�);)07;D@;V\E;�#H;�jI;(�I;s�I;�I;L�I;�vI;�YI;�BI;�0I;g"I;CI;�I;EI;�I;N I;�H;�H;�H;N I;�I;EI;�I;CI;g"I;�0I;�BI;�YI;�vI;L�I;�I;s�I;(�I;�jI;�#H;V\E;D@;)07;�);�;ij�:���:�m�9�#�%���T�;❻#�ԻG"��� ���7���I�,}U�      "�ü�l������S��cߓ���{�f�M�҉ ����S�����B�$찺��o���u:���:�Q;D�';)07;ք@;�E;�kH;N�I;��I;��I;+�I;��I;�kI;�PI;D;I;�*I;�I;�I;|I;�I;[I;CI;� I;CI;[I;�I;|I;�I;�I;�*I;D;I;�PI;�kI;��I;+�I;��I;��I;N�I;�kH;�E;ք@;)07;D�';�Q;���:��u:��o�$찺��B�S������҉ �f�M���{�cߓ�S�������l��      �'��-$�r��l�,���.?ټ-w��`����yY�-l���Ի���	[������ R:���:�Q;�);��8;��A;�F;R�H;I�I;��I;��I;ȨI;$�I;�_I;GI;�3I;�$I;cI;�I;�
I;�I;*I;]I;*I;�I;�
I;�I;cI;�$I;�3I;GI;�_I;$�I;ȨI;��I;��I;I�I;R�H;�F;��A;��8;�);�Q;���: R:����	[�������Ի-l��yY�`���-w��.?ټ,���l�r���-$�      b+����k̀�?l��Q�8�2�T����7����@����>��2���V���2���� R:���:�;�[,;P;;;C;�dG;w8I;��I;U�I;��I;^�I;�pI;�SI;=I;W,I;KI;�I;�I;�	I;+I;'I;+I;�	I;�I;�I;KI;W,I;=I;�SI;�pI;^�I;��I;U�I;��I;w8I;�dG;;C;P;;�[,;�;���: R:���2��V���2����>��@��7������T�8�2��Q�?l�k̀���      s�ཾhܽw�нfy��h什Y ��-l��n<�`���>ټ�𛼞|U����H᝻�2�������u:ij�:�;}61;j(>;rE;+IH;p�I;��I;��I;�I;��I;zaI;�GI;G4I;~%I;�I;�I;XI;<
I;6	I;<
I;XI;�I;�I;~%I;G4I;�GI;zaI;��I;�I;��I;��I;p�I;+IH;rE;j(>;}61;�;ij�:��u:�����2�H᝻����|U����>ټ`���n<�-l�Y ��h什fy��w�н�hܽ      ��4�j1�	�&������q�ཌྷ�������`��'�-��yR����]�����V��	[����o����:{�;=~#;/�6;nsA;r�F;�I;��I;��I;��I;6�I;�oI;�RI;�<I;�+I;�I;�I;�I;`I;VI;`I;�I;�I;�I;�+I;�<I;�RI;�oI;6�I;��I;��I;��I;�I;r�F;nsA;/�6;=~#;{�;���:��o�	[���V�������]�yR��-��'��`��������q�������	�&�j1�      �x���o��ń�KUo���O�-�-�{��hܽd什�x��2��b��yR���|U��2�����$찺�m�9��:C;��,;�g<;�qD;g$H;�I;��I;��I;&�I;&I;�]I;(EI;r2I;�$I;�I;}I;�I;PI;�I;}I;�I;�$I;r2I;(EI;�]I;&I;&�I;��I;��I;�I;g$H;�qD;�g<;��,;C;��:�m�9$찺����2���|U�yR���b���2��x�d什�hܽ{�-�-���O�KUo�ń��o��      v���ྃ�Ѿ(����נ�	ń�<�S�
�#�gO���n��R̀��2�-������>���Ի��B��#�Ym:�E�:o ;��5;�EA;��F;�I;r�I;p�I;ŽI;��I;�iI;�MI;.9I;�)I;I;�I;�I;iI;�I;�I;I;�)I;.9I;�MI;�iI;��I;ŽI;p�I;r�I;�I;��F;�EA;��5;o ;�E�:Ym:�#���B���Ի��>���-���2�R̀��n��gO��
�#�<�S�	ń��נ�(�����Ѿ��      �3���/��X#��	��A��ՌȾ�f��JUo�`1�Ӱ���n���x��'��>ټ�@��-l�S���%���39�!�:;Q; d-;�.=;�E;~wH;��I;,�I;��I; �I;6uI;�VI;�?I;/I;B#I;_I;�I;TI;�I;_I;B#I;/I;�?I;�VI;6uI; �I;��I;,�I;��I;~wH;�E;�.=; d-;;Q;�!�:�39%��S���-l��@���>ټ�'��x��n��Ӱ��`1�JUo��f��ՌȾ�A���	��X#���/�      ���S���Q�v��RZ�Z58�˂�p��d���hoy�`1�gO��d什�`�`��7����yY���컟�T��1���u:��:\~#;.88;�B;��G;lI;-�I;!�I;L�I;��I;�^I;!FI;4I;C'I;�I;�I;)I;�I;�I;C'I;4I;!FI;�^I;��I;L�I;!�I;-�I;lI;��G;�B;.88;\~#;��:��u:�1���T���컷yY�7���`���`�d什gO��`1�hoy�d���p��˂�Z58��RZ�Q�v�S���      Ŀ3g��$ﱿ���R����U��X#�r��d���JUo�
�#��hܽ����n<����`���҉ �;❻J�Ժ�l�9q��:�U;�2;�@;t�F;�I;�I;b�I;K�I;��I;%gI;.LI;�8I;+I;�!I;�I;�I;�I;�!I;+I;�8I;.LI;%gI;��I;K�I;b�I;�I;�I;t�F;�@;�2;�U;q��:�l�9J�Ժ;❻҉ �`�������n<�����hܽ
�#�JUo�d���r���X#��U�R������$ﱿ3g��      |x�N9�M��pؿkQ��c_��4�_��X#�p���f��<�S�{�����-l�T�-w��f�M�#�Ի �+��LT���:�d;�[,;/=;�AE;|�H;��I;��I;��I;֕I;�nI;�QI;/=I;|.I;�$I;I;cI;I;�$I;|.I;/=I;�QI;�nI;֕I;��I;��I;��I;|�H;�AE;/=;�[,;�d;��:�LT� �+�#�Իf�M�-w��T�-l�����{�<�S��f��p���X#�4�_�c_��kQ��pؿM��N9�      �X1���,�e���<���2g��c_���U�˂�ՌȾ	ń�-�-�q��Y ��8�2�.?ټ��{�G"��n��O���u:�O ;�&;5":;[�C;!%H;0�I;C�I;��I;�I;�uI;�VI;AI;�1I;3'I;c!I;}I;c!I;3'I;�1I;AI;�VI;�uI;�I;��I;C�I;0�I;!%H;[�C;5":;�&;�O ;��u:�O��n�G"���{�.?ټ8�2�Y ��q��-�-�	ń�ՌȾ˂��U�c_��2g���<�e����,�      d��]]�1K��X1�Xf���kQ��R���Z58��A���נ���O���h什�Q�,���cߓ��� �W��}谺�":��:# ;�/7;�B;`�G;{I;�I;��I;ԦI;]{I;Z[I;hDI;;4I;X)I;Q#I;G!I;Q#I;X)I;;4I;hDI;Z[I;]{I;ԦI;��I;�I;{I;`�G;�B;�/7;# ;��:�":}谺W���� �cߓ�,����Q�h什����O��נ��A��Z58�R���kQ����Xf��X1�1K��]]�      L������4z���V��X1��<�pؿ����RZ��	�(���KUo����fy��?l�l�S����7������𺢽�9��:��;\�4;�sA;�1G;�WI;��I;r�I;)�I;�I;�^I;GI;A6I;+I;�$I;�"I;�$I;+I;A6I;GI;�^I;�I;)�I;r�I;��I;�WI;�1G;�sA;\�4;��;��:���9�𺙼����7�S��l�?l�fy�����KUo�(����	��RZ����pؿ�<��X1���V��4z�����      �o��c^���ē��4z�1K�e��M��$ﱿQ�v��X#���Ѿń�	�&�w�нk̀�r��������I� ǻ�5��9�
�:W�;!�2;��@;�F;:I;�I;�I;��I;��I;qaI;II;�7I;~,I;�%I;�#I;�%I;~,I;�7I;II;qaI;��I;��I;�I;�I;:I;�F;��@;!�2;W�;�
�:�9�5� ǻ��I�����r��k̀�w�н	�&�ń���Ѿ�X#�Q�v�$ﱿM��e��1K��4z��ē�c^��      o'���X��c^�������]]���,�N9�3g��S�����/����o��j1��hܽ���-$��l��,}U��Ի~!� �-���:;�41;��?;m�F;N&I;��I;7�I;Y�I;ąI;�bI;\JI;�8I;E-I;�&I;�$I;�&I;E-I;�8I;\JI;�bI;ąI;Y�I;7�I;��I;N&I;m�F;��?;�41;;��: �-�~!��Ի,}U��l���-$����hܽj1��o���྘�/�S���3g��N9���,��]]�����c^���X��      j����������΢��+�j��5���	���ȿ%8����7�D�꾂S���7�3但L��-�)��ƼE�\���ݻ�+�4wɸ��:>w;��0;��?;}�F;+I;��I;�I;�I;H�I;�gI;NI;�;I;�/I;�(I;�&I;�(I;�/I;�;I;NI;�gI;H�I;�I;�I;��I;+I;}�F;��?;��0;>w;��:4wɸ�+���ݻE�\��Ƽ-�)��L��3��7��S��D�꾧�7�%8����ȿ��	��5�+�j�΢����������      ��������B��Z�����c�321�#X��ÿhڇ�q�3��s��7��74�i�Gى���&�-Nür�X�>�ػ��%���J�ρ�:�a;z�0;��?;8�F;�1I;�I;c�I;
�I;m�I;xgI;�MI;R;I;�/I;~(I;�&I;~(I;�/I;R;I;�MI;xgI;m�I;
�I;c�I;�I;�1I;8�F;��?;z�0;�a;ρ�:��J���%�>�ػr�X�-Nü��&�Gى�i�74��7���s�q�3�hڇ��ÿ#X�321���c�Z����B�����      �����B����C��s�P���#�I�������x|��'�YD־�X��s�)�&Խ�Ă�\<�]_���-M�j ˻^��	�8Б�:�;J2;/u@;��F;�EI;��I;+�I;F�I;%�I;�eI;YLI;c:I;�.I;�'I;�%I;�'I;�.I;c:I;YLI;�eI;%�I;F�I;+�I;��I;�EI;��F;/u@;J2;�;Б�:	�8^��j ˻�-M�]_��\<��Ă�&Խs�)��X��YD־�'��x|����I�����#�s�P�C�����B��      ΢��Z���C���/]��5�L���,ݿ)8��nm_��K��t��Y�s�'>�����J�o��3��۩��:��T�������9�d�:�;;�^4;&gA;:7G;�cI;%�I;P�I;w�I;��I;KcI;7JI;�8I;m-I;�&I;�$I;�&I;m-I;�8I;7JI;KcI;��I;w�I;P�I;%�I;�cI;:7G;&gA;�^4;�;;�d�:��9����T���:��۩��3�J�o�����'>�Y�s��t���K�nm_�)8���,ݿL���5��/]�C��Z���      +�j���c�s�P��5���o��E���gڇ�Dv<�&���q���_S��������+T��� �P$��+H#�W���p3����:ǯ�:Q�;67;��B;��G;׆I;6�I;��I;�I;��I;�_I;fGI;�6I;�+I;*%I;#I;*%I;�+I;�6I;fGI;�_I;��I;�I;��I;6�I;׆I;��G;��B;67;Q�;ǯ�:��:p3��W���+H#�P$���� �+T���������_S�q��&���Dv<�gڇ�E���o�����5�s�P���c�      �5�321���#�L��o���ÿ�ҕ�Z������̾�X����0�3�8W����5��zܼ������l�s��Y\�]�n:���:��%;��9;��C;.H;1�I;1�I;%�I;��I;�zI;-[I;�CI;�3I;L)I;8#I;8!I;8#I;L)I;�3I;�CI;-[I;�zI;��I;%�I;1�I;1�I;.H;��C;��9;��%;���:]�n:�Y\�l�s��������zܼ��5�8W��3佃�0��X����̾���Z��ҕ��ÿo��L����#�321�      ��	�#X�I����,ݿE����ҕ� �d��'�?��#���{�W����t���C�o��G��*���Q�'�ػ�0�4�~���:��;N,;q=;WAE;��H;��I;��I;h�I;�I;�sI;�UI;�?I;�0I;�&I;� I;�I;� I;�&I;�0I;�?I;�UI;�sI;�I;h�I;��I;��I;��H;WAE;q=;N,;��;��:4�~��0�'�ػ�Q��*���G�C�o�t������{�W�#���?�꾊'� �d��ҕ�E����,ݿI���#X�      ��ȿ�ÿ���)8��gڇ�Z��'�����l8��Y�s�0�&�`�9{??�W�A琼�G#��7���Vܺ��9U�:��;8K2;c@;��F;I;��I;��I;p�I;d�I;�kI;�OI;u;I;-I;�#I;CI;dI;CI;�#I;-I;u;I;�OI;�kI;d�I;p�I;��I;��I;I;��F;c@;8K2;��;U�:��9�Vܺ�7���G#�A琼W�{??�9`�0�&�Y�s�l8�������'�Z�gڇ�)8������ÿ      %8��hڇ��x|�nm_�Dv<����?��l8��'6~�r74��l������Inc�G��_��2�\�A:�UZ�� >���n:[��:#;�8;ܿB;��G;�wI;��I;��I;��I;��I;ZcI;�II;�6I;5)I;W I;lI;�I;lI;W I;5)I;�6I;�II;ZcI;��I;��I;��I;��I;�wI;��G;ܿB;�8;#;[��:��n:� >�UZ�A:�2�\�_��G��Inc������l��r74�'6~�l8��?�꾎��Dv<�nm_��x|�hڇ�      ��7�q�3��'��K�&�����̾#���Y�s�r74����*N���|��)�^zܼZ��� � ��P���D9ꇹ:-�;-;%=;�E;!�H;o�I;M�I;��I;ǤI;<zI;�ZI;�BI;q1I;2%I;�I;II;�I;II;�I;2%I;q1I;�BI;�ZI;<zI;ǤI;��I;M�I;o�I;!�H;�E;%=;-;-�;ꇹ:D9P��� ��� �Z��^zܼ�)��|�*N�����r74�Y�s�#�����̾&����K��'�q�3�      D���s�YD־�t��q���X��{�W�0�&��l��*N���Ă�|�5�׃���Q��#�A���ػ��G�!&/�8f:`�:Õ;x�5;�8A;]�F;�)I;��I;��I;+�I;}�I;QnI;�QI;�;I;4,I;� I;aI;I;�I;I;aI;� I;4,I;�;I;�QI;QnI;}�I;+�I;��I;��I;�)I;]�F;�8A;x�5;Õ;`�:8f:!&/���G���ػ#�A��Q��׃��|�5��Ă�*N���l��0�&�{�W��X��q���t��YD־�s�      �S���7���X��Y�s��_S���0����`ང����|�|�5����۩��X�fc �����5����9"��:��;�,;�K<;vnD;'-H;�I;��I;��I;u�I;q�I;ZbI;|HI;�4I;�&I;eI;�I;�I;�I;�I;�I;eI;�&I;�4I;|HI;ZbI;q�I;u�I;��I;��I;�I;'-H;vnD;�K<;�,;��;"��:��9�5�����fc ��X�۩����|�5��|�����`ས����0��_S�Y�s��X���7��      �7�74�s�)�'>����3�t���9Inc��)�׃��۩��a�2R�ݒ��%O�v�ȸ%��:��;�#;��6;gA;��F;�I;Y�I;��I;0�I;��I;�tI;�VI;�?I;%.I;|!I;2I;I;�I;xI;�I;I;2I;|!I;%.I;�?I;�VI;�tI;��I;0�I;��I;Y�I;�I;��F;gA;��6;�#;��;%��:v�ȸ%O�ݒ��2R��a�۩�׃���)�Inc�9t���3����'>�s�)�74�      3�i�&Խ��������8W��C�o�{??�G��^zܼ�Q���X�2R�/7�������Ϲ��n:�k�:!=;��0;�>;KE;rRH;d�I;��I;�I;[�I;y�I;�eI;DKI;�6I;'I;$I;I;{I;8I;Y
I;8I;{I;I;$I;'I;�6I;DKI;�eI;y�I;[�I;�I;��I;d�I;rRH;KE;�>;��0;!=;�k�:��n:��Ϲ���/7��2R��X��Q��^zܼG��{??�C�o�8W����������&Խi�      �L��Gى��Ă�J�o�+T���5��G�W�_��Z��#�A�fc �ݒ��������8�J:tj�:�d;3,;��:;"4C;+kG;DI;�I;��I;��I;��I;�uI;�WI;b@I;�.I;,!I;�I;�I;�
I;I;eI;I;�
I;�I;�I;,!I;�.I;b@I;�WI;�uI;��I;��I;��I;�I;DI;+kG;"4C;��:;3,;�d;tj�:8�J:������ݒ��fc �#�A�Z��_��W��G���5�+T�J�o��Ă�Gى�      -�)���&�\<��3��� ��zܼ�*��A琼2�\�� ���ػ���%O���Ϲ8�J:yh�:v�;��(;�d8;��A;*�F;��H;=�I;��I;!�I;�I;}�I;zdI;�JI;36I;�&I;I;&I;�I;{I;�I;@I;�I;{I;�I;&I;I;�&I;36I;�JI;zdI;}�I;�I;!�I;��I;=�I;��H;*�F;��A;�d8;��(;v�;yh�:8�J:��Ϲ%O������ػ� �2�\�A琼�*���zܼ�� ��3�\<���&�      �Ƽ-Nü]_���۩�P$������Q��G#�A:� ����G��5��v�ȸ��n:tj�:v�;*�';�7;�u@;<�E;.uH;�I;��I;��I;]�I;��I;�pI;�TI;I>I;�,I;�I;,I;�I;�I;YI;I;7I;I;YI;�I;�I;,I;�I;�,I;I>I;�TI;�pI;��I;]�I;��I;��I;�I;.uH;<�E;�u@;�7;*�';v�;tj�:��n:v�ȸ�5����G� ��A:�G#��Q����P$���۩�]_��-Nü      E�\�r�X��-M��:�+H#����'�ػ�7��UZ�P���!&/���9%��:�k�:�d;��(;�7;�@;;\E;�,H;OvI;��I;��I;��I;ܡI;�{I;�]I;�EI;3I;b$I;�I;�I;[	I;UI;7I;@�H;��H;@�H;7I;UI;[	I;�I;�I;b$I;3I;�EI;�]I;�{I;ܡI;��I;��I;��I;OvI;�,H;;\E;�@;�7;��(;�d;�k�:%��:��9!&/�P���UZ��7��'�ػ���+H#��:��-M�r�X�      ��ݻ>�ػj ˻�T��W���l�s��0��Vܺ� >�D98f:"��:��;!=;3,;�d8;�u@;;\E;IH;aI;*�I;��I;X�I;��I;y�I;fI;MI;�8I;)I;~I;�I;I;II;I;Y�H;��H;��H;��H;Y�H;I;II;I;�I;~I;)I;�8I;MI;fI;y�I;��I;X�I;��I;*�I;aI;IH;;\E;�u@;�d8;3,;!=;��;"��:8f:D9� >��Vܺ�0�l�s�W����T��j ˻>�ػ      �+���%�^�����p3���Y\�4�~���9��n:ꇹ:`�:��;�#;��0;��:;��A;<�E;�,H;aI;��I;��I;��I;!�I;͌I;�lI;SI; >I;I-I;�I;kI;I;tI;�I;�H;��H;�H;��H;�H;��H;�H;�I;tI;I;kI;�I;I-I; >I;SI;�lI;͌I;!�I;��I;��I;��I;aI;�,H;<�E;��A;��:;��0;�#;��;`�:ꇹ:��n:��94�~��Y\�p3�����^����%�      4wɸ��J�	�8��9��:]�n:��:U�:[��:-�;Õ;�,;��6;�>;"4C;*�F;.uH;OvI;*�I;��I;O�I;޷I;n�I;�qI;�WI;JBI;1I;<#I;�I;�I;�I;XI;Q�H;@�H;��H;��H;��H;��H;��H;@�H;Q�H;XI;�I;�I;�I;<#I;1I;JBI;�WI;�qI;n�I;޷I;O�I;��I;*�I;OvI;.uH;*�F;"4C;�>;��6;�,;Õ;-�;[��:U�:��:]�n:��:��9	�8��J�      ��:ρ�:Б�:�d�:ǯ�:���:��;��;#;-;x�5;�K<;gA;KE;+kG;��H;�I;��I;��I;��I;޷I;	�I;tI;�ZI;gEI;�3I;�%I;FI;�I;b	I;~I;��H;�H;��H;��H;��H;x�H;��H;��H;��H;�H;��H;~I;b	I;�I;FI;�%I;�3I;gEI;�ZI;tI;	�I;޷I;��I;��I;��I;�I;��H;+kG;KE;gA;�K<;x�5;-;#;��;��;���:ǯ�:�d�:Б�:ρ�:      >w;�a;�;�;;Q�;��%;N,;8K2;�8;%=;�8A;vnD;��F;rRH;DI;=�I;��I;��I;X�I;!�I;n�I;tI;u[I;�FI;�5I;�'I;�I;TI;�
I;]I;V�H;��H;]�H;�H;��H;��H;��H;��H;��H;�H;]�H;��H;V�H;]I;�
I;TI;�I;�'I;�5I;�FI;u[I;tI;n�I;!�I;X�I;��I;��I;=�I;DI;rRH;��F;vnD;�8A;%=;�8;8K2;N,;��%;Q�;�;;�;�a;      ��0;z�0;J2;�^4;67;��9;q=;c@;ܿB;�E;]�F;'-H;�I;d�I;�I;��I;��I;��I;��I;͌I;�qI;�ZI;�FI;36I;�(I;I;hI;�I;@I;��H;��H;��H;
�H; �H;��H;�H;��H;�H;��H; �H;
�H;��H;��H;��H;@I;�I;hI;I;�(I;36I;�FI;�ZI;�qI;͌I;��I;��I;��I;��I;�I;d�I;�I;'-H;]�F;�E;ܿB;c@;q=;��9;67;�^4;J2;z�0;      ��?;��?;/u@;&gA;��B;��C;WAE;��F;��G;!�H;�)I;�I;Y�I;��I;��I;!�I;]�I;ܡI;y�I;�lI;�WI;gEI;�5I;�(I;qI;�I;HI;�I;� I;D�H;��H;��H;��H;7�H;�H;v�H;=�H;v�H;�H;7�H;��H;��H;��H;D�H;� I;�I;HI;�I;qI;�(I;�5I;gEI;�WI;�lI;y�I;ܡI;]�I;!�I;��I;��I;Y�I;�I;�)I;!�H;��G;��F;WAE;��C;��B;&gA;/u@;��?;      }�F;8�F;��F;:7G;��G;.H;��H;I;�wI;o�I;��I;��I;��I;�I;��I;�I;��I;�{I;fI;SI;JBI;�3I;�'I;I;�I;�I;CI;� I;{�H;��H;�H;��H;��H;��H;��H; �H;��H; �H;��H;��H;��H;��H;�H;��H;{�H;� I;CI;�I;�I;I;�'I;�3I;JBI;SI;fI;�{I;��I;�I;��I;�I;��I;��I;��I;o�I;�wI;I;��H;.H;��G;:7G;��F;8�F;      +I;�1I;�EI;�cI;׆I;1�I;��I;��I;��I;M�I;��I;��I;0�I;[�I;��I;}�I;�pI;�]I;MI; >I;1I;�%I;�I;hI;HI;CI;� I;��H;�H;	�H;��H;��H;E�H;(�H;3�H;��H;��H;��H;3�H;(�H;E�H;��H;��H;	�H;�H;��H;� I;CI;HI;hI;�I;�%I;1I; >I;MI;�]I;�pI;}�I;��I;[�I;0�I;��I;��I;M�I;��I;��I;��I;1�I;׆I;�cI;�EI;�1I;      ��I;�I;��I;%�I;6�I;1�I;��I;��I;��I;��I;+�I;u�I;��I;y�I;�uI;zdI;�TI;�EI;�8I;I-I;<#I;FI;TI;�I;�I;� I;��H;?�H;'�H;��H;��H;�H;��H;��H;(�H;��H;��H;��H;(�H;��H;��H;�H;��H;��H;'�H;?�H;��H;� I;�I;�I;TI;FI;<#I;I-I;�8I;�EI;�TI;zdI;�uI;y�I;��I;u�I;+�I;��I;��I;��I;��I;1�I;6�I;%�I;��I;�I;      �I;c�I;+�I;P�I;��I;%�I;h�I;p�I;��I;ǤI;}�I;q�I;�tI;�eI;�WI;�JI;I>I;3I;)I;�I;�I;�I;�
I;@I;� I;{�H;�H;'�H;��H;��H;��H;��H;[�H;��H;A�H;��H;��H;��H;A�H;��H;[�H;��H;��H;��H;��H;'�H;�H;{�H;� I;@I;�
I;�I;�I;�I;)I;3I;I>I;�JI;�WI;�eI;�tI;q�I;}�I;ǤI;��I;p�I;h�I;%�I;��I;P�I;+�I;c�I;      �I;
�I;F�I;w�I;�I;��I;�I;d�I;��I;<zI;QnI;ZbI;�VI;DKI;b@I;36I;�,I;b$I;~I;kI;�I;b	I;]I;��H;D�H;��H;	�H;��H;��H;��H;��H;O�H;e�H;��H;'�H;��H;��H;��H;'�H;��H;e�H;O�H;��H;��H;��H;��H;	�H;��H;D�H;��H;]I;b	I;�I;kI;~I;b$I;�,I;36I;b@I;DKI;�VI;ZbI;QnI;<zI;��I;d�I;�I;��I;�I;w�I;F�I;
�I;      H�I;m�I;%�I;��I;��I;�zI;�sI;�kI;ZcI;�ZI;�QI;|HI;�?I;�6I;�.I;�&I;�I;�I;�I;I;�I;~I;V�H;��H;��H;�H;��H;��H;��H;��H;C�H;>�H;��H;��H;p�H;N�H;5�H;N�H;p�H;��H;��H;>�H;C�H;��H;��H;��H;��H;�H;��H;��H;V�H;~I;�I;I;�I;�I;�I;�&I;�.I;�6I;�?I;|HI;�QI;�ZI;ZcI;�kI;�sI;�zI;��I;��I;%�I;m�I;      �gI;xgI;�eI;KcI;�_I;-[I;�UI;�OI;�II;�BI;�;I;�4I;%.I;'I;,!I;I;,I;�I;I;tI;XI;��H;��H;��H;��H;��H;��H;�H;��H;O�H;>�H;��H;��H;8�H;��H;��H;��H;��H;��H;8�H;��H;��H;>�H;O�H;��H;�H;��H;��H;��H;��H;��H;��H;XI;tI;I;�I;,I;I;,!I;'I;%.I;�4I;�;I;�BI;�II;�OI;�UI;-[I;�_I;KcI;�eI;xgI;      NI;�MI;YLI;7JI;fGI;�CI;�?I;u;I;�6I;q1I;4,I;�&I;|!I;$I;�I;&I;�I;[	I;II;�I;Q�H;�H;]�H;
�H;��H;��H;E�H;��H;[�H;e�H;��H;��H;�H;��H;{�H;;�H;2�H;;�H;{�H;��H;�H;��H;��H;e�H;[�H;��H;E�H;��H;��H;
�H;]�H;�H;Q�H;�I;II;[	I;�I;&I;�I;$I;|!I;�&I;4,I;q1I;�6I;u;I;�?I;�CI;fGI;7JI;YLI;�MI;      �;I;R;I;c:I;�8I;�6I;�3I;�0I;-I;5)I;2%I;� I;eI;2I;I;�I;�I;�I;UI;I;�H;@�H;��H;�H; �H;7�H;��H;(�H;��H;��H;��H;��H;8�H;��H;W�H;�H;��H;��H;��H;�H;W�H;��H;8�H;��H;��H;��H;��H;(�H;��H;7�H; �H;�H;��H;@�H;�H;I;UI;�I;�I;�I;I;2I;eI;� I;2%I;5)I;-I;�0I;�3I;�6I;�8I;c:I;R;I;      �/I;�/I;�.I;m-I;�+I;L)I;�&I;�#I;W I;�I;aI;�I;I;{I;�
I;{I;YI;7I;Y�H;��H;��H;��H;��H;��H;�H;��H;3�H;(�H;A�H;'�H;p�H;��H;{�H;�H;��H;��H;��H;��H;��H;�H;{�H;��H;p�H;'�H;A�H;(�H;3�H;��H;�H;��H;��H;��H;��H;��H;Y�H;7I;YI;{I;�
I;{I;I;�I;aI;�I;W I;�#I;�&I;L)I;�+I;m-I;�.I;�/I;      �(I;~(I;�'I;�&I;*%I;8#I;� I;CI;lI;II;I;�I;�I;8I;I;�I;I;@�H;��H;�H;��H;��H;��H;�H;v�H; �H;��H;��H;��H;��H;N�H;��H;;�H;��H;��H;o�H;i�H;o�H;��H;��H;;�H;��H;N�H;��H;��H;��H;��H; �H;v�H;�H;��H;��H;��H;�H;��H;@�H;I;�I;I;8I;�I;�I;I;II;lI;CI;� I;8#I;*%I;�&I;�'I;~(I;      �&I;�&I;�%I;�$I;#I;8!I;�I;dI;�I;�I;�I;�I;xI;Y
I;eI;@I;7I;��H;��H;��H;��H;x�H;��H;��H;=�H;��H;��H;��H;��H;��H;5�H;��H;2�H;��H;��H;i�H;L�H;i�H;��H;��H;2�H;��H;5�H;��H;��H;��H;��H;��H;=�H;��H;��H;x�H;��H;��H;��H;��H;7I;@I;eI;Y
I;xI;�I;�I;�I;�I;dI;�I;8!I;#I;�$I;�%I;�&I;      �(I;~(I;�'I;�&I;*%I;8#I;� I;CI;lI;II;I;�I;�I;8I;I;�I;I;@�H;��H;�H;��H;��H;��H;�H;v�H; �H;��H;��H;��H;��H;N�H;��H;;�H;��H;��H;o�H;i�H;o�H;��H;��H;;�H;��H;N�H;��H;��H;��H;��H; �H;v�H;�H;��H;��H;��H;�H;��H;@�H;I;�I;I;8I;�I;�I;I;II;lI;CI;� I;8#I;*%I;�&I;�'I;~(I;      �/I;�/I;�.I;m-I;�+I;L)I;�&I;�#I;W I;�I;aI;�I;I;{I;�
I;{I;YI;7I;Y�H;��H;��H;��H;��H;��H;�H;��H;3�H;(�H;A�H;'�H;p�H;��H;{�H;�H;��H;��H;��H;��H;��H;�H;{�H;��H;p�H;'�H;A�H;(�H;3�H;��H;�H;��H;��H;��H;��H;��H;Y�H;7I;YI;{I;�
I;{I;I;�I;aI;�I;W I;�#I;�&I;L)I;�+I;m-I;�.I;�/I;      �;I;R;I;c:I;�8I;�6I;�3I;�0I;-I;5)I;2%I;� I;eI;2I;I;�I;�I;�I;UI;I;�H;@�H;��H;�H; �H;7�H;��H;(�H;��H;��H;��H;��H;8�H;��H;W�H;�H;��H;��H;��H;�H;W�H;��H;8�H;��H;��H;��H;��H;(�H;��H;7�H; �H;�H;��H;@�H;�H;I;UI;�I;�I;�I;I;2I;eI;� I;2%I;5)I;-I;�0I;�3I;�6I;�8I;c:I;R;I;      NI;�MI;YLI;7JI;fGI;�CI;�?I;u;I;�6I;q1I;4,I;�&I;|!I;$I;�I;&I;�I;[	I;II;�I;Q�H;�H;]�H;
�H;��H;��H;E�H;��H;[�H;e�H;��H;��H;�H;��H;{�H;;�H;2�H;;�H;{�H;��H;�H;��H;��H;e�H;[�H;��H;E�H;��H;��H;
�H;]�H;�H;Q�H;�I;II;[	I;�I;&I;�I;$I;|!I;�&I;4,I;q1I;�6I;u;I;�?I;�CI;fGI;7JI;YLI;�MI;      �gI;xgI;�eI;KcI;�_I;-[I;�UI;�OI;�II;�BI;�;I;�4I;%.I;'I;,!I;I;,I;�I;I;tI;XI;��H;��H;��H;��H;��H;��H;�H;��H;O�H;>�H;��H;��H;8�H;��H;��H;��H;��H;��H;8�H;��H;��H;>�H;O�H;��H;�H;��H;��H;��H;��H;��H;��H;XI;tI;I;�I;,I;I;,!I;'I;%.I;�4I;�;I;�BI;�II;�OI;�UI;-[I;�_I;KcI;�eI;xgI;      H�I;m�I;%�I;��I;��I;�zI;�sI;�kI;ZcI;�ZI;�QI;|HI;�?I;�6I;�.I;�&I;�I;�I;�I;I;�I;~I;V�H;��H;��H;�H;��H;��H;��H;��H;C�H;>�H;��H;��H;p�H;N�H;5�H;N�H;p�H;��H;��H;>�H;C�H;��H;��H;��H;��H;�H;��H;��H;V�H;~I;�I;I;�I;�I;�I;�&I;�.I;�6I;�?I;|HI;�QI;�ZI;ZcI;�kI;�sI;�zI;��I;��I;%�I;m�I;      �I;
�I;F�I;w�I;�I;��I;�I;d�I;��I;<zI;QnI;ZbI;�VI;DKI;b@I;36I;�,I;b$I;~I;kI;�I;b	I;]I;��H;D�H;��H;	�H;��H;��H;��H;��H;O�H;e�H;��H;'�H;��H;��H;��H;'�H;��H;e�H;O�H;��H;��H;��H;��H;	�H;��H;D�H;��H;]I;b	I;�I;kI;~I;b$I;�,I;36I;b@I;DKI;�VI;ZbI;QnI;<zI;��I;d�I;�I;��I;�I;w�I;F�I;
�I;      �I;c�I;+�I;P�I;��I;%�I;h�I;p�I;��I;ǤI;}�I;q�I;�tI;�eI;�WI;�JI;I>I;3I;)I;�I;�I;�I;�
I;@I;� I;{�H;�H;'�H;��H;��H;��H;��H;[�H;��H;A�H;��H;��H;��H;A�H;��H;[�H;��H;��H;��H;��H;'�H;�H;{�H;� I;@I;�
I;�I;�I;�I;)I;3I;I>I;�JI;�WI;�eI;�tI;q�I;}�I;ǤI;��I;p�I;h�I;%�I;��I;P�I;+�I;c�I;      ��I;�I;��I;%�I;6�I;1�I;��I;��I;��I;��I;+�I;u�I;��I;y�I;�uI;zdI;�TI;�EI;�8I;I-I;<#I;FI;TI;�I;�I;� I;��H;?�H;'�H;��H;��H;�H;��H;��H;(�H;��H;��H;��H;(�H;��H;��H;�H;��H;��H;'�H;?�H;��H;� I;�I;�I;TI;FI;<#I;I-I;�8I;�EI;�TI;zdI;�uI;y�I;��I;u�I;+�I;��I;��I;��I;��I;1�I;6�I;%�I;��I;�I;      +I;�1I;�EI;�cI;׆I;1�I;��I;��I;��I;M�I;��I;��I;0�I;[�I;��I;}�I;�pI;�]I;MI; >I;1I;�%I;�I;hI;HI;CI;� I;��H;�H;	�H;��H;��H;E�H;(�H;3�H;��H;��H;��H;3�H;(�H;E�H;��H;��H;	�H;�H;��H;� I;CI;HI;hI;�I;�%I;1I; >I;MI;�]I;�pI;}�I;��I;[�I;0�I;��I;��I;M�I;��I;��I;��I;1�I;׆I;�cI;�EI;�1I;      }�F;8�F;��F;:7G;��G;.H;��H;I;�wI;o�I;��I;��I;��I;�I;��I;�I;��I;�{I;fI;SI;JBI;�3I;�'I;I;�I;�I;CI;� I;{�H;��H;�H;��H;��H;��H;��H; �H;��H; �H;��H;��H;��H;��H;�H;��H;{�H;� I;CI;�I;�I;I;�'I;�3I;JBI;SI;fI;�{I;��I;�I;��I;�I;��I;��I;��I;o�I;�wI;I;��H;.H;��G;:7G;��F;8�F;      ��?;��?;/u@;&gA;��B;��C;WAE;��F;��G;!�H;�)I;�I;Y�I;��I;��I;!�I;]�I;ܡI;y�I;�lI;�WI;gEI;�5I;�(I;qI;�I;HI;�I;� I;D�H;��H;��H;��H;7�H;�H;v�H;=�H;v�H;�H;7�H;��H;��H;��H;D�H;� I;�I;HI;�I;qI;�(I;�5I;gEI;�WI;�lI;y�I;ܡI;]�I;!�I;��I;��I;Y�I;�I;�)I;!�H;��G;��F;WAE;��C;��B;&gA;/u@;��?;      ��0;z�0;J2;�^4;67;��9;q=;c@;ܿB;�E;]�F;'-H;�I;d�I;�I;��I;��I;��I;��I;͌I;�qI;�ZI;�FI;36I;�(I;I;hI;�I;@I;��H;��H;��H;
�H; �H;��H;�H;��H;�H;��H; �H;
�H;��H;��H;��H;@I;�I;hI;I;�(I;36I;�FI;�ZI;�qI;͌I;��I;��I;��I;��I;�I;d�I;�I;'-H;]�F;�E;ܿB;c@;q=;��9;67;�^4;J2;z�0;      >w;�a;�;�;;Q�;��%;N,;8K2;�8;%=;�8A;vnD;��F;rRH;DI;=�I;��I;��I;X�I;!�I;n�I;tI;u[I;�FI;�5I;�'I;�I;TI;�
I;]I;V�H;��H;]�H;�H;��H;��H;��H;��H;��H;�H;]�H;��H;V�H;]I;�
I;TI;�I;�'I;�5I;�FI;u[I;tI;n�I;!�I;X�I;��I;��I;=�I;DI;rRH;��F;vnD;�8A;%=;�8;8K2;N,;��%;Q�;�;;�;�a;      ��:ρ�:Б�:�d�:ǯ�:���:��;��;#;-;x�5;�K<;gA;KE;+kG;��H;�I;��I;��I;��I;޷I;	�I;tI;�ZI;gEI;�3I;�%I;FI;�I;b	I;~I;��H;�H;��H;��H;��H;x�H;��H;��H;��H;�H;��H;~I;b	I;�I;FI;�%I;�3I;gEI;�ZI;tI;	�I;޷I;��I;��I;��I;�I;��H;+kG;KE;gA;�K<;x�5;-;#;��;��;���:ǯ�:�d�:Б�:ρ�:      4wɸ��J�	�8��9��:]�n:��:U�:[��:-�;Õ;�,;��6;�>;"4C;*�F;.uH;OvI;*�I;��I;O�I;޷I;n�I;�qI;�WI;JBI;1I;<#I;�I;�I;�I;XI;Q�H;@�H;��H;��H;��H;��H;��H;@�H;Q�H;XI;�I;�I;�I;<#I;1I;JBI;�WI;�qI;n�I;޷I;O�I;��I;*�I;OvI;.uH;*�F;"4C;�>;��6;�,;Õ;-�;[��:U�:��:]�n:��:��9	�8��J�      �+���%�^�����p3���Y\�4�~���9��n:ꇹ:`�:��;�#;��0;��:;��A;<�E;�,H;aI;��I;��I;��I;!�I;͌I;�lI;SI; >I;I-I;�I;kI;I;tI;�I;�H;��H;�H;��H;�H;��H;�H;�I;tI;I;kI;�I;I-I; >I;SI;�lI;͌I;!�I;��I;��I;��I;aI;�,H;<�E;��A;��:;��0;�#;��;`�:ꇹ:��n:��94�~��Y\�p3�����^����%�      ��ݻ>�ػj ˻�T��W���l�s��0��Vܺ� >�D98f:"��:��;!=;3,;�d8;�u@;;\E;IH;aI;*�I;��I;X�I;��I;y�I;fI;MI;�8I;)I;~I;�I;I;II;I;Y�H;��H;��H;��H;Y�H;I;II;I;�I;~I;)I;�8I;MI;fI;y�I;��I;X�I;��I;*�I;aI;IH;;\E;�u@;�d8;3,;!=;��;"��:8f:D9� >��Vܺ�0�l�s�W����T��j ˻>�ػ      E�\�r�X��-M��:�+H#����'�ػ�7��UZ�P���!&/���9%��:�k�:�d;��(;�7;�@;;\E;�,H;OvI;��I;��I;��I;ܡI;�{I;�]I;�EI;3I;b$I;�I;�I;[	I;UI;7I;@�H;��H;@�H;7I;UI;[	I;�I;�I;b$I;3I;�EI;�]I;�{I;ܡI;��I;��I;��I;OvI;�,H;;\E;�@;�7;��(;�d;�k�:%��:��9!&/�P���UZ��7��'�ػ���+H#��:��-M�r�X�      �Ƽ-Nü]_���۩�P$������Q��G#�A:� ����G��5��v�ȸ��n:tj�:v�;*�';�7;�u@;<�E;.uH;�I;��I;��I;]�I;��I;�pI;�TI;I>I;�,I;�I;,I;�I;�I;YI;I;7I;I;YI;�I;�I;,I;�I;�,I;I>I;�TI;�pI;��I;]�I;��I;��I;�I;.uH;<�E;�u@;�7;*�';v�;tj�:��n:v�ȸ�5����G� ��A:�G#��Q����P$���۩�]_��-Nü      -�)���&�\<��3��� ��zܼ�*��A琼2�\�� ���ػ���%O���Ϲ8�J:yh�:v�;��(;�d8;��A;*�F;��H;=�I;��I;!�I;�I;}�I;zdI;�JI;36I;�&I;I;&I;�I;{I;�I;@I;�I;{I;�I;&I;I;�&I;36I;�JI;zdI;}�I;�I;!�I;��I;=�I;��H;*�F;��A;�d8;��(;v�;yh�:8�J:��Ϲ%O������ػ� �2�\�A琼�*���zܼ�� ��3�\<���&�      �L��Gى��Ă�J�o�+T���5��G�W�_��Z��#�A�fc �ݒ��������8�J:tj�:�d;3,;��:;"4C;+kG;DI;�I;��I;��I;��I;�uI;�WI;b@I;�.I;,!I;�I;�I;�
I;I;eI;I;�
I;�I;�I;,!I;�.I;b@I;�WI;�uI;��I;��I;��I;�I;DI;+kG;"4C;��:;3,;�d;tj�:8�J:������ݒ��fc �#�A�Z��_��W��G���5�+T�J�o��Ă�Gى�      3�i�&Խ��������8W��C�o�{??�G��^zܼ�Q���X�2R�/7�������Ϲ��n:�k�:!=;��0;�>;KE;rRH;d�I;��I;�I;[�I;y�I;�eI;DKI;�6I;'I;$I;I;{I;8I;Y
I;8I;{I;I;$I;'I;�6I;DKI;�eI;y�I;[�I;�I;��I;d�I;rRH;KE;�>;��0;!=;�k�:��n:��Ϲ���/7��2R��X��Q��^zܼG��{??�C�o�8W����������&Խi�      �7�74�s�)�'>����3�t���9Inc��)�׃��۩��a�2R�ݒ��%O�v�ȸ%��:��;�#;��6;gA;��F;�I;Y�I;��I;0�I;��I;�tI;�VI;�?I;%.I;|!I;2I;I;�I;xI;�I;I;2I;|!I;%.I;�?I;�VI;�tI;��I;0�I;��I;Y�I;�I;��F;gA;��6;�#;��;%��:v�ȸ%O�ݒ��2R��a�۩�׃���)�Inc�9t���3����'>�s�)�74�      �S���7���X��Y�s��_S���0����`ང����|�|�5����۩��X�fc �����5����9"��:��;�,;�K<;vnD;'-H;�I;��I;��I;u�I;q�I;ZbI;|HI;�4I;�&I;eI;�I;�I;�I;�I;�I;eI;�&I;�4I;|HI;ZbI;q�I;u�I;��I;��I;�I;'-H;vnD;�K<;�,;��;"��:��9�5�����fc ��X�۩����|�5��|�����`ས����0��_S�Y�s��X���7��      D���s�YD־�t��q���X��{�W�0�&��l��*N���Ă�|�5�׃���Q��#�A���ػ��G�!&/�8f:`�:Õ;x�5;�8A;]�F;�)I;��I;��I;+�I;}�I;QnI;�QI;�;I;4,I;� I;aI;I;�I;I;aI;� I;4,I;�;I;�QI;QnI;}�I;+�I;��I;��I;�)I;]�F;�8A;x�5;Õ;`�:8f:!&/���G���ػ#�A��Q��׃��|�5��Ă�*N���l��0�&�{�W��X��q���t��YD־�s�      ��7�q�3��'��K�&�����̾#���Y�s�r74����*N���|��)�^zܼZ��� � ��P���D9ꇹ:-�;-;%=;�E;!�H;o�I;M�I;��I;ǤI;<zI;�ZI;�BI;q1I;2%I;�I;II;�I;II;�I;2%I;q1I;�BI;�ZI;<zI;ǤI;��I;M�I;o�I;!�H;�E;%=;-;-�;ꇹ:D9P��� ��� �Z��^zܼ�)��|�*N�����r74�Y�s�#�����̾&����K��'�q�3�      %8��hڇ��x|�nm_�Dv<����?��l8��'6~�r74��l������Inc�G��_��2�\�A:�UZ�� >���n:[��:#;�8;ܿB;��G;�wI;��I;��I;��I;��I;ZcI;�II;�6I;5)I;W I;lI;�I;lI;W I;5)I;�6I;�II;ZcI;��I;��I;��I;��I;�wI;��G;ܿB;�8;#;[��:��n:� >�UZ�A:�2�\�_��G��Inc������l��r74�'6~�l8��?�꾎��Dv<�nm_��x|�hڇ�      ��ȿ�ÿ���)8��gڇ�Z��'�����l8��Y�s�0�&�`�9{??�W�A琼�G#��7���Vܺ��9U�:��;8K2;c@;��F;I;��I;��I;p�I;d�I;�kI;�OI;u;I;-I;�#I;CI;dI;CI;�#I;-I;u;I;�OI;�kI;d�I;p�I;��I;��I;I;��F;c@;8K2;��;U�:��9�Vܺ�7���G#�A琼W�{??�9`�0�&�Y�s�l8�������'�Z�gڇ�)8������ÿ      ��	�#X�I����,ݿE����ҕ� �d��'�?��#���{�W����t���C�o��G��*���Q�'�ػ�0�4�~���:��;N,;q=;WAE;��H;��I;��I;h�I;�I;�sI;�UI;�?I;�0I;�&I;� I;�I;� I;�&I;�0I;�?I;�UI;�sI;�I;h�I;��I;��I;��H;WAE;q=;N,;��;��:4�~��0�'�ػ�Q��*���G�C�o�t������{�W�#���?�꾊'� �d��ҕ�E����,ݿI���#X�      �5�321���#�L��o���ÿ�ҕ�Z������̾�X����0�3�8W����5��zܼ������l�s��Y\�]�n:���:��%;��9;��C;.H;1�I;1�I;%�I;��I;�zI;-[I;�CI;�3I;L)I;8#I;8!I;8#I;L)I;�3I;�CI;-[I;�zI;��I;%�I;1�I;1�I;.H;��C;��9;��%;���:]�n:�Y\�l�s��������zܼ��5�8W��3佃�0��X����̾���Z��ҕ��ÿo��L����#�321�      +�j���c�s�P��5���o��E���gڇ�Dv<�&���q���_S��������+T��� �P$��+H#�W���p3����:ǯ�:Q�;67;��B;��G;׆I;6�I;��I;�I;��I;�_I;fGI;�6I;�+I;*%I;#I;*%I;�+I;�6I;fGI;�_I;��I;�I;��I;6�I;׆I;��G;��B;67;Q�;ǯ�:��:p3��W���+H#�P$���� �+T���������_S�q��&���Dv<�gڇ�E���o�����5�s�P���c�      ΢��Z���C���/]��5�L���,ݿ)8��nm_��K��t��Y�s�'>�����J�o��3��۩��:��T�������9�d�:�;;�^4;&gA;:7G;�cI;%�I;P�I;w�I;��I;KcI;7JI;�8I;m-I;�&I;�$I;�&I;m-I;�8I;7JI;KcI;��I;w�I;P�I;%�I;�cI;:7G;&gA;�^4;�;;�d�:��9����T���:��۩��3�J�o�����'>�Y�s��t���K�nm_�)8���,ݿL���5��/]�C��Z���      �����B����C��s�P���#�I�������x|��'�YD־�X��s�)�&Խ�Ă�\<�]_���-M�j ˻^��	�8Б�:�;J2;/u@;��F;�EI;��I;+�I;F�I;%�I;�eI;YLI;c:I;�.I;�'I;�%I;�'I;�.I;c:I;YLI;�eI;%�I;F�I;+�I;��I;�EI;��F;/u@;J2;�;Б�:	�8^��j ˻�-M�]_��\<��Ă�&Խs�)��X��YD־�'��x|����I�����#�s�P�C�����B��      ��������B��Z�����c�321�#X��ÿhڇ�q�3��s��7��74�i�Gى���&�-Nür�X�>�ػ��%���J�ρ�:�a;z�0;��?;8�F;�1I;�I;c�I;
�I;m�I;xgI;�MI;R;I;�/I;~(I;�&I;~(I;�/I;R;I;�MI;xgI;m�I;
�I;c�I;�I;�1I;8�F;��?;z�0;�a;ρ�:��J���%�>�ػr�X�-Nü��&�Gى�i�74��7���s�q�3�hڇ��ÿ#X�321���c�Z����B�����      A(��o'���o��L�d��X1�|x�Ŀ����3�v���x����4�s��b+���'�"�ü�yY�llٻq&�`�p�X��:_;��0;��?;�F;tI;�I;��I;H�I;��I;ucI;�JI;�8I;�-I;�&I;�$I;�&I;�-I;�8I;�JI;ucI;��I;H�I;��I;�I;tI;�F;��?;��0;_;X��:`�p�q&�llٻ�yY�"�ü�'�b+��s����4��x��v���3����Ŀ|x��X1�d�L��o��o'��      o'���X��c^�������]]���,�N9�3g��S�����/����o��j1��hܽ���-$��l��,}U��Ի~!�
�-���:;�41;��?;m�F;N&I;��I;7�I;Y�I;ąI;�bI;\JI;�8I;E-I;�&I;�$I;�&I;E-I;�8I;\JI;�bI;ąI;Y�I;7�I;��I;N&I;m�F;��?;�41;;��:
�-�~!��Ի,}U��l���-$����hܽj1��o���྘�/�S���3g��N9���,��]]�����c^���X��      �o��c^���ē��4z�1K�e��M��$ﱿQ�v��X#���Ѿń�	�&�w�нk̀�r��������I� ǻ�5��9�
�:W�;!�2;��@;�F;:I;�I;�I;��I;��I;qaI;II;�7I;~,I;�%I;�#I;�%I;~,I;�7I;II;qaI;��I;��I;�I;�I;:I;�F;��@;!�2;W�;�
�:�9�5� ǻ��I�����r��k̀�w�н	�&�ń���Ѿ�X#�Q�v�$ﱿM��e��1K��4z��ē�c^��      L������4z���V��X1��<�pؿ����RZ��	�(���KUo����fy��?l�l�S����7������𺣽�9��:��;]�4;�sA;�1G;�WI;��I;r�I;)�I;�I;�^I;GI;A6I;+I;�$I;�"I;�$I;+I;A6I;GI;�^I;�I;)�I;r�I;��I;�WI;�1G;�sA;]�4;��;��:���9�𺙼����7�S��l�?l�fy�����KUo�(����	��RZ����pؿ�<��X1���V��4z�����      d��]]�1K��X1�Xf���kQ��R���Z58��A���נ���O���h什�Q�,���cߓ��� �W��}谺�":��:# ;�/7;�B;`�G;{I;�I;��I;ԦI;]{I;Z[I;hDI;;4I;X)I;Q#I;G!I;Q#I;X)I;;4I;hDI;Z[I;]{I;ԦI;��I;�I;{I;`�G;�B;�/7;# ;��:�":}谺W���� �cߓ�,����Q�h什����O��נ��A��Z58�R���kQ����Xf��X1�1K��]]�      �X1���,�e���<���2g��c_���U�˂�ՌȾ	ń�-�-�q��Y ��8�2�.?ټ��{�G"��n��O���u:�O ;�&;5":;[�C;!%H;0�I;D�I;��I;�I;�uI;�VI;AI;�1I;3'I;c!I;}I;c!I;3'I;�1I;AI;�VI;�uI;�I;��I;D�I;0�I;!%H;[�C;5":;�&;�O ;��u:�O��n�G"���{�.?ټ8�2�Y ��q��-�-�	ń�ՌȾ˂��U�c_��2g���<�e����,�      |x�N9�M��pؿkQ��c_��4�_��X#�p���f��<�S�{�����-l�T�-w��f�M�#�Ի �+��LT���:�d;�[,;/=;�AE;|�H;��I;��I;��I;֕I;�nI;�QI;/=I;|.I;�$I;I;cI;I;�$I;|.I;/=I;�QI;�nI;֕I;��I;��I;��I;|�H;�AE;/=;�[,;�d;��:�LT� �+�#�Իf�M�-w��T�-l�����{�<�S��f��p���X#�4�_�c_��kQ��pؿM��N9�      Ŀ3g��$ﱿ���R����U��X#�r��d���JUo�
�#��hܽ����n<����`���҉ �;❻J�Ժ�l�9r��:�U;�2;�@;t�F;�I;�I;b�I;K�I;��I;%gI;.LI;�8I;+I;�!I;�I;�I;�I;�!I;+I;�8I;.LI;%gI;��I;K�I;b�I;�I;�I;t�F;�@;�2;�U;r��:�l�9J�Ժ;❻҉ �`�������n<�����hܽ
�#�JUo�d���r���X#��U�R������$ﱿ3g��      ���S���Q�v��RZ�Z58�˂�p��d���hoy�`1�gO��d什�`�`��7����yY���컟�T��1���u:��:\~#;.88;�B;��G;lI;-�I;!�I;L�I;��I;�^I;!FI;4I;C'I;�I;�I;)I;�I;�I;C'I;4I;!FI;�^I;��I;L�I;!�I;-�I;lI;��G;�B;.88;\~#;��:��u:�1���T���컷yY�7���`���`�d什gO��`1�hoy�d���p��˂�Z58��RZ�Q�v�S���      �3���/��X#��	��A��ՌȾ�f��JUo�`1�Ӱ���n���x��'��>ټ�@��-l�S���%���39�!�:;Q; d-;�.=;�E;~wH;��I;,�I;��I; �I;6uI;�VI;�?I;/I;B#I;_I;�I;TI;�I;_I;B#I;/I;�?I;�VI;6uI; �I;��I;,�I;��I;~wH;�E;�.=; d-;;Q;�!�:�39%��S���-l��@���>ټ�'��x��n��Ӱ��`1�JUo��f��ՌȾ�A���	��X#���/�      v���ྃ�Ѿ(����נ�	ń�<�S�
�#�gO���n��R̀��2�-������>���Ի��B��#�Zm:�E�:o ;��5;�EA;��F;�I;r�I;p�I;ŽI;��I;�iI;�MI;.9I;�)I;I;�I;�I;iI;�I;�I;I;�)I;.9I;�MI;�iI;��I;ŽI;p�I;r�I;�I;��F;�EA;��5;o ;�E�:Zm:�#���B���Ի��>���-���2�R̀��n��gO��
�#�<�S�	ń��נ�(�����Ѿ��      �x���o��ń�KUo���O�-�-�{��hܽd什�x��2��b��yR���|U��2�����$찺�m�9��:C;��,;�g<;�qD;g$H;�I;��I;��I;&�I;&I;�]I;(EI;r2I;�$I;�I;}I;�I;PI;�I;}I;�I;�$I;r2I;(EI;�]I;&I;&�I;��I;��I;�I;g$H;�qD;�g<;��,;C;��:�m�9$찺����2���|U�yR���b���2��x�d什�hܽ{�-�-���O�KUo�ń��o��      ��4�j1�	�&������q�ཌྷ�������`��'�-��yR����]�����V��[����o����:{�;=~#;/�6;nsA;r�F;�I;��I;��I;��I;6�I;�oI;�RI;�<I;�+I;�I;�I;�I;`I;VI;`I;�I;�I;�I;�+I;�<I;�RI;�oI;6�I;��I;��I;��I;�I;r�F;nsA;/�6;=~#;{�;���:��o�[���V�������]�yR��-��'��`��������q�������	�&�j1�      s�ཾhܽw�нfy��h什Y ��-l��n<�`���>ټ�𛼝|U����H᝻�2�������u:ij�:�;}61;j(>;rE;+IH;p�I;��I;��I;�I;��I;zaI;�GI;G4I;~%I;�I;�I;XI;<
I;6	I;<
I;XI;�I;�I;~%I;G4I;�GI;zaI;��I;�I;��I;��I;p�I;+IH;rE;j(>;}61;�;ij�:��u:�����2�H᝻����|U����>ټ`���n<�-l�Y ��h什fy��w�н�hܽ      b+����k̀�?l��Q�8�2�T����7����@����>��2���V���2���� R:���:�;�[,;P;;;C;�dG;w8I;��I;U�I;��I;^�I;�pI;�SI;=I;W,I;KI;�I;�I;�	I;+I;'I;+I;�	I;�I;�I;KI;W,I;=I;�SI;�pI;^�I;��I;U�I;��I;w8I;�dG;;C;P;;�[,;�;���: R:���2��V���2����>��@��7������T�8�2��Q�?l�k̀���      �'��-$�r��l�,���.?ټ-w��`����yY�-l���Ի���[������ R:���:�Q;�);��8;��A;�F;R�H;I�I;��I;��I;ȨI;$�I;�_I;GI;�3I;�$I;cI;�I;�
I;�I;*I;]I;*I;�I;�
I;�I;cI;�$I;�3I;GI;�_I;$�I;ȨI;��I;��I;I�I;R�H;�F;��A;��8;�);�Q;���: R:����[�������Ի-l��yY�`���-w��.?ټ,���l�r���-$�      "�ü�l������S��cߓ���{�f�M�҉ ����S�����B�$찺��o���u:���:�Q;D�';)07;ք@;�E;�kH;N�I;��I;��I;+�I;��I;�kI;�PI;D;I;�*I;�I;�I;|I;�I;[I;CI;� I;CI;[I;�I;|I;�I;�I;�*I;D;I;�PI;�kI;��I;+�I;��I;��I;N�I;�kH;�E;ք@;)07;D�';�Q;���:��u:��o�$찺��B�S������҉ �f�M���{�cߓ�S�������l��      �yY�,}U���I���7��� �G"�#�Ի;❻��T�%���#��m�9���:ij�:�;�);)07;D@;V\E;�#H;�jI;(�I;s�I;�I;L�I;�vI;�YI;�BI;�0I;g"I;DI;�I;EI;�I;N I;�H;�H;�H;N I;�I;EI;�I;DI;g"I;�0I;�BI;�YI;�vI;L�I;�I;s�I;(�I;�jI;�#H;V\E;D@;)07;�);�;ij�:���:�m�9�#�%���T�;❻#�ԻG"��� ���7���I�,}U�      llٻ�Ի ǻ����W���n� �+�J�Ժ�1��39Zm:��:{�;�;�[,;��8;ք@;V\E;�	H;jUI;��I;	�I;�I;}�I;#�I;�aI;}II;>6I;�&I;�I;GI;�	I;NI;O I;{�H;��H;��H;��H;{�H;O I;NI;�	I;GI;�I;�&I;>6I;}II;�aI;#�I;}�I;�I;	�I;��I;jUI;�	H;V\E;ք@;��8;�[,;�;{�;��:Zm:�39�1�J�Ժ �+��n�W������ ǻ�Ի      q&�~!��5���}谺�O��LT��l�9��u:�!�:�E�:C;=~#;}61;P;;��A;�E;�#H;jUI;,�I;��I;0�I;��I;�I;-hI;BOI;6;I;+I;3I;�I;�I;�I;� I;F�H;��H;��H;�H;��H;��H;F�H;� I;�I;�I;�I;3I;+I;6;I;BOI;-hI;�I;��I;0�I;��I;,�I;jUI;�#H;�E;��A;P;;}61;=~#;C;�E�:�!�:��u:�l�9�LT��O�}谺���5�~!�      `�p�
�-��9���9�":��u:��:r��:��:;Q;o ;��,;/�6;j(>;;C;�F;�kH;�jI;��I;��I;��I;4�I;��I;�lI;�SI;??I;�.I;8!I;nI;�I;�I;�I;��H;��H;��H;c�H;��H;c�H;��H;��H;��H;�I;�I;�I;nI;8!I;�.I;??I;�SI;�lI;��I;4�I;��I;��I;��I;�jI;�kH;�F;;C;j(>;/�6;��,;o ;;Q;��:r��:��:��u:�":���9�9
�-�      X��:��:�
�:��:��:�O ;�d;�U;\~#; d-;��5;�g<;nsA;rE;�dG;R�H;N�I;(�I;	�I;0�I;4�I;�I;!oI;aVI;BI;X1I;�#I;�I;�I;VI;�I;�H;��H;�H;f�H;>�H;��H;>�H;f�H;�H;��H;�H;�I;VI;�I;�I;�#I;X1I;BI;aVI;!oI;�I;4�I;0�I;	�I;(�I;N�I;R�H;�dG;rE;nsA;�g<;��5; d-;\~#;�U;�d;�O ;��:��:�
�:��:      _;;W�;��;# ;�&;�[,;�2;.88;�.=;�EA;�qD;r�F;+IH;w8I;I�I;��I;s�I;�I;��I;��I;!oI;bWI;�CI;3I;r%I;7I;�I;�	I;�I;��H;��H;��H;��H;H�H;V�H;�H;V�H;H�H;��H;��H;��H;��H;�I;�	I;�I;7I;r%I;3I;�CI;bWI;!oI;��I;��I;�I;s�I;��I;I�I;w8I;+IH;r�F;�qD;�EA;�.=;.88;�2;�[,;�&;# ;��;W�;;      ��0;�41;!�2;]�4;�/7;5":;/=;�@;�B;�E;��F;g$H;�I;p�I;��I;��I;��I;�I;}�I;�I;�lI;aVI;�CI;�3I;Y&I;DI;I;�
I;II;>�H;A�H;��H;��H;��H;o�H;��H;w�H;��H;o�H;��H;��H;��H;A�H;>�H;II;�
I;I;DI;Y&I;�3I;�CI;aVI;�lI;�I;}�I;�I;��I;��I;��I;p�I;�I;g$H;��F;�E;�B;�@;/=;5":;�/7;]�4;!�2;�41;      ��?;��?;��@;�sA;�B;[�C;�AE;t�F;��G;~wH;�I;�I;��I;��I;U�I;��I;+�I;L�I;#�I;-hI;�SI;BI;3I;Y&I;�I;�I;)I;�I;��H;��H;&�H;z�H;p�H;��H;��H;5�H;�H;5�H;��H;��H;p�H;z�H;&�H;��H;��H;�I;)I;�I;�I;Y&I;3I;BI;�SI;-hI;#�I;L�I;+�I;��I;U�I;��I;��I;�I;�I;~wH;��G;t�F;�AE;[�C;�B;�sA;��@;��?;      �F;m�F;�F;�1G;`�G;!%H;|�H;�I;lI;��I;r�I;��I;��I;��I;��I;ȨI;��I;�vI;�aI;BOI;??I;X1I;r%I;DI;�I;OI;1I; I;��H;U�H;��H;c�H;��H;4�H;e�H;��H;��H;��H;e�H;4�H;��H;c�H;��H;U�H;��H; I;1I;OI;�I;DI;r%I;X1I;??I;BOI;�aI;�vI;��I;ȨI;��I;��I;��I;��I;r�I;��I;lI;�I;|�H;!%H;`�G;�1G;�F;m�F;      tI;N&I;:I;�WI;{I;0�I;��I;�I;-�I;,�I;p�I;��I;��I;�I;^�I;$�I;�kI;�YI;}II;6;I;�.I;�#I;7I;I;)I;1I; I;��H;}�H;��H;\�H;`�H;��H;��H;�H;��H;w�H;��H;�H;��H;��H;`�H;\�H;��H;}�H;��H; I;1I;)I;I;7I;�#I;�.I;6;I;}II;�YI;�kI;$�I;^�I;�I;��I;��I;p�I;,�I;-�I;�I;��I;0�I;{I;�WI;:I;N&I;      �I;��I;�I;��I;�I;D�I;��I;b�I;!�I;��I;ŽI;&�I;6�I;��I;�pI;�_I;�PI;�BI;>6I;+I;8!I;�I;�I;�
I;�I; I;��H;y�H;��H;c�H;a�H;��H;��H;��H;��H;��H;y�H;��H;��H;��H;��H;��H;a�H;c�H;��H;y�H;��H; I;�I;�
I;�I;�I;8!I;+I;>6I;�BI;�PI;�_I;�pI;��I;6�I;&�I;ŽI;��I;!�I;b�I;��I;D�I;�I;��I;�I;��I;      ��I;7�I;�I;r�I;��I;��I;��I;K�I;L�I; �I;��I;&I;�oI;zaI;�SI;GI;D;I;�0I;�&I;3I;nI;�I;�	I;II;��H;��H;}�H;��H;X�H;[�H;��H;Z�H;K�H;��H;��H;��H;��H;��H;��H;��H;K�H;Z�H;��H;[�H;X�H;��H;}�H;��H;��H;II;�	I;�I;nI;3I;�&I;�0I;D;I;GI;�SI;zaI;�oI;&I;��I; �I;L�I;K�I;��I;��I;��I;r�I;�I;7�I;      H�I;Y�I;��I;)�I;ԦI;�I;֕I;��I;��I;6uI;�iI;�]I;�RI;�GI;=I;�3I;�*I;g"I;�I;�I;�I;VI;�I;>�H;��H;U�H;��H;c�H;[�H;��H;6�H;�H;B�H;��H;�H;��H;��H;��H;�H;��H;B�H;�H;6�H;��H;[�H;c�H;��H;U�H;��H;>�H;�I;VI;�I;�I;�I;g"I;�*I;�3I;=I;�GI;�RI;�]I;�iI;6uI;��I;��I;֕I;�I;ԦI;)�I;��I;Y�I;      ��I;ąI;��I;�I;]{I;�uI;�nI;%gI;�^I;�VI;�MI;(EI;�<I;G4I;W,I;�$I;�I;DI;GI;�I;�I;�I;��H;A�H;&�H;��H;\�H;a�H;��H;6�H;�H;�H;\�H;��H;z�H;7�H;��H;7�H;z�H;��H;\�H;�H;�H;6�H;��H;a�H;\�H;��H;&�H;A�H;��H;�I;�I;�I;GI;DI;�I;�$I;W,I;G4I;�<I;(EI;�MI;�VI;�^I;%gI;�nI;�uI;]{I;�I;��I;ąI;      ucI;�bI;qaI;�^I;Z[I;�VI;�QI;.LI;!FI;�?I;.9I;r2I;�+I;~%I;KI;cI;�I;�I;�	I;�I;�I;�H;��H;��H;z�H;c�H;`�H;��H;Z�H;�H;�H;U�H;��H;,�H;��H;��H;��H;��H;��H;,�H;��H;U�H;�H;�H;Z�H;��H;`�H;c�H;z�H;��H;��H;�H;�I;�I;�	I;�I;�I;cI;KI;~%I;�+I;r2I;.9I;�?I;!FI;.LI;�QI;�VI;Z[I;�^I;qaI;�bI;      �JI;\JI;II;GI;hDI;AI;/=I;�8I;4I;/I;�)I;�$I;�I;�I;�I;�I;|I;EI;NI;� I;��H;��H;��H;��H;p�H;��H;��H;��H;K�H;B�H;\�H;��H;�H;��H;M�H;!�H;3�H;!�H;M�H;��H;�H;��H;\�H;B�H;K�H;��H;��H;��H;p�H;��H;��H;��H;��H;� I;NI;EI;|I;�I;�I;�I;�I;�$I;�)I;/I;4I;�8I;/=I;AI;hDI;GI;II;\JI;      �8I;�8I;�7I;A6I;;4I;�1I;|.I;+I;C'I;B#I;I;�I;�I;�I;�I;�
I;�I;�I;O I;F�H;��H;�H;��H;��H;��H;4�H;��H;��H;��H;��H;��H;,�H;��H;<�H;��H;��H;��H;��H;��H;<�H;��H;,�H;��H;��H;��H;��H;��H;4�H;��H;��H;��H;�H;��H;F�H;O I;�I;�I;�
I;�I;�I;�I;�I;I;B#I;C'I;+I;|.I;�1I;;4I;A6I;�7I;�8I;      �-I;E-I;~,I;+I;X)I;3'I;�$I;�!I;�I;_I;�I;}I;�I;XI;�	I;�I;[I;N I;{�H;��H;��H;f�H;H�H;o�H;��H;e�H;�H;��H;��H;�H;z�H;��H;M�H;��H;��H;��H;�H;��H;��H;��H;M�H;��H;z�H;�H;��H;��H;�H;e�H;��H;o�H;H�H;f�H;��H;��H;{�H;N I;[I;�I;�	I;XI;�I;}I;�I;_I;�I;�!I;�$I;3'I;X)I;+I;~,I;E-I;      �&I;�&I;�%I;�$I;Q#I;c!I;I;�I;�I;�I;�I;�I;`I;<
I;+I;*I;CI;�H;��H;��H;c�H;>�H;V�H;��H;5�H;��H;��H;��H;��H;��H;7�H;��H;!�H;��H;��H;k�H;r�H;k�H;��H;��H;!�H;��H;7�H;��H;��H;��H;��H;��H;5�H;��H;V�H;>�H;c�H;��H;��H;�H;CI;*I;+I;<
I;`I;�I;�I;�I;�I;�I;I;c!I;Q#I;�$I;�%I;�&I;      �$I;�$I;�#I;�"I;G!I;}I;cI;�I;)I;TI;iI;PI;VI;6	I;'I;]I;� I;�H;��H;�H;��H;��H;�H;w�H;�H;��H;w�H;y�H;��H;��H;��H;��H;3�H;��H;�H;r�H;w�H;r�H;�H;��H;3�H;��H;��H;��H;��H;y�H;w�H;��H;�H;w�H;�H;��H;��H;�H;��H;�H;� I;]I;'I;6	I;VI;PI;iI;TI;)I;�I;cI;}I;G!I;�"I;�#I;�$I;      �&I;�&I;�%I;�$I;Q#I;c!I;I;�I;�I;�I;�I;�I;`I;<
I;+I;*I;CI;�H;��H;��H;c�H;>�H;V�H;��H;5�H;��H;��H;��H;��H;��H;7�H;��H;!�H;��H;��H;k�H;r�H;k�H;��H;��H;!�H;��H;7�H;��H;��H;��H;��H;��H;5�H;��H;V�H;>�H;c�H;��H;��H;�H;CI;*I;+I;<
I;`I;�I;�I;�I;�I;�I;I;c!I;Q#I;�$I;�%I;�&I;      �-I;E-I;~,I;+I;X)I;3'I;�$I;�!I;�I;_I;�I;}I;�I;XI;�	I;�I;[I;N I;{�H;��H;��H;f�H;H�H;o�H;��H;e�H;�H;��H;��H;�H;z�H;��H;M�H;��H;��H;��H;�H;��H;��H;��H;M�H;��H;z�H;�H;��H;��H;�H;e�H;��H;o�H;H�H;f�H;��H;��H;{�H;N I;[I;�I;�	I;XI;�I;}I;�I;_I;�I;�!I;�$I;3'I;X)I;+I;~,I;E-I;      �8I;�8I;�7I;A6I;;4I;�1I;|.I;+I;C'I;B#I;I;�I;�I;�I;�I;�
I;�I;�I;O I;F�H;��H;�H;��H;��H;��H;4�H;��H;��H;��H;��H;��H;,�H;��H;<�H;��H;��H;��H;��H;��H;<�H;��H;,�H;��H;��H;��H;��H;��H;4�H;��H;��H;��H;�H;��H;F�H;O I;�I;�I;�
I;�I;�I;�I;�I;I;B#I;C'I;+I;|.I;�1I;;4I;A6I;�7I;�8I;      �JI;\JI;II;GI;hDI;AI;/=I;�8I;4I;/I;�)I;�$I;�I;�I;�I;�I;|I;EI;NI;� I;��H;��H;��H;��H;p�H;��H;��H;��H;K�H;B�H;\�H;��H;�H;��H;M�H;!�H;3�H;!�H;M�H;��H;�H;��H;\�H;B�H;K�H;��H;��H;��H;p�H;��H;��H;��H;��H;� I;NI;EI;|I;�I;�I;�I;�I;�$I;�)I;/I;4I;�8I;/=I;AI;hDI;GI;II;\JI;      ucI;�bI;qaI;�^I;Z[I;�VI;�QI;.LI;!FI;�?I;.9I;r2I;�+I;~%I;KI;cI;�I;�I;�	I;�I;�I;�H;��H;��H;z�H;c�H;`�H;��H;Z�H;�H;�H;U�H;��H;,�H;��H;��H;��H;��H;��H;,�H;��H;U�H;�H;�H;Z�H;��H;`�H;c�H;z�H;��H;��H;�H;�I;�I;�	I;�I;�I;cI;KI;~%I;�+I;r2I;.9I;�?I;!FI;.LI;�QI;�VI;Z[I;�^I;qaI;�bI;      ��I;ąI;��I;�I;]{I;�uI;�nI;%gI;�^I;�VI;�MI;(EI;�<I;G4I;W,I;�$I;�I;DI;GI;�I;�I;�I;��H;A�H;&�H;��H;\�H;a�H;��H;6�H;�H;�H;\�H;��H;z�H;7�H;��H;7�H;z�H;��H;\�H;�H;�H;6�H;��H;a�H;\�H;��H;&�H;A�H;��H;�I;�I;�I;GI;DI;�I;�$I;W,I;G4I;�<I;(EI;�MI;�VI;�^I;%gI;�nI;�uI;]{I;�I;��I;ąI;      H�I;Y�I;��I;)�I;ԦI;�I;֕I;��I;��I;6uI;�iI;�]I;�RI;�GI;=I;�3I;�*I;g"I;�I;�I;�I;VI;�I;>�H;��H;U�H;��H;c�H;[�H;��H;6�H;�H;B�H;��H;�H;��H;��H;��H;�H;��H;B�H;�H;6�H;��H;[�H;c�H;��H;U�H;��H;>�H;�I;VI;�I;�I;�I;g"I;�*I;�3I;=I;�GI;�RI;�]I;�iI;6uI;��I;��I;֕I;�I;ԦI;)�I;��I;Y�I;      ��I;7�I;�I;r�I;��I;��I;��I;K�I;L�I; �I;��I;&I;�oI;zaI;�SI;GI;D;I;�0I;�&I;3I;nI;�I;�	I;II;��H;��H;}�H;��H;X�H;[�H;��H;Z�H;K�H;��H;��H;��H;��H;��H;��H;��H;K�H;Z�H;��H;[�H;X�H;��H;}�H;��H;��H;II;�	I;�I;nI;3I;�&I;�0I;D;I;GI;�SI;zaI;�oI;&I;��I; �I;L�I;K�I;��I;��I;��I;r�I;�I;7�I;      �I;��I;�I;��I;�I;D�I;��I;b�I;!�I;��I;ŽI;&�I;6�I;��I;�pI;�_I;�PI;�BI;>6I;+I;8!I;�I;�I;�
I;�I; I;��H;y�H;��H;c�H;a�H;��H;��H;��H;��H;��H;y�H;��H;��H;��H;��H;��H;a�H;c�H;��H;y�H;��H; I;�I;�
I;�I;�I;8!I;+I;>6I;�BI;�PI;�_I;�pI;��I;6�I;&�I;ŽI;��I;!�I;b�I;��I;D�I;�I;��I;�I;��I;      tI;N&I;:I;�WI;{I;0�I;��I;�I;-�I;,�I;p�I;��I;��I;�I;^�I;$�I;�kI;�YI;}II;6;I;�.I;�#I;7I;I;)I;1I; I;��H;}�H;��H;\�H;`�H;��H;��H;�H;��H;w�H;��H;�H;��H;��H;`�H;\�H;��H;}�H;��H; I;1I;)I;I;7I;�#I;�.I;6;I;}II;�YI;�kI;$�I;^�I;�I;��I;��I;p�I;,�I;-�I;�I;��I;0�I;{I;�WI;:I;N&I;      �F;m�F;�F;�1G;`�G;!%H;|�H;�I;lI;��I;r�I;��I;��I;��I;��I;ȨI;��I;�vI;�aI;BOI;??I;X1I;r%I;DI;�I;OI;1I; I;��H;U�H;��H;c�H;��H;4�H;e�H;��H;��H;��H;e�H;4�H;��H;c�H;��H;U�H;��H; I;1I;OI;�I;DI;r%I;X1I;??I;BOI;�aI;�vI;��I;ȨI;��I;��I;��I;��I;r�I;��I;lI;�I;|�H;!%H;`�G;�1G;�F;m�F;      ��?;��?;��@;�sA;�B;[�C;�AE;t�F;��G;~wH;�I;�I;��I;��I;U�I;��I;+�I;L�I;#�I;-hI;�SI;BI;3I;Y&I;�I;�I;)I;�I;��H;��H;&�H;z�H;p�H;��H;��H;5�H;�H;5�H;��H;��H;p�H;z�H;&�H;��H;��H;�I;)I;�I;�I;Y&I;3I;BI;�SI;-hI;#�I;L�I;+�I;��I;U�I;��I;��I;�I;�I;~wH;��G;t�F;�AE;[�C;�B;�sA;��@;��?;      ��0;�41;!�2;]�4;�/7;5":;/=;�@;�B;�E;��F;g$H;�I;p�I;��I;��I;��I;�I;}�I;�I;�lI;aVI;�CI;�3I;Y&I;DI;I;�
I;II;>�H;A�H;��H;��H;��H;o�H;��H;w�H;��H;o�H;��H;��H;��H;A�H;>�H;II;�
I;I;DI;Y&I;�3I;�CI;aVI;�lI;�I;}�I;�I;��I;��I;��I;p�I;�I;g$H;��F;�E;�B;�@;/=;5":;�/7;]�4;!�2;�41;      _;;W�;��;# ;�&;�[,;�2;.88;�.=;�EA;�qD;r�F;+IH;w8I;I�I;��I;s�I;�I;��I;��I;!oI;bWI;�CI;3I;r%I;7I;�I;�	I;�I;��H;��H;��H;��H;H�H;V�H;�H;V�H;H�H;��H;��H;��H;��H;�I;�	I;�I;7I;r%I;3I;�CI;bWI;!oI;��I;��I;�I;s�I;��I;I�I;w8I;+IH;r�F;�qD;�EA;�.=;.88;�2;�[,;�&;# ;��;W�;;      X��:��:�
�:��:��:�O ;�d;�U;\~#; d-;��5;�g<;nsA;rE;�dG;R�H;N�I;(�I;	�I;0�I;4�I;�I;!oI;aVI;BI;X1I;�#I;�I;�I;VI;�I;�H;��H;�H;f�H;>�H;��H;>�H;f�H;�H;��H;�H;�I;VI;�I;�I;�#I;X1I;BI;aVI;!oI;�I;4�I;0�I;	�I;(�I;N�I;R�H;�dG;rE;nsA;�g<;��5; d-;\~#;�U;�d;�O ;��:��:�
�:��:      `�p�
�-��9���9�":��u:��:r��:��:;Q;o ;��,;/�6;j(>;;C;�F;�kH;�jI;��I;��I;��I;4�I;��I;�lI;�SI;??I;�.I;8!I;nI;�I;�I;�I;��H;��H;��H;c�H;��H;c�H;��H;��H;��H;�I;�I;�I;nI;8!I;�.I;??I;�SI;�lI;��I;4�I;��I;��I;��I;�jI;�kH;�F;;C;j(>;/�6;��,;o ;;Q;��:r��:��:��u:�":���9�9
�-�      q&�~!��5���}谺�O��LT��l�9��u:�!�:�E�:C;=~#;}61;P;;��A;�E;�#H;jUI;,�I;��I;0�I;��I;�I;-hI;BOI;6;I;+I;3I;�I;�I;�I;� I;F�H;��H;��H;�H;��H;��H;F�H;� I;�I;�I;�I;3I;+I;6;I;BOI;-hI;�I;��I;0�I;��I;,�I;jUI;�#H;�E;��A;P;;}61;=~#;C;�E�:�!�:��u:�l�9�LT��O�}谺���5�~!�      llٻ�Ի ǻ����W���n� �+�J�Ժ�1��39Zm:��:{�;�;�[,;��8;ք@;V\E;�	H;jUI;��I;	�I;�I;}�I;#�I;�aI;}II;>6I;�&I;�I;GI;�	I;NI;O I;{�H;��H;��H;��H;{�H;O I;NI;�	I;GI;�I;�&I;>6I;}II;�aI;#�I;}�I;�I;	�I;��I;jUI;�	H;V\E;ք@;��8;�[,;�;{�;��:Zm:�39�1�J�Ժ �+��n�W������ ǻ�Ի      �yY�,}U���I���7��� �G"�#�Ի;❻��T�%���#��m�9���:ij�:�;�);)07;D@;V\E;�#H;�jI;(�I;s�I;�I;L�I;�vI;�YI;�BI;�0I;g"I;DI;�I;EI;�I;N I;�H;�H;�H;N I;�I;EI;�I;DI;g"I;�0I;�BI;�YI;�vI;L�I;�I;s�I;(�I;�jI;�#H;V\E;D@;)07;�);�;ij�:���:�m�9�#�%���T�;❻#�ԻG"��� ���7���I�,}U�      "�ü�l������S��cߓ���{�f�M�҉ ����S�����B�$찺��o���u:���:�Q;D�';)07;ք@;�E;�kH;N�I;��I;��I;+�I;��I;�kI;�PI;D;I;�*I;�I;�I;|I;�I;[I;CI;� I;CI;[I;�I;|I;�I;�I;�*I;D;I;�PI;�kI;��I;+�I;��I;��I;N�I;�kH;�E;ք@;)07;D�';�Q;���:��u:��o�$찺��B�S������҉ �f�M���{�cߓ�S�������l��      �'��-$�r��l�,���.?ټ-w��`����yY�-l���Ի���[������ R:���:�Q;�);��8;��A;�F;R�H;I�I;��I;��I;ȨI;$�I;�_I;GI;�3I;�$I;cI;�I;�
I;�I;*I;]I;*I;�I;�
I;�I;cI;�$I;�3I;GI;�_I;$�I;ȨI;��I;��I;I�I;R�H;�F;��A;��8;�);�Q;���: R:����[�������Ի-l��yY�`���-w��.?ټ,���l�r���-$�      b+����k̀�?l��Q�8�2�T����7����@����>��2���V���2���� R:���:�;�[,;P;;;C;�dG;w8I;��I;U�I;��I;^�I;�pI;�SI;=I;W,I;KI;�I;�I;�	I;+I;'I;+I;�	I;�I;�I;KI;W,I;=I;�SI;�pI;^�I;��I;U�I;��I;w8I;�dG;;C;P;;�[,;�;���: R:���2��V���2����>��@��7������T�8�2��Q�?l�k̀���      s�ཾhܽw�нfy��h什Y ��-l��n<�`���>ټ�𛼝|U����H᝻�2�������u:ij�:�;}61;j(>;rE;+IH;p�I;��I;��I;�I;��I;zaI;�GI;G4I;~%I;�I;�I;XI;<
I;6	I;<
I;XI;�I;�I;~%I;G4I;�GI;zaI;��I;�I;��I;��I;p�I;+IH;rE;j(>;}61;�;ij�:��u:�����2�H᝻����|U����>ټ`���n<�-l�Y ��h什fy��w�н�hܽ      ��4�j1�	�&������q�ཌྷ�������`��'�-��yR����]�����V��[����o����:{�;=~#;/�6;nsA;r�F;�I;��I;��I;��I;6�I;�oI;�RI;�<I;�+I;�I;�I;�I;`I;VI;`I;�I;�I;�I;�+I;�<I;�RI;�oI;6�I;��I;��I;��I;�I;r�F;nsA;/�6;=~#;{�;���:��o�[���V�������]�yR��-��'��`��������q�������	�&�j1�      �x���o��ń�KUo���O�-�-�{��hܽd什�x��2��b��yR���|U��2�����$찺�m�9��:C;��,;�g<;�qD;g$H;�I;��I;��I;&�I;&I;�]I;(EI;r2I;�$I;�I;}I;�I;PI;�I;}I;�I;�$I;r2I;(EI;�]I;&I;&�I;��I;��I;�I;g$H;�qD;�g<;��,;C;��:�m�9$찺����2���|U�yR���b���2��x�d什�hܽ{�-�-���O�KUo�ń��o��      v���ྃ�Ѿ(����נ�	ń�<�S�
�#�gO���n��R̀��2�-������>���Ի��B��#�Zm:�E�:o ;��5;�EA;��F;�I;r�I;p�I;ŽI;��I;�iI;�MI;.9I;�)I;I;�I;�I;iI;�I;�I;I;�)I;.9I;�MI;�iI;��I;ŽI;p�I;r�I;�I;��F;�EA;��5;o ;�E�:Zm:�#���B���Ի��>���-���2�R̀��n��gO��
�#�<�S�	ń��נ�(�����Ѿ��      �3���/��X#��	��A��ՌȾ�f��JUo�`1�Ӱ���n���x��'��>ټ�@��-l�S���%���39�!�:;Q; d-;�.=;�E;~wH;��I;,�I;��I; �I;6uI;�VI;�?I;/I;B#I;_I;�I;TI;�I;_I;B#I;/I;�?I;�VI;6uI; �I;��I;,�I;��I;~wH;�E;�.=; d-;;Q;�!�:�39%��S���-l��@���>ټ�'��x��n��Ӱ��`1�JUo��f��ՌȾ�A���	��X#���/�      ���S���Q�v��RZ�Z58�˂�p��d���hoy�`1�gO��d什�`�`��7����yY���컟�T��1���u:��:\~#;.88;�B;��G;lI;-�I;!�I;L�I;��I;�^I;!FI;4I;C'I;�I;�I;)I;�I;�I;C'I;4I;!FI;�^I;��I;L�I;!�I;-�I;lI;��G;�B;.88;\~#;��:��u:�1���T���컷yY�7���`���`�d什gO��`1�hoy�d���p��˂�Z58��RZ�Q�v�S���      Ŀ3g��$ﱿ���R����U��X#�r��d���JUo�
�#��hܽ����n<����`���҉ �;❻J�Ժ�l�9r��:�U;�2;�@;t�F;�I;�I;b�I;K�I;��I;%gI;.LI;�8I;+I;�!I;�I;�I;�I;�!I;+I;�8I;.LI;%gI;��I;K�I;b�I;�I;�I;t�F;�@;�2;�U;r��:�l�9J�Ժ;❻҉ �`�������n<�����hܽ
�#�JUo�d���r���X#��U�R������$ﱿ3g��      |x�N9�M��pؿkQ��c_��4�_��X#�p���f��<�S�{�����-l�T�-w��f�M�#�Ի �+��LT���:�d;�[,;/=;�AE;|�H;��I;��I;��I;֕I;�nI;�QI;/=I;|.I;�$I;I;cI;I;�$I;|.I;/=I;�QI;�nI;֕I;��I;��I;��I;|�H;�AE;/=;�[,;�d;��:�LT� �+�#�Իf�M�-w��T�-l�����{�<�S��f��p���X#�4�_�c_��kQ��pؿM��N9�      �X1���,�e���<���2g��c_���U�˂�ՌȾ	ń�-�-�q��Y ��8�2�.?ټ��{�G"��n��O���u:�O ;�&;5":;[�C;!%H;0�I;D�I;��I;�I;�uI;�VI;AI;�1I;3'I;c!I;}I;c!I;3'I;�1I;AI;�VI;�uI;�I;��I;D�I;0�I;!%H;[�C;5":;�&;�O ;��u:�O��n�G"���{�.?ټ8�2�Y ��q��-�-�	ń�ՌȾ˂��U�c_��2g���<�e����,�      d��]]�1K��X1�Xf���kQ��R���Z58��A���נ���O���h什�Q�,���cߓ��� �W��}谺�":��:# ;�/7;�B;`�G;{I;�I;��I;ԦI;]{I;Z[I;hDI;;4I;X)I;Q#I;G!I;Q#I;X)I;;4I;hDI;Z[I;]{I;ԦI;��I;�I;{I;`�G;�B;�/7;# ;��:�":}谺W���� �cߓ�,����Q�h什����O��נ��A��Z58�R���kQ����Xf��X1�1K��]]�      L������4z���V��X1��<�pؿ����RZ��	�(���KUo����fy��?l�l�S����7������𺣽�9��:��;]�4;�sA;�1G;�WI;��I;r�I;)�I;�I;�^I;GI;A6I;+I;�$I;�"I;�$I;+I;A6I;GI;�^I;�I;)�I;r�I;��I;�WI;�1G;�sA;]�4;��;��:���9�𺙼����7�S��l�?l�fy�����KUo�(����	��RZ����pؿ�<��X1���V��4z�����      �o��c^���ē��4z�1K�e��M��$ﱿQ�v��X#���Ѿń�	�&�w�нk̀�r��������I� ǻ�5��9�
�:W�;!�2;��@;�F;:I;�I;�I;��I;��I;qaI;II;�7I;~,I;�%I;�#I;�%I;~,I;�7I;II;qaI;��I;��I;�I;�I;:I;�F;��@;!�2;W�;�
�:�9�5� ǻ��I�����r��k̀�w�н	�&�ń���Ѿ�X#�Q�v�$ﱿM��e��1K��4z��ē�c^��      o'���X��c^�������]]���,�N9�3g��S�����/����o��j1��hܽ���-$��l��,}U��Ի~!�
�-���:;�41;��?;m�F;N&I;��I;7�I;Y�I;ąI;�bI;\JI;�8I;E-I;�&I;�$I;�&I;E-I;�8I;\JI;�bI;ąI;Y�I;7�I;��I;N&I;m�F;��?;�41;;��:
�-�~!��Ի,}U��l���-$����hܽj1��o���྘�/�S���3g��N9���,��]]�����c^���X��      ����,������Q���F�Q�Ù$�.���~�7�}�E(�>�׾�T���L+���սr����@L��jO�9�ͻ�����l8�m�:��;T�1;��?;uF;s�H;��I;��I;��I;�uI;�VI;�@I;1I;�&I;� I;I;� I;�&I;1I;�@I;�VI;�uI;��I;��I;��I;s�H;uF;��?;T�1;��;�m�:��l8���9�ͻjO�@L����r����ս�L+��T��>�׾E(�7�}�~�.���Ù$�F�Q�Q��������,��      �,��^�� P���{��K��x �����n�����w��$���Ҿf��� (���ѽٷ��7����$�K��ɻ����8���:��;��1;@;��F;.I;�I;4�I;ĝI;�tI;NVI;�@I;�0I;�&I;� I;�I;� I;�&I;�0I;�@I;NVI;�tI;ĝI;4�I;�I;.I;��F;@;��1;��;���:��8���ɻ$�K����7�ٷ����ѽ (�f�����Ҿ�$���w�n��������x ��K��{� P��^��      ���� P�������d���;� ����㿰���#f�b��ž��z���C�ƽ40v�e5�R����o@����pj��Pu9^I�:=\;�63;@�@;�F;WI;��I;{�I;o�I;�rI;�TI;^?I;0I;&I;, I;MI;, I;&I;0I;^?I;�TI;�rI;o�I;{�I;��I;WI;�F;@�@;�63;=\;^I�:�Pu9pj�����o@�R���e5�40v�C�ƽ����z�žb��#f�������� ����;���d���� P��      Q����{���d��F�Ù$�7����ɿ,蒿��K�O���j�� Zb�H�8�����a����`���%�.� e��W�غǨ�9�W�:VW;�15;?�A;� G;Z6I;��I;k�I;m�I;�oI;�RI;�=I;�.I;�$I;AI;OI;AI;�$I;�.I;�=I;�RI;�oI;m�I;k�I;��I;Z6I;� G;?�A;�15;VW;�W�:Ǩ�9W�غ e��%�.�`��������a�8���H� Zb��j��O����K�,蒿��ɿ7��Ù$��F���d��{�      F�Q��K���;�Ù$��;
��޿�����w�o,���澝���(�D������I��3�G�����N��Ǩ�2��:�����9:���:�m!;��7;۸B;}�G;
YI;L�I;��I;ّI;�kI;�OI;4;I;�,I;3#I;�I;�I;�I;3#I;�,I;4;I;�OI;�kI;ّI;��I;L�I;
YI;}�G;۸B;��7;�m!;���:��9::���2��Ǩ��N�����3�G��I������(�D��������o,���w�����޿�;
�Ù$���;��K�      Ù$��x � ��7���޿m���ǅ����F�{�
��~����z��$���ս$���P2+���ϼXPp����J�]��*�"��:,�;�7';��:;�C;,H;�|I;?�I;��I;��I;�fI;�KI;98I;V*I;E!I;I;GI;I;E!I;V*I;98I;�KI;�fI;��I;��I;?�I;�|I;,H;�C;��:;�7';,�;"��:�*�J�]����XPp���ϼP2+�$�����ս�$���z��~��{�
���F�ǅ��m����޿7�� ���x �      .���������㿆�ɿ���ǅ����P�b��:�׾�`��U�H����@��a�a�!����!D�Hɻ�!������U�:�~;�H-;H{=;ABE;ȄH;)�I; �I;��I;ւI;�`I;BGI;�4I;�'I;�I; I;pI; I;�I;�'I;�4I;BGI;�`I;ւI;��I; �I;)�I;ȄH;ABE;H{=;�H-;�~;�U�:�����!�Hɻ!D���!��a�a��@����U�H��`��:�׾b����P�ǅ�������ɿ��㿯���      ~�n�������,蒿��w���F�b��Ȱ�����Yb�+����ѽ�%��'D4����@X��ʨ��H���轺L��9bp�:�; 93;;P@;�uF;9�H;%�I;��I;��I;�yI;�YI;3BI;�0I;�$I;eI;�I;@I;�I;eI;�$I;�0I;3BI;�YI;�yI;��I;��I;%�I;9�H;�uF;;P@; 93;�;bp�:L��9�轺�H��ʨ�@X�����'D4��%����ѽ+���Yb����Ȱ�b����F���w�,蒿����n���      7�}���w�#f���K�o,�{�
�:�׾�����k���'�lz꽥I���;V�LM�*����iO��G�npE����b�:T� ;��$;˳8;q�B;�G;VJI;1�I;:�I;a�I;*pI;�RI;�<I;�,I;%!I;�I;9I;�I;9I;�I;%!I;�,I;�<I;�RI;*pI;a�I;:�I;1�I;VJI;�G;q�B;˳8;��$;T� ;b�:���npE��G��iO�*���LM��;V��I��lz���'���k����:�׾{�
�o,���K�#f���w�      E(��$�b��O������~���`���Yb���'��U�N$��S�m�5����ϼ0�����_�����غ�0�9c��:F;�F.;3{=;aE;�[H;B�I;��I;��I;�I;%fI;&KI;7I;&(I;�I;�I;�I;DI;�I;�I;�I;&(I;7I;&KI;%fI;�I;��I;��I;B�I;�[H;aE;3{=;�F.;F;c��:�0�9��غ_������0����ϼ5��S�m�N$���U���'��Yb��`���~�����O��b���$�      >�׾��Ҿž�j��������z�U�H�+��lz�N$��0v�!2+����9���5�-ɻ44�0�����:���:Nn!;*O6;)kA;��F;��H;��I;��I;�I;k|I;�[I;~CI;%1I;�#I;�I;jI;�I;�I;�I;jI;�I;�#I;%1I;~CI;�[I;k|I;�I;��I;��I;��H;��F;)kA;*O6;Nn!;���:���:0��44�-ɻ�5�9�����!2+�0v�N$��lz�+��U�H���z������j��ž��Ҿ      �T��f�����z� Zb�(�D��$�����ѽ�I��S�m�!2+��������K��ﻙ�p�;��� ��9LR�:�.;��-;��<;iyD;uH;�lI;�I;��I;��I;�nI;�QI;�;I;!+I;�I;*I;OI;�I;�I;�I;OI;*I;�I;!+I;�;I;�QI;�nI;��I;��I;�I;�lI;uH;iyD;��<;��-;�.;LR�: ��9;�����p��ﻍ�K������!2+�S�m��I����ѽ���$�(�D� Zb���z�f���      �L+� (���H�������ս�@���%���;V�5���������MS�������zF��n8o�:�;��$;^7;K�A;��F;�H;��I;��I;��I;��I;uaI;�GI;-4I;A%I;II;ZI;I;�	I; 	I;�	I;I;ZI;II;A%I;-4I;�GI;uaI;��I;��I;��I;��I;�H;��F;K�A;^7;��$;�;o�:�n8zF⺧������MS�������5���;V��%���@����ս����H��� (�      ��ս��ѽC�ƽ8����I��$���a�a�'D4�LM���ϼ9����K�����G��]g�m�o���:�@�:�X;��1;jk>;�
E;/H;;pI;"�I;	�I;��I;!rI;�TI;>I;�,I;~I;�I;�I;�	I;/I;MI;/I;�	I;�I;�I;~I;�,I;>I;�TI;!rI;��I;	�I;"�I;;pI;/H;�
E;jk>;��1;�X;�@�:��:m�o�]g��G�������K�9����ϼLM�'D4�a�a�$����I��8���C�ƽ��ѽ      r��ٷ��40v���a�3�G�P2+�!�����*���0���5��ﻧ��]g��ହ�g:^�:�;1H-;3f;;NC;)RG;�I;�I;@�I;�I;%�I;+bI;�HI;�4I;�%I;�I;PI;�
I;�I;eI;sI;eI;�I;�
I;PI;�I;�%I;�4I;�HI;+bI;%�I;�I;@�I;�I;�I;)RG;NC;3f;;1H-;�;^�:�g:�ହ]g�������5�0��*������!��P2+�3�G���a�40v�ٷ��      ��7�e5���������ϼ��@X���iO����-ɻ��p�zF�m�o��g:^�:ZF;�*;�9;��A;�tF;;�H;�I;��I;ɺI;e�I;�oI;SSI;n=I;9,I;�I;�I;I;pI;�I;�I;� I;�I;�I;pI;I;�I;�I;9,I;n=I;SSI;�oI;e�I;ɺI;��I;�I;;�H;�tF;��A;�9;�*;ZF;^�:�g:m�o�zF⺙�p�-ɻ����iO�@X������ϼ������e5�7�      @L�����R���`����N��XPp�!D�ʨ��G�_���44�;����n8��:^�:ZF;�(;��7;v�@;��E;mPH;5lI;��I;�I;��I;C|I;�]I;�EI;�2I;�#I;zI;�I;		I;(I;� I; �H;h�H; �H;� I;(I;		I;�I;zI;�#I;�2I;�EI;�]I;C|I;��I;�I;��I;5lI;mPH;��E;v�@;��7;�(;ZF;^�:��:�n8;���44�_����G�ʨ�!D�XPp��N��`���R������      jO�$�K��o@�%�.�Ǩ����Hɻ�H��npE���غ0�� ��9o�:�@�:�;�*;��7;�O@;�[E;H;�HI;��I;��I;)�I;|�I;ZgI;�MI;z9I;W)I;�I;�I;�
I;,I;'I;G�H;s�H;��H;s�H;G�H;'I;,I;�
I;�I;�I;W)I;z9I;�MI;ZgI;|�I;)�I;��I;��I;�HI;H;�[E;�O@;��7;�*;�;�@�:o�: ��90����غnpE��H��Hɻ���Ǩ�%�.��o@�$�K�      9�ͻ�ɻ��� e��2��J�]��!��轺����0�9���:LR�:�;�X;1H-;�9;v�@;�[E;��G;Q4I;ճI;d�I;��I;m�I;�oI;�TI;q?I;M.I;� I;�I;YI;�I;�I;6�H;��H;,�H;��H;,�H;��H;6�H;�I;�I;YI;�I;� I;M.I;q?I;�TI;�oI;m�I;��I;d�I;ճI;Q4I;��G;�[E;v�@;�9;1H-;�X;�;LR�:���:�0�9����轺�!�J�]�2�� e������ɻ      �����pj�W�غ:����*�����L��9b�:c��:���:�.;��$;��1;3f;;��A;��E;H;Q4I;X�I;��I;m�I;��I;�uI;tZI;xDI;�2I;K$I;�I;�I;hI;�I;��H;s�H;7�H;��H;��H;��H;7�H;s�H;��H;�I;hI;�I;�I;K$I;�2I;xDI;tZI;�uI;��I;m�I;��I;X�I;Q4I;H;��E;��A;3f;;��1;��$;�.;���:c��:b�:L��9�����*�:���W�غpj���      ��l8��8�Pu9Ǩ�9��9:"��:�U�:bp�:T� ;F;Nn!;��-;^7;jk>;NC;�tF;mPH;�HI;ճI;��I;ϺI;әI;�yI;�^I;aHI;d6I;}'I;vI;�I;1
I;�I;>�H;��H;��H;�H;��H;��H;��H;�H;��H;��H;>�H;�I;1
I;�I;vI;}'I;d6I;aHI;�^I;�yI;әI;ϺI;��I;ճI;�HI;mPH;�tF;NC;jk>;^7;��-;Nn!;F;T� ;bp�:�U�:"��:��9:Ǩ�9�Pu9��8      �m�:���:^I�:�W�:���:,�;�~;�;��$;�F.;*O6;��<;K�A;�
E;)RG;;�H;5lI;��I;d�I;m�I;әI;�zI;�`I;�JI;�8I;�)I;�I;�I;�I;9I; I;�H;��H;{�H; �H;�H;��H;�H; �H;{�H;��H;�H; I;9I;�I;�I;�I;�)I;�8I;�JI;�`I;�zI;әI;m�I;d�I;��I;5lI;;�H;)RG;�
E;K�A;��<;*O6;�F.;��$;�;�~;,�;���:�W�:^I�:���:      ��;��;=\;VW;�m!;�7';�H-; 93;˳8;3{=;)kA;iyD;��F;/H;�I;�I;��I;��I;��I;��I;�yI;�`I;�KI;4:I;+I;EI;8I;I;MI;� I;��H;�H;w�H;�H;�H;a�H;2�H;a�H;�H;�H;w�H;�H;��H;� I;MI;I;8I;EI;+I;4:I;�KI;�`I;�yI;��I;��I;��I;��I;�I;�I;/H;��F;iyD;)kA;3{=;˳8; 93;�H-;�7';�m!;VW;=\;��;      T�1;��1;�63;�15;��7;��:;H{=;;P@;q�B;aE;��F;uH;�H;;pI;�I;��I;�I;)�I;m�I;�uI;�^I;�JI;4:I;�+I; I;+I;�I;*I;�I;�H;��H;~�H;4�H;��H;{�H;��H;��H;��H;{�H;��H;4�H;~�H;��H;�H;�I;*I;�I;+I; I;�+I;4:I;�JI;�^I;�uI;m�I;)�I;�I;��I;�I;;pI;�H;uH;��F;aE;q�B;;P@;H{=;��:;��7;�15;�63;��1;      ��?;@;@�@;?�A;۸B;�C;ABE;�uF;�G;�[H;��H;�lI;��I;"�I;@�I;ɺI;��I;|�I;�oI;tZI;aHI;�8I;+I; I;�I;sI;�I;I;t�H;��H;��H;;�H;d�H;��H;��H;f�H;=�H;f�H;��H;��H;d�H;;�H;��H;��H;t�H;I;�I;sI;�I; I;+I;�8I;aHI;tZI;�oI;|�I;��I;ɺI;@�I;"�I;��I;�lI;��H;�[H;�G;�uF;ABE;�C;۸B;?�A;@�@;@;      uF;��F;�F;� G;}�G;,H;ȄH;9�H;VJI;B�I;��I;�I;��I;	�I;�I;e�I;C|I;ZgI;�TI;xDI;d6I;�)I;EI;+I;sI;�I;ZI;��H;��H;��H;6�H;I�H;��H;j�H;��H;$�H;��H;$�H;��H;j�H;��H;I�H;6�H;��H;��H;��H;ZI;�I;sI;+I;EI;�)I;d6I;xDI;�TI;ZgI;C|I;e�I;�I;	�I;��I;�I;��I;B�I;VJI;9�H;ȄH;,H;}�G;� G;�F;��F;      s�H;.I;WI;Z6I;
YI;�|I;)�I;%�I;1�I;��I;��I;��I;��I;��I;%�I;�oI;�]I;�MI;q?I;�2I;}'I;�I;8I;�I;�I;ZI;��H;2�H;��H;@�H;1�H;s�H;%�H;#�H;��H;�H;��H;�H;��H;#�H;%�H;s�H;1�H;@�H;��H;2�H;��H;ZI;�I;�I;8I;�I;}'I;�2I;q?I;�MI;�]I;�oI;%�I;��I;��I;��I;��I;��I;1�I;%�I;)�I;�|I;
YI;Z6I;WI;.I;      ��I;�I;��I;��I;L�I;?�I; �I;��I;:�I;��I;�I;��I;��I;!rI;+bI;SSI;�EI;z9I;M.I;K$I;vI;�I;I;*I;I;��H;2�H;�H;M�H;-�H;d�H;��H;��H;�H;b�H;�H;��H;�H;b�H;�H;��H;��H;d�H;-�H;M�H;�H;2�H;��H;I;*I;I;�I;vI;K$I;M.I;z9I;�EI;SSI;+bI;!rI;��I;��I;�I;��I;:�I;��I; �I;?�I;L�I;��I;��I;�I;      ��I;4�I;{�I;k�I;��I;��I;��I;��I;a�I;�I;k|I;�nI;uaI;�TI;�HI;n=I;�2I;W)I;� I;�I;�I;�I;MI;�I;t�H;��H;��H;M�H;8�H;a�H;��H;��H;��H;�H;��H;<�H;5�H;<�H;��H;�H;��H;��H;��H;a�H;8�H;M�H;��H;��H;t�H;�I;MI;�I;�I;�I;� I;W)I;�2I;n=I;�HI;�TI;uaI;�nI;k|I;�I;a�I;��I;��I;��I;��I;k�I;{�I;4�I;      ��I;ĝI;o�I;m�I;ّI;��I;ւI;�yI;*pI;%fI;�[I;�QI;�GI;>I;�4I;9,I;�#I;�I;�I;�I;1
I;9I;� I;�H;��H;��H;@�H;-�H;a�H;��H;��H;��H;��H;"�H;��H;��H;c�H;��H;��H;"�H;��H;��H;��H;��H;a�H;-�H;@�H;��H;��H;�H;� I;9I;1
I;�I;�I;�I;�#I;9,I;�4I;>I;�GI;�QI;�[I;%fI;*pI;�yI;ւI;��I;ّI;m�I;o�I;ĝI;      �uI;�tI;�rI;�oI;�kI;�fI;�`I;�YI;�RI;&KI;~CI;�;I;-4I;�,I;�%I;�I;zI;�I;YI;hI;�I; I;��H;��H;��H;6�H;1�H;d�H;��H;��H;��H;��H;��H;c�H;�H;��H;��H;��H;�H;c�H;��H;��H;��H;��H;��H;d�H;1�H;6�H;��H;��H;��H; I;�I;hI;YI;�I;zI;�I;�%I;�,I;-4I;�;I;~CI;&KI;�RI;�YI;�`I;�fI;�kI;�oI;�rI;�tI;      �VI;NVI;�TI;�RI;�OI;�KI;BGI;3BI;�<I;7I;%1I;!+I;A%I;~I;�I;�I;�I;�
I;�I;�I;>�H;�H;�H;~�H;;�H;I�H;s�H;��H;��H;��H;��H;��H;K�H;��H;��H;J�H;P�H;J�H;��H;��H;K�H;��H;��H;��H;��H;��H;s�H;I�H;;�H;~�H;�H;�H;>�H;�I;�I;�
I;�I;�I;�I;~I;A%I;!+I;%1I;7I;�<I;3BI;BGI;�KI;�OI;�RI;�TI;NVI;      �@I;�@I;^?I;�=I;4;I;98I;�4I;�0I;�,I;&(I;�#I;�I;II;�I;PI;I;		I;,I;�I;��H;��H;��H;w�H;4�H;d�H;��H;%�H;��H;��H;��H;��H;K�H;��H;d�H;�H;��H;��H;��H;�H;d�H;��H;K�H;��H;��H;��H;��H;%�H;��H;d�H;4�H;w�H;��H;��H;��H;�I;,I;		I;I;PI;�I;II;�I;�#I;&(I;�,I;�0I;�4I;98I;4;I;�=I;^?I;�@I;      1I;�0I;0I;�.I;�,I;V*I;�'I;�$I;%!I;�I;�I;*I;ZI;�I;�
I;pI;(I;'I;6�H;s�H;��H;{�H;�H;��H;��H;j�H;#�H;�H;�H;"�H;c�H;��H;d�H;��H;��H;��H;��H;��H;��H;��H;d�H;��H;c�H;"�H;�H;�H;#�H;j�H;��H;��H;�H;{�H;��H;s�H;6�H;'I;(I;pI;�
I;�I;ZI;*I;�I;�I;%!I;�$I;�'I;V*I;�,I;�.I;0I;�0I;      �&I;�&I;&I;�$I;3#I;E!I;�I;eI;�I;�I;jI;OI;I;�	I;�I;�I;� I;G�H;��H;7�H;�H; �H;�H;{�H;��H;��H;��H;b�H;��H;��H;�H;��H;�H;��H;��H;d�H;[�H;d�H;��H;��H;�H;��H;�H;��H;��H;b�H;��H;��H;��H;{�H;�H; �H;�H;7�H;��H;G�H;� I;�I;�I;�	I;I;OI;jI;�I;�I;eI;�I;E!I;3#I;�$I;&I;�&I;      � I;� I;, I;AI;�I;I; I;�I;9I;�I;�I;�I;�	I;/I;eI;�I; �H;s�H;,�H;��H;��H;�H;a�H;��H;f�H;$�H;�H;�H;<�H;��H;��H;J�H;��H;��H;d�H;2�H;/�H;2�H;d�H;��H;��H;J�H;��H;��H;<�H;�H;�H;$�H;f�H;��H;a�H;�H;��H;��H;,�H;s�H; �H;�I;eI;/I;�	I;�I;�I;�I;9I;�I; I;I;�I;AI;, I;� I;      I;�I;MI;OI;�I;GI;pI;@I;�I;DI;�I;�I; 	I;MI;sI;� I;h�H;��H;��H;��H;��H;��H;2�H;��H;=�H;��H;��H;��H;5�H;c�H;��H;P�H;��H;��H;[�H;/�H;�H;/�H;[�H;��H;��H;P�H;��H;c�H;5�H;��H;��H;��H;=�H;��H;2�H;��H;��H;��H;��H;��H;h�H;� I;sI;MI; 	I;�I;�I;DI;�I;@I;pI;GI;�I;OI;MI;�I;      � I;� I;, I;AI;�I;I; I;�I;9I;�I;�I;�I;�	I;/I;eI;�I; �H;s�H;,�H;��H;��H;�H;a�H;��H;f�H;$�H;�H;�H;<�H;��H;��H;J�H;��H;��H;d�H;2�H;/�H;2�H;d�H;��H;��H;J�H;��H;��H;<�H;�H;�H;$�H;f�H;��H;a�H;�H;��H;��H;,�H;s�H; �H;�I;eI;/I;�	I;�I;�I;�I;9I;�I; I;I;�I;AI;, I;� I;      �&I;�&I;&I;�$I;3#I;E!I;�I;eI;�I;�I;jI;OI;I;�	I;�I;�I;� I;G�H;��H;7�H;�H; �H;�H;{�H;��H;��H;��H;b�H;��H;��H;�H;��H;�H;��H;��H;d�H;[�H;d�H;��H;��H;�H;��H;�H;��H;��H;b�H;��H;��H;��H;{�H;�H; �H;�H;7�H;��H;G�H;� I;�I;�I;�	I;I;OI;jI;�I;�I;eI;�I;E!I;3#I;�$I;&I;�&I;      1I;�0I;0I;�.I;�,I;V*I;�'I;�$I;%!I;�I;�I;*I;ZI;�I;�
I;pI;(I;'I;6�H;s�H;��H;{�H;�H;��H;��H;j�H;#�H;�H;�H;"�H;c�H;��H;d�H;��H;��H;��H;��H;��H;��H;��H;d�H;��H;c�H;"�H;�H;�H;#�H;j�H;��H;��H;�H;{�H;��H;s�H;6�H;'I;(I;pI;�
I;�I;ZI;*I;�I;�I;%!I;�$I;�'I;V*I;�,I;�.I;0I;�0I;      �@I;�@I;^?I;�=I;4;I;98I;�4I;�0I;�,I;&(I;�#I;�I;II;�I;PI;I;		I;,I;�I;��H;��H;��H;w�H;4�H;d�H;��H;%�H;��H;��H;��H;��H;K�H;��H;d�H;�H;��H;��H;��H;�H;d�H;��H;K�H;��H;��H;��H;��H;%�H;��H;d�H;4�H;w�H;��H;��H;��H;�I;,I;		I;I;PI;�I;II;�I;�#I;&(I;�,I;�0I;�4I;98I;4;I;�=I;^?I;�@I;      �VI;NVI;�TI;�RI;�OI;�KI;BGI;3BI;�<I;7I;%1I;!+I;A%I;~I;�I;�I;�I;�
I;�I;�I;>�H;�H;�H;~�H;;�H;I�H;s�H;��H;��H;��H;��H;��H;K�H;��H;��H;J�H;P�H;J�H;��H;��H;K�H;��H;��H;��H;��H;��H;s�H;I�H;;�H;~�H;�H;�H;>�H;�I;�I;�
I;�I;�I;�I;~I;A%I;!+I;%1I;7I;�<I;3BI;BGI;�KI;�OI;�RI;�TI;NVI;      �uI;�tI;�rI;�oI;�kI;�fI;�`I;�YI;�RI;&KI;~CI;�;I;-4I;�,I;�%I;�I;zI;�I;YI;hI;�I; I;��H;��H;��H;6�H;1�H;d�H;��H;��H;��H;��H;��H;c�H;�H;��H;��H;��H;�H;c�H;��H;��H;��H;��H;��H;d�H;1�H;6�H;��H;��H;��H; I;�I;hI;YI;�I;zI;�I;�%I;�,I;-4I;�;I;~CI;&KI;�RI;�YI;�`I;�fI;�kI;�oI;�rI;�tI;      ��I;ĝI;o�I;m�I;ّI;��I;ւI;�yI;*pI;%fI;�[I;�QI;�GI;>I;�4I;9,I;�#I;�I;�I;�I;1
I;9I;� I;�H;��H;��H;@�H;-�H;a�H;��H;��H;��H;��H;"�H;��H;��H;c�H;��H;��H;"�H;��H;��H;��H;��H;a�H;-�H;@�H;��H;��H;�H;� I;9I;1
I;�I;�I;�I;�#I;9,I;�4I;>I;�GI;�QI;�[I;%fI;*pI;�yI;ւI;��I;ّI;m�I;o�I;ĝI;      ��I;4�I;{�I;k�I;��I;��I;��I;��I;a�I;�I;k|I;�nI;uaI;�TI;�HI;n=I;�2I;W)I;� I;�I;�I;�I;MI;�I;t�H;��H;��H;M�H;8�H;a�H;��H;��H;��H;�H;��H;<�H;5�H;<�H;��H;�H;��H;��H;��H;a�H;8�H;M�H;��H;��H;t�H;�I;MI;�I;�I;�I;� I;W)I;�2I;n=I;�HI;�TI;uaI;�nI;k|I;�I;a�I;��I;��I;��I;��I;k�I;{�I;4�I;      ��I;�I;��I;��I;L�I;?�I; �I;��I;:�I;��I;�I;��I;��I;!rI;+bI;SSI;�EI;z9I;M.I;K$I;vI;�I;I;*I;I;��H;2�H;�H;M�H;-�H;d�H;��H;��H;�H;b�H;�H;��H;�H;b�H;�H;��H;��H;d�H;-�H;M�H;�H;2�H;��H;I;*I;I;�I;vI;K$I;M.I;z9I;�EI;SSI;+bI;!rI;��I;��I;�I;��I;:�I;��I; �I;?�I;L�I;��I;��I;�I;      s�H;.I;WI;Z6I;
YI;�|I;)�I;%�I;1�I;��I;��I;��I;��I;��I;%�I;�oI;�]I;�MI;q?I;�2I;}'I;�I;8I;�I;�I;ZI;��H;2�H;��H;@�H;1�H;s�H;%�H;#�H;��H;�H;��H;�H;��H;#�H;%�H;s�H;1�H;@�H;��H;2�H;��H;ZI;�I;�I;8I;�I;}'I;�2I;q?I;�MI;�]I;�oI;%�I;��I;��I;��I;��I;��I;1�I;%�I;)�I;�|I;
YI;Z6I;WI;.I;      uF;��F;�F;� G;}�G;,H;ȄH;9�H;VJI;B�I;��I;�I;��I;	�I;�I;e�I;C|I;ZgI;�TI;xDI;d6I;�)I;EI;+I;sI;�I;ZI;��H;��H;��H;6�H;I�H;��H;j�H;��H;$�H;��H;$�H;��H;j�H;��H;I�H;6�H;��H;��H;��H;ZI;�I;sI;+I;EI;�)I;d6I;xDI;�TI;ZgI;C|I;e�I;�I;	�I;��I;�I;��I;B�I;VJI;9�H;ȄH;,H;}�G;� G;�F;��F;      ��?;@;@�@;?�A;۸B;�C;ABE;�uF;�G;�[H;��H;�lI;��I;"�I;@�I;ɺI;��I;|�I;�oI;tZI;aHI;�8I;+I; I;�I;sI;�I;I;t�H;��H;��H;;�H;d�H;��H;��H;f�H;=�H;f�H;��H;��H;d�H;;�H;��H;��H;t�H;I;�I;sI;�I; I;+I;�8I;aHI;tZI;�oI;|�I;��I;ɺI;@�I;"�I;��I;�lI;��H;�[H;�G;�uF;ABE;�C;۸B;?�A;@�@;@;      T�1;��1;�63;�15;��7;��:;H{=;;P@;q�B;aE;��F;uH;�H;;pI;�I;��I;�I;)�I;m�I;�uI;�^I;�JI;4:I;�+I; I;+I;�I;*I;�I;�H;��H;~�H;4�H;��H;{�H;��H;��H;��H;{�H;��H;4�H;~�H;��H;�H;�I;*I;�I;+I; I;�+I;4:I;�JI;�^I;�uI;m�I;)�I;�I;��I;�I;;pI;�H;uH;��F;aE;q�B;;P@;H{=;��:;��7;�15;�63;��1;      ��;��;=\;VW;�m!;�7';�H-; 93;˳8;3{=;)kA;iyD;��F;/H;�I;�I;��I;��I;��I;��I;�yI;�`I;�KI;4:I;+I;EI;8I;I;MI;� I;��H;�H;w�H;�H;�H;a�H;2�H;a�H;�H;�H;w�H;�H;��H;� I;MI;I;8I;EI;+I;4:I;�KI;�`I;�yI;��I;��I;��I;��I;�I;�I;/H;��F;iyD;)kA;3{=;˳8; 93;�H-;�7';�m!;VW;=\;��;      �m�:���:^I�:�W�:���:,�;�~;�;��$;�F.;*O6;��<;K�A;�
E;)RG;;�H;5lI;��I;d�I;m�I;әI;�zI;�`I;�JI;�8I;�)I;�I;�I;�I;9I; I;�H;��H;{�H; �H;�H;��H;�H; �H;{�H;��H;�H; I;9I;�I;�I;�I;�)I;�8I;�JI;�`I;�zI;әI;m�I;d�I;��I;5lI;;�H;)RG;�
E;K�A;��<;*O6;�F.;��$;�;�~;,�;���:�W�:^I�:���:      ��l8��8�Pu9Ǩ�9��9:"��:�U�:bp�:T� ;F;Nn!;��-;^7;jk>;NC;�tF;mPH;�HI;ճI;��I;ϺI;әI;�yI;�^I;aHI;d6I;}'I;vI;�I;1
I;�I;>�H;��H;��H;�H;��H;��H;��H;�H;��H;��H;>�H;�I;1
I;�I;vI;}'I;d6I;aHI;�^I;�yI;әI;ϺI;��I;ճI;�HI;mPH;�tF;NC;jk>;^7;��-;Nn!;F;T� ;bp�:�U�:"��:��9:Ǩ�9�Pu9��8      �����pj�W�غ:����*�����L��9b�:c��:���:�.;��$;��1;3f;;��A;��E;H;Q4I;X�I;��I;m�I;��I;�uI;tZI;xDI;�2I;K$I;�I;�I;hI;�I;��H;s�H;7�H;��H;��H;��H;7�H;s�H;��H;�I;hI;�I;�I;K$I;�2I;xDI;tZI;�uI;��I;m�I;��I;X�I;Q4I;H;��E;��A;3f;;��1;��$;�.;���:c��:b�:L��9�����*�:���W�غpj���      9�ͻ�ɻ��� e��2��J�]��!��轺����0�9���:LR�:�;�X;1H-;�9;v�@;�[E;��G;Q4I;ճI;d�I;��I;m�I;�oI;�TI;q?I;M.I;� I;�I;YI;�I;�I;6�H;��H;,�H;��H;,�H;��H;6�H;�I;�I;YI;�I;� I;M.I;q?I;�TI;�oI;m�I;��I;d�I;ճI;Q4I;��G;�[E;v�@;�9;1H-;�X;�;LR�:���:�0�9����轺�!�J�]�2�� e������ɻ      jO�$�K��o@�%�.�Ǩ����Hɻ�H��npE���غ0�� ��9o�:�@�:�;�*;��7;�O@;�[E;H;�HI;��I;��I;)�I;|�I;ZgI;�MI;z9I;W)I;�I;�I;�
I;,I;'I;G�H;s�H;��H;s�H;G�H;'I;,I;�
I;�I;�I;W)I;z9I;�MI;ZgI;|�I;)�I;��I;��I;�HI;H;�[E;�O@;��7;�*;�;�@�:o�: ��90����غnpE��H��Hɻ���Ǩ�%�.��o@�$�K�      @L�����R���`����N��XPp�!D�ʨ��G�_���44�;����n8��:^�:ZF;�(;��7;v�@;��E;mPH;5lI;��I;�I;��I;C|I;�]I;�EI;�2I;�#I;zI;�I;		I;(I;� I; �H;h�H; �H;� I;(I;		I;�I;zI;�#I;�2I;�EI;�]I;C|I;��I;�I;��I;5lI;mPH;��E;v�@;��7;�(;ZF;^�:��:�n8;���44�_����G�ʨ�!D�XPp��N��`���R������      ��7�e5���������ϼ��@X���iO����-ɻ��p�zF�m�o��g:^�:ZF;�*;�9;��A;�tF;;�H;�I;��I;ɺI;e�I;�oI;SSI;n=I;9,I;�I;�I;I;pI;�I;�I;� I;�I;�I;pI;I;�I;�I;9,I;n=I;SSI;�oI;e�I;ɺI;��I;�I;;�H;�tF;��A;�9;�*;ZF;^�:�g:m�o�zF⺙�p�-ɻ����iO�@X������ϼ������e5�7�      r��ٷ��40v���a�3�G�P2+�!�����*���0���5��ﻧ��]g��ହ�g:^�:�;1H-;3f;;NC;)RG;�I;�I;@�I;�I;%�I;+bI;�HI;�4I;�%I;�I;PI;�
I;�I;eI;sI;eI;�I;�
I;PI;�I;�%I;�4I;�HI;+bI;%�I;�I;@�I;�I;�I;)RG;NC;3f;;1H-;�;^�:�g:�ହ]g�������5�0��*������!��P2+�3�G���a�40v�ٷ��      ��ս��ѽC�ƽ8����I��$���a�a�'D4�LM���ϼ9����K�����G��]g�m�o���:�@�:�X;��1;jk>;�
E;/H;;pI;"�I;	�I;��I;!rI;�TI;>I;�,I;~I;�I;�I;�	I;/I;MI;/I;�	I;�I;�I;~I;�,I;>I;�TI;!rI;��I;	�I;"�I;;pI;/H;�
E;jk>;��1;�X;�@�:��:m�o�]g��G�������K�9����ϼLM�'D4�a�a�$����I��8���C�ƽ��ѽ      �L+� (���H�������ս�@���%���;V�5���������MS�������zF��n8o�:�;��$;^7;K�A;��F;�H;��I;��I;��I;��I;uaI;�GI;-4I;A%I;II;ZI;I;�	I; 	I;�	I;I;ZI;II;A%I;-4I;�GI;uaI;��I;��I;��I;��I;�H;��F;K�A;^7;��$;�;o�:�n8zF⺧������MS�������5���;V��%���@����ս����H��� (�      �T��f�����z� Zb�(�D��$�����ѽ�I��S�m�!2+��������K��ﻙ�p�;��� ��9LR�:�.;��-;��<;iyD;uH;�lI;�I;��I;��I;�nI;�QI;�;I;!+I;�I;*I;OI;�I;�I;�I;OI;*I;�I;!+I;�;I;�QI;�nI;��I;��I;�I;�lI;uH;iyD;��<;��-;�.;LR�: ��9;�����p��ﻍ�K������!2+�S�m��I����ѽ���$�(�D� Zb���z�f���      >�׾��Ҿž�j��������z�U�H�+��lz�N$��0v�!2+����9���5�-ɻ44�0�����:���:Nn!;*O6;)kA;��F;��H;��I;��I;�I;k|I;�[I;~CI;%1I;�#I;�I;jI;�I;�I;�I;jI;�I;�#I;%1I;~CI;�[I;k|I;�I;��I;��I;��H;��F;)kA;*O6;Nn!;���:���:0��44�-ɻ�5�9�����!2+�0v�N$��lz�+��U�H���z������j��ž��Ҿ      E(��$�b��O������~���`���Yb���'��U�N$��S�m�5����ϼ0�����_�����غ�0�9c��:F;�F.;3{=;aE;�[H;B�I;��I;��I;�I;%fI;&KI;7I;&(I;�I;�I;�I;DI;�I;�I;�I;&(I;7I;&KI;%fI;�I;��I;��I;B�I;�[H;aE;3{=;�F.;F;c��:�0�9��غ_������0����ϼ5��S�m�N$���U���'��Yb��`���~�����O��b���$�      7�}���w�#f���K�o,�{�
�:�׾�����k���'�lz꽥I���;V�LM�*����iO��G�npE����b�:T� ;��$;˳8;q�B;�G;VJI;1�I;:�I;a�I;*pI;�RI;�<I;�,I;%!I;�I;9I;�I;9I;�I;%!I;�,I;�<I;�RI;*pI;a�I;:�I;1�I;VJI;�G;q�B;˳8;��$;T� ;b�:���npE��G��iO�*���LM��;V��I��lz���'���k����:�׾{�
�o,���K�#f���w�      ~�n�������,蒿��w���F�b��Ȱ�����Yb�+����ѽ�%��'D4����@X��ʨ��H���轺L��9bp�:�; 93;;P@;�uF;9�H;%�I;��I;��I;�yI;�YI;3BI;�0I;�$I;eI;�I;@I;�I;eI;�$I;�0I;3BI;�YI;�yI;��I;��I;%�I;9�H;�uF;;P@; 93;�;bp�:L��9�轺�H��ʨ�@X�����'D4��%����ѽ+���Yb����Ȱ�b����F���w�,蒿����n���      .���������㿆�ɿ���ǅ����P�b��:�׾�`��U�H����@��a�a�!����!D�Hɻ�!������U�:�~;�H-;H{=;ABE;ȄH;)�I; �I;��I;ւI;�`I;BGI;�4I;�'I;�I; I;pI; I;�I;�'I;�4I;BGI;�`I;ւI;��I; �I;)�I;ȄH;ABE;H{=;�H-;�~;�U�:�����!�Hɻ!D���!��a�a��@����U�H��`��:�׾b����P�ǅ�������ɿ��㿯���      Ù$��x � ��7���޿m���ǅ����F�{�
��~����z��$���ս$���P2+���ϼXPp����J�]��*�"��:,�;�7';��:;�C;,H;�|I;?�I;��I;��I;�fI;�KI;98I;V*I;E!I;I;GI;I;E!I;V*I;98I;�KI;�fI;��I;��I;?�I;�|I;,H;�C;��:;�7';,�;"��:�*�J�]����XPp���ϼP2+�$�����ս�$���z��~��{�
���F�ǅ��m����޿7�� ���x �      F�Q��K���;�Ù$��;
��޿�����w�o,���澝���(�D������I��3�G�����N��Ǩ�2��:�����9:���:�m!;��7;۸B;}�G;
YI;L�I;��I;ّI;�kI;�OI;4;I;�,I;3#I;�I;�I;�I;3#I;�,I;4;I;�OI;�kI;ّI;��I;L�I;
YI;}�G;۸B;��7;�m!;���:��9::���2��Ǩ��N�����3�G��I������(�D��������o,���w�����޿�;
�Ù$���;��K�      Q����{���d��F�Ù$�7����ɿ,蒿��K�O���j�� Zb�H�8�����a����`���%�.� e��W�غǨ�9�W�:VW;�15;?�A;� G;Z6I;��I;k�I;m�I;�oI;�RI;�=I;�.I;�$I;AI;OI;AI;�$I;�.I;�=I;�RI;�oI;m�I;k�I;��I;Z6I;� G;?�A;�15;VW;�W�:Ǩ�9W�غ e��%�.�`��������a�8���H� Zb��j��O����K�,蒿��ɿ7��Ù$��F���d��{�      ���� P�������d���;� ����㿰���#f�b��ž��z���C�ƽ40v�e5�R����o@����pj��Pu9^I�:=\;�63;@�@;�F;WI;��I;{�I;o�I;�rI;�TI;^?I;0I;&I;, I;MI;, I;&I;0I;^?I;�TI;�rI;o�I;{�I;��I;WI;�F;@�@;�63;=\;^I�:�Pu9pj�����o@�R���e5�40v�C�ƽ����z�žb��#f�������� ����;���d���� P��      �,��^�� P���{��K��x �����n�����w��$���Ҿf��� (���ѽٷ��7����$�K��ɻ����8���:��;��1;@;��F;.I;�I;4�I;ĝI;�tI;NVI;�@I;�0I;�&I;� I;�I;� I;�&I;�0I;�@I;NVI;�tI;ĝI;4�I;�I;.I;��F;@;��1;��;���:��8���ɻ$�K����7�ٷ����ѽ (�f�����Ҿ�$���w�n��������x ��K��{� P��^��      ݶ��O���ά��(�_���7�w�}߿���~,b��V�*l¾Fx�c.���Ž��t�6�����*�?��N�����sx9���:��;��2;T?@;�eF;D�H;��I;��I;9{I;�ZI;�BI;#1I;�$I;�I;�I;NI;�I;�I;�$I;#1I;�BI;�ZI;9{I;��I;��I;D�H;�eF;T?@;��2;��;���:�sx9���N��*�?����6����t���Žc.�Fx�*l¾�V�~,b����}߿w���7�(�_�ά��O���      O���A���}��+Y��3�����$ڿ"����\����(���s��3�9�����p�p�p���<<����e������9|��:�;V$3;io@;yF;��H;�I;�I;�zI;sZI;yBI;�0I;t$I;EI;tI; I;tI;EI;t$I;�0I;yBI;sZI;�zI;�I;�I;��H;yF;io@;V$3;�;|��:���9e�������<<�p��p���p�9����3��s�(�������\�"���$ڿ����3��+Y�}�A���      ά��}�8tf��lG�Ң%��p�*�ʿV����>M����S����d�ɤ�̷�9�d��
��I��@�1���������9���:N;�T4;��@;�F;@�H;�I;ܙI;�xI;�XI;bAI;�/I;�#I;�I;�I;�I;�I;�I;�#I;�/I;bAI;�XI;�xI;ܙI;�I;@�H;�F;��@;�T4;N;���:��9������@�1��I���
�9�d�̷�ɤ��d�S�������>M�V���*�ʿ�p�Ң%��lG�8tf�}�      (�_��+Y��lG�f.�w���꿭���J䂿��5���󾋰��M�N�W��V��-�Q�*�������;i!��g��+󳺐:��:�;e06;��A;uG;I;Z�I;��I;�uI;qVI;�?I;�.I;�"I;�I;'I;�I;'I;�I;�"I;�.I;�?I;qVI;�uI;��I;Z�I;I;uG;��A;e06;�;��:�:+��g��;i!�����*���-�Q�V��W��M�N���������5�J䂿�������w�f.��lG��+Y�      ��7��3�Ң%�w��<����ſ�����\�9����Ͼ����`�3����z����9�z�ἷ���z��8}�ht�I�^:�)�:Ϣ#;��8;��B;ArG;�$I;јI;�I;$qI;7SI;=I;�,I;1!I;oI;I;�I;I;oI;1!I;�,I;=I;7SI;$qI;�I;јI;�$I;ArG;��B;��8;Ϣ#;�)�:I�^:ht��8}��z����z�Ἁ�9��z����`�3�������Ͼ9����\������ſ�<��w�Ң%��3�      w�����p������ſ!��{Ps���1�-r���d���d�}I�҈Ž��}�l*�fC��W�^�RC�f�D�&N๪��:��;�);.6;;KD;e�G;kGI;ΜI;ȎI;�kI;OI;�9I;3*I;9I;�I;�I;KI;�I;�I;9I;3*I;�9I;OI;�kI;ȎI;ΜI;kGI;e�G;KD;.6;;�);��;���:&N�f�D�RC�W�^�fC��l*���}�҈Ž}I��d��d��-r����1�{Ps�!����ſ��꿀p����      }߿�$ڿ*�ʿ�������{Ps�MX:����#l¾�ǆ���7����<5��$�Q�����t��85�������*��8 ȼ:��;��.;��=;�DE;�XH;�gI;G�I;ڇI;GeI;@JI;E6I;a'I;�I;I;�I;�I;�I;I;�I;a'I;E6I;@JI;GeI;ڇI;G�I;�gI;�XH;�DE;��=;��.;��; ȼ:*��8������85��t�����$�Q�<5�������7��ǆ�#l¾���MX:�{Ps��������*�ʿ�$ڿ      ���"��V���J䂿��\���1�����J˾睒�C�N�y��L������c�'���Ҽ �|��z�ko��z��(�&:�N�:˧;�V4;�@;HfF;��H;.�I;A�I;UI;=^I;�DI;&2I;<$I;cI;�I;I;�I;I;�I;cI;<$I;&2I;�DI;=^I;UI;A�I;.�I;��H;HfF;�@;�V4;˧;�N�:(�&:z��ko���z� �|���Ҽc�'����L���y��C�N�睒��J˾�����1���\�J䂿V���"��      ~,b���\��>M���5�9��-r��#l¾睒�"&W��3�<Sؽ�z��fG�����I���?��̻{�-����L��:��;Ͽ&;C{9;�C;�cG;sI;]�I;r�I;ruI;�VI;O?I;�-I;� I;�I;yI;�I;�I;�I;yI;�I;� I;�-I;O?I;�VI;ruI;r�I;]�I;sI;�cG;�C;C{9;Ͽ&;��;L��:���{�-��̻�?��I�����fG��z��<Sؽ�3�"&W�睒�#l¾-r��9����5��>M���\�      �V������������Ͼ�d���ǆ�C�N��3��c�[����\�@��EC��N�o�Ъ	�t숻0�N��9J��:�g;o�/;\�=;bE;2H;�VI;ٜI;�I;�jI;�NI;G9I;)I;=I;�I;I;�I;�
I;�I;I;�I;=I;)I;G9I;�NI;�jI;�I;ٜI;�VI;2H;bE;\�=;o�/;�g;J��:N��90�t숻Ъ	�N�o�EC��@����\�[���cཱ3�C�N��ǆ��d����Ͼ���������      *l¾(��S������������d���7�y��<Sؽ[�� �d�P*�kּI\����'�����S������
�:�Y;�#;Y<7;M�A;2�F;|�H;��I;	�I;րI;	`I;�FI;3I;C$I;�I;�I;vI;i	I;iI;i	I;vI;�I;�I;C$I;3I;�FI;	`I;րI;	�I;��I;|�H;2�F;M�A;Y<7;�#;�Y;�
�:�����S������'�I\��kּP*� �d�[��<Sؽy����7��d���������S���(��      Fx��s��d�M�N�`�3�}I����L����z����\�P*�'�ݼe���j<<��ڻ��V��gt�s�&:���:\B;�;/;oC=;��D;��G;8I;�I;ÓI;4sI;IUI;}>I;�,I;�I;�I;yI;�	I;I;.I;I;�	I;yI;�I;�I;�,I;}>I;IUI;4sI;ÓI;�I;8I;��G;��D;oC=;�;/;\B;���:s�&:�gt���V��ڻj<<�e���'�ݼP*���\��z��L������}I�`�3�M�N��d��s�      c.��3�ɤ�W����҈Ž<5�����fG�@��kּe���:yC�?�W7}�𮼺O�x9���:&	;O�&;�:8;��A;F;ϸH;WxI;��I;�I;PeI;�JI;m6I;�&I;�I;�I;uI;/I;�I;�I;�I;/I;uI;�I;�I;�&I;m6I;�JI;PeI;�I;��I;WxI;ϸH;F;��A;�:8;O�&;&	;���:O�x9𮼺W7}�?�:yC�e���kּ@��fG����<5��҈Ž��W��ɤ��3�      ��Ž9���̷�V���z����}�$�Q�c�'����EC��I\��j<<�?��n����IU�c��:Z��:-�;�&3;��>;�E;�H;};I;�I;ÔI;�uI;�WI;�@I;�.I;� I;�I;I;oI;�I;<I;�I;<I;�I;oI;I;�I;� I;�.I;�@I;�WI;�uI;ÔI;�I;};I;�H;�E;��>;�&3;-�;Z��:c��:IU����n��?�j<<�I\��EC�����c�'�$�Q���}��z��V��̷�9���      ��t���p�9�d�-�Q���9�l*������Ҽ�I��N�o���'��ڻW7}���lH��߄:�k�:��;�.;5<;�nC;^6G;��H;�I;��I;�I;;eI;^KI;7I;�&I;�I;�I;i
I;cI;�I;��H;l�H;��H;�I;cI;i
I;�I;�I;�&I;7I;^KI;;eI;�I;��I;�I;��H;^6G;�nC;5<;�.;��;�k�:�߄:lH���W7}��ڻ��'�N�o��I����Ҽ���l*���9�-�Q�9�d���p�      6��p��
�*���z��fC���t�� �|��?�Ъ	������V�𮼺IU��߄:��:�g;6�+;�9;��A;�eF;w�H;�^I;��I;��I; rI;�UI;�?I;�-I; I;uI;(I;�I;�I;i�H;��H;�H;��H;i�H;�I;�I;(I;uI; I;�-I;�?I;�UI; rI;��I;��I;�^I;w�H;�eF;��A;�9;6�+;�g;��:�߄:IU�𮼺��V����Ъ	��?� �|��t��fC��z��*����
�p�      ���p���I���������W�^�85��z��̻t숻�S��gt�O�x9c��:�k�:�g;z�*;�8;�@; �E;W'H;�7I;ߒI;3�I;o}I;�_I;�GI;�4I;y%I;�I;RI;	I;�I;��H;�H;i�H;��H;i�H;�H;��H;�I;	I;RI;�I;y%I;�4I;�GI;�_I;o}I;3�I;ߒI;�7I;W'H; �E;�@;�8;z�*;�g;�k�:c��:O�x9�gt��S�t숻�̻�z�85�W�^���������I��p��      *�?��<<�@�1�;i!��z�RC����ko��{�-�0򳺯���s�&:���:Z��:��;6�+;�8;W�@;]E;��G;eI;	�I;l�I;P�I;�hI;UOI;";I;�*I;�I;�I;nI;EI;� I;��H;��H;d�H;��H;d�H;��H;��H;� I;EI;nI;�I;�I;�*I;";I;UOI;�hI;P�I;l�I;	�I;eI;��G;]E;W�@;�8;6�+;��;Z��:���:s�&:����0�{�-�ko�����RC��z�;i!�@�1��<<�      �N����������g���8}�f�D����z�����N��9�
�:���:&	;-�;�.;�9;�@;]E;��G;]I;�~I;#�I;g�I;�oI;�UI;�@I;�/I;�!I;�I;I;I;�I;��H;s�H;��H;r�H;��H;r�H;��H;s�H;��H;�I;I;I;�I;�!I;�/I;�@I;�UI;�oI;g�I;#�I;�~I;]I;��G;]E;�@;�9;�.;-�;&	;���:�
�:N��9���z�����f�D��8}��g���������      ��e�����+�ht�&N�*��8(�&:L��:J��:�Y;\B;O�&;�&3;5<;��A; �E;��G;]I;w{I;��I;��I;�tI;�ZI;*EI;�3I;E%I;�I;bI;�I;I;O�H;��H;I�H;��H;��H;1�H;��H;��H;I�H;��H;O�H;I;�I;bI;�I;E%I;�3I;*EI;�ZI;�tI;��I;��I;w{I;]I;��G; �E;��A;5<;�&3;O�&;\B;�Y;J��:L��:(�&:*��8&N�ht�+���e���      �sx9���9��9�:I�^:���: ȼ:�N�:��;�g;�#;�;/;�:8;��>;�nC;�eF;W'H;eI;�~I;��I;ːI;wI;�]I;QHI;�6I;(I;#I;�I;�
I;\I;b�H;]�H;h�H;L�H;��H;��H;��H;��H;��H;L�H;h�H;]�H;b�H;\I;�
I;�I;#I;(I;�6I;QHI;�]I;wI;ːI;��I;�~I;eI;W'H;�eF;�nC;��>;�:8;�;/;�#;�g;��;�N�: ȼ:���:I�^:�:��9���9      ���:|��:���:��:�)�:��;��;˧;Ͽ&;o�/;Y<7;oC=;��A;�E;^6G;w�H;�7I;	�I;#�I;��I;wI;�^I;�II;�8I;*I;I;LI;QI;�I;L I;�H;��H;*�H;M�H;��H;�H;��H;�H;��H;M�H;*�H;��H;�H;L I;�I;QI;LI;I;*I;�8I;�II;�^I;wI;��I;#�I;	�I;�7I;w�H;^6G;�E;��A;oC=;Y<7;o�/;Ͽ&;˧;��;��;�)�:��:���:|��:      ��;�;N;�;Ϣ#;�);��.;�V4;C{9;\�=;M�A;��D;F;�H;��H;�^I;ߒI;l�I;g�I;�tI;�]I;�II;>9I;6+I;VI;�I;gI;�I;4I;��H;�H;F�H;�H;{�H;p�H;��H;b�H;��H;p�H;{�H;�H;F�H;�H;��H;4I;�I;gI;�I;VI;6+I;>9I;�II;�]I;�tI;g�I;l�I;ߒI;�^I;��H;�H;F;��D;M�A;\�=;C{9;�V4;��.;�);Ϣ#;�;N;�;      ��2;V$3;�T4;e06;��8;.6;;��=;�@;�C;bE;2�F;��G;ϸH;};I;�I;��I;3�I;P�I;�oI;�ZI;QHI;�8I;6+I;�I;5I;2I;iI;�I;Y�H;t�H;q�H;:�H;L�H;��H;��H;i�H;�H;i�H;��H;��H;L�H;:�H;q�H;t�H;Y�H;�I;iI;2I;5I;�I;6+I;�8I;QHI;�ZI;�oI;P�I;3�I;��I;�I;};I;ϸH;��G;2�F;bE;�C;�@;��=;.6;;��8;e06;�T4;V$3;      T?@;io@;��@;��A;��B;KD;�DE;HfF;�cG;2H;|�H;8I;WxI;�I;��I;��I;o}I;�hI;�UI;*EI;�6I;*I;VI;5I;tI;�I;QI;��H;��H;��H;.�H;0�H;��H;}�H;��H;,�H;	�H;,�H;��H;}�H;��H;0�H;.�H;��H;��H;��H;QI;�I;tI;5I;VI;*I;�6I;*EI;�UI;�hI;o}I;��I;��I;�I;WxI;8I;|�H;2H;�cG;HfF;�DE;KD;��B;��A;��@;io@;      �eF;yF;�F;uG;ArG;e�G;�XH;��H;sI;�VI;��I;�I;��I;ÔI;�I; rI;�_I;UOI;�@I;�3I;(I;I;�I;2I;�I;jI;��H;�H;��H;b�H;?�H;q�H;#�H;9�H;|�H;�H;�H;�H;|�H;9�H;#�H;q�H;?�H;b�H;��H;�H;��H;jI;�I;2I;�I;I;(I;�3I;�@I;UOI;�_I; rI;�I;ÔI;��I;�I;��I;�VI;sI;��H;�XH;e�G;ArG;uG;�F;yF;      D�H;��H;@�H;I;�$I;kGI;�gI;.�I;]�I;ٜI;	�I;ÓI;�I;�uI;;eI;�UI;�GI;";I;�/I;E%I;#I;LI;gI;iI;QI;��H;�H;��H;s�H;@�H;{�H; �H;��H;�H;q�H;�H;�H;�H;q�H;�H;��H; �H;{�H;@�H;s�H;��H;�H;��H;QI;iI;gI;LI;#I;E%I;�/I;";I;�GI;�UI;;eI;�uI;�I;ÓI;	�I;ٜI;]�I;.�I;�gI;kGI;�$I;I;@�H;��H;      ��I;�I;�I;Z�I;јI;ΜI;G�I;A�I;r�I;�I;րI;4sI;PeI;�WI;^KI;�?I;�4I;�*I;�!I;�I;�I;QI;�I;�I;��H;�H;��H;k�H;Q�H;j�H;��H;��H;��H;�H;��H;H�H;1�H;H�H;��H;�H;��H;��H;��H;j�H;Q�H;k�H;��H;�H;��H;�I;�I;QI;�I;�I;�!I;�*I;�4I;�?I;^KI;�WI;PeI;4sI;րI;�I;r�I;A�I;G�I;ΜI;јI;Z�I;�I;�I;      ��I;�I;ܙI;��I;�I;ȎI;ڇI;UI;ruI;�jI;	`I;IUI;�JI;�@I;7I;�-I;y%I;�I;�I;bI;�
I;�I;4I;Y�H;��H;��H;s�H;Q�H;j�H;��H;��H;��H;��H;-�H;��H;��H;Y�H;��H;��H;-�H;��H;��H;��H;��H;j�H;Q�H;s�H;��H;��H;Y�H;4I;�I;�
I;bI;�I;�I;y%I;�-I;7I;�@I;�JI;IUI;	`I;�jI;ruI;UI;ڇI;ȎI;�I;��I;ܙI;�I;      9{I;�zI;�xI;�uI;$qI;�kI;GeI;=^I;�VI;�NI;�FI;}>I;m6I;�.I;�&I; I;�I;�I;I;�I;\I;L I;��H;t�H;��H;b�H;@�H;j�H;��H;��H;��H;��H;�H;��H;�H;��H;��H;��H;�H;��H;�H;��H;��H;��H;��H;j�H;@�H;b�H;��H;t�H;��H;L I;\I;�I;I;�I;�I; I;�&I;�.I;m6I;}>I;�FI;�NI;�VI;=^I;GeI;�kI;$qI;�uI;�xI;�zI;      �ZI;sZI;�XI;qVI;7SI;OI;@JI;�DI;O?I;G9I;3I;�,I;�&I;� I;�I;uI;RI;nI;I;I;b�H;�H;�H;q�H;.�H;?�H;{�H;��H;��H;��H;��H;��H;_�H;��H;|�H;c�H;Z�H;c�H;|�H;��H;_�H;��H;��H;��H;��H;��H;{�H;?�H;.�H;q�H;�H;�H;b�H;I;I;nI;RI;uI;�I;� I;�&I;�,I;3I;G9I;O?I;�DI;@JI;OI;7SI;qVI;�XI;sZI;      �BI;yBI;bAI;�?I;=I;�9I;E6I;&2I;�-I;)I;C$I;�I;�I;�I;�I;(I;	I;EI;�I;O�H;]�H;��H;F�H;:�H;0�H;q�H; �H;��H;��H;��H;��H;I�H;��H;U�H;�H;��H;��H;��H;�H;U�H;��H;I�H;��H;��H;��H;��H; �H;q�H;0�H;:�H;F�H;��H;]�H;O�H;�I;EI;	I;(I;�I;�I;�I;�I;C$I;)I;�-I;&2I;E6I;�9I;=I;�?I;bAI;yBI;      #1I;�0I;�/I;�.I;�,I;3*I;a'I;<$I;� I;=I;�I;�I;�I;I;i
I;�I;�I;� I;��H;��H;h�H;*�H;�H;L�H;��H;#�H;��H;��H;��H;�H;_�H;��H;9�H;��H;��H;��H;t�H;��H;��H;��H;9�H;��H;_�H;�H;��H;��H;��H;#�H;��H;L�H;�H;*�H;h�H;��H;��H;� I;�I;�I;i
I;I;�I;�I;�I;=I;� I;<$I;a'I;3*I;�,I;�.I;�/I;�0I;      �$I;t$I;�#I;�"I;1!I;9I;�I;cI;�I;�I;�I;yI;uI;oI;cI;�I;��H;��H;s�H;I�H;L�H;M�H;{�H;��H;}�H;9�H;�H;�H;-�H;��H;��H;U�H;��H;��H;b�H;@�H;)�H;@�H;b�H;��H;��H;U�H;��H;��H;-�H;�H;�H;9�H;}�H;��H;{�H;M�H;L�H;I�H;s�H;��H;��H;�I;cI;oI;uI;yI;�I;�I;�I;cI;�I;9I;1!I;�"I;�#I;t$I;      �I;EI;�I;�I;oI;�I;I;�I;yI;I;vI;�	I;/I;�I;�I;i�H;�H;��H;��H;��H;��H;��H;p�H;��H;��H;|�H;q�H;��H;��H;�H;|�H;�H;��H;b�H;�H;�H;�H;�H;�H;b�H;��H;�H;|�H;�H;��H;��H;q�H;|�H;��H;��H;p�H;��H;��H;��H;��H;��H;�H;i�H;�I;�I;/I;�	I;vI;I;yI;�I;I;�I;oI;�I;�I;EI;      �I;tI;�I;'I;I;�I;�I;I;�I;�I;i	I;I;�I;<I;��H;��H;i�H;d�H;r�H;��H;��H;�H;��H;i�H;,�H;�H;�H;H�H;��H;��H;c�H;��H;��H;@�H;�H;��H;��H;��H;�H;@�H;��H;��H;c�H;��H;��H;H�H;�H;�H;,�H;i�H;��H;�H;��H;��H;r�H;d�H;i�H;��H;��H;<I;�I;I;i	I;�I;�I;I;�I;�I;I;'I;�I;tI;      NI; I;�I;�I;�I;KI;�I;�I;�I;�
I;iI;.I;�I;�I;l�H;�H;��H;��H;��H;1�H;��H;��H;b�H;�H;	�H;�H;�H;1�H;Y�H;��H;Z�H;��H;t�H;)�H;�H;��H;��H;��H;�H;)�H;t�H;��H;Z�H;��H;Y�H;1�H;�H;�H;	�H;�H;b�H;��H;��H;1�H;��H;��H;��H;�H;l�H;�I;�I;.I;iI;�
I;�I;�I;�I;KI;�I;�I;�I; I;      �I;tI;�I;'I;I;�I;�I;I;�I;�I;i	I;I;�I;<I;��H;��H;i�H;d�H;r�H;��H;��H;�H;��H;i�H;,�H;�H;�H;H�H;��H;��H;c�H;��H;��H;@�H;�H;��H;��H;��H;�H;@�H;��H;��H;c�H;��H;��H;H�H;�H;�H;,�H;i�H;��H;�H;��H;��H;r�H;d�H;i�H;��H;��H;<I;�I;I;i	I;�I;�I;I;�I;�I;I;'I;�I;tI;      �I;EI;�I;�I;oI;�I;I;�I;yI;I;vI;�	I;/I;�I;�I;i�H;�H;��H;��H;��H;��H;��H;p�H;��H;��H;|�H;q�H;��H;��H;�H;|�H;�H;��H;b�H;�H;�H;�H;�H;�H;b�H;��H;�H;|�H;�H;��H;��H;q�H;|�H;��H;��H;p�H;��H;��H;��H;��H;��H;�H;i�H;�I;�I;/I;�	I;vI;I;yI;�I;I;�I;oI;�I;�I;EI;      �$I;t$I;�#I;�"I;1!I;9I;�I;cI;�I;�I;�I;yI;uI;oI;cI;�I;��H;��H;s�H;I�H;L�H;M�H;{�H;��H;}�H;9�H;�H;�H;-�H;��H;��H;U�H;��H;��H;b�H;@�H;)�H;@�H;b�H;��H;��H;U�H;��H;��H;-�H;�H;�H;9�H;}�H;��H;{�H;M�H;L�H;I�H;s�H;��H;��H;�I;cI;oI;uI;yI;�I;�I;�I;cI;�I;9I;1!I;�"I;�#I;t$I;      #1I;�0I;�/I;�.I;�,I;3*I;a'I;<$I;� I;=I;�I;�I;�I;I;i
I;�I;�I;� I;��H;��H;h�H;*�H;�H;L�H;��H;#�H;��H;��H;��H;�H;_�H;��H;9�H;��H;��H;��H;t�H;��H;��H;��H;9�H;��H;_�H;�H;��H;��H;��H;#�H;��H;L�H;�H;*�H;h�H;��H;��H;� I;�I;�I;i
I;I;�I;�I;�I;=I;� I;<$I;a'I;3*I;�,I;�.I;�/I;�0I;      �BI;yBI;bAI;�?I;=I;�9I;E6I;&2I;�-I;)I;C$I;�I;�I;�I;�I;(I;	I;EI;�I;O�H;]�H;��H;F�H;:�H;0�H;q�H; �H;��H;��H;��H;��H;I�H;��H;U�H;�H;��H;��H;��H;�H;U�H;��H;I�H;��H;��H;��H;��H; �H;q�H;0�H;:�H;F�H;��H;]�H;O�H;�I;EI;	I;(I;�I;�I;�I;�I;C$I;)I;�-I;&2I;E6I;�9I;=I;�?I;bAI;yBI;      �ZI;sZI;�XI;qVI;7SI;OI;@JI;�DI;O?I;G9I;3I;�,I;�&I;� I;�I;uI;RI;nI;I;I;b�H;�H;�H;q�H;.�H;?�H;{�H;��H;��H;��H;��H;��H;_�H;��H;|�H;c�H;Z�H;c�H;|�H;��H;_�H;��H;��H;��H;��H;��H;{�H;?�H;.�H;q�H;�H;�H;b�H;I;I;nI;RI;uI;�I;� I;�&I;�,I;3I;G9I;O?I;�DI;@JI;OI;7SI;qVI;�XI;sZI;      9{I;�zI;�xI;�uI;$qI;�kI;GeI;=^I;�VI;�NI;�FI;}>I;m6I;�.I;�&I; I;�I;�I;I;�I;\I;L I;��H;t�H;��H;b�H;@�H;j�H;��H;��H;��H;��H;�H;��H;�H;��H;��H;��H;�H;��H;�H;��H;��H;��H;��H;j�H;@�H;b�H;��H;t�H;��H;L I;\I;�I;I;�I;�I; I;�&I;�.I;m6I;}>I;�FI;�NI;�VI;=^I;GeI;�kI;$qI;�uI;�xI;�zI;      ��I;�I;ܙI;��I;�I;ȎI;ڇI;UI;ruI;�jI;	`I;IUI;�JI;�@I;7I;�-I;y%I;�I;�I;bI;�
I;�I;4I;Y�H;��H;��H;s�H;Q�H;j�H;��H;��H;��H;��H;-�H;��H;��H;Y�H;��H;��H;-�H;��H;��H;��H;��H;j�H;Q�H;s�H;��H;��H;Y�H;4I;�I;�
I;bI;�I;�I;y%I;�-I;7I;�@I;�JI;IUI;	`I;�jI;ruI;UI;ڇI;ȎI;�I;��I;ܙI;�I;      ��I;�I;�I;Z�I;јI;ΜI;G�I;A�I;r�I;�I;րI;4sI;PeI;�WI;^KI;�?I;�4I;�*I;�!I;�I;�I;QI;�I;�I;��H;�H;��H;k�H;Q�H;j�H;��H;��H;��H;�H;��H;H�H;1�H;H�H;��H;�H;��H;��H;��H;j�H;Q�H;k�H;��H;�H;��H;�I;�I;QI;�I;�I;�!I;�*I;�4I;�?I;^KI;�WI;PeI;4sI;րI;�I;r�I;A�I;G�I;ΜI;јI;Z�I;�I;�I;      D�H;��H;@�H;I;�$I;kGI;�gI;.�I;]�I;ٜI;	�I;ÓI;�I;�uI;;eI;�UI;�GI;";I;�/I;E%I;#I;LI;gI;iI;QI;��H;�H;��H;s�H;@�H;{�H; �H;��H;�H;q�H;�H;�H;�H;q�H;�H;��H; �H;{�H;@�H;s�H;��H;�H;��H;QI;iI;gI;LI;#I;E%I;�/I;";I;�GI;�UI;;eI;�uI;�I;ÓI;	�I;ٜI;]�I;.�I;�gI;kGI;�$I;I;@�H;��H;      �eF;yF;�F;uG;ArG;e�G;�XH;��H;sI;�VI;��I;�I;��I;ÔI;�I; rI;�_I;UOI;�@I;�3I;(I;I;�I;2I;�I;jI;��H;�H;��H;b�H;?�H;q�H;#�H;9�H;|�H;�H;�H;�H;|�H;9�H;#�H;q�H;?�H;b�H;��H;�H;��H;jI;�I;2I;�I;I;(I;�3I;�@I;UOI;�_I; rI;�I;ÔI;��I;�I;��I;�VI;sI;��H;�XH;e�G;ArG;uG;�F;yF;      T?@;io@;��@;��A;��B;KD;�DE;HfF;�cG;2H;|�H;8I;WxI;�I;��I;��I;o}I;�hI;�UI;*EI;�6I;*I;VI;5I;tI;�I;QI;��H;��H;��H;.�H;0�H;��H;}�H;��H;,�H;	�H;,�H;��H;}�H;��H;0�H;.�H;��H;��H;��H;QI;�I;tI;5I;VI;*I;�6I;*EI;�UI;�hI;o}I;��I;��I;�I;WxI;8I;|�H;2H;�cG;HfF;�DE;KD;��B;��A;��@;io@;      ��2;V$3;�T4;e06;��8;.6;;��=;�@;�C;bE;2�F;��G;ϸH;};I;�I;��I;3�I;P�I;�oI;�ZI;QHI;�8I;6+I;�I;5I;2I;iI;�I;Y�H;t�H;q�H;:�H;L�H;��H;��H;i�H;�H;i�H;��H;��H;L�H;:�H;q�H;t�H;Y�H;�I;iI;2I;5I;�I;6+I;�8I;QHI;�ZI;�oI;P�I;3�I;��I;�I;};I;ϸH;��G;2�F;bE;�C;�@;��=;.6;;��8;e06;�T4;V$3;      ��;�;N;�;Ϣ#;�);��.;�V4;C{9;\�=;M�A;��D;F;�H;��H;�^I;ߒI;l�I;g�I;�tI;�]I;�II;>9I;6+I;VI;�I;gI;�I;4I;��H;�H;F�H;�H;{�H;p�H;��H;b�H;��H;p�H;{�H;�H;F�H;�H;��H;4I;�I;gI;�I;VI;6+I;>9I;�II;�]I;�tI;g�I;l�I;ߒI;�^I;��H;�H;F;��D;M�A;\�=;C{9;�V4;��.;�);Ϣ#;�;N;�;      ���:|��:���:��:�)�:��;��;˧;Ͽ&;o�/;Y<7;oC=;��A;�E;^6G;w�H;�7I;	�I;#�I;��I;wI;�^I;�II;�8I;*I;I;LI;QI;�I;L I;�H;��H;*�H;M�H;��H;�H;��H;�H;��H;M�H;*�H;��H;�H;L I;�I;QI;LI;I;*I;�8I;�II;�^I;wI;��I;#�I;	�I;�7I;w�H;^6G;�E;��A;oC=;Y<7;o�/;Ͽ&;˧;��;��;�)�:��:���:|��:      �sx9���9��9�:I�^:���: ȼ:�N�:��;�g;�#;�;/;�:8;��>;�nC;�eF;W'H;eI;�~I;��I;ːI;wI;�]I;QHI;�6I;(I;#I;�I;�
I;\I;b�H;]�H;h�H;L�H;��H;��H;��H;��H;��H;L�H;h�H;]�H;b�H;\I;�
I;�I;#I;(I;�6I;QHI;�]I;wI;ːI;��I;�~I;eI;W'H;�eF;�nC;��>;�:8;�;/;�#;�g;��;�N�: ȼ:���:I�^:�:��9���9      ��e�����+�ht�&N�*��8(�&:L��:J��:�Y;\B;O�&;�&3;5<;��A; �E;��G;]I;w{I;��I;��I;�tI;�ZI;*EI;�3I;E%I;�I;bI;�I;I;O�H;��H;I�H;��H;��H;1�H;��H;��H;I�H;��H;O�H;I;�I;bI;�I;E%I;�3I;*EI;�ZI;�tI;��I;��I;w{I;]I;��G; �E;��A;5<;�&3;O�&;\B;�Y;J��:L��:(�&:*��8&N�ht�+���e���      �N����������g���8}�f�D����z�����N��9�
�:���:&	;-�;�.;�9;�@;]E;��G;]I;�~I;#�I;g�I;�oI;�UI;�@I;�/I;�!I;�I;I;I;�I;��H;s�H;��H;r�H;��H;r�H;��H;s�H;��H;�I;I;I;�I;�!I;�/I;�@I;�UI;�oI;g�I;#�I;�~I;]I;��G;]E;�@;�9;�.;-�;&	;���:�
�:N��9���z�����f�D��8}��g���������      *�?��<<�@�1�;i!��z�RC����ko��{�-�0򳺯���s�&:���:Z��:��;6�+;�8;W�@;]E;��G;eI;	�I;l�I;P�I;�hI;UOI;";I;�*I;�I;�I;nI;EI;� I;��H;��H;d�H;��H;d�H;��H;��H;� I;EI;nI;�I;�I;�*I;";I;UOI;�hI;P�I;l�I;	�I;eI;��G;]E;W�@;�8;6�+;��;Z��:���:s�&:����0�{�-�ko�����RC��z�;i!�@�1��<<�      ���p���I���������W�^�85��z��̻t숻�S��gt�O�x9c��:�k�:�g;z�*;�8;�@; �E;W'H;�7I;ߒI;3�I;o}I;�_I;�GI;�4I;y%I;�I;RI;	I;�I;��H;�H;i�H;��H;i�H;�H;��H;�I;	I;RI;�I;y%I;�4I;�GI;�_I;o}I;3�I;ߒI;�7I;W'H; �E;�@;�8;z�*;�g;�k�:c��:O�x9�gt��S�t숻�̻�z�85�W�^���������I��p��      6��p��
�*���z��fC���t�� �|��?�Ъ	������V�𮼺IU��߄:��:�g;6�+;�9;��A;�eF;w�H;�^I;��I;��I; rI;�UI;�?I;�-I; I;uI;(I;�I;�I;i�H;��H;�H;��H;i�H;�I;�I;(I;uI; I;�-I;�?I;�UI; rI;��I;��I;�^I;w�H;�eF;��A;�9;6�+;�g;��:�߄:IU�𮼺��V����Ъ	��?� �|��t��fC��z��*����
�p�      ��t���p�9�d�-�Q���9�l*������Ҽ�I��N�o���'��ڻW7}���lH��߄:�k�:��;�.;5<;�nC;^6G;��H;�I;��I;�I;;eI;^KI;7I;�&I;�I;�I;i
I;cI;�I;��H;l�H;��H;�I;cI;i
I;�I;�I;�&I;7I;^KI;;eI;�I;��I;�I;��H;^6G;�nC;5<;�.;��;�k�:�߄:lH���W7}��ڻ��'�N�o��I����Ҽ���l*���9�-�Q�9�d���p�      ��Ž9���̷�V���z����}�$�Q�c�'����EC��I\��j<<�?��n����IU�c��:Z��:-�;�&3;��>;�E;�H;};I;�I;ÔI;�uI;�WI;�@I;�.I;� I;�I;I;oI;�I;<I;�I;<I;�I;oI;I;�I;� I;�.I;�@I;�WI;�uI;ÔI;�I;};I;�H;�E;��>;�&3;-�;Z��:c��:IU����n��?�j<<�I\��EC�����c�'�$�Q���}��z��V��̷�9���      c.��3�ɤ�W����҈Ž<5�����fG�@��kּe���:yC�?�W7}�𮼺O�x9���:&	;O�&;�:8;��A;F;ϸH;WxI;��I;�I;PeI;�JI;m6I;�&I;�I;�I;uI;/I;�I;�I;�I;/I;uI;�I;�I;�&I;m6I;�JI;PeI;�I;��I;WxI;ϸH;F;��A;�:8;O�&;&	;���:O�x9𮼺W7}�?�:yC�e���kּ@��fG����<5��҈Ž��W��ɤ��3�      Fx��s��d�M�N�`�3�}I����L����z����\�P*�'�ݼe���j<<��ڻ��V��gt�s�&:���:\B;�;/;oC=;��D;��G;8I;�I;ÓI;4sI;IUI;}>I;�,I;�I;�I;yI;�	I;I;.I;I;�	I;yI;�I;�I;�,I;}>I;IUI;4sI;ÓI;�I;8I;��G;��D;oC=;�;/;\B;���:s�&:�gt���V��ڻj<<�e���'�ݼP*���\��z��L������}I�`�3�M�N��d��s�      *l¾(��S������������d���7�y��<Sؽ[�� �d�P*�kּI\����'�����S������
�:�Y;�#;Y<7;M�A;2�F;|�H;��I;	�I;րI;	`I;�FI;3I;C$I;�I;�I;vI;i	I;iI;i	I;vI;�I;�I;C$I;3I;�FI;	`I;րI;	�I;��I;|�H;2�F;M�A;Y<7;�#;�Y;�
�:�����S������'�I\��kּP*� �d�[��<Sؽy����7��d���������S���(��      �V������������Ͼ�d���ǆ�C�N��3��c�[����\�@��EC��N�o�Ъ	�t숻0�N��9J��:�g;o�/;\�=;bE;2H;�VI;ٜI;�I;�jI;�NI;G9I;)I;=I;�I;I;�I;�
I;�I;I;�I;=I;)I;G9I;�NI;�jI;�I;ٜI;�VI;2H;bE;\�=;o�/;�g;J��:N��90�t숻Ъ	�N�o�EC��@����\�[���cཱ3�C�N��ǆ��d����Ͼ���������      ~,b���\��>M���5�9��-r��#l¾睒�"&W��3�<Sؽ�z��fG�����I���?��̻{�-����L��:��;Ͽ&;C{9;�C;�cG;sI;]�I;r�I;ruI;�VI;O?I;�-I;� I;�I;yI;�I;�I;�I;yI;�I;� I;�-I;O?I;�VI;ruI;r�I;]�I;sI;�cG;�C;C{9;Ͽ&;��;L��:���{�-��̻�?��I�����fG��z��<Sؽ�3�"&W�睒�#l¾-r��9����5��>M���\�      ���"��V���J䂿��\���1�����J˾睒�C�N�y��L������c�'���Ҽ �|��z�ko��z��(�&:�N�:˧;�V4;�@;HfF;��H;.�I;A�I;UI;=^I;�DI;&2I;<$I;cI;�I;I;�I;I;�I;cI;<$I;&2I;�DI;=^I;UI;A�I;.�I;��H;HfF;�@;�V4;˧;�N�:(�&:z��ko���z� �|���Ҽc�'����L���y��C�N�睒��J˾�����1���\�J䂿V���"��      }߿�$ڿ*�ʿ�������{Ps�MX:����#l¾�ǆ���7����<5��$�Q�����t��85�������*��8 ȼ:��;��.;��=;�DE;�XH;�gI;G�I;ڇI;GeI;@JI;E6I;a'I;�I;I;�I;�I;�I;I;�I;a'I;E6I;@JI;GeI;ڇI;G�I;�gI;�XH;�DE;��=;��.;��; ȼ:*��8������85��t�����$�Q�<5�������7��ǆ�#l¾���MX:�{Ps��������*�ʿ�$ڿ      w�����p������ſ!��{Ps���1�-r���d���d�}I�҈Ž��}�l*�fC��W�^�RC�f�D�&N๪��:��;�);.6;;KD;e�G;kGI;ΜI;ȎI;�kI;OI;�9I;3*I;9I;�I;�I;KI;�I;�I;9I;3*I;�9I;OI;�kI;ȎI;ΜI;kGI;e�G;KD;.6;;�);��;���:&N�f�D�RC�W�^�fC��l*���}�҈Ž}I��d��d��-r����1�{Ps�!����ſ��꿀p����      ��7��3�Ң%�w��<����ſ�����\�9����Ͼ����`�3����z����9�z�ἷ���z��8}�ht�I�^:�)�:Ϣ#;��8;��B;ArG;�$I;јI;�I;$qI;7SI;=I;�,I;1!I;oI;I;�I;I;oI;1!I;�,I;=I;7SI;$qI;�I;јI;�$I;ArG;��B;��8;Ϣ#;�)�:I�^:ht��8}��z����z�Ἁ�9��z����`�3�������Ͼ9����\������ſ�<��w�Ң%��3�      (�_��+Y��lG�f.�w���꿭���J䂿��5���󾋰��M�N�W��V��-�Q�*�������;i!��g��+󳺐:��:�;e06;��A;uG;I;Z�I;��I;�uI;qVI;�?I;�.I;�"I;�I;'I;�I;'I;�I;�"I;�.I;�?I;qVI;�uI;��I;Z�I;I;uG;��A;e06;�;��:�:+��g��;i!�����*���-�Q�V��W��M�N���������5�J䂿�������w�f.��lG��+Y�      ά��}�8tf��lG�Ң%��p�*�ʿV����>M����S����d�ɤ�̷�9�d��
��I��@�1���������9���:N;�T4;��@;�F;@�H;�I;ܙI;�xI;�XI;bAI;�/I;�#I;�I;�I;�I;�I;�I;�#I;�/I;bAI;�XI;�xI;ܙI;�I;@�H;�F;��@;�T4;N;���:��9������@�1��I���
�9�d�̷�ɤ��d�S�������>M�V���*�ʿ�p�Ң%��lG�8tf�}�      O���A���}��+Y��3�����$ڿ"����\����(���s��3�9�����p�p�p���<<����e������9|��:�;V$3;io@;yF;��H;�I;�I;�zI;sZI;yBI;�0I;t$I;EI;tI; I;tI;EI;t$I;�0I;yBI;sZI;�zI;�I;�I;��H;yF;io@;V$3;�;|��:���9e�������<<�p��p���p�9����3��s�(�������\�"���$ڿ����3��+Y�}�A���      �Aq���i���U�A:�@�����6���q���uA�a5�� ��y^Z�����A���]�����d��|",�6��9�Ѻ���9(��:e�;eX4;p�@;�UF;��H;�FI;�aI;2NI;B9I;�(I;=I;�I;�I;�I;�
I;�I;�I;�I;=I;�(I;B9I;2NI;�aI;�FI;��H;�UF;p�@;eX4;e�;(��:���99�Ѻ6��|",��d������]��A�����y^Z�� ��a5�uA�q���6�������@�A:���U���i�      ��i���b�T�O�.5�-i������������q<�����e��[
V�FE	�!���IY�s9�Z����(� S����Ⱥ��:���:(�;L�4;h�@;kgF;��H;4HI;�aI;�MI;�8I;�(I;I;~I;�I;{I;x
I;{I;�I;~I;I;�(I;�8I;�MI;�aI;4HI;��H;kgF;h�@;L�4;(�;���:��:��Ⱥ S���(�Z���s9��IY�!��FE	�[
V��e������q<������������-i�.5�T�O���b�      ��U�T�O�B-?�(�'���F�`欿Y�{�aa/���뾙���I����e���ZN�o5��Ǩ��nH�� ��􊮺ާ":��:��;��5;�_A;ٚF;Z�H;<LI;aI;�LI;�7I;(I;aI;I;`I;&I;&
I;&I;`I;I;aI;(I;�7I;�LI;aI;<LI;Z�H;ٚF;�_A;��5;��;��:ާ":􊮺� ��nH�Ǩ��o5���ZN�e������I�������aa/�Y�{��欿F����(�'�B-?�T�O�      A:�.5�(�'��������dȿ���e$_���Q�Ҿؕ��
�6�����*���`=�P���)��{G��6��A����Q:�:/";�7;�%B;�F;��H;RI;�_I;�JI;C6I;�&I;ZI;7I;�I;�
I;�	I;�
I;�I;7I;ZI;�&I;C6I;�JI;�_I;RI;��H;�F;�%B;�7;/";�:��Q:A���6��{G��)��P���`=��*�����
�6�ؕ��Q�Ҿ��e$_����dȿ�������(�'�.5�      @�-i�������B�ѿf�������q<��:��a����q����Wн齅���'�ib̼�zl�/���X�x��!�:��;
�&;٪9;LC;wLG;�H;]XI;�]I;�GI;4I;�$I;I;(I;�I;�	I;�I;�	I;�I;(I;I;�$I;4I;�GI;�]I;]XI;�H;wLG;LC;٪9;
�&;��;!�:x���X�/���zl�ib̼��'�齅��Wн����q��a���:��q<����f���B�ѿ������-i�      �������F��dȿf���������O���u]׾w���	�I�����A��C�d�v��֮�<RH�Kkλ�$�m5����:mM;˅+;�<;"3D;�G;�I;�]I;�ZI;	DI;I1I;�"I;aI;�I;�I;�I;�I;�I;�I;�I;aI;�"I;I1I;	DI;�ZI;�]I;�I;�G;"3D;�<;˅+;mM;���:m5��$�Kkλ<RH��֮�v�C�d��A�����	�I�w���u]׾����O�����f���dȿF�ῢ��      6��������欿��������O�}x����� ���l���"��ܽ���`=�Ý��l"��R���ۺR��9�=�:�K;��0;͞>;�LE;}"H;�$I;�`I;(VI;�?I;.I;` I;[I;"I;/
I;mI;�I;mI;/
I;"I;[I;` I;.I;�?I;(VI;�`I;�$I;}"H;�LE;͞>;��0;�K;�=�:R��9�ۺ�R��l"����Ý��`=����ܽ��"��l�� �����}x���O��������欿����      q�������Y�{�e$_��q<�������}��w���6�����!��!�h��������� d��.��g_e�SL[���Z:���:�+ ;��5;�A;�UF;̃H;@I;�aI;�PI;;I;e*I;�I;+I;WI;�I;I;LI;I;�I;WI;+I;�I;e*I;;I;�PI;�aI;@I;̃H;�UF;�A;��5;�+ ;���:��Z:SL[�g_e��.��� d��������!�h�!�������6�w���}��������q<�e$_�Y�{�����      uA��q<�aa/����:�u]׾� ��w��>�BE	�����ܽ����3�r�꼰���>",�X��3��6AQ�ٮ�:�L
;�e);ބ:;D?C;?G;|�H;gSI;�^I;KJI;6I;t&I;�I;�I;ZI;�I;�I;�I;�I;�I;ZI;�I;�I;t&I;6I;KJI;�^I;gSI;|�H;?G;D?C;ބ:;�e);�L
;ٮ�:6AQ�3��X��>",�����r�꼠�3�ܽ������BE	�>�w��� ��u]׾�:���aa/��q<�      a5�������Q�Ҿ�a��w����l��6�BE	���Ƚk���aG����z֮�C�W����9�k����V`,:���:�;��1;m�>;^E;L�G;CI;G^I;hYI;ZCI;�0I;V"I;cI;I;#	I;,I;�I;=I;�I;,I;#	I;I;cI;V"I;�0I;ZCI;hYI;G^I;CI;L�G;^E;m�>;��1;�;���:V`,:���9�k����C�W�z֮�����aG�k����ȽBE	��6��l�w����a��Q�Ҿ������      � ���e�����ؕ����q�	�I���"���������k���ZN�c�6¼~�y��$�PR��\� �D�[��:G/;J�&;w8;��A;��F;��H;?I;aI;�QI;;<I;7+I;�I;I;vI;�I;WI;9I;� I;9I;WI;�I;vI;I;�I;7+I;;<I;�QI;aI;?I;��H;��F;��A;w8;J�&;G/;�:D�[�\� �PR���$�~�y�6¼c��ZN�k������������"�	�I���q�ؕ������e��      y^Z�[
V��I�
�6�������ܽ!��ܽ���aG�c��ȼ�)����(����H5� ��/�Z:k�:8R;/&1;��=;ПD;P�G;�H;�WI;:]I;�HI;5I;�%I;�I;�I;�	I;�I;mI;|�H;��H;|�H;mI;�I;�	I;�I;�I;�%I;5I;�HI;:]I;�WI;�H;P�G;ПD;��=;/&1;8R;k�:/�Z: ��H5������(��)���ȼc��aG�ܽ��!���ܽ�����
�6��I�[
V�      ���FE	��������Wн�A����!�h���3����6¼�)��ax/�u�һC�X�%����9���:�=;[e);�_9;�%B;ډF;�|H;�5I;v`I;�TI;�?I;�-I; I;jI;DI;�I;jI;q�H;��H;�H;��H;q�H;jI;�I;DI;jI; I;�-I;�?I;�TI;v`I;�5I;�|H;ډF;�%B;�_9;[e);�=;���:��9%��C�X�u�һax/��)��6¼�����3�!�h��󑽢A���Wн��콹��FE	�      �A��!��e���*��齅�C�d��`=����r��z֮�~�y���(�u�һj^e������f9���:Y�;m0";B�4;�l?;E;��G;��H;�VI;�]I;(JI;�6I;'I;�I;FI;�	I;>I;7 I;��H;��H;V�H;��H;��H;7 I;>I;�	I;FI;�I;'I;�6I;(JI;�]I;�VI;��H;��G;E;�l?;B�4;m0";Y�;���:�f9����j^e�u�һ��(�~�y�z֮�r�꼠���`=�C�d�齅��*��e��!��      �]��IY��ZN��`=���'�v�Ý���������C�W��$����C�X������9�ޚ:���:��;˷0;�<;v�C;HG;�H;�>I;P`I;�SI;^?I;2.I;z I;�I;.I;�I;�I;��H;��H;&�H;��H;&�H;��H;��H;�I;�I;.I;�I;z I;2.I;^?I;�SI;P`I;�>I;�H;HG;v�C;�<;˷0;��;���:�ޚ:�9����C�X�����$�C�W���������Ý�v���'��`=��ZN��IY�      ���s9�o5��P��ib̼�֮����� d�>",����PR��H5�%���f9�ޚ:��:6�;��-;��:;KB;_UF;;JH; I;�[I;G[I;�GI;%5I;<&I;7I;�I;9	I;^I;�H;��H;��H;n�H;�H;n�H;��H;��H;�H;^I;9	I;�I;7I;<&I;%5I;�GI;G[I;�[I; I;;JH;_UF;KB;��:;��-;6�;��:�ޚ:�f9%��H5�PR�����>",�� d�����֮�ib̼P��o5��s9�      �d��Z���Ǩ���)���zl�<RH�l"��.��X��9�k�\� � ����9���:���:6�;�-;�9;j`A;۹E;J�G;��H;#RI;4_I;OI;�;I;�+I;�I;MI;*I;�I;p I;��H;��H;��H;��H;|�H;��H;��H;��H;��H;p I;�I;*I;MI;�I;�+I;�;I;OI;4_I;#RI;��H;J�G;۹E;j`A;�9;�-;6�;���:���:��9 ��\� �9�k�X���.��l"�<RH��zl��)��Ǩ��Z���      |",��(�nH�{G�/��Kkλ�R��g_e�3�����D�[�/�Z:���:Y�;��;��-;�9;�A;�bE;E�G;��H;tFI;`I;�TI;bAI;�0I;#I;�I;I;�I;I;��H;b�H;��H;!�H;,�H;��H;,�H;!�H;��H;b�H;��H;I;�I;I;�I;#I;�0I;bAI;�TI;`I;tFI;��H;E�G;�bE;�A;�9;��-;��;Y�;���:/�Z:D�[����3��g_e��R��Kkλ/��{G�nH��(�      6�� S��� ���6���X��$��ۺSL[�6AQ�V`,:�:k�:�=;m0";˷0;��:;j`A;�bE;�G;��H;�<I;N_I;�XI;FI;5I;�&I;I;�I;
I;�I;��H;�H;6�H;�H;��H;��H;S�H;��H;��H;�H;6�H;�H;��H;�I;
I;�I;I;�&I;5I;FI;�XI;N_I;�<I;��H;�G;�bE;j`A;��:;˷0;m0";�=;k�:�:V`,:6AQ�SL[��ۺ�$��X��6��� �� S��      9�Ѻ��Ⱥ􊮺A��x��m5�R��9��Z:ٮ�:���:G/;8R;[e);B�4;�<;KB;۹E;E�G;��H;�9I;q^I;�ZI;?II;8I;�)I;�I;I;I;vI;$ I;��H;��H;%�H;C�H;�H;F�H;��H;F�H;�H;C�H;%�H;��H;��H;$ I;vI;I;I;�I;�)I;8I;?II;�ZI;q^I;�9I;��H;E�G;۹E;KB;�<;B�4;[e);8R;G/;���:ٮ�:��Z:R��9m5�x��A��􊮺��Ⱥ      ���9��:ާ":��Q:!�:���:�=�:���:�L
;�;J�&;/&1;�_9;�l?;v�C;_UF;J�G;��H;�<I;q^I;1[I;�JI;1:I;�+I;�I;I;�I;�I;`I;��H;L�H;��H;K�H;��H;��H;��H;��H;��H;��H;��H;K�H;��H;L�H;��H;`I;�I;�I;I;�I;�+I;1:I;�JI;1[I;q^I;�<I;��H;J�G;_UF;v�C;�l?;�_9;/&1;J�&;�;�L
;���:�=�:���:!�:��Q:ާ":��:      (��:���:��:�:��;mM;�K;�+ ;�e);��1;w8;��=;�%B;E;HG;;JH;��H;tFI;N_I;�ZI;�JI;�:I;-I;H!I;QI;+I;0I;xI;��H;��H;��H;}�H;��H;.�H;R�H;��H;y�H;��H;R�H;.�H;��H;}�H;��H;��H;��H;xI;0I;+I;QI;H!I;-I;�:I;�JI;�ZI;N_I;tFI;��H;;JH;HG;E;�%B;��=;w8;��1;�e);�+ ;�K;mM;��;�:��:���:      e�;(�;��;/";
�&;˅+;��0;��5;ބ:;m�>;��A;ПD;ډF;��G;�H; I;#RI;`I;�XI;?II;1:I;-I;�!I;I;�I;	I;BI;]�H;��H;j�H;��H;��H;�H;��H; �H;��H;p�H;��H; �H;��H;�H;��H;��H;j�H;��H;]�H;BI;	I;�I;I;�!I;-I;1:I;?II;�XI;`I;#RI; I;�H;��G;ډF;ПD;��A;m�>;ބ:;��5;��0;˅+;
�&;/";��;(�;      eX4;L�4;��5;�7;٪9;�<;͞>;�A;D?C;^E;��F;P�G;�|H;��H;�>I;�[I;4_I;�TI;FI;8I;�+I;H!I;I;9I;v	I;�I; �H;��H;��H;��H;��H;�H;��H;��H;��H;��H;u�H;��H;��H;��H;��H;�H;��H;��H;��H;��H; �H;�I;v	I;9I;I;H!I;�+I;8I;FI;�TI;4_I;�[I;�>I;��H;�|H;P�G;��F;^E;D?C;�A;͞>;�<;٪9;�7;��5;L�4;      p�@;h�@;�_A;�%B;LC;"3D;�LE;�UF;?G;L�G;��H;�H;�5I;�VI;P`I;G[I;OI;bAI;5I;�)I;�I;QI;�I;v	I;I;.�H;D�H;��H;0�H;��H;�H;��H;[�H;��H;��H;��H;r�H;��H;��H;��H;[�H;��H;�H;��H;0�H;��H;D�H;.�H;I;v	I;�I;QI;�I;�)I;5I;bAI;OI;G[I;P`I;�VI;�5I;�H;��H;L�G;?G;�UF;�LE;"3D;LC;�%B;�_A;h�@;      �UF;kgF;ٚF;�F;wLG;�G;}"H;̃H;|�H;CI;?I;�WI;v`I;�]I;�SI;�GI;�;I;�0I;�&I;�I;I;+I;	I;�I;.�H;W�H;'�H;j�H;��H;�H;��H;V�H;L�H;��H;�H;��H;��H;��H;�H;��H;L�H;V�H;��H;�H;��H;j�H;'�H;W�H;.�H;�I;	I;+I;I;�I;�&I;�0I;�;I;�GI;�SI;�]I;v`I;�WI;?I;CI;|�H;̃H;}"H;�G;wLG;�F;ٚF;kgF;      ��H;��H;Z�H;��H;�H;�I;�$I;@I;gSI;G^I;aI;:]I;�TI;(JI;^?I;%5I;�+I;#I;I;I;�I;0I;BI; �H;D�H;'�H;\�H;�H;7�H;|�H;7�H;�H;F�H;��H;@�H;��H;��H;��H;@�H;��H;F�H;�H;7�H;|�H;7�H;�H;\�H;'�H;D�H; �H;BI;0I;�I;I;I;#I;�+I;%5I;^?I;(JI;�TI;:]I;aI;G^I;gSI;@I;�$I;�I;�H;��H;Z�H;��H;      �FI;4HI;<LI;RI;]XI;�]I;�`I;�aI;�^I;hYI;�QI;�HI;�?I;�6I;2.I;<&I;�I;�I;�I;I;�I;xI;]�H;��H;��H;j�H;�H;�H;��H;3�H;�H;�H;p�H;��H;|�H;F�H;@�H;F�H;|�H;��H;p�H;�H;�H;3�H;��H;�H;�H;j�H;��H;��H;]�H;xI;�I;I;�I;�I;�I;<&I;2.I;�6I;�?I;�HI;�QI;hYI;�^I;�aI;�`I;�]I;]XI;RI;<LI;4HI;      �aI;�aI;aI;�_I;�]I;�ZI;(VI;�PI;KJI;ZCI;;<I;5I;�-I;'I;z I;7I;MI;I;
I;vI;`I;��H;��H;��H;0�H;��H;7�H;��H;*�H;�H; �H;B�H;��H;2�H;��H;��H;��H;��H;��H;2�H;��H;B�H; �H;�H;*�H;��H;7�H;��H;0�H;��H;��H;��H;`I;vI;
I;I;MI;7I;z I;'I;�-I;5I;;<I;ZCI;KJI;�PI;(VI;�ZI;�]I;�_I;aI;�aI;      2NI;�MI;�LI;�JI;�GI;	DI;�?I;;I;6I;�0I;7+I;�%I; I;�I;�I;�I;*I;�I;�I;$ I;��H;��H;j�H;��H;��H;�H;|�H;3�H;�H;�H;1�H;��H;��H;��H;H�H;(�H;%�H;(�H;H�H;��H;��H;��H;1�H;�H;�H;3�H;|�H;�H;��H;��H;j�H;��H;��H;$ I;�I;�I;*I;�I;�I;�I; I;�%I;7+I;�0I;6I;;I;�?I;	DI;�GI;�JI;�LI;�MI;      B9I;�8I;�7I;C6I;4I;I1I;.I;e*I;t&I;V"I;�I;�I;jI;FI;.I;9	I;�I;I;��H;��H;L�H;��H;��H;��H;�H;��H;7�H;�H; �H;1�H;��H;��H;d�H;�H;��H;��H;��H;��H;��H;�H;d�H;��H;��H;1�H; �H;�H;7�H;��H;�H;��H;��H;��H;L�H;��H;��H;I;�I;9	I;.I;FI;jI;�I;�I;V"I;t&I;e*I;.I;I1I;4I;C6I;�7I;�8I;      �(I;�(I;(I;�&I;�$I;�"I;` I;�I;�I;cI;I;�I;DI;�	I;�I;^I;p I;��H;�H;��H;��H;}�H;��H;�H;��H;V�H;�H;�H;B�H;��H;��H;{�H;��H;��H;z�H;T�H;>�H;T�H;z�H;��H;��H;{�H;��H;��H;B�H;�H;�H;V�H;��H;�H;��H;}�H;��H;��H;�H;��H;p I;^I;�I;�	I;DI;�I;I;cI;�I;�I;` I;�"I;�$I;�&I;(I;�(I;      =I;I;aI;ZI;I;aI;[I;+I;�I;I;vI;�	I;�I;>I;�I;�H;��H;b�H;6�H;%�H;K�H;��H;�H;��H;[�H;L�H;F�H;p�H;��H;��H;d�H;��H;��H;\�H;�H;�H;�H;�H;�H;\�H;��H;��H;d�H;��H;��H;p�H;F�H;L�H;[�H;��H;�H;��H;K�H;%�H;6�H;b�H;��H;�H;�I;>I;�I;�	I;vI;I;�I;+I;[I;aI;I;ZI;aI;I;      �I;~I;I;7I;(I;�I;"I;WI;ZI;#	I;�I;�I;jI;7 I;��H;��H;��H;��H;�H;C�H;��H;.�H;��H;��H;��H;��H;��H;��H;2�H;��H;�H;��H;\�H; �H;��H;��H;��H;��H;��H; �H;\�H;��H;�H;��H;2�H;��H;��H;��H;��H;��H;��H;.�H;��H;C�H;�H;��H;��H;��H;��H;7 I;jI;�I;�I;#	I;ZI;WI;"I;�I;(I;7I;I;~I;      �I;�I;`I;�I;�I;�I;/
I;�I;�I;,I;WI;mI;q�H;��H;��H;��H;��H;!�H;��H;�H;��H;R�H; �H;��H;��H;�H;@�H;|�H;��H;H�H;��H;z�H;�H;��H;��H;��H;��H;��H;��H;��H;�H;z�H;��H;H�H;��H;|�H;@�H;�H;��H;��H; �H;R�H;��H;�H;��H;!�H;��H;��H;��H;��H;q�H;mI;WI;,I;�I;�I;/
I;�I;�I;�I;`I;�I;      �I;{I;&I;�
I;�	I;�I;mI;I;�I;�I;9I;|�H;��H;��H;&�H;n�H;��H;,�H;��H;F�H;��H;��H;��H;��H;��H;��H;��H;F�H;��H;(�H;��H;T�H;�H;��H;��H;��H;}�H;��H;��H;��H;�H;T�H;��H;(�H;��H;F�H;��H;��H;��H;��H;��H;��H;��H;F�H;��H;,�H;��H;n�H;&�H;��H;��H;|�H;9I;�I;�I;I;mI;�I;�	I;�
I;&I;{I;      �
I;x
I;&
I;�	I;�I;�I;�I;LI;�I;=I;� I;��H;�H;V�H;��H;�H;|�H;��H;S�H;��H;��H;y�H;p�H;u�H;r�H;��H;��H;@�H;��H;%�H;��H;>�H;�H;��H;��H;}�H;��H;}�H;��H;��H;�H;>�H;��H;%�H;��H;@�H;��H;��H;r�H;u�H;p�H;y�H;��H;��H;S�H;��H;|�H;�H;��H;V�H;�H;��H;� I;=I;�I;LI;�I;�I;�I;�	I;&
I;x
I;      �I;{I;&I;�
I;�	I;�I;mI;I;�I;�I;9I;|�H;��H;��H;&�H;n�H;��H;,�H;��H;F�H;��H;��H;��H;��H;��H;��H;��H;F�H;��H;(�H;��H;T�H;�H;��H;��H;��H;}�H;��H;��H;��H;�H;T�H;��H;(�H;��H;F�H;��H;��H;��H;��H;��H;��H;��H;F�H;��H;,�H;��H;n�H;&�H;��H;��H;|�H;9I;�I;�I;I;mI;�I;�	I;�
I;&I;{I;      �I;�I;`I;�I;�I;�I;/
I;�I;�I;,I;WI;mI;q�H;��H;��H;��H;��H;!�H;��H;�H;��H;R�H; �H;��H;��H;�H;@�H;|�H;��H;H�H;��H;z�H;�H;��H;��H;��H;��H;��H;��H;��H;�H;z�H;��H;H�H;��H;|�H;@�H;�H;��H;��H; �H;R�H;��H;�H;��H;!�H;��H;��H;��H;��H;q�H;mI;WI;,I;�I;�I;/
I;�I;�I;�I;`I;�I;      �I;~I;I;7I;(I;�I;"I;WI;ZI;#	I;�I;�I;jI;7 I;��H;��H;��H;��H;�H;C�H;��H;.�H;��H;��H;��H;��H;��H;��H;2�H;��H;�H;��H;\�H; �H;��H;��H;��H;��H;��H; �H;\�H;��H;�H;��H;2�H;��H;��H;��H;��H;��H;��H;.�H;��H;C�H;�H;��H;��H;��H;��H;7 I;jI;�I;�I;#	I;ZI;WI;"I;�I;(I;7I;I;~I;      =I;I;aI;ZI;I;aI;[I;+I;�I;I;vI;�	I;�I;>I;�I;�H;��H;b�H;6�H;%�H;K�H;��H;�H;��H;[�H;L�H;F�H;p�H;��H;��H;d�H;��H;��H;\�H;�H;�H;�H;�H;�H;\�H;��H;��H;d�H;��H;��H;p�H;F�H;L�H;[�H;��H;�H;��H;K�H;%�H;6�H;b�H;��H;�H;�I;>I;�I;�	I;vI;I;�I;+I;[I;aI;I;ZI;aI;I;      �(I;�(I;(I;�&I;�$I;�"I;` I;�I;�I;cI;I;�I;DI;�	I;�I;^I;p I;��H;�H;��H;��H;}�H;��H;�H;��H;V�H;�H;�H;B�H;��H;��H;{�H;��H;��H;z�H;T�H;>�H;T�H;z�H;��H;��H;{�H;��H;��H;B�H;�H;�H;V�H;��H;�H;��H;}�H;��H;��H;�H;��H;p I;^I;�I;�	I;DI;�I;I;cI;�I;�I;` I;�"I;�$I;�&I;(I;�(I;      B9I;�8I;�7I;C6I;4I;I1I;.I;e*I;t&I;V"I;�I;�I;jI;FI;.I;9	I;�I;I;��H;��H;L�H;��H;��H;��H;�H;��H;7�H;�H; �H;1�H;��H;��H;d�H;�H;��H;��H;��H;��H;��H;�H;d�H;��H;��H;1�H; �H;�H;7�H;��H;�H;��H;��H;��H;L�H;��H;��H;I;�I;9	I;.I;FI;jI;�I;�I;V"I;t&I;e*I;.I;I1I;4I;C6I;�7I;�8I;      2NI;�MI;�LI;�JI;�GI;	DI;�?I;;I;6I;�0I;7+I;�%I; I;�I;�I;�I;*I;�I;�I;$ I;��H;��H;j�H;��H;��H;�H;|�H;3�H;�H;�H;1�H;��H;��H;��H;H�H;(�H;%�H;(�H;H�H;��H;��H;��H;1�H;�H;�H;3�H;|�H;�H;��H;��H;j�H;��H;��H;$ I;�I;�I;*I;�I;�I;�I; I;�%I;7+I;�0I;6I;;I;�?I;	DI;�GI;�JI;�LI;�MI;      �aI;�aI;aI;�_I;�]I;�ZI;(VI;�PI;KJI;ZCI;;<I;5I;�-I;'I;z I;7I;MI;I;
I;vI;`I;��H;��H;��H;0�H;��H;7�H;��H;*�H;�H; �H;B�H;��H;2�H;��H;��H;��H;��H;��H;2�H;��H;B�H; �H;�H;*�H;��H;7�H;��H;0�H;��H;��H;��H;`I;vI;
I;I;MI;7I;z I;'I;�-I;5I;;<I;ZCI;KJI;�PI;(VI;�ZI;�]I;�_I;aI;�aI;      �FI;4HI;<LI;RI;]XI;�]I;�`I;�aI;�^I;hYI;�QI;�HI;�?I;�6I;2.I;<&I;�I;�I;�I;I;�I;xI;]�H;��H;��H;j�H;�H;�H;��H;3�H;�H;�H;p�H;��H;|�H;F�H;@�H;F�H;|�H;��H;p�H;�H;�H;3�H;��H;�H;�H;j�H;��H;��H;]�H;xI;�I;I;�I;�I;�I;<&I;2.I;�6I;�?I;�HI;�QI;hYI;�^I;�aI;�`I;�]I;]XI;RI;<LI;4HI;      ��H;��H;Z�H;��H;�H;�I;�$I;@I;gSI;G^I;aI;:]I;�TI;(JI;^?I;%5I;�+I;#I;I;I;�I;0I;BI; �H;D�H;'�H;\�H;�H;7�H;|�H;7�H;�H;F�H;��H;@�H;��H;��H;��H;@�H;��H;F�H;�H;7�H;|�H;7�H;�H;\�H;'�H;D�H; �H;BI;0I;�I;I;I;#I;�+I;%5I;^?I;(JI;�TI;:]I;aI;G^I;gSI;@I;�$I;�I;�H;��H;Z�H;��H;      �UF;kgF;ٚF;�F;wLG;�G;}"H;̃H;|�H;CI;?I;�WI;v`I;�]I;�SI;�GI;�;I;�0I;�&I;�I;I;+I;	I;�I;.�H;W�H;'�H;j�H;��H;�H;��H;V�H;L�H;��H;�H;��H;��H;��H;�H;��H;L�H;V�H;��H;�H;��H;j�H;'�H;W�H;.�H;�I;	I;+I;I;�I;�&I;�0I;�;I;�GI;�SI;�]I;v`I;�WI;?I;CI;|�H;̃H;}"H;�G;wLG;�F;ٚF;kgF;      p�@;h�@;�_A;�%B;LC;"3D;�LE;�UF;?G;L�G;��H;�H;�5I;�VI;P`I;G[I;OI;bAI;5I;�)I;�I;QI;�I;v	I;I;.�H;D�H;��H;0�H;��H;�H;��H;[�H;��H;��H;��H;r�H;��H;��H;��H;[�H;��H;�H;��H;0�H;��H;D�H;.�H;I;v	I;�I;QI;�I;�)I;5I;bAI;OI;G[I;P`I;�VI;�5I;�H;��H;L�G;?G;�UF;�LE;"3D;LC;�%B;�_A;h�@;      eX4;L�4;��5;�7;٪9;�<;͞>;�A;D?C;^E;��F;P�G;�|H;��H;�>I;�[I;4_I;�TI;FI;8I;�+I;H!I;I;9I;v	I;�I; �H;��H;��H;��H;��H;�H;��H;��H;��H;��H;u�H;��H;��H;��H;��H;�H;��H;��H;��H;��H; �H;�I;v	I;9I;I;H!I;�+I;8I;FI;�TI;4_I;�[I;�>I;��H;�|H;P�G;��F;^E;D?C;�A;͞>;�<;٪9;�7;��5;L�4;      e�;(�;��;/";
�&;˅+;��0;��5;ބ:;m�>;��A;ПD;ډF;��G;�H; I;#RI;`I;�XI;?II;1:I;-I;�!I;I;�I;	I;BI;]�H;��H;j�H;��H;��H;�H;��H; �H;��H;p�H;��H; �H;��H;�H;��H;��H;j�H;��H;]�H;BI;	I;�I;I;�!I;-I;1:I;?II;�XI;`I;#RI; I;�H;��G;ډF;ПD;��A;m�>;ބ:;��5;��0;˅+;
�&;/";��;(�;      (��:���:��:�:��;mM;�K;�+ ;�e);��1;w8;��=;�%B;E;HG;;JH;��H;tFI;N_I;�ZI;�JI;�:I;-I;H!I;QI;+I;0I;xI;��H;��H;��H;}�H;��H;.�H;R�H;��H;y�H;��H;R�H;.�H;��H;}�H;��H;��H;��H;xI;0I;+I;QI;H!I;-I;�:I;�JI;�ZI;N_I;tFI;��H;;JH;HG;E;�%B;��=;w8;��1;�e);�+ ;�K;mM;��;�:��:���:      ���9��:ާ":��Q:!�:���:�=�:���:�L
;�;J�&;/&1;�_9;�l?;v�C;_UF;J�G;��H;�<I;q^I;1[I;�JI;1:I;�+I;�I;I;�I;�I;`I;��H;L�H;��H;K�H;��H;��H;��H;��H;��H;��H;��H;K�H;��H;L�H;��H;`I;�I;�I;I;�I;�+I;1:I;�JI;1[I;q^I;�<I;��H;J�G;_UF;v�C;�l?;�_9;/&1;J�&;�;�L
;���:�=�:���:!�:��Q:ާ":��:      9�Ѻ��Ⱥ􊮺A��x��m5�R��9��Z:ٮ�:���:G/;8R;[e);B�4;�<;KB;۹E;E�G;��H;�9I;q^I;�ZI;?II;8I;�)I;�I;I;I;vI;$ I;��H;��H;%�H;C�H;�H;F�H;��H;F�H;�H;C�H;%�H;��H;��H;$ I;vI;I;I;�I;�)I;8I;?II;�ZI;q^I;�9I;��H;E�G;۹E;KB;�<;B�4;[e);8R;G/;���:ٮ�:��Z:R��9m5�x��A��􊮺��Ⱥ      6�� S��� ���6���X��$��ۺSL[�6AQ�V`,:�:k�:�=;m0";˷0;��:;j`A;�bE;�G;��H;�<I;N_I;�XI;FI;5I;�&I;I;�I;
I;�I;��H;�H;6�H;�H;��H;��H;S�H;��H;��H;�H;6�H;�H;��H;�I;
I;�I;I;�&I;5I;FI;�XI;N_I;�<I;��H;�G;�bE;j`A;��:;˷0;m0";�=;k�:�:V`,:6AQ�SL[��ۺ�$��X��6��� �� S��      |",��(�nH�{G�/��Kkλ�R��g_e�3�����D�[�/�Z:���:Y�;��;��-;�9;�A;�bE;E�G;��H;tFI;`I;�TI;bAI;�0I;#I;�I;I;�I;I;��H;b�H;��H;!�H;,�H;��H;,�H;!�H;��H;b�H;��H;I;�I;I;�I;#I;�0I;bAI;�TI;`I;tFI;��H;E�G;�bE;�A;�9;��-;��;Y�;���:/�Z:D�[����3��g_e��R��Kkλ/��{G�nH��(�      �d��Z���Ǩ���)���zl�<RH�l"��.��X��9�k�\� � ����9���:���:6�;�-;�9;j`A;۹E;J�G;��H;#RI;4_I;OI;�;I;�+I;�I;MI;*I;�I;p I;��H;��H;��H;��H;|�H;��H;��H;��H;��H;p I;�I;*I;MI;�I;�+I;�;I;OI;4_I;#RI;��H;J�G;۹E;j`A;�9;�-;6�;���:���:��9 ��\� �9�k�X���.��l"�<RH��zl��)��Ǩ��Z���      ���s9�o5��P��ib̼�֮����� d�>",����PR��H5�%���f9�ޚ:��:6�;��-;��:;KB;_UF;;JH; I;�[I;G[I;�GI;%5I;<&I;7I;�I;9	I;^I;�H;��H;��H;n�H;�H;n�H;��H;��H;�H;^I;9	I;�I;7I;<&I;%5I;�GI;G[I;�[I; I;;JH;_UF;KB;��:;��-;6�;��:�ޚ:�f9%��H5�PR�����>",�� d�����֮�ib̼P��o5��s9�      �]��IY��ZN��`=���'�v�Ý���������C�W��$����C�X������9�ޚ:���:��;˷0;�<;v�C;HG;�H;�>I;P`I;�SI;^?I;2.I;z I;�I;.I;�I;�I;��H;��H;&�H;��H;&�H;��H;��H;�I;�I;.I;�I;z I;2.I;^?I;�SI;P`I;�>I;�H;HG;v�C;�<;˷0;��;���:�ޚ:�9����C�X�����$�C�W���������Ý�v���'��`=��ZN��IY�      �A��!��e���*��齅�C�d��`=����r��z֮�~�y���(�u�һj^e������f9���:Y�;m0";B�4;�l?;E;��G;��H;�VI;�]I;(JI;�6I;'I;�I;FI;�	I;>I;7 I;��H;��H;V�H;��H;��H;7 I;>I;�	I;FI;�I;'I;�6I;(JI;�]I;�VI;��H;��G;E;�l?;B�4;m0";Y�;���:�f9����j^e�u�һ��(�~�y�z֮�r�꼠���`=�C�d�齅��*��e��!��      ���FE	��������Wн�A����!�h���3����6¼�)��ax/�u�һC�X�%����9���:�=;[e);�_9;�%B;ډF;�|H;�5I;v`I;�TI;�?I;�-I; I;jI;DI;�I;jI;q�H;��H;�H;��H;q�H;jI;�I;DI;jI; I;�-I;�?I;�TI;v`I;�5I;�|H;ډF;�%B;�_9;[e);�=;���:��9%��C�X�u�һax/��)��6¼�����3�!�h��󑽢A���Wн��콹��FE	�      y^Z�[
V��I�
�6�������ܽ!��ܽ���aG�c��ȼ�)����(����H5� ��/�Z:k�:8R;/&1;��=;ПD;P�G;�H;�WI;:]I;�HI;5I;�%I;�I;�I;�	I;�I;mI;|�H;��H;|�H;mI;�I;�	I;�I;�I;�%I;5I;�HI;:]I;�WI;�H;P�G;ПD;��=;/&1;8R;k�:/�Z: ��H5������(��)���ȼc��aG�ܽ��!���ܽ�����
�6��I�[
V�      � ���e�����ؕ����q�	�I���"���������k���ZN�c�6¼~�y��$�PR��\� �D�[��:G/;J�&;w8;��A;��F;��H;?I;aI;�QI;;<I;7+I;�I;I;vI;�I;WI;9I;� I;9I;WI;�I;vI;I;�I;7+I;;<I;�QI;aI;?I;��H;��F;��A;w8;J�&;G/;�:D�[�\� �PR���$�~�y�6¼c��ZN�k������������"�	�I���q�ؕ������e��      a5�������Q�Ҿ�a��w����l��6�BE	���Ƚk���aG����z֮�C�W����9�k����V`,:���:�;��1;m�>;^E;L�G;CI;G^I;hYI;ZCI;�0I;V"I;cI;I;#	I;,I;�I;=I;�I;,I;#	I;I;cI;V"I;�0I;ZCI;hYI;G^I;CI;L�G;^E;m�>;��1;�;���:V`,:���9�k����C�W�z֮�����aG�k����ȽBE	��6��l�w����a��Q�Ҿ������      uA��q<�aa/����:�u]׾� ��w��>�BE	�����ܽ����3�r�꼰���>",�X��3��6AQ�ٮ�:�L
;�e);ބ:;D?C;?G;|�H;gSI;�^I;KJI;6I;t&I;�I;�I;ZI;�I;�I;�I;�I;�I;ZI;�I;�I;t&I;6I;KJI;�^I;gSI;|�H;?G;D?C;ބ:;�e);�L
;ٮ�:6AQ�3��X��>",�����r�꼠�3�ܽ������BE	�>�w��� ��u]׾�:���aa/��q<�      q�������Y�{�e$_��q<�������}��w���6�����!��!�h��������� d��.��g_e�SL[���Z:���:�+ ;��5;�A;�UF;̃H;@I;�aI;�PI;;I;e*I;�I;+I;WI;�I;I;LI;I;�I;WI;+I;�I;e*I;;I;�PI;�aI;@I;̃H;�UF;�A;��5;�+ ;���:��Z:SL[�g_e��.��� d��������!�h�!�������6�w���}��������q<�e$_�Y�{�����      6��������欿��������O�}x����� ���l���"��ܽ���`=�Ý��l"��R���ۺR��9�=�:�K;��0;͞>;�LE;}"H;�$I;�`I;(VI;�?I;.I;` I;[I;"I;/
I;mI;�I;mI;/
I;"I;[I;` I;.I;�?I;(VI;�`I;�$I;}"H;�LE;͞>;��0;�K;�=�:R��9�ۺ�R��l"����Ý��`=����ܽ��"��l�� �����}x���O��������欿����      �������F��dȿf���������O���u]׾w���	�I�����A��C�d�v��֮�<RH�Kkλ�$�m5����:mM;˅+;�<;"3D;�G;�I;�]I;�ZI;	DI;I1I;�"I;aI;�I;�I;�I;�I;�I;�I;�I;aI;�"I;I1I;	DI;�ZI;�]I;�I;�G;"3D;�<;˅+;mM;���:m5��$�Kkλ<RH��֮�v�C�d��A�����	�I�w���u]׾����O�����f���dȿF�ῢ��      @�-i�������B�ѿf�������q<��:��a����q����Wн齅���'�ib̼�zl�/���X�x��!�:��;
�&;٪9;LC;wLG;�H;]XI;�]I;�GI;4I;�$I;I;(I;�I;�	I;�I;�	I;�I;(I;I;�$I;4I;�GI;�]I;]XI;�H;wLG;LC;٪9;
�&;��;!�:x���X�/���zl�ib̼��'�齅��Wн����q��a���:��q<����f���B�ѿ������-i�      A:�.5�(�'��������dȿ���e$_���Q�Ҿؕ��
�6�����*���`=�P���)��{G��6��A����Q:�:/";�7;�%B;�F;��H;RI;�_I;�JI;C6I;�&I;ZI;7I;�I;�
I;�	I;�
I;�I;7I;ZI;�&I;C6I;�JI;�_I;RI;��H;�F;�%B;�7;/";�:��Q:A���6��{G��)��P���`=��*�����
�6�ؕ��Q�Ҿ��e$_����dȿ�������(�'�.5�      ��U�T�O�B-?�(�'���F�`欿Y�{�aa/���뾙���I����e���ZN�o5��Ǩ��nH�� ��􊮺ާ":��:��;��5;�_A;ٚF;Z�H;<LI;aI;�LI;�7I;(I;aI;I;`I;&I;&
I;&I;`I;I;aI;(I;�7I;�LI;aI;<LI;Z�H;ٚF;�_A;��5;��;��:ާ":􊮺� ��nH�Ǩ��o5���ZN�e������I�������aa/�Y�{��欿F����(�'�B-?�T�O�      ��i���b�T�O�.5�-i������������q<�����e��[
V�FE	�!���IY�s9�Z����(� S����Ⱥ��:���:(�;L�4;h�@;kgF;��H;4HI;�aI;�MI;�8I;�(I;I;~I;�I;{I;x
I;{I;�I;~I;I;�(I;�8I;�MI;�aI;4HI;��H;kgF;h�@;L�4;(�;���:��:��Ⱥ S���(�Z���s9��IY�!��FE	�[
V��e������q<������������-i�.5�T�O���b�      �>���8���*�O������˿�o��<�b�=\�+m־^��K�:��J�&��F�B�F���������/��������>:�r�:eo ;�I6;DA;�HF;�MH;�H;!I;�I;I;�I;mI;I;q�H;��H;+�H;��H;q�H;I;mI;�I;I;�I;!I;�H;�MH;�HF;DA;�I6;eo ;�r�:��>:�����/���������F��F�B�&���J�K�:�^��+m־=\�<�b��o���˿����O���*���8�      ��8��4��g&�0��2����<ƿ벗��>]����G�Ѿ�p���*7����"W��MR?�	}�8����s������9�G:���: !;&�6;(kA;�XF;�SH;s�H;!I;�I;�I;�I;FI;�I;e�H;��H;�H;��H;e�H;�I;FI;�I;�I;�I;!I;s�H;�SH;�XF;(kA;&�6; !;���:9�G:���s�����8��	}�MR?�"W�����*7��p��G�Ѿ����>]�벗��<ƿ2���0���g&��4�      ��*��g&��#�o�K[�jL�������M�l5��>ľ
����,��D�撐��5�;�ݼ���q
���x��wk���b:�j�:#;ۖ7;��A;�F;�cH;�I;\!I;I;oI;BI;�I;�I;!�H;x�H;��H;x�H;!�H;�I;�I;BI;oI;I;\!I;�I;�cH;�F;��A;ۖ7;#;�j�:��b:�wk���x��q
���;�ݼ�5�撐��Dὤ�,�
���>ľl5���M����jL��K[�o��#��g&�      O�0��o����˿:1��-�y���6��z �����)�l�+��ͽ!�����&���˼_�k�q���k�X��� �г�:p�;)&;�9;��B;�F;�|H;�I;f!I;5I;�I;�
I;qI;FI;��H;"�H;��H;"�H;��H;FI;qI;�
I;�I;5I;f!I;�I;�|H;�F;��B;�9;)&;p�;г�:�� �k�X�q���_�k���˼��&�!����ͽ+�)�l������z ���6�-�y�:1���˿���o�0��      ����2���K[忭˿�T��蟉�s�R�����E۾̗����M�~�	������j��3�"d��ɆO���׻c�/��
�����:��	;%*;l;;�iC;�&G;�H;�I;
!I;�I;�I;�	I;�I;� I;I�H;��H; �H;��H;I�H;� I;�I;�	I;�I;�I;
!I;�I;�H;�&G;�iC;l;;%*;��	;���:�
��c�/���׻ɆO�"d���3���j����~�	���M�̗���E۾���s�R�蟉��T���˿K[�2���      �˿�<ƿjL��:1��蟉��>]���)��$���ճ���{���,�j��$��Q`I��J��-��4/�S,��˻ ��!69
3�:�;o.;0-=;o`D;�G;o�H;�I;? I;aI;TI;�I;�I;��H;��H;�H;d�H;�H;��H;��H;�I;�I;TI;aI;? I;�I;o�H;�G;o`D;0-=;o.;�;
3�:�!69˻ �S,��4/�-���J��Q`I�$��j�齞�,���{��ճ��$����)��>]�蟉�:1��jL���<ƿ      �o��벗����-�y�s�R���)�iv��>ľ�]����I�Tl�~��������&�߮Ҽ	�}�VB�"���������!:?)�:Vy;�3;li?;�[E;��G;��H;tI;�I;�I;�I;|I;�I;�H;��H;c�H;��H;c�H;��H;�H;�I;|I;�I;�I;�I;tI;��H;��G;�[E;li?;�3;Vy;?)�:��!:����"���VB�	�}�߮Ҽ��&����~���Tl���I��]���>ľiv���)�s�R�-�y����벗�      <�b��>]���M���6�����$���>ľq��q�Z�+�K9ݽW����L����/F��&�G�\�׻�;�u�Ǌ:�h;6O$;�7;y�A;IF;:BH;��H;�I;mI;xI;I;-I;�I;�H;��H;��H;�H;��H;��H;�H;�I;-I;I;xI;mI;�I;��H;:BH;IF;y�A;�7;6O$;�h;Ǌ:u칹;�\�׻&�G�/F�������L�W��K9ݽ+�q�Z�q���>ľ�$�������6���M��>]�      =\����l5��z ��E۾�ճ��]��q�Z�F?#����A����j�(��Oϼ��������Rnۺo3�9�2�:p�;y�,;��;;C�C;�G;Q�H;�
I;� I;�I;GI;.
I;�I;? I;�H;�H;��H;!�H;��H;�H;�H;? I;�I;.
I;GI;�I;� I;�
I;Q�H;�G;C�C;��;;y�,;p�;�2�:o3�9Rnۺ��������Oϼ(����j��A�����F?#�q�Z��]���ճ��E۾�z �l5����      +m־G�Ѿ�>ľ����̗����{���I�+����V���{�?�/�.���,��c=���һ�@�:� ���k:C�:$a;��3;Ai?;w1E;��G;p�H;7I;wI;�I;�I;%I;�I;��H;��H;��H;��H;V�H;��H;��H;��H;��H;�I;%I;�I;�I;wI;7I;p�H;��G;w1E;Ai?;��3;$a;C�:��k::� ��@���һc=��,��.��?�/��{��V�����+���I���{�̗�������>ľG�Ѿ      ^���p��
��)�l���M���,�Tl�K9ݽ�A���{���5��J��;���T[�I?������Q��J�9�:��;:*;5�9;jjB;ۆF;�MH;��H; I;�I;�I;"I;I;@I;_�H;��H;��H;��H;j�H;��H;��H;��H;_�H;@I;I;"I;�I;�I; I;��H;�MH;ۆF;jjB;5�9;:*;��;�:J�9�Q������I?��T[�;���J����5��{��A��K9ݽTl���,���M�)�l�
���p��      K�:��*7���,�+�~�	�j��~���W����j�?�/��J���I��%�k���b.���� ��<Ǌ:�m�:(;nq3;1�>;8�D;t�G;S�H;I;/ I;�I;�I;�	I;�I;`�H;��H;��H;��H;��H;_�H;��H;��H;��H;��H;`�H;�I;�	I;�I;�I;/ I;I;S�H;t�G;8�D;1�>;nq3;(;�m�:<Ǌ: ����b.����%�k��I���J��?�/���j�W��~���j��~�	�+���,��*7�      �J���D��ͽ���$�������L�(��.��;��%�k����I����/��"/�*�>:���:�A;w�,;��:;>�B;�wF;�;H;��H;
I;�I;�I;AI;�I;�I;��H;s�H;5�H;o�H;��H;l�H;��H;o�H;5�H;s�H;��H;�I;�I;AI;�I;�I;
I;��H;�;H;�wF;>�B;��:;w�,;�A;���:*�>:�"/���/��I����%�k�;��.��(����L����$������ͽ�Dὼ��      &��"W��撐�!�����j�Q`I���&����Oϼ�,���T[����I��;��qk�m:i3�:� ;!&;�6;� @;D1E;�G;��H;�I;�I;OI;I;�	I;;I;u�H;��H;�H;��H;^�H;��H;D�H;��H;^�H;��H;�H;��H;u�H;;I;�	I;I;OI;�I;�I;��H;�G;D1E;� @;�6;!&;� ;i3�:m:�qk�;��I�����T[��,��Oϼ�����&�Q`I���j�!���撐�"W��      F�B�MR?��5���&��3��J��߮Ҽ/F����c=�I?�b.����/��qk����9�ճ:�;K!;l3;��=;��C;*�F;cH;��H;�I;I;�I;$I;�I;�I;D�H;��H;��H;|�H;?�H;|�H;3�H;|�H;?�H;|�H;��H;��H;D�H;�I;�I;$I;�I;I;�I;��H;cH;*�F;��C;��=;l3;K!;�;�ճ:���9�qk���/�b.��I?�c=���/F��߮Ҽ�J���3���&��5�MR?�      F��	}�;�ݼ��˼"d��-��	�}�&�G������һ�������"/�m:�ճ:#�;�a;Ģ0;�<;��B;�HF;vH;,�H;�I;yI;I;8I;Y	I;�I;�H;/�H;T�H;�H;#�H;�H;r�H;5�H;r�H;�H;#�H;�H;T�H;/�H;�H;�I;Y	I;8I;I;yI;�I;,�H;vH;�HF;��B;�<;Ģ0;�a;#�;�ճ:m:�"/���������һ���&�G�	�}�-��"d����˼;�ݼ	}�      ����8����_�k�ɆO�4/�VB�\�׻����@��Q�� ��*�>:i3�:�;�a;��/;=;;J�A;��E;ʾG;��H;�	I;hI;I;�I;�I;�I;� I;��H;;�H;��H;��H;��H;�H;d�H;)�H;d�H;�H;��H;��H;��H;;�H;��H;� I;�I;�I;�I;I;hI;�	I;��H;ʾG;��E;J�A;=;;��/;�a;�;i3�:*�>: ���Q���@����\�׻VB�4/�ɆO�_�k���8��      ������q
�q�����׻S,��"����;�Rnۺ:� �J�9<Ǌ:���:� ;K!;Ģ0;=;;͒A;�oE;}�G;ԍH;��H;�I;9I;ZI; I;�I;oI;��H;=�H;x�H;�H;�H;��H;��H;[�H;1�H;[�H;��H;��H;�H;�H;x�H;=�H;��H;oI;�I; I;ZI;9I;�I;��H;ԍH;}�G;�oE;͒A;=;;Ģ0;K!;� ;���:<Ǌ:J�9:� �Rnۺ�;�"���S,����׻q����q
���      �/��s�����x�k�X�c�/�˻ �����u�o3�9��k:�:�m�:�A;!&;l3;�<;J�A;�oE;isG;�{H;.�H;,I;rI;CI;�I;i	I;�I;L�H;I�H;�H;��H;x�H;��H;��H;��H;l�H;\�H;l�H;��H;��H;��H;x�H;��H;�H;I�H;L�H;�I;i	I;�I;CI;rI;,I;.�H;�{H;isG;�oE;J�A;�<;l3;!&;�A;�m�:�:��k:o3�9u칊���˻ �c�/�k�X���x�s���      ��������wk��� ��
���!69��!:Ǌ:�2�:C�:��;(;w�,;�6;��=;��B;��E;}�G;�{H;��H;zI;I;�I;WI;�
I;"I;� I;A�H;��H;4�H;��H;�H;��H;��H;��H;~�H;l�H;~�H;��H;��H;��H;�H;��H;4�H;��H;A�H;� I;"I;�
I;WI;�I;I;zI;��H;�{H;}�G;��E;��B;��=;�6;w�,;(;��;C�:�2�:Ǌ:��!:�!69�
���� ��wk����      ��>:9�G:��b:г�:���:
3�:?)�:�h;p�;$a;:*;nq3;��:;� @;��C;�HF;ʾG;ԍH;.�H;zI;I;CI;9I;�I;I;VI;�H;��H;��H;o�H;B�H;��H;��H;��H;	�H;��H;y�H;��H;	�H;��H;��H;��H;B�H;o�H;��H;��H;�H;VI;I;�I;9I;CI;I;zI;.�H;ԍH;ʾG;�HF;��C;� @;��:;nq3;:*;$a;p�;�h;?)�:
3�:���:г�:��b:9�G:      �r�:���:�j�:p�;��	;�;Vy;6O$;y�,;��3;5�9;1�>;>�B;D1E;*�F;vH;��H;��H;,I;I;CI;�I;6I;�I;�I;��H;�H;G�H;��H;��H;��H;��H;��H;��H;)�H;��H;��H;��H;)�H;��H;��H;��H;��H;��H;��H;G�H;�H;��H;�I;�I;6I;�I;CI;I;,I;��H;��H;vH;*�F;D1E;>�B;1�>;5�9;��3;y�,;6O$;Vy;�;��	;p�;�j�:���:      eo ; !;#;)&;%*;o.;�3;�7;��;;Ai?;jjB;8�D;�wF;�G;cH;,�H;�	I;�I;rI;�I;9I;6I;�I;RI;4�H;��H;��H; �H;��H;�H;��H;x�H;��H;��H;E�H;�H;��H;�H;E�H;��H;��H;x�H;��H;�H;��H; �H;��H;��H;4�H;RI;�I;6I;9I;�I;rI;�I;�	I;,�H;cH;�G;�wF;8�D;jjB;Ai?;��;;�7;�3;o.;%*;)&;#; !;      �I6;&�6;ۖ7;�9;l;;0-=;li?;y�A;C�C;w1E;ۆF;t�G;�;H;��H;��H;�I;hI;9I;CI;WI;�I;�I;RI;E�H;��H;��H;Y�H;$�H;1�H;��H;~�H;e�H;��H;�H;��H;]�H;:�H;]�H;��H;�H;��H;e�H;~�H;��H;1�H;$�H;Y�H;��H;��H;E�H;RI;�I;�I;WI;CI;9I;hI;�I;��H;��H;�;H;t�G;ۆF;w1E;C�C;y�A;li?;0-=;l;;�9;ۖ7;&�6;      DA;(kA;��A;��B;�iC;o`D;�[E;IF;�G;��G;�MH;S�H;��H;�I;�I;yI;I;ZI;�I;�
I;I;�I;4�H;��H;��H;w�H;-�H;@�H;��H;��H;`�H;u�H;��H;O�H;��H;��H;��H;��H;��H;O�H;��H;u�H;`�H;��H;��H;@�H;-�H;w�H;��H;��H;4�H;�I;I;�
I;�I;ZI;I;yI;�I;�I;��H;S�H;�MH;��G;�G;IF;�[E;o`D;�iC;��B;��A;(kA;      �HF;�XF;�F;�F;�&G;�G;��G;:BH;Q�H;p�H;��H;I;
I;�I;I;I;�I; I;i	I;"I;VI;��H;��H;��H;w�H;S�H;Z�H;��H;��H;i�H;X�H;��H;&�H;��H;@�H;"�H;�H;"�H;@�H;��H;&�H;��H;X�H;i�H;��H;��H;Z�H;S�H;w�H;��H;��H;��H;VI;"I;i	I; I;�I;I;I;�I;
I;I;��H;p�H;Q�H;:BH;��G;�G;�&G;�F;�F;�XF;      �MH;�SH;�cH;�|H;�H;o�H;��H;��H;�
I;7I; I;/ I;�I;OI;�I;8I;�I;�I;�I;� I;�H;�H;��H;Y�H;-�H;Z�H;��H;��H;X�H;[�H;��H;��H;d�H;��H;��H;��H;��H;��H;��H;��H;d�H;��H;��H;[�H;X�H;��H;��H;Z�H;-�H;Y�H;��H;�H;�H;� I;�I;�I;�I;8I;�I;OI;�I;/ I; I;7I;�
I;��H;��H;o�H;�H;�|H;�cH;�SH;      �H;s�H;�I;�I;�I;�I;tI;�I;� I;wI;�I;�I;�I;I;$I;Y	I;�I;oI;L�H;A�H;��H;G�H; �H;$�H;@�H;��H;��H;k�H;O�H;��H;��H;;�H;��H;|�H;9�H;
�H;�H;
�H;9�H;|�H;��H;;�H;��H;��H;O�H;k�H;��H;��H;@�H;$�H; �H;G�H;��H;A�H;L�H;oI;�I;Y	I;$I;I;�I;�I;�I;wI;� I;�I;tI;�I;�I;�I;�I;s�H;      !I;!I;\!I;f!I;
!I;? I;�I;mI;�I;�I;�I;�I;AI;�	I;�I;�I;� I;��H;I�H;��H;��H;��H;��H;1�H;��H;��H;X�H;O�H;��H;��H;/�H;��H;M�H;��H;��H;��H;��H;��H;��H;��H;M�H;��H;/�H;��H;��H;O�H;X�H;��H;��H;1�H;��H;��H;��H;��H;I�H;��H;� I;�I;�I;�	I;AI;�I;�I;�I;�I;mI;�I;? I;
!I;f!I;\!I;!I;      �I;�I;I;5I;�I;aI;�I;xI;GI;�I;"I;�	I;�I;;I;�I;�H;��H;=�H;�H;4�H;o�H;��H;�H;��H;��H;i�H;[�H;��H;��H;�H;��H;C�H;��H;��H;g�H;J�H;:�H;J�H;g�H;��H;��H;C�H;��H;�H;��H;��H;[�H;i�H;��H;��H;�H;��H;o�H;4�H;�H;=�H;��H;�H;�I;;I;�I;�	I;"I;�I;GI;xI;�I;aI;�I;5I;I;�I;      I;�I;oI;�I;�I;TI;�I;I;.
I;%I;I;�I;�I;u�H;D�H;/�H;;�H;x�H;��H;��H;B�H;��H;��H;~�H;`�H;X�H;��H;��H;/�H;��H;'�H;��H;v�H;<�H;	�H;��H;��H;��H;	�H;<�H;v�H;��H;'�H;��H;/�H;��H;��H;X�H;`�H;~�H;��H;��H;B�H;��H;��H;x�H;;�H;/�H;D�H;u�H;�I;�I;I;%I;.
I;I;�I;TI;�I;�I;oI;�I;      �I;�I;BI;�
I;�	I;�I;|I;-I;�I;�I;@I;`�H;��H;��H;��H;T�H;��H;�H;x�H;�H;��H;��H;x�H;e�H;u�H;��H;��H;;�H;��H;C�H;��H;R�H;!�H;��H;��H;��H;��H;��H;��H;��H;!�H;R�H;��H;C�H;��H;;�H;��H;��H;u�H;e�H;x�H;��H;��H;�H;x�H;�H;��H;T�H;��H;��H;��H;`�H;@I;�I;�I;-I;|I;�I;�	I;�
I;BI;�I;      mI;FI;�I;qI;�I;�I;�I;�I;? I;��H;_�H;��H;s�H;�H;��H;�H;��H;�H;��H;��H;��H;��H;��H;��H;��H;&�H;d�H;��H;M�H;��H;v�H;!�H;��H;��H;��H;m�H;f�H;m�H;��H;��H;��H;!�H;v�H;��H;M�H;��H;d�H;&�H;��H;��H;��H;��H;��H;��H;��H;�H;��H;�H;��H;�H;s�H;��H;_�H;��H;? I;�I;�I;�I;�I;qI;�I;FI;      I;�I;�I;FI;� I;��H;�H;�H;�H;��H;��H;��H;5�H;��H;|�H;#�H;��H;��H;��H;��H;��H;��H;��H;�H;O�H;��H;��H;|�H;��H;��H;<�H;��H;��H;n�H;V�H;J�H;9�H;J�H;V�H;n�H;��H;��H;<�H;��H;��H;|�H;��H;��H;O�H;�H;��H;��H;��H;��H;��H;��H;��H;#�H;|�H;��H;5�H;��H;��H;��H;�H;�H;�H;��H;� I;FI;�I;�I;      q�H;e�H;!�H;��H;I�H;��H;��H;��H;�H;��H;��H;��H;o�H;^�H;?�H;�H;�H;��H;��H;��H;	�H;)�H;E�H;��H;��H;@�H;��H;9�H;��H;g�H;	�H;��H;��H;V�H;1�H;&�H;(�H;&�H;1�H;V�H;��H;��H;	�H;g�H;��H;9�H;��H;@�H;��H;��H;E�H;)�H;	�H;��H;��H;��H;�H;�H;?�H;^�H;o�H;��H;��H;��H;�H;��H;��H;��H;I�H;��H;!�H;e�H;      ��H;��H;x�H;"�H;��H;�H;c�H;��H;��H;��H;��H;��H;��H;��H;|�H;r�H;d�H;[�H;l�H;~�H;��H;��H;�H;]�H;��H;"�H;��H;
�H;��H;J�H;��H;��H;m�H;J�H;&�H;
�H;�H;
�H;&�H;J�H;m�H;��H;��H;J�H;��H;
�H;��H;"�H;��H;]�H;�H;��H;��H;~�H;l�H;[�H;d�H;r�H;|�H;��H;��H;��H;��H;��H;��H;��H;c�H;�H;��H;"�H;x�H;��H;      +�H;�H;��H;��H; �H;d�H;��H;�H;!�H;V�H;j�H;_�H;l�H;D�H;3�H;5�H;)�H;1�H;\�H;l�H;y�H;��H;��H;:�H;��H;�H;��H;�H;��H;:�H;��H;��H;f�H;9�H;(�H;�H;	�H;�H;(�H;9�H;f�H;��H;��H;:�H;��H;�H;��H;�H;��H;:�H;��H;��H;y�H;l�H;\�H;1�H;)�H;5�H;3�H;D�H;l�H;_�H;j�H;V�H;!�H;�H;��H;d�H; �H;��H;��H;�H;      ��H;��H;x�H;"�H;��H;�H;c�H;��H;��H;��H;��H;��H;��H;��H;|�H;r�H;d�H;[�H;l�H;~�H;��H;��H;�H;]�H;��H;"�H;��H;
�H;��H;J�H;��H;��H;m�H;J�H;&�H;
�H;�H;
�H;&�H;J�H;m�H;��H;��H;J�H;��H;
�H;��H;"�H;��H;]�H;�H;��H;��H;~�H;l�H;[�H;d�H;r�H;|�H;��H;��H;��H;��H;��H;��H;��H;c�H;�H;��H;"�H;x�H;��H;      q�H;e�H;!�H;��H;I�H;��H;��H;��H;�H;��H;��H;��H;o�H;^�H;?�H;�H;�H;��H;��H;��H;	�H;)�H;E�H;��H;��H;@�H;��H;9�H;��H;g�H;	�H;��H;��H;V�H;1�H;&�H;(�H;&�H;1�H;V�H;��H;��H;	�H;g�H;��H;9�H;��H;@�H;��H;��H;E�H;)�H;	�H;��H;��H;��H;�H;�H;?�H;^�H;o�H;��H;��H;��H;�H;��H;��H;��H;I�H;��H;!�H;e�H;      I;�I;�I;FI;� I;��H;�H;�H;�H;��H;��H;��H;5�H;��H;|�H;#�H;��H;��H;��H;��H;��H;��H;��H;�H;O�H;��H;��H;|�H;��H;��H;<�H;��H;��H;n�H;V�H;J�H;9�H;J�H;V�H;n�H;��H;��H;<�H;��H;��H;|�H;��H;��H;O�H;�H;��H;��H;��H;��H;��H;��H;��H;#�H;|�H;��H;5�H;��H;��H;��H;�H;�H;�H;��H;� I;FI;�I;�I;      mI;FI;�I;qI;�I;�I;�I;�I;? I;��H;_�H;��H;s�H;�H;��H;�H;��H;�H;��H;��H;��H;��H;��H;��H;��H;&�H;d�H;��H;M�H;��H;v�H;!�H;��H;��H;��H;m�H;f�H;m�H;��H;��H;��H;!�H;v�H;��H;M�H;��H;d�H;&�H;��H;��H;��H;��H;��H;��H;��H;�H;��H;�H;��H;�H;s�H;��H;_�H;��H;? I;�I;�I;�I;�I;qI;�I;FI;      �I;�I;BI;�
I;�	I;�I;|I;-I;�I;�I;@I;`�H;��H;��H;��H;T�H;��H;�H;x�H;�H;��H;��H;x�H;e�H;u�H;��H;��H;;�H;��H;C�H;��H;R�H;!�H;��H;��H;��H;��H;��H;��H;��H;!�H;R�H;��H;C�H;��H;;�H;��H;��H;u�H;e�H;x�H;��H;��H;�H;x�H;�H;��H;T�H;��H;��H;��H;`�H;@I;�I;�I;-I;|I;�I;�	I;�
I;BI;�I;      I;�I;oI;�I;�I;TI;�I;I;.
I;%I;I;�I;�I;u�H;D�H;/�H;;�H;x�H;��H;��H;B�H;��H;��H;~�H;`�H;X�H;��H;��H;/�H;��H;'�H;��H;v�H;<�H;	�H;��H;��H;��H;	�H;<�H;v�H;��H;'�H;��H;/�H;��H;��H;X�H;`�H;~�H;��H;��H;B�H;��H;��H;x�H;;�H;/�H;D�H;u�H;�I;�I;I;%I;.
I;I;�I;TI;�I;�I;oI;�I;      �I;�I;I;5I;�I;aI;�I;xI;GI;�I;"I;�	I;�I;;I;�I;�H;��H;=�H;�H;4�H;o�H;��H;�H;��H;��H;i�H;[�H;��H;��H;�H;��H;C�H;��H;��H;g�H;J�H;:�H;J�H;g�H;��H;��H;C�H;��H;�H;��H;��H;[�H;i�H;��H;��H;�H;��H;o�H;4�H;�H;=�H;��H;�H;�I;;I;�I;�	I;"I;�I;GI;xI;�I;aI;�I;5I;I;�I;      !I;!I;\!I;f!I;
!I;? I;�I;mI;�I;�I;�I;�I;AI;�	I;�I;�I;� I;��H;I�H;��H;��H;��H;��H;1�H;��H;��H;X�H;O�H;��H;��H;/�H;��H;M�H;��H;��H;��H;��H;��H;��H;��H;M�H;��H;/�H;��H;��H;O�H;X�H;��H;��H;1�H;��H;��H;��H;��H;I�H;��H;� I;�I;�I;�	I;AI;�I;�I;�I;�I;mI;�I;? I;
!I;f!I;\!I;!I;      �H;s�H;�I;�I;�I;�I;tI;�I;� I;wI;�I;�I;�I;I;$I;Y	I;�I;oI;L�H;A�H;��H;G�H; �H;$�H;@�H;��H;��H;k�H;O�H;��H;��H;;�H;��H;|�H;9�H;
�H;�H;
�H;9�H;|�H;��H;;�H;��H;��H;O�H;k�H;��H;��H;@�H;$�H; �H;G�H;��H;A�H;L�H;oI;�I;Y	I;$I;I;�I;�I;�I;wI;� I;�I;tI;�I;�I;�I;�I;s�H;      �MH;�SH;�cH;�|H;�H;o�H;��H;��H;�
I;7I; I;/ I;�I;OI;�I;8I;�I;�I;�I;� I;�H;�H;��H;Y�H;-�H;Z�H;��H;��H;X�H;[�H;��H;��H;d�H;��H;��H;��H;��H;��H;��H;��H;d�H;��H;��H;[�H;X�H;��H;��H;Z�H;-�H;Y�H;��H;�H;�H;� I;�I;�I;�I;8I;�I;OI;�I;/ I; I;7I;�
I;��H;��H;o�H;�H;�|H;�cH;�SH;      �HF;�XF;�F;�F;�&G;�G;��G;:BH;Q�H;p�H;��H;I;
I;�I;I;I;�I; I;i	I;"I;VI;��H;��H;��H;w�H;S�H;Z�H;��H;��H;i�H;X�H;��H;&�H;��H;@�H;"�H;�H;"�H;@�H;��H;&�H;��H;X�H;i�H;��H;��H;Z�H;S�H;w�H;��H;��H;��H;VI;"I;i	I; I;�I;I;I;�I;
I;I;��H;p�H;Q�H;:BH;��G;�G;�&G;�F;�F;�XF;      DA;(kA;��A;��B;�iC;o`D;�[E;IF;�G;��G;�MH;S�H;��H;�I;�I;yI;I;ZI;�I;�
I;I;�I;4�H;��H;��H;w�H;-�H;@�H;��H;��H;`�H;u�H;��H;O�H;��H;��H;��H;��H;��H;O�H;��H;u�H;`�H;��H;��H;@�H;-�H;w�H;��H;��H;4�H;�I;I;�
I;�I;ZI;I;yI;�I;�I;��H;S�H;�MH;��G;�G;IF;�[E;o`D;�iC;��B;��A;(kA;      �I6;&�6;ۖ7;�9;l;;0-=;li?;y�A;C�C;w1E;ۆF;t�G;�;H;��H;��H;�I;hI;9I;CI;WI;�I;�I;RI;E�H;��H;��H;Y�H;$�H;1�H;��H;~�H;e�H;��H;�H;��H;]�H;:�H;]�H;��H;�H;��H;e�H;~�H;��H;1�H;$�H;Y�H;��H;��H;E�H;RI;�I;�I;WI;CI;9I;hI;�I;��H;��H;�;H;t�G;ۆF;w1E;C�C;y�A;li?;0-=;l;;�9;ۖ7;&�6;      eo ; !;#;)&;%*;o.;�3;�7;��;;Ai?;jjB;8�D;�wF;�G;cH;,�H;�	I;�I;rI;�I;9I;6I;�I;RI;4�H;��H;��H; �H;��H;�H;��H;x�H;��H;��H;E�H;�H;��H;�H;E�H;��H;��H;x�H;��H;�H;��H; �H;��H;��H;4�H;RI;�I;6I;9I;�I;rI;�I;�	I;,�H;cH;�G;�wF;8�D;jjB;Ai?;��;;�7;�3;o.;%*;)&;#; !;      �r�:���:�j�:p�;��	;�;Vy;6O$;y�,;��3;5�9;1�>;>�B;D1E;*�F;vH;��H;��H;,I;I;CI;�I;6I;�I;�I;��H;�H;G�H;��H;��H;��H;��H;��H;��H;)�H;��H;��H;��H;)�H;��H;��H;��H;��H;��H;��H;G�H;�H;��H;�I;�I;6I;�I;CI;I;,I;��H;��H;vH;*�F;D1E;>�B;1�>;5�9;��3;y�,;6O$;Vy;�;��	;p�;�j�:���:      ��>:9�G:��b:г�:���:
3�:?)�:�h;p�;$a;:*;nq3;��:;� @;��C;�HF;ʾG;ԍH;.�H;zI;I;CI;9I;�I;I;VI;�H;��H;��H;o�H;B�H;��H;��H;��H;	�H;��H;y�H;��H;	�H;��H;��H;��H;B�H;o�H;��H;��H;�H;VI;I;�I;9I;CI;I;zI;.�H;ԍH;ʾG;�HF;��C;� @;��:;nq3;:*;$a;p�;�h;?)�:
3�:���:г�:��b:9�G:      ��������wk��� ��
���!69��!:Ǌ:�2�:C�:��;(;w�,;�6;��=;��B;��E;}�G;�{H;��H;zI;I;�I;WI;�
I;"I;� I;A�H;��H;4�H;��H;�H;��H;��H;��H;~�H;l�H;~�H;��H;��H;��H;�H;��H;4�H;��H;A�H;� I;"I;�
I;WI;�I;I;zI;��H;�{H;}�G;��E;��B;��=;�6;w�,;(;��;C�:�2�:Ǌ:��!:�!69�
���� ��wk����      �/��s�����x�k�X�c�/�˻ �����u�o3�9��k:�:�m�:�A;!&;l3;�<;J�A;�oE;isG;�{H;.�H;,I;rI;CI;�I;i	I;�I;L�H;I�H;�H;��H;x�H;��H;��H;��H;l�H;\�H;l�H;��H;��H;��H;x�H;��H;�H;I�H;L�H;�I;i	I;�I;CI;rI;,I;.�H;�{H;isG;�oE;J�A;�<;l3;!&;�A;�m�:�:��k:o3�9u칊���˻ �c�/�k�X���x�s���      ������q
�q�����׻S,��"����;�Rnۺ:� �J�9<Ǌ:���:� ;K!;Ģ0;=;;͒A;�oE;}�G;ԍH;��H;�I;9I;ZI; I;�I;oI;��H;=�H;x�H;�H;�H;��H;��H;[�H;1�H;[�H;��H;��H;�H;�H;x�H;=�H;��H;oI;�I; I;ZI;9I;�I;��H;ԍH;}�G;�oE;͒A;=;;Ģ0;K!;� ;���:<Ǌ:J�9:� �Rnۺ�;�"���S,����׻q����q
���      ����8����_�k�ɆO�4/�VB�\�׻����@��Q�� ��*�>:i3�:�;�a;��/;=;;J�A;��E;ʾG;��H;�	I;hI;I;�I;�I;�I;� I;��H;;�H;��H;��H;��H;�H;d�H;)�H;d�H;�H;��H;��H;��H;;�H;��H;� I;�I;�I;�I;I;hI;�	I;��H;ʾG;��E;J�A;=;;��/;�a;�;i3�:*�>: ���Q���@����\�׻VB�4/�ɆO�_�k���8��      F��	}�;�ݼ��˼"d��-��	�}�&�G������һ�������"/�m:�ճ:#�;�a;Ģ0;�<;��B;�HF;vH;,�H;�I;yI;I;8I;Y	I;�I;�H;/�H;T�H;�H;#�H;�H;r�H;5�H;r�H;�H;#�H;�H;T�H;/�H;�H;�I;Y	I;8I;I;yI;�I;,�H;vH;�HF;��B;�<;Ģ0;�a;#�;�ճ:m:�"/���������һ���&�G�	�}�-��"d����˼;�ݼ	}�      F�B�MR?��5���&��3��J��߮Ҽ/F����c=�I?�b.����/��qk����9�ճ:�;K!;l3;��=;��C;*�F;cH;��H;�I;I;�I;$I;�I;�I;D�H;��H;��H;|�H;?�H;|�H;3�H;|�H;?�H;|�H;��H;��H;D�H;�I;�I;$I;�I;I;�I;��H;cH;*�F;��C;��=;l3;K!;�;�ճ:���9�qk���/�b.��I?�c=���/F��߮Ҽ�J���3���&��5�MR?�      &��"W��撐�!�����j�Q`I���&����Oϼ�,���T[����I��;��qk�m:i3�:� ;!&;�6;� @;D1E;�G;��H;�I;�I;OI;I;�	I;;I;u�H;��H;�H;��H;^�H;��H;D�H;��H;^�H;��H;�H;��H;u�H;;I;�	I;I;OI;�I;�I;��H;�G;D1E;� @;�6;!&;� ;i3�:m:�qk�;��I�����T[��,��Oϼ�����&�Q`I���j�!���撐�"W��      �J���D��ͽ���$�������L�(��.��;��%�k����I����/��"/�*�>:���:�A;w�,;��:;>�B;�wF;�;H;��H;
I;�I;�I;AI;�I;�I;��H;s�H;5�H;o�H;��H;l�H;��H;o�H;5�H;s�H;��H;�I;�I;AI;�I;�I;
I;��H;�;H;�wF;>�B;��:;w�,;�A;���:*�>:�"/���/��I����%�k�;��.��(����L����$������ͽ�Dὼ��      K�:��*7���,�+�~�	�j��~���W����j�?�/��J���I��%�k���b.���� ��<Ǌ:�m�:(;nq3;1�>;8�D;t�G;S�H;I;/ I;�I;�I;�	I;�I;`�H;��H;��H;��H;��H;_�H;��H;��H;��H;��H;`�H;�I;�	I;�I;�I;/ I;I;S�H;t�G;8�D;1�>;nq3;(;�m�:<Ǌ: ����b.����%�k��I���J��?�/���j�W��~���j��~�	�+���,��*7�      ^���p��
��)�l���M���,�Tl�K9ݽ�A���{���5��J��;���T[�I?������Q��J�9�:��;:*;5�9;jjB;ۆF;�MH;��H; I;�I;�I;"I;I;@I;_�H;��H;��H;��H;j�H;��H;��H;��H;_�H;@I;I;"I;�I;�I; I;��H;�MH;ۆF;jjB;5�9;:*;��;�:J�9�Q������I?��T[�;���J����5��{��A��K9ݽTl���,���M�)�l�
���p��      +m־G�Ѿ�>ľ����̗����{���I�+����V���{�?�/�.���,��c=���һ�@�:� ���k:C�:$a;��3;Ai?;w1E;��G;p�H;7I;wI;�I;�I;%I;�I;��H;��H;��H;��H;V�H;��H;��H;��H;��H;�I;%I;�I;�I;wI;7I;p�H;��G;w1E;Ai?;��3;$a;C�:��k::� ��@���һc=��,��.��?�/��{��V�����+���I���{�̗�������>ľG�Ѿ      =\����l5��z ��E۾�ճ��]��q�Z�F?#����A����j�(��Oϼ��������Rnۺo3�9�2�:p�;y�,;��;;C�C;�G;Q�H;�
I;� I;�I;GI;.
I;�I;? I;�H;�H;��H;!�H;��H;�H;�H;? I;�I;.
I;GI;�I;� I;�
I;Q�H;�G;C�C;��;;y�,;p�;�2�:o3�9Rnۺ��������Oϼ(����j��A�����F?#�q�Z��]���ճ��E۾�z �l5����      <�b��>]���M���6�����$���>ľq��q�Z�+�K9ݽW����L����/F��&�G�\�׻�;�u�Ǌ:�h;6O$;�7;y�A;IF;:BH;��H;�I;mI;xI;I;-I;�I;�H;��H;��H;�H;��H;��H;�H;�I;-I;I;xI;mI;�I;��H;:BH;IF;y�A;�7;6O$;�h;Ǌ:u칹;�\�׻&�G�/F�������L�W��K9ݽ+�q�Z�q���>ľ�$�������6���M��>]�      �o��벗����-�y�s�R���)�iv��>ľ�]����I�Tl�~��������&�߮Ҽ	�}�VB�"���������!:?)�:Vy;�3;li?;�[E;��G;��H;tI;�I;�I;�I;|I;�I;�H;��H;c�H;��H;c�H;��H;�H;�I;|I;�I;�I;�I;tI;��H;��G;�[E;li?;�3;Vy;?)�:��!:����"���VB�	�}�߮Ҽ��&����~���Tl���I��]���>ľiv���)�s�R�-�y����벗�      �˿�<ƿjL��:1��蟉��>]���)��$���ճ���{���,�j��$��Q`I��J��-��4/�S,��˻ ��!69
3�:�;o.;0-=;o`D;�G;o�H;�I;? I;aI;TI;�I;�I;��H;��H;�H;d�H;�H;��H;��H;�I;�I;TI;aI;? I;�I;o�H;�G;o`D;0-=;o.;�;
3�:�!69˻ �S,��4/�-���J��Q`I�$��j�齞�,���{��ճ��$����)��>]�蟉�:1��jL���<ƿ      ����2���K[忭˿�T��蟉�s�R�����E۾̗����M�~�	������j��3�"d��ɆO���׻c�/��
�����:��	;%*;l;;�iC;�&G;�H;�I;
!I;�I;�I;�	I;�I;� I;I�H;��H; �H;��H;I�H;� I;�I;�	I;�I;�I;
!I;�I;�H;�&G;�iC;l;;%*;��	;���:�
��c�/���׻ɆO�"d���3���j����~�	���M�̗���E۾���s�R�蟉��T���˿K[�2���      O�0��o����˿:1��-�y���6��z �����)�l�+��ͽ!�����&���˼_�k�q���k�X��� �г�:p�;)&;�9;��B;�F;�|H;�I;f!I;5I;�I;�
I;qI;FI;��H;"�H;��H;"�H;��H;FI;qI;�
I;�I;5I;f!I;�I;�|H;�F;��B;�9;)&;p�;г�:�� �k�X�q���_�k���˼��&�!����ͽ+�)�l������z ���6�-�y�:1���˿���o�0��      ��*��g&��#�o�K[�jL�������M�l5��>ľ
����,��D�撐��5�;�ݼ���q
���x��wk���b:�j�:#;ۖ7;��A;�F;�cH;�I;\!I;I;oI;BI;�I;�I;!�H;x�H;��H;x�H;!�H;�I;�I;BI;oI;I;\!I;�I;�cH;�F;��A;ۖ7;#;�j�:��b:�wk���x��q
���;�ݼ�5�撐��Dὤ�,�
���>ľl5���M����jL��K[�o��#��g&�      ��8��4��g&�0��2����<ƿ벗��>]����G�Ѿ�p���*7����"W��MR?�	}�8����s������9�G:���: !;&�6;(kA;�XF;�SH;s�H;!I;�I;�I;�I;FI;�I;e�H;��H;�H;��H;e�H;�I;FI;�I;�I;�I;!I;s�H;�SH;�XF;(kA;&�6; !;���:9�G:���s�����8��	}�MR?�"W�����*7��p��G�Ѿ����>]�벗��<ƿ2���0���g&��4�      ���$������꿥�ſ�ޞ�3s��2�/����� j���nHͽ������'�B<ͼ��n������Q^�0.��:�V;�R%;~n8;��A;nCF;�H;��H;��H;��H;L�H;>�H;C�H;��H;��H;��H;+�H;��H;��H;��H;C�H;>�H;L�H;��H;��H;��H;�H;nCF;��A;~n8;�R%;�V;�:0.��Q^�������n�B<ͼ��'�����nHͽ�� j���/����2�3s��ޞ���ſ������$�      $��������~�����cm�L�-�����Fh��Ide�-�̪ɽ�v��#�$���ɼ�mj�o����X�5��nĆ:�w;i�%;M�8;B;{QF;H;5�H;U�H;	�H;p�H;B�H;6�H;��H;��H;��H;$�H;��H;��H;��H;6�H;B�H;p�H;	�H;U�H;5�H;H;{QF;B;M�8;i�%;�w;nĆ:5���X�o����mj���ɼ#�$��v��̪ɽ-�Ide�Fh������L�-�cm����~���忖����      ������{���ԿBw�����/�\��"����b��M0X�}���;����w����������]�X��UF�,��oȒ:1�;_�';؎9;2oB;�yF;� H;��H;7�H;�H;��H;F�H;:�H;��H;��H;��H;�H;��H;��H;��H;:�H;F�H;��H;�H;7�H;��H;� H;�yF;2oB;؎9;_�';1�;oȒ:,��UF�X�黼�]����������w��;��}��M0X�b������"�/�\����Bw���Կ{�𿖏�      ������Կp���ޞ�RF�]�C�$E��;�I��sD�|�"��]�c�y��֯���J�P�ѻ\�)���K����:Q�
;M*;��:;�C;�F;�7H;Z�H;��H;w�H;��H;>�H;:�H;��H;��H;��H;��H;��H;��H;��H;:�H;>�H;��H;w�H;��H;Z�H;�7H;�F;�C;��:;M*;Q�
;���:��K�\�)�P�ѻ��J��֯�y�]�c�"��|�sD��I���;$E�]�C�RF��ޞ�p���Կ��      ��ſ~��Bw���ޞ�|���3�W�,�%�����^ɰ��|x�\{+�ű����J��  �Ҷ��n�1�f����+�
9r�:�;4�-;��<;��C;�G;�SH;Q�H;��H;��H;��H;V�H;3�H;��H;��H;��H;��H;��H;��H;��H;3�H;V�H;��H;��H;��H;Q�H;�SH;�G;��C;��<;4�-;�;r�:
9�+�f���n�1�Ҷ���  ��J���ű�\{+��|x�^ɰ�����,�%�3�W�|����ޞ�Bw��~��      �ޞ�������RF�3�W�M�-���4Kɾ�G����O�z��ƽ����Ȅ-���ۼㄼL4�[ǐ�,ж��Z:o��:�;ʕ1;
c>;|�D;�[G;KrH;��H;i�H;e�H;'�H;u�H;)�H;h�H;��H;|�H;��H;|�H;��H;h�H;)�H;u�H;'�H;e�H;i�H;��H;KrH;�[G;|�D;
c>;ʕ1;�;o��:�Z:,ж�[ǐ�L4�ㄼ��ۼȄ-�����ƽz����O��G��4Kɾ��M�-�3�W�RF�������      3s�cm�/�\�]�C�,�%����TҾa����i��C(����UP����[�x������Y�k���X���<���k:���:)� ;�5;ZQ@;otE;�G;9�H;L�H;��H;�H;I�H;l�H;$�H;c�H;s�H;X�H;��H;X�H;s�H;c�H;$�H;l�H;I�H;�H;��H;L�H;9�H;�G;otE;ZQ@;�5;)� ;���:��k:��<��X�k����Y����x���[�UP����콡C(���i�a���TҾ��,�%�]�C�/�\�cm�      �2�L�-��"�$E�����4Kɾa��w�s�.�5�y�k㻽�v��z0��;��+��-�*�S����6�"jS�L�:��	;��(;6�9;�.B;�CF;YH;ժH;��H;��H;��H;w�H;��H;�H;0�H;C�H;<�H;Y�H;<�H;C�H;0�H;�H;��H;w�H;��H;��H;��H;ժH;YH;�CF;�.B;6�9;��(;��	;L�:"jS��6�S���-�*��+���;�z0��v��k㻽y�.�5�w�s�a��4Kɾ����$E��"�L�-�      /�����������;^ɰ��G����i�.�5��	�ĪɽR����J�p���沼��]�I���U
x��
���k:5��:v;��/;�,=;��C;N�F;#HH;��H;(�H;��H;#�H;��H;��H;��H;�H;�H;�H;$�H;�H;�H;�H;��H;��H;��H;#�H;��H;(�H;��H;#HH;N�F;��C;�,=;��/;v;5��:�k:�
��U
x�I�����]��沼p���J�R���Īɽ�	�.�5���i��G��^ɰ��;��徨���      ��Fh��b���I���|x���O��C(�y�Īɽ����IDX�D��'<ͼㄼ�X!�t��hX��K����:�x;7�#;$H6;IQ@;�OE;��G;��H;��H;2�H;��H;��H;��H;v�H;��H;��H;��H;��H;��H;��H;��H;��H;��H;v�H;��H;��H;��H;2�H;��H;��H;��G;�OE;IQ@;$H6;7�#;�x;���:�K�hX�t���X!�ㄼ'<ͼD��IDX�����Īɽy��C(���O��|x��I��b��Fh��       j�Ide�M0X�sD�\{+�z�����k㻽R���IDX������ۼо����;�>ۻ�X���y�><":J��:��;��-;��;;�B;�yF;�H;��H;|�H;&�H;��H;��H;��H;n�H;��H;��H;��H;��H;z�H;��H;��H;��H;��H;n�H;��H;��H;��H;&�H;|�H;��H;�H;�yF;�B;��;;��-;��;J��:><":��y��X�>ۻ��;�о����ۼ���IDX�R���k㻽���z��\{+�sD�M0X�Ide�      ��-�}��|�ű�ƽUP���v���J�D����ۼ��u�J������+���sѺ.
9fL�:�;�$;#�5;�?;��D;j[G;eH;��H;��H;��H;��H;!�H;��H;T�H;n�H;Y�H;T�H;a�H;7�H;a�H;T�H;Y�H;n�H;T�H;��H;!�H;��H;��H;��H;��H;eH;j[G;��D;�?;#�5;�$;�;fL�:.
9�sѺ�+������u�J�����ۼD���J��v��UP��ƽű�|�}��-�      nHͽ̪ɽ�;��"����������[�z0�p��'<ͼо��u�J���k��+��(����:�`�:|�;�/;�K<;!C;9lF;��G;�H;�H;�H;�H;A�H;T�H;��H;%�H;/�H;�H;�H;�H;��H;�H;�H;�H;/�H;%�H;��H;T�H;A�H;�H;�H;�H;�H;��G;9lF;!C;�K<;�/;|�;�`�:���:�(�+�k����u�J�о��'<ͼp��z0���[�������"���;��̪ɽ      �����v����w�]�c��J�Ȅ-�x��;缈沼ㄼ��;�����k��56�d��M<Q:֣�:�h;M*;��8;��@;�OE;�tG;DhH;��H;��H;�H;#�H;��H;y�H;��H;��H;��H;��H;��H;��H;��H;��H;��H;��H;��H;��H;��H;y�H;��H;#�H;�H;��H;��H;DhH;�tG;�OE;��@;��8;M*;�h;֣�:M<Q:d��56�k��������;�ㄼ�沼�;�x�Ȅ-��J�]�c���w��v��      ��'�#�$����y��  ���ۼ����+����]��X!�>ۻ�+��+�d���>:]��:@�;Z�%;	�5;��>;�'D;�F;� H;8�H;[�H;��H;��H;��H;��H;k�H;��H;��H;��H;��H;h�H;K�H;m�H;K�H;h�H;��H;��H;��H;��H;k�H;��H;��H;��H;��H;[�H;8�H;� H;�F;�'D;��>;	�5;Z�%;@�;]��:�>:d��+��+��>ۻ�X!���]��+�������ۼ�  �y����#�$�      B<ͼ��ɼ�����֯�Ҷ��ㄼ��Y�-�*�I���t���X��sѺ�(�M<Q:]��:��
;v�#;��3;�b=;#C;3CF;�G;�H;��H;�H;9�H;��H;X�H;!�H;d�H;��H;b�H;5�H;O�H;	�H;��H;�H;��H;	�H;O�H;5�H;b�H;��H;d�H;!�H;X�H;��H;9�H;�H;��H;�H;�G;3CF;#C;�b=;��3;v�#;��
;]��:M<Q:�(��sѺ�X�t��I���-�*���Y�ㄼҶ���֯�������ɼ      ��n��mj���]���J�n�1�L4�k��S���U
x�hX���y�.
9���:֣�:@�;v�#;w�2;�<;�oB;7�E;��G;�dH;��H;8�H;��H;��H;��H;��H;9�H;F�H;8�H;�H;��H;��H;��H;��H;��H;��H;��H;��H;��H;�H;8�H;F�H;9�H;��H;��H;��H;��H;8�H;��H;�dH;��G;7�E;�oB;�<;w�2;v�#;@�;֣�:���:.
9��y�hX�U
x�S���k��L4�n�1���J���]��mj�      ����o���X��P�ѻf���[ǐ��X��6��
���K�><":fL�:�`�:�h;Z�%;��3;�<;Y/B;��E;�[G;�GH;N�H;��H;a�H;�H;7�H;=�H;��H;�H;�H;��H;��H;��H;]�H;O�H;K�H;'�H;K�H;O�H;]�H;��H;��H;��H;�H;�H;��H;=�H;7�H;�H;a�H;��H;N�H;�GH;�[G;��E;Y/B;�<;��3;Z�%;�h;�`�:fL�:><":�K��
���6��X�[ǐ�f���P�ѻX��o���      �Q^��X�UF�\�)��+�,ж���<�"jS��k:���:J��:�;|�;M*;	�5;�b=;�oB;��E;�IG;]7H;s�H;��H;�H;-�H;��H;��H;��H;��H;��H;��H;��H;u�H;P�H;��H;��H;��H;��H;��H;��H;��H;P�H;u�H;��H;��H;��H;��H;��H;��H;��H;-�H;�H;��H;s�H;]7H;�IG;��E;�oB;�b=;	�5;M*;|�;�;J��:���:�k:"jS���<�,ж��+�\�)�UF��X�      0.�5��,�깜�K�
9�Z:��k:L�:5��:�x;��;�$;�/;��8;��>;#C;7�E;�[G;]7H;ͤH;�H;&�H;��H;5�H;��H;P�H;��H;��H;��H;z�H;5�H;�H;��H;��H;��H;��H;u�H;��H;��H;��H;��H;�H;5�H;z�H;��H;��H;��H;P�H;��H;5�H;��H;&�H;�H;ͤH;]7H;�[G;7�E;#C;��>;��8;�/;�$;��;�x;5��:L�:��k:�Z:
9��K�,��5��      �:nĆ:oȒ:���:r�:o��:���:��	;v;7�#;��-;#�5;�K<;��@;�'D;3CF;��G;�GH;s�H;�H;��H;P�H;��H;\�H;#�H;��H;��H;��H;[�H;�H;��H;��H;m�H;[�H;*�H;�H;�H;�H;*�H;[�H;m�H;��H;��H;�H;[�H;��H;��H;��H;#�H;\�H;��H;P�H;��H;�H;s�H;�GH;��G;3CF;�'D;��@;�K<;#�5;��-;7�#;v;��	;���:o��:r�:���:oȒ:nĆ:      �V;�w;1�;Q�
;�;�;)� ;��(;��/;$H6;��;;�?;!C;�OE;�F;�G;�dH;N�H;��H;&�H;P�H;��H;1�H;��H;f�H;�H;��H;b�H;��H;��H;��H;B�H;�H;�H;��H;��H;��H;��H;��H;�H;�H;B�H;��H;��H;��H;b�H;��H;�H;f�H;��H;1�H;��H;P�H;&�H;��H;N�H;�dH;�G;�F;�OE;!C;�?;��;;$H6;��/;��(;)� ;�;�;Q�
;1�;�w;      �R%;i�%;_�';M*;4�-;ʕ1;�5;6�9;�,=;IQ@;�B;��D;9lF;�tG;� H;�H;��H;��H;�H;��H;��H;1�H;�H;b�H;��H;r�H;5�H;��H;��H;��H;�H;��H;��H;��H;}�H;e�H;L�H;e�H;}�H;��H;��H;��H;�H;��H;��H;��H;5�H;r�H;��H;b�H;�H;1�H;��H;��H;�H;��H;��H;�H;� H;�tG;9lF;��D;�B;IQ@;�,=;6�9;�5;ʕ1;4�-;M*;_�';i�%;      ~n8;M�8;؎9;��:;��<;
c>;ZQ@;�.B;��C;�OE;�yF;j[G;��G;DhH;8�H;��H;8�H;a�H;-�H;5�H;\�H;��H;b�H;k�H;j�H;D�H;��H;��H;e�H;	�H;��H;��H;Y�H;(�H;"�H;�H;��H;�H;"�H;(�H;Y�H;��H;��H;	�H;e�H;��H;��H;D�H;j�H;k�H;b�H;��H;\�H;5�H;-�H;a�H;8�H;��H;8�H;DhH;��G;j[G;�yF;�OE;��C;�.B;ZQ@;
c>;��<;��:;؎9;M�8;      ��A;B;2oB;�C;��C;|�D;otE;�CF;N�F;��G;�H;eH;�H;��H;[�H;�H;��H;�H;��H;��H;#�H;f�H;��H;j�H;-�H;��H;��H;i�H; �H;��H;r�H;@�H;�H;��H;��H;��H;��H;��H;��H;��H;�H;@�H;r�H;��H; �H;i�H;��H;��H;-�H;j�H;��H;f�H;#�H;��H;��H;�H;��H;�H;[�H;��H;�H;eH;�H;��G;N�F;�CF;otE;|�D;��C;�C;2oB;B;      nCF;{QF;�yF;�F;�G;�[G;�G;YH;#HH;��H;��H;��H;�H;��H;��H;9�H;��H;7�H;��H;P�H;��H;�H;r�H;D�H;��H;��H;_�H;��H;��H;a�H;�H;��H;��H;��H;o�H;\�H;n�H;\�H;o�H;��H;��H;��H;�H;a�H;��H;��H;_�H;��H;��H;D�H;r�H;�H;��H;P�H;��H;7�H;��H;9�H;��H;��H;�H;��H;��H;��H;#HH;YH;�G;�[G;�G;�F;�yF;{QF;      �H;H;� H;�7H;�SH;KrH;9�H;ժH;��H;��H;|�H;��H;�H;�H;��H;��H;��H;=�H;��H;��H;��H;��H;5�H;��H;��H;_�H;��H;��H;H�H;�H;��H;��H;b�H;D�H;(�H;�H;�H;�H;(�H;D�H;b�H;��H;��H;�H;H�H;��H;��H;_�H;��H;��H;5�H;��H;��H;��H;��H;=�H;��H;��H;��H;�H;�H;��H;|�H;��H;��H;ժH;9�H;KrH;�SH;�7H;� H;H;      ��H;5�H;��H;Z�H;Q�H;��H;L�H;��H;(�H;2�H;&�H;��H;�H;#�H;��H;X�H;��H;��H;��H;��H;��H;b�H;��H;��H;i�H;��H;��H;W�H;�H;��H;u�H;F�H;!�H;��H;��H;��H;��H;��H;��H;��H;!�H;F�H;u�H;��H;�H;W�H;��H;��H;i�H;��H;��H;b�H;��H;��H;��H;��H;��H;X�H;��H;#�H;�H;��H;&�H;2�H;(�H;��H;L�H;��H;Q�H;Z�H;��H;5�H;      ��H;U�H;7�H;��H;��H;i�H;��H;��H;��H;��H;��H;��H;A�H;��H;��H;!�H;9�H;�H;��H;��H;[�H;��H;��H;e�H; �H;��H;H�H;�H;��H;k�H;7�H;��H;��H;��H;��H;��H;�H;��H;��H;��H;��H;��H;7�H;k�H;��H;�H;H�H;��H; �H;e�H;��H;��H;[�H;��H;��H;�H;9�H;!�H;��H;��H;A�H;��H;��H;��H;��H;��H;��H;i�H;��H;��H;7�H;U�H;      ��H;	�H;�H;w�H;��H;e�H;�H;��H;#�H;��H;��H;!�H;T�H;y�H;k�H;d�H;F�H;�H;��H;z�H;�H;��H;��H;	�H;��H;a�H;�H;��H;k�H;-�H;��H;��H;��H;��H;d�H;K�H;A�H;K�H;d�H;��H;��H;��H;��H;-�H;k�H;��H;�H;a�H;��H;	�H;��H;��H;�H;z�H;��H;�H;F�H;d�H;k�H;y�H;T�H;!�H;��H;��H;#�H;��H;�H;e�H;��H;w�H;�H;	�H;      L�H;p�H;��H;��H;��H;'�H;I�H;w�H;��H;��H;��H;��H;��H;��H;��H;��H;8�H;��H;��H;5�H;��H;��H;�H;��H;r�H;�H;��H;u�H;7�H;��H;��H;��H;w�H;?�H;�H;'�H;(�H;'�H;�H;?�H;w�H;��H;��H;��H;7�H;u�H;��H;�H;r�H;��H;�H;��H;��H;5�H;��H;��H;8�H;��H;��H;��H;��H;��H;��H;��H;��H;w�H;I�H;'�H;��H;��H;��H;p�H;      >�H;B�H;F�H;>�H;V�H;u�H;l�H;��H;��H;v�H;n�H;T�H;%�H;��H;��H;b�H;�H;��H;u�H;�H;��H;B�H;��H;��H;@�H;��H;��H;F�H;��H;��H;��H;_�H;A�H;�H;��H;��H;��H;��H;��H;�H;A�H;_�H;��H;��H;��H;F�H;��H;��H;@�H;��H;��H;B�H;��H;�H;u�H;��H;�H;b�H;��H;��H;%�H;T�H;n�H;v�H;��H;��H;l�H;u�H;V�H;>�H;F�H;B�H;      C�H;6�H;:�H;:�H;3�H;)�H;$�H;�H;��H;��H;��H;n�H;/�H;��H;��H;5�H;��H;��H;P�H;��H;m�H;�H;��H;Y�H;�H;��H;b�H;!�H;��H;��H;w�H;A�H;��H;��H;��H;��H;��H;��H;��H;��H;��H;A�H;w�H;��H;��H;!�H;b�H;��H;�H;Y�H;��H;�H;m�H;��H;P�H;��H;��H;5�H;��H;��H;/�H;n�H;��H;��H;��H;�H;$�H;)�H;3�H;:�H;:�H;6�H;      ��H;��H;��H;��H;��H;h�H;c�H;0�H;�H;��H;��H;Y�H;�H;��H;��H;O�H;��H;]�H;��H;��H;[�H;�H;��H;(�H;��H;��H;D�H;��H;��H;��H;?�H;�H;��H;��H;��H;��H;��H;��H;��H;��H;��H;�H;?�H;��H;��H;��H;D�H;��H;��H;(�H;��H;�H;[�H;��H;��H;]�H;��H;O�H;��H;��H;�H;Y�H;��H;��H;�H;0�H;c�H;h�H;��H;��H;��H;��H;      ��H;��H;��H;��H;��H;��H;s�H;C�H;�H;��H;��H;T�H;�H;��H;h�H;	�H;��H;O�H;��H;��H;*�H;��H;}�H;"�H;��H;o�H;(�H;��H;��H;d�H;�H;��H;��H;��H;��H;��H;��H;��H;��H;��H;��H;��H;�H;d�H;��H;��H;(�H;o�H;��H;"�H;}�H;��H;*�H;��H;��H;O�H;��H;	�H;h�H;��H;�H;T�H;��H;��H;�H;C�H;s�H;��H;��H;��H;��H;��H;      ��H;��H;��H;��H;��H;|�H;X�H;<�H;�H;��H;��H;a�H;�H;��H;K�H;��H;��H;K�H;��H;��H;�H;��H;e�H;�H;��H;\�H;�H;��H;��H;K�H;'�H;��H;��H;��H;��H;��H;��H;��H;��H;��H;��H;��H;'�H;K�H;��H;��H;�H;\�H;��H;�H;e�H;��H;�H;��H;��H;K�H;��H;��H;K�H;��H;�H;a�H;��H;��H;�H;<�H;X�H;|�H;��H;��H;��H;��H;      +�H;$�H;�H;��H;��H;��H;��H;Y�H;$�H;��H;z�H;7�H;��H;��H;m�H;�H;��H;'�H;��H;u�H;�H;��H;L�H;��H;��H;n�H;�H;��H;�H;A�H;(�H;��H;��H;��H;��H;��H;~�H;��H;��H;��H;��H;��H;(�H;A�H;�H;��H;�H;n�H;��H;��H;L�H;��H;�H;u�H;��H;'�H;��H;�H;m�H;��H;��H;7�H;z�H;��H;$�H;Y�H;��H;��H;��H;��H;�H;$�H;      ��H;��H;��H;��H;��H;|�H;X�H;<�H;�H;��H;��H;a�H;�H;��H;K�H;��H;��H;K�H;��H;��H;�H;��H;e�H;�H;��H;\�H;�H;��H;��H;K�H;'�H;��H;��H;��H;��H;��H;��H;��H;��H;��H;��H;��H;'�H;K�H;��H;��H;�H;\�H;��H;�H;e�H;��H;�H;��H;��H;K�H;��H;��H;K�H;��H;�H;a�H;��H;��H;�H;<�H;X�H;|�H;��H;��H;��H;��H;      ��H;��H;��H;��H;��H;��H;s�H;C�H;�H;��H;��H;T�H;�H;��H;h�H;	�H;��H;O�H;��H;��H;*�H;��H;}�H;"�H;��H;o�H;(�H;��H;��H;d�H;�H;��H;��H;��H;��H;��H;��H;��H;��H;��H;��H;��H;�H;d�H;��H;��H;(�H;o�H;��H;"�H;}�H;��H;*�H;��H;��H;O�H;��H;	�H;h�H;��H;�H;T�H;��H;��H;�H;C�H;s�H;��H;��H;��H;��H;��H;      ��H;��H;��H;��H;��H;h�H;c�H;0�H;�H;��H;��H;Y�H;�H;��H;��H;O�H;��H;]�H;��H;��H;[�H;�H;��H;(�H;��H;��H;D�H;��H;��H;��H;?�H;�H;��H;��H;��H;��H;��H;��H;��H;��H;��H;�H;?�H;��H;��H;��H;D�H;��H;��H;(�H;��H;�H;[�H;��H;��H;]�H;��H;O�H;��H;��H;�H;Y�H;��H;��H;�H;0�H;c�H;h�H;��H;��H;��H;��H;      C�H;6�H;:�H;:�H;3�H;)�H;$�H;�H;��H;��H;��H;n�H;/�H;��H;��H;5�H;��H;��H;P�H;��H;m�H;�H;��H;Y�H;�H;��H;b�H;!�H;��H;��H;w�H;A�H;��H;��H;��H;��H;��H;��H;��H;��H;��H;A�H;w�H;��H;��H;!�H;b�H;��H;�H;Y�H;��H;�H;m�H;��H;P�H;��H;��H;5�H;��H;��H;/�H;n�H;��H;��H;��H;�H;$�H;)�H;3�H;:�H;:�H;6�H;      >�H;B�H;F�H;>�H;V�H;u�H;l�H;��H;��H;v�H;n�H;T�H;%�H;��H;��H;b�H;�H;��H;u�H;�H;��H;B�H;��H;��H;@�H;��H;��H;F�H;��H;��H;��H;_�H;A�H;�H;��H;��H;��H;��H;��H;�H;A�H;_�H;��H;��H;��H;F�H;��H;��H;@�H;��H;��H;B�H;��H;�H;u�H;��H;�H;b�H;��H;��H;%�H;T�H;n�H;v�H;��H;��H;l�H;u�H;V�H;>�H;F�H;B�H;      L�H;p�H;��H;��H;��H;'�H;I�H;w�H;��H;��H;��H;��H;��H;��H;��H;��H;8�H;��H;��H;5�H;��H;��H;�H;��H;r�H;�H;��H;u�H;7�H;��H;��H;��H;w�H;?�H;�H;'�H;(�H;'�H;�H;?�H;w�H;��H;��H;��H;7�H;u�H;��H;�H;r�H;��H;�H;��H;��H;5�H;��H;��H;8�H;��H;��H;��H;��H;��H;��H;��H;��H;w�H;I�H;'�H;��H;��H;��H;p�H;      ��H;	�H;�H;w�H;��H;e�H;�H;��H;#�H;��H;��H;!�H;T�H;y�H;k�H;d�H;F�H;�H;��H;z�H;�H;��H;��H;	�H;��H;a�H;�H;��H;k�H;-�H;��H;��H;��H;��H;d�H;K�H;A�H;K�H;d�H;��H;��H;��H;��H;-�H;k�H;��H;�H;a�H;��H;	�H;��H;��H;�H;z�H;��H;�H;F�H;d�H;k�H;y�H;T�H;!�H;��H;��H;#�H;��H;�H;e�H;��H;w�H;�H;	�H;      ��H;U�H;7�H;��H;��H;i�H;��H;��H;��H;��H;��H;��H;A�H;��H;��H;!�H;9�H;�H;��H;��H;[�H;��H;��H;e�H; �H;��H;H�H;�H;��H;k�H;7�H;��H;��H;��H;��H;��H;�H;��H;��H;��H;��H;��H;7�H;k�H;��H;�H;H�H;��H; �H;e�H;��H;��H;[�H;��H;��H;�H;9�H;!�H;��H;��H;A�H;��H;��H;��H;��H;��H;��H;i�H;��H;��H;7�H;U�H;      ��H;5�H;��H;Z�H;Q�H;��H;L�H;��H;(�H;2�H;&�H;��H;�H;#�H;��H;X�H;��H;��H;��H;��H;��H;b�H;��H;��H;i�H;��H;��H;W�H;�H;��H;u�H;F�H;!�H;��H;��H;��H;��H;��H;��H;��H;!�H;F�H;u�H;��H;�H;W�H;��H;��H;i�H;��H;��H;b�H;��H;��H;��H;��H;��H;X�H;��H;#�H;�H;��H;&�H;2�H;(�H;��H;L�H;��H;Q�H;Z�H;��H;5�H;      �H;H;� H;�7H;�SH;KrH;9�H;ժH;��H;��H;|�H;��H;�H;�H;��H;��H;��H;=�H;��H;��H;��H;��H;5�H;��H;��H;_�H;��H;��H;H�H;�H;��H;��H;b�H;D�H;(�H;�H;�H;�H;(�H;D�H;b�H;��H;��H;�H;H�H;��H;��H;_�H;��H;��H;5�H;��H;��H;��H;��H;=�H;��H;��H;��H;�H;�H;��H;|�H;��H;��H;ժH;9�H;KrH;�SH;�7H;� H;H;      nCF;{QF;�yF;�F;�G;�[G;�G;YH;#HH;��H;��H;��H;�H;��H;��H;9�H;��H;7�H;��H;P�H;��H;�H;r�H;D�H;��H;��H;_�H;��H;��H;a�H;�H;��H;��H;��H;o�H;\�H;n�H;\�H;o�H;��H;��H;��H;�H;a�H;��H;��H;_�H;��H;��H;D�H;r�H;�H;��H;P�H;��H;7�H;��H;9�H;��H;��H;�H;��H;��H;��H;#HH;YH;�G;�[G;�G;�F;�yF;{QF;      ��A;B;2oB;�C;��C;|�D;otE;�CF;N�F;��G;�H;eH;�H;��H;[�H;�H;��H;�H;��H;��H;#�H;f�H;��H;j�H;-�H;��H;��H;i�H; �H;��H;r�H;@�H;�H;��H;��H;��H;��H;��H;��H;��H;�H;@�H;r�H;��H; �H;i�H;��H;��H;-�H;j�H;��H;f�H;#�H;��H;��H;�H;��H;�H;[�H;��H;�H;eH;�H;��G;N�F;�CF;otE;|�D;��C;�C;2oB;B;      ~n8;M�8;؎9;��:;��<;
c>;ZQ@;�.B;��C;�OE;�yF;j[G;��G;DhH;8�H;��H;8�H;a�H;-�H;5�H;\�H;��H;b�H;k�H;j�H;D�H;��H;��H;e�H;	�H;��H;��H;Y�H;(�H;"�H;�H;��H;�H;"�H;(�H;Y�H;��H;��H;	�H;e�H;��H;��H;D�H;j�H;k�H;b�H;��H;\�H;5�H;-�H;a�H;8�H;��H;8�H;DhH;��G;j[G;�yF;�OE;��C;�.B;ZQ@;
c>;��<;��:;؎9;M�8;      �R%;i�%;_�';M*;4�-;ʕ1;�5;6�9;�,=;IQ@;�B;��D;9lF;�tG;� H;�H;��H;��H;�H;��H;��H;1�H;�H;b�H;��H;r�H;5�H;��H;��H;��H;�H;��H;��H;��H;}�H;e�H;L�H;e�H;}�H;��H;��H;��H;�H;��H;��H;��H;5�H;r�H;��H;b�H;�H;1�H;��H;��H;�H;��H;��H;�H;� H;�tG;9lF;��D;�B;IQ@;�,=;6�9;�5;ʕ1;4�-;M*;_�';i�%;      �V;�w;1�;Q�
;�;�;)� ;��(;��/;$H6;��;;�?;!C;�OE;�F;�G;�dH;N�H;��H;&�H;P�H;��H;1�H;��H;f�H;�H;��H;b�H;��H;��H;��H;B�H;�H;�H;��H;��H;��H;��H;��H;�H;�H;B�H;��H;��H;��H;b�H;��H;�H;f�H;��H;1�H;��H;P�H;&�H;��H;N�H;�dH;�G;�F;�OE;!C;�?;��;;$H6;��/;��(;)� ;�;�;Q�
;1�;�w;      �:nĆ:oȒ:���:r�:o��:���:��	;v;7�#;��-;#�5;�K<;��@;�'D;3CF;��G;�GH;s�H;�H;��H;P�H;��H;\�H;#�H;��H;��H;��H;[�H;�H;��H;��H;m�H;[�H;*�H;�H;�H;�H;*�H;[�H;m�H;��H;��H;�H;[�H;��H;��H;��H;#�H;\�H;��H;P�H;��H;�H;s�H;�GH;��G;3CF;�'D;��@;�K<;#�5;��-;7�#;v;��	;���:o��:r�:���:oȒ:nĆ:      0.�5��,�깜�K�
9�Z:��k:L�:5��:�x;��;�$;�/;��8;��>;#C;7�E;�[G;]7H;ͤH;�H;&�H;��H;5�H;��H;P�H;��H;��H;��H;z�H;5�H;�H;��H;��H;��H;��H;u�H;��H;��H;��H;��H;�H;5�H;z�H;��H;��H;��H;P�H;��H;5�H;��H;&�H;�H;ͤH;]7H;�[G;7�E;#C;��>;��8;�/;�$;��;�x;5��:L�:��k:�Z:
9��K�,��5��      �Q^��X�UF�\�)��+�,ж���<�"jS��k:���:J��:�;|�;M*;	�5;�b=;�oB;��E;�IG;]7H;s�H;��H;�H;-�H;��H;��H;��H;��H;��H;��H;��H;u�H;P�H;��H;��H;��H;��H;��H;��H;��H;P�H;u�H;��H;��H;��H;��H;��H;��H;��H;-�H;�H;��H;s�H;]7H;�IG;��E;�oB;�b=;	�5;M*;|�;�;J��:���:�k:"jS���<�,ж��+�\�)�UF��X�      ����o���X��P�ѻf���[ǐ��X��6��
���K�><":fL�:�`�:�h;Z�%;��3;�<;Y/B;��E;�[G;�GH;N�H;��H;a�H;�H;7�H;=�H;��H;�H;�H;��H;��H;��H;]�H;O�H;K�H;'�H;K�H;O�H;]�H;��H;��H;��H;�H;�H;��H;=�H;7�H;�H;a�H;��H;N�H;�GH;�[G;��E;Y/B;�<;��3;Z�%;�h;�`�:fL�:><":�K��
���6��X�[ǐ�f���P�ѻX��o���      ��n��mj���]���J�n�1�L4�k��S���U
x�hX���y�.
9���:֣�:@�;v�#;w�2;�<;�oB;7�E;��G;�dH;��H;8�H;��H;��H;��H;��H;9�H;F�H;8�H;�H;��H;��H;��H;��H;��H;��H;��H;��H;��H;�H;8�H;F�H;9�H;��H;��H;��H;��H;8�H;��H;�dH;��G;7�E;�oB;�<;w�2;v�#;@�;֣�:���:.
9��y�hX�U
x�S���k��L4�n�1���J���]��mj�      B<ͼ��ɼ�����֯�Ҷ��ㄼ��Y�-�*�I���t���X��sѺ�(�M<Q:]��:��
;v�#;��3;�b=;#C;3CF;�G;�H;��H;�H;9�H;��H;X�H;!�H;d�H;��H;b�H;5�H;O�H;	�H;��H;�H;��H;	�H;O�H;5�H;b�H;��H;d�H;!�H;X�H;��H;9�H;�H;��H;�H;�G;3CF;#C;�b=;��3;v�#;��
;]��:M<Q:�(��sѺ�X�t��I���-�*���Y�ㄼҶ���֯�������ɼ      ��'�#�$����y��  ���ۼ����+����]��X!�>ۻ�+��+�d���>:]��:@�;Z�%;	�5;��>;�'D;�F;� H;8�H;[�H;��H;��H;��H;��H;k�H;��H;��H;��H;��H;h�H;K�H;m�H;K�H;h�H;��H;��H;��H;��H;k�H;��H;��H;��H;��H;[�H;8�H;� H;�F;�'D;��>;	�5;Z�%;@�;]��:�>:d��+��+��>ۻ�X!���]��+�������ۼ�  �y����#�$�      �����v����w�]�c��J�Ȅ-�x��;缈沼ㄼ��;�����k��56�d��M<Q:֣�:�h;M*;��8;��@;�OE;�tG;DhH;��H;��H;�H;#�H;��H;y�H;��H;��H;��H;��H;��H;��H;��H;��H;��H;��H;��H;��H;��H;y�H;��H;#�H;�H;��H;��H;DhH;�tG;�OE;��@;��8;M*;�h;֣�:M<Q:d��56�k��������;�ㄼ�沼�;�x�Ȅ-��J�]�c���w��v��      nHͽ̪ɽ�;��"����������[�z0�p��'<ͼо��u�J���k��+��(����:�`�:|�;�/;�K<;!C;9lF;��G;�H;�H;�H;�H;A�H;T�H;��H;%�H;/�H;�H;�H;�H;��H;�H;�H;�H;/�H;%�H;��H;T�H;A�H;�H;�H;�H;�H;��G;9lF;!C;�K<;�/;|�;�`�:���:�(�+�k����u�J�о��'<ͼp��z0���[�������"���;��̪ɽ      ��-�}��|�ű�ƽUP���v���J�D����ۼ��u�J������+���sѺ.
9fL�:�;�$;#�5;�?;��D;j[G;eH;��H;��H;��H;��H;!�H;��H;T�H;n�H;Y�H;T�H;a�H;7�H;a�H;T�H;Y�H;n�H;T�H;��H;!�H;��H;��H;��H;��H;eH;j[G;��D;�?;#�5;�$;�;fL�:.
9�sѺ�+������u�J�����ۼD���J��v��UP��ƽű�|�}��-�       j�Ide�M0X�sD�\{+�z�����k㻽R���IDX������ۼо����;�>ۻ�X���y�><":J��:��;��-;��;;�B;�yF;�H;��H;|�H;&�H;��H;��H;��H;n�H;��H;��H;��H;��H;z�H;��H;��H;��H;��H;n�H;��H;��H;��H;&�H;|�H;��H;�H;�yF;�B;��;;��-;��;J��:><":��y��X�>ۻ��;�о����ۼ���IDX�R���k㻽���z��\{+�sD�M0X�Ide�      ��Fh��b���I���|x���O��C(�y�Īɽ����IDX�D��'<ͼㄼ�X!�t��hX��K����:�x;7�#;$H6;IQ@;�OE;��G;��H;��H;2�H;��H;��H;��H;v�H;��H;��H;��H;��H;��H;��H;��H;��H;��H;v�H;��H;��H;��H;2�H;��H;��H;��G;�OE;IQ@;$H6;7�#;�x;���:�K�hX�t���X!�ㄼ'<ͼD��IDX�����Īɽy��C(���O��|x��I��b��Fh��      /�����������;^ɰ��G����i�.�5��	�ĪɽR����J�p���沼��]�I���U
x��
���k:5��:v;��/;�,=;��C;N�F;#HH;��H;(�H;��H;#�H;��H;��H;��H;�H;�H;�H;$�H;�H;�H;�H;��H;��H;��H;#�H;��H;(�H;��H;#HH;N�F;��C;�,=;��/;v;5��:�k:�
��U
x�I�����]��沼p���J�R���Īɽ�	�.�5���i��G��^ɰ��;��徨���      �2�L�-��"�$E�����4Kɾa��w�s�.�5�y�k㻽�v��z0��;��+��-�*�S����6�"jS�L�:��	;��(;6�9;�.B;�CF;YH;ժH;��H;��H;��H;w�H;��H;�H;0�H;C�H;<�H;Y�H;<�H;C�H;0�H;�H;��H;w�H;��H;��H;��H;ժH;YH;�CF;�.B;6�9;��(;��	;L�:"jS��6�S���-�*��+���;�z0��v��k㻽y�.�5�w�s�a��4Kɾ����$E��"�L�-�      3s�cm�/�\�]�C�,�%����TҾa����i��C(����UP����[�x������Y�k���X���<���k:���:)� ;�5;ZQ@;otE;�G;9�H;L�H;��H;�H;I�H;l�H;$�H;c�H;s�H;X�H;��H;X�H;s�H;c�H;$�H;l�H;I�H;�H;��H;L�H;9�H;�G;otE;ZQ@;�5;)� ;���:��k:��<��X�k����Y����x���[�UP����콡C(���i�a���TҾ��,�%�]�C�/�\�cm�      �ޞ�������RF�3�W�M�-���4Kɾ�G����O�z��ƽ����Ȅ-���ۼㄼL4�[ǐ�,ж��Z:o��:�;ʕ1;
c>;|�D;�[G;KrH;��H;i�H;e�H;'�H;u�H;)�H;h�H;��H;|�H;��H;|�H;��H;h�H;)�H;u�H;'�H;e�H;i�H;��H;KrH;�[G;|�D;
c>;ʕ1;�;o��:�Z:,ж�[ǐ�L4�ㄼ��ۼȄ-�����ƽz����O��G��4Kɾ��M�-�3�W�RF�������      ��ſ~��Bw���ޞ�|���3�W�,�%�����^ɰ��|x�\{+�ű����J��  �Ҷ��n�1�f����+�
9r�:�;4�-;��<;��C;�G;�SH;Q�H;��H;��H;��H;V�H;3�H;��H;��H;��H;��H;��H;��H;��H;3�H;V�H;��H;��H;��H;Q�H;�SH;�G;��C;��<;4�-;�;r�:
9�+�f���n�1�Ҷ���  ��J���ű�\{+��|x�^ɰ�����,�%�3�W�|����ޞ�Bw��~��      ������Կp���ޞ�RF�]�C�$E��;�I��sD�|�"��]�c�y��֯���J�P�ѻ\�)���K����:Q�
;M*;��:;�C;�F;�7H;Z�H;��H;w�H;��H;>�H;:�H;��H;��H;��H;��H;��H;��H;��H;:�H;>�H;��H;w�H;��H;Z�H;�7H;�F;�C;��:;M*;Q�
;���:��K�\�)�P�ѻ��J��֯�y�]�c�"��|�sD��I���;$E�]�C�RF��ޞ�p���Կ��      ������{���ԿBw�����/�\��"����b��M0X�}���;����w����������]�X��UF�,��oȒ:1�;_�';؎9;2oB;�yF;� H;��H;7�H;�H;��H;F�H;:�H;��H;��H;��H;�H;��H;��H;��H;:�H;F�H;��H;�H;7�H;��H;� H;�yF;2oB;؎9;_�';1�;oȒ:,��UF�X�黼�]����������w��;��}��M0X�b������"�/�\����Bw���Կ{�𿖏�      $��������~�����cm�L�-�����Fh��Ide�-�̪ɽ�v��#�$���ɼ�mj�o����X�5��nĆ:�w;i�%;M�8;B;{QF;H;5�H;U�H;	�H;p�H;B�H;6�H;��H;��H;��H;$�H;��H;��H;��H;6�H;B�H;p�H;	�H;U�H;5�H;H;{QF;B;M�8;i�%;�w;nĆ:5���X�o����mj���ɼ#�$��v��̪ɽ-�Ide�Fh������L�-�cm����~���忖����      Vܿ%�ֿ�aǿ2^��&���Io���7����iþ�(���-=��` ��@����_�&]�&p����I�q�ѻ��)��R�\�:��
;*;D�:;�B;UHF;=�G;�kH;3�H;��H;i�H;��H;��H;p�H;��H;(�H;��H;(�H;��H;p�H;��H;��H;i�H;��H;3�H;�kH;=�G;UHF;�B;D�:;*;��
;\�:�R���)�q�ѻ��I�&p��&]���_��@���` ��-=��(���iþ����7�Io�&���2^���aǿ%�ֿ      %�ֿ5pѿ֊¿������PXi�Õ3��
�GD��;l��1�9�j.���R��\� �\x��1�E��ͻ��$�� ����:��;��*;\�:;.�B;3TF;��G;[mH;ϠH;ݶH;��H;��H;��H;�H;��H;<�H;��H;<�H;��H;�H;��H;��H;��H;ݶH;ϠH;[mH;��G;3TF;.�B;\�:;��*;��;���:� ���$��ͻ1�E�\x�� �\��R��j.��1�9�;l��GD���
�Õ3�PXi�������֊¿5pѿ      �aǿ֊¿���������s"Y��f'�����)o���.}��k/�m��ڟ�<Q�%#�ע��(;�P��������7���:J�;�,;��;;�C;RvF;/�G;�qH;[�H;��H;=�H;�H;�H;��H;��H;j�H;��H;j�H;��H;��H;�H;�H;=�H;��H;[�H;�qH;/�G;RvF;�C;��;;�,;J�;��:��7����P����(;�ע�%#�<Q�ڟ�m���k/��.}�)o�������f'�s"Y����������֊¿      2^������b���Io���@���޾����&ce�"����ڽ绒��f@������R���O*�mG�����<^9Ҳ�:[;�c.;'�<;ՏC;G�F;��G;�xH;ĤH;8�H;I�H;��H;��H;��H;�H;��H;7�H;��H;�H;��H;��H;��H;I�H;8�H;ĤH;�xH;��G;G�F;ՏC;'�<;�c.;[;Ҳ�:<^9���mG���O*��R�������f@�绒���ڽ"��&ce������޾���@�Io�b�������      &����������Io��!J�@�#��\��HD������jPH�����b��C��t +�u�ټ%��������������:���:��;�X1;3>;�/D;��F;�H;r�H;��H;*�H;��H;��H;)�H;��H;p�H;��H;�H;��H;p�H;��H;)�H;��H;��H;*�H;��H;r�H;�H;��F;�/D;3>;�X1;��;���:��:����������%��u�ټt +�C���b�����jPH�����HD���\��@�#��!J�Io��������      Io�PXi�s"Y���@�@�#��
��о�A�� �i���(�i��gr����_��5��ɺ�n�`��<����d�=�\�P�X:PO�:7`;#�4;�?;��D;�7G;�/H;ȊH;��H;��H;.�H;��H;��H;�H;��H;-�H;��H;-�H;��H;�H;��H;��H;.�H;��H;��H;ȊH;�/H;�7G;��D;�?;#�4;7`;PO�:P�X:=�\���d��<��n�`��ɺ��5���_�gr��i����(� �i��A���о�
�@�#���@�s"Y�PXi�      ��7�Õ3��f'���\���о�����.}��-=�o
�y�ĽO��:����������7�?GĻ*�$�
S�����:�z;�C&;E+8;FIA;1�E;��G;�KH;�H;��H;S�H;�H;(�H;��H;��H;A�H;��H;5�H;��H;A�H;��H;��H;(�H;�H;S�H;��H;�H;�KH;��G;1�E;FIA;E+8;�C&;�z;���:
S��*�$�?GĻ�7���������:�O��y�Ľo
��-=��.}������о�\����f'�Õ3�      ���
������޾HD���A���.}��D�[t���ڽ�!��\����P�ļ�
v�F�����Jɺ�N�9���:i';�-;ӊ;;��B;�HF;��G;?eH;ʜH;�H;N�H;��H;��H;��H;{�H;��H;�H;��H;�H;��H;{�H;��H;��H;��H;N�H;�H;ʜH;?eH;��G;�HF;��B;ӊ;;�-;i';���:�N�9�Jɺ��F���
v�P�ļ���\��!����ڽ[t��D��.}��A��HD���޾�����
�      �iþGD��)o���������� �i��-=�[t����R��Tys�m +����s񗼗(;�G�ѻt@�͇!��1j:�O�:4�;�C3;~�>;DED;��F;�H;_{H;��H;��H;W�H;�H;�H;��H;9�H;R�H;��H;�H;��H;R�H;9�H;��H;�H;�H;W�H;��H;��H;_{H;�H;��F;DED;~�>;�C3;4�;�O�:�1j:͇!�t@�G�ѻ�(;�s����m +�Tys��R����[t��-=� �i���������)o��GD��      �(��;l���.}�&ce�jPH���(�o
���ڽ�R����{�4�6�� �$p��\�`�ר�-��JҺ�C^9a��:=�;�}(;t�8;IA;6{E;GiG;�<H;i�H; �H;H�H;��H;N�H;��H;��H;��H;��H;�H;i�H;�H;��H;��H;��H;��H;N�H;��H;H�H; �H;i�H;�<H;GiG;6{E;IA;t�8;�}(;=�;a��:�C^9JҺ-��ר�\�`�$p��� �4�6���{��R����ڽo
���(�jPH�&ce��.}�;l��      �-=�1�9��k/�"�����i��y�Ľ�!��Tys�4�6�#��ɺ��vz����c^��˃$�{����r:���:7�;�X1;?H=;jwC;WvF;R�G;/eH;m�H;��H;��H;��H;v�H;�H;��H;��H;��H;��H;��H;��H;��H;��H;��H;�H;v�H;��H;��H;��H;m�H;/eH;R�G;WvF;jwC;?H=;�X1;7�;���:��r:{��˃$�c^������vz��ɺ�#�4�6�Tys��!��y�Ľi���"���k/�1�9�      �` �j.��m��ڽ�b��gr��O��\�m +�� ��ɺ�<��O*�bͻP6R��ǅ���:���:ڃ;�);6t8;��@;�)E;�7G;t#H;p�H;d�H;�H;J�H;��H;��H;��H;�H;n�H;�H; �H;?�H; �H;�H;n�H;�H;��H;��H;��H;J�H;�H;d�H;p�H;t#H;�7G;�)E;��@;6t8;�);ڃ;���:��:�ǅ�P6R�bͻ�O*�<��ɺ�� �m +�\�O��gr���b����ڽm��j.��      �@���R��ڟ�绒�C����_�:�������$p���vz��O*�5ֻfk������09�:`0;�� ;�C3;��=;�C;kF;��G;�[H;ÖH;o�H;&�H;b�H;��H;��H;��H;�H;'�H;��H;o�H;��H;o�H;��H;'�H;�H;��H;��H;��H;b�H;&�H;o�H;ÖH;�[H;��G;kF;�C;��=;�C3;�� ;`0;�:��09���fk�5ֻ�O*��vz�$p����輙��:���_�C��绒�ڟ��R��      ��_�\�<Q��f@�t +��5�����P�ļs�\�`����bͻfk��Iɺ�	7��:�O�:y�;%d.;��:;Z�A;c{E;�MG;q&H;/�H;�H;��H;��H;J�H;n�H;|�H;S�H;�H;��H;*�H;��H;�H;��H;*�H;��H;�H;S�H;|�H;n�H;J�H;��H;��H;�H;/�H;q&H;�MG;c{E;Z�A;��:;%d.;y�;�O�:�:�	7��Iɺfk�bͻ���\�`�s�P�ļ�����5�t +��f@�<Q�\�      &]� �%#�����u�ټ�ɺ������
v��(;�ר�c^��P6R�����	7����:���:O�;l�*;+8;� @;��D;��F;'�G; eH;��H;��H;žH;��H;�H;��H;B�H;��H;��H;��H;��H;B�H;u�H;B�H;��H;��H;��H;��H;B�H;��H;�H;��H;žH;��H;��H; eH;'�G;��F;��D;� @;+8;l�*;O�;���:���:�	7����P6R�c^��ר��(;��
v������ɺ�u�ټ����%#� �      &p��\x��ע��R��%��n�`��7�F��G�ѻ-��˃$��ǅ���09�:���:�; ~(;�Y6;��>;�C;&HF;�G;DH;s�H;�H;ϸH;3�H;K�H;2�H;�H;��H;��H;��H;,�H;�H;��H;��H;��H;�H;,�H;��H;��H;��H;�H;2�H;K�H;3�H;ϸH;�H;s�H;DH;�G;&HF;�C;��>;�Y6; ~(;�;���:�:��09�ǅ�˃$�-��G�ѻF���7�n�`�%���R��ע�\x��      ��I�1�E��(;��O*�����<��?GĻ��t@�JҺ{��:�:�O�:O�; ~(;S�5;>;qC;k�E;�bG;k#H;"{H;_�H;I�H;��H;��H;Y�H;��H;;�H;x�H;��H;h�H;��H;Y�H;��H;�H;��H;Y�H;��H;h�H;��H;x�H;;�H;��H;Y�H;��H;��H;I�H;_�H;"{H;k#H;�bG;k�E;qC;>;S�5; ~(;O�;�O�:�:��:{��JҺt@���?GĻ�<������O*��(;�1�E�      q�ѻ�ͻP���mG�������d�*�$��Jɺ͇!��C^9��r:���:`0;y�;l�*;�Y6;>;n�B;��E;8G;�H;,mH;A�H;m�H;μH;��H;��H;��H;h�H;�H;��H;��H;�H;�H;��H;�H;<�H;�H;��H;�H;�H;��H;��H;�H;h�H;��H;��H;��H;μH;m�H;A�H;,mH;�H;8G;��E;n�B;>;�Y6;l�*;y�;`0;���:��r:�C^9͇!��Jɺ*�$���d����mG��P����ͻ      ��)���$�����������=�\�
S���N�9�1j:a��:���:ڃ;�� ;%d.;+8;��>;qC;��E;�(G;��G;>cH;��H;��H;��H;��H;T�H;��H;��H;��H;��H;��H;b�H;��H;w�H;�H;I�H;c�H;I�H;�H;w�H;��H;b�H;��H;��H;��H;��H;��H;T�H;��H;��H;��H;��H;>cH;��G;�(G;��E;qC;��>;+8;%d.;�� ;ڃ;���:a��:�1j:�N�9
S��=�\�������������$�      �R�� ���7�<^9��:P�X:���:���:�O�:=�;7�;�);�C3;��:;� @;�C;k�E;8G;��G;�_H;��H;?�H;@�H;��H;d�H;Q�H;i�H;w�H;��H;��H;��H;$�H; �H;��H;@�H;{�H;{�H;{�H;@�H;��H; �H;$�H;��H;��H;��H;w�H;i�H;Q�H;d�H;��H;@�H;?�H;��H;�_H;��G;8G;k�E;�C;� @;��:;�C3;�);7�;=�;�O�:���:���:P�X:��:<^9��7�� �      \�:���:��:Ҳ�:���:PO�:�z;i';4�;�}(;�X1;6t8;��=;Z�A;��D;&HF;�bG;�H;>cH;��H;m�H;��H;S�H;�H;��H;Y�H;d�H;��H;<�H;��H;��H;��H;m�H;��H;Y�H;��H;��H;��H;Y�H;��H;m�H;��H;��H;��H;<�H;��H;d�H;Y�H;��H;�H;S�H;��H;m�H;��H;>cH;�H;�bG;&HF;��D;Z�A;��=;6t8;�X1;�}(;4�;i';�z;PO�:���:Ҳ�:��:���:      ��
;��;J�;[;��;7`;�C&;�-;�C3;t�8;?H=;��@;�C;c{E;��F;�G;k#H;,mH;��H;?�H;��H;��H;Y�H;:�H;��H;��H;��H;��H;�H;�H;4�H;�H;��H;1�H;r�H;��H;��H;��H;r�H;1�H;��H;�H;4�H;�H;�H;��H;��H;��H;��H;:�H;Y�H;��H;��H;?�H;��H;,mH;k#H;�G;��F;c{E;�C;��@;?H=;t�8;�C3;�-;�C&;7`;��;[;J�;��;      *;��*;�,;�c.;�X1;#�4;E+8;ӊ;;~�>;IA;jwC;�)E;kF;�MG;'�G;DH;"{H;A�H;��H;@�H;S�H;Y�H;��H;�H;�H;w�H;#�H;�H;��H;��H;��H;��H;��H;L�H;��H;��H;��H;��H;��H;L�H;��H;��H;��H;��H;��H;�H;#�H;w�H;�H;�H;��H;Y�H;S�H;@�H;��H;A�H;"{H;DH;'�G;�MG;kF;�)E;jwC;IA;~�>;ӊ;;E+8;#�4;�X1;�c.;�,;��*;      D�:;\�:;��;;'�<;3>;�?;FIA;��B;DED;6{E;WvF;�7G;��G;q&H; eH;s�H;_�H;m�H;��H;��H;�H;:�H;�H;��H;5�H;��H;��H;G�H;��H;~�H;(�H;��H;,�H;l�H;��H;��H;��H;��H;��H;l�H;,�H;��H;(�H;~�H;��H;G�H;��H;��H;5�H;��H;�H;:�H;�H;��H;��H;m�H;_�H;s�H; eH;q&H;��G;�7G;WvF;6{E;DED;��B;FIA;�?;3>;'�<;��;;\�:;      �B;.�B;�C;ՏC;�/D;��D;1�E;�HF;��F;GiG;R�G;t#H;�[H;/�H;��H;�H;I�H;μH;��H;d�H;��H;��H;�H;5�H;��H;��H;�H;T�H;8�H;�H;��H;��H;=�H;��H;��H;��H;��H;��H;��H;��H;=�H;��H;��H;�H;8�H;T�H;�H;��H;��H;5�H;�H;��H;��H;d�H;��H;μH;I�H;�H;��H;/�H;�[H;t#H;R�G;GiG;��F;�HF;1�E;��D;�/D;ՏC;�C;.�B;      UHF;3TF;RvF;G�F;��F;�7G;��G;��G;�H;�<H;/eH;p�H;ÖH;�H;��H;ϸH;��H;��H;T�H;Q�H;Y�H;��H;w�H;��H;��H;	�H;9�H;�H;��H;R�H;��H;.�H;C�H;}�H;��H;��H;��H;��H;��H;}�H;C�H;.�H;��H;R�H;��H;�H;9�H;	�H;��H;��H;w�H;��H;Y�H;Q�H;T�H;��H;��H;ϸH;��H;�H;ÖH;p�H;/eH;�<H;�H;��G;��G;�7G;��F;G�F;RvF;3TF;      =�G;��G;/�G;��G;�H;�/H;�KH;?eH;_{H;i�H;m�H;d�H;o�H;��H;žH;3�H;��H;��H;��H;i�H;d�H;��H;#�H;��H;�H;9�H;�H;��H;[�H;��H;��H;<�H;\�H;�H;��H;��H;��H;��H;��H;�H;\�H;<�H;��H;��H;[�H;��H;�H;9�H;�H;��H;#�H;��H;d�H;i�H;��H;��H;��H;3�H;žH;��H;o�H;d�H;m�H;i�H;_{H;?eH;�KH;�/H;�H;��G;/�G;��G;      �kH;[mH;�qH;�xH;r�H;ȊH;�H;ʜH;��H; �H;��H;�H;&�H;��H;��H;K�H;Y�H;��H;��H;w�H;��H;��H;�H;G�H;T�H;�H;��H;B�H;��H;��H;�H;B�H;k�H;l�H;��H;��H;��H;��H;��H;l�H;k�H;B�H;�H;��H;��H;B�H;��H;�H;T�H;G�H;�H;��H;��H;w�H;��H;��H;Y�H;K�H;��H;��H;&�H;�H;��H; �H;��H;ʜH;�H;ȊH;r�H;�xH;�qH;[mH;      3�H;ϠH;[�H;ĤH;��H;��H;��H;�H;��H;H�H;��H;J�H;b�H;J�H;�H;2�H;��H;h�H;��H;��H;<�H;�H;��H;��H;8�H;��H;[�H;��H;��H;�H;6�H;S�H;j�H;l�H;j�H;u�H;u�H;u�H;j�H;l�H;j�H;S�H;6�H;�H;��H;��H;[�H;��H;8�H;��H;��H;�H;<�H;��H;��H;h�H;��H;2�H;�H;J�H;b�H;J�H;��H;H�H;��H;�H;��H;��H;��H;ĤH;[�H;ϠH;      ��H;ݶH;��H;8�H;*�H;��H;S�H;N�H;W�H;��H;��H;��H;��H;n�H;��H;�H;;�H;�H;��H;��H;��H;�H;��H;~�H;�H;R�H;��H;��H;�H;+�H;J�H;I�H;Y�H;h�H;P�H;b�H;{�H;b�H;P�H;h�H;Y�H;I�H;J�H;+�H;�H;��H;��H;R�H;�H;~�H;��H;�H;��H;��H;��H;�H;;�H;�H;��H;n�H;��H;��H;��H;��H;W�H;N�H;S�H;��H;*�H;8�H;��H;ݶH;      i�H;��H;=�H;I�H;��H;.�H;�H;��H;�H;N�H;v�H;��H;��H;|�H;B�H;��H;x�H;��H;��H;��H;��H;4�H;��H;(�H;��H;��H;��H;�H;6�H;J�H;a�H;T�H;E�H;E�H;c�H;U�H;6�H;U�H;c�H;E�H;E�H;T�H;a�H;J�H;6�H;�H;��H;��H;��H;(�H;��H;4�H;��H;��H;��H;��H;x�H;��H;B�H;|�H;��H;��H;v�H;N�H;�H;��H;�H;.�H;��H;I�H;=�H;��H;      ��H;��H;�H;��H;��H;��H;(�H;��H;�H;��H;�H;��H;��H;S�H;��H;��H;��H;��H;b�H;$�H;��H;�H;��H;��H;��H;.�H;<�H;B�H;S�H;I�H;T�H;Z�H;C�H;=�H;O�H;4�H;+�H;4�H;O�H;=�H;C�H;Z�H;T�H;I�H;S�H;B�H;<�H;.�H;��H;��H;��H;�H;��H;$�H;b�H;��H;��H;��H;��H;S�H;��H;��H;�H;��H;�H;��H;(�H;��H;��H;��H;�H;��H;      ��H;��H;�H;��H;)�H;��H;��H;��H;��H;��H;��H;�H;�H;�H;��H;��H;h�H;�H;��H; �H;m�H;��H;��H;,�H;=�H;C�H;\�H;k�H;j�H;Y�H;E�H;C�H;H�H;C�H;#�H;#�H;S�H;#�H;#�H;C�H;H�H;C�H;E�H;Y�H;j�H;k�H;\�H;C�H;=�H;,�H;��H;��H;m�H; �H;��H;�H;h�H;��H;��H;�H;�H;�H;��H;��H;��H;��H;��H;��H;)�H;��H;�H;��H;      p�H;�H;��H;��H;��H;�H;��H;{�H;9�H;��H;��H;n�H;'�H;��H;��H;,�H;��H;�H;w�H;��H;��H;1�H;L�H;l�H;��H;}�H;�H;l�H;l�H;h�H;E�H;=�H;C�H;-�H;�H;$�H;)�H;$�H;�H;-�H;C�H;=�H;E�H;h�H;l�H;l�H;�H;}�H;��H;l�H;L�H;1�H;��H;��H;w�H;�H;��H;,�H;��H;��H;'�H;n�H;��H;��H;9�H;{�H;��H;�H;��H;��H;��H;�H;      ��H;��H;��H;�H;p�H;��H;A�H;��H;R�H;��H;��H;�H;��H;*�H;��H;�H;Y�H;��H;�H;@�H;Y�H;r�H;��H;��H;��H;��H;��H;��H;j�H;P�H;c�H;O�H;#�H;�H;'�H;�H;�H;�H;'�H;�H;#�H;O�H;c�H;P�H;j�H;��H;��H;��H;��H;��H;��H;r�H;Y�H;@�H;�H;��H;Y�H;�H;��H;*�H;��H;�H;��H;��H;R�H;��H;A�H;��H;p�H;�H;��H;��H;      (�H;<�H;j�H;��H;��H;-�H;��H;�H;��H;�H;��H; �H;o�H;��H;B�H;��H;��H;�H;I�H;{�H;��H;��H;��H;��H;��H;��H;��H;��H;u�H;b�H;U�H;4�H;#�H;$�H;�H;�H;�H;�H;�H;$�H;#�H;4�H;U�H;b�H;u�H;��H;��H;��H;��H;��H;��H;��H;��H;{�H;I�H;�H;��H;��H;B�H;��H;o�H; �H;��H;�H;��H;�H;��H;-�H;��H;��H;j�H;<�H;      ��H;��H;��H;7�H;�H;��H;5�H;��H;�H;i�H;��H;?�H;��H;�H;u�H;��H;�H;<�H;c�H;{�H;��H;��H;��H;��H;��H;��H;��H;��H;u�H;{�H;6�H;+�H;S�H;)�H;�H;�H;�H;�H;�H;)�H;S�H;+�H;6�H;{�H;u�H;��H;��H;��H;��H;��H;��H;��H;��H;{�H;c�H;<�H;�H;��H;u�H;�H;��H;?�H;��H;i�H;�H;��H;5�H;��H;�H;7�H;��H;��H;      (�H;<�H;j�H;��H;��H;-�H;��H;�H;��H;�H;��H; �H;o�H;��H;B�H;��H;��H;�H;I�H;{�H;��H;��H;��H;��H;��H;��H;��H;��H;u�H;b�H;U�H;4�H;#�H;$�H;�H;�H;�H;�H;�H;$�H;#�H;4�H;U�H;b�H;u�H;��H;��H;��H;��H;��H;��H;��H;��H;{�H;I�H;�H;��H;��H;B�H;��H;o�H; �H;��H;�H;��H;�H;��H;-�H;��H;��H;j�H;<�H;      ��H;��H;��H;�H;p�H;��H;A�H;��H;R�H;��H;��H;�H;��H;*�H;��H;�H;Y�H;��H;�H;@�H;Y�H;r�H;��H;��H;��H;��H;��H;��H;j�H;P�H;c�H;O�H;#�H;�H;'�H;�H;�H;�H;'�H;�H;#�H;O�H;c�H;P�H;j�H;��H;��H;��H;��H;��H;��H;r�H;Y�H;@�H;�H;��H;Y�H;�H;��H;*�H;��H;�H;��H;��H;R�H;��H;A�H;��H;p�H;�H;��H;��H;      p�H;�H;��H;��H;��H;�H;��H;{�H;9�H;��H;��H;n�H;'�H;��H;��H;,�H;��H;�H;w�H;��H;��H;1�H;L�H;l�H;��H;}�H;�H;l�H;l�H;h�H;E�H;=�H;C�H;-�H;�H;$�H;)�H;$�H;�H;-�H;C�H;=�H;E�H;h�H;l�H;l�H;�H;}�H;��H;l�H;L�H;1�H;��H;��H;w�H;�H;��H;,�H;��H;��H;'�H;n�H;��H;��H;9�H;{�H;��H;�H;��H;��H;��H;�H;      ��H;��H;�H;��H;)�H;��H;��H;��H;��H;��H;��H;�H;�H;�H;��H;��H;h�H;�H;��H; �H;m�H;��H;��H;,�H;=�H;C�H;\�H;k�H;j�H;Y�H;E�H;C�H;H�H;C�H;#�H;#�H;S�H;#�H;#�H;C�H;H�H;C�H;E�H;Y�H;j�H;k�H;\�H;C�H;=�H;,�H;��H;��H;m�H; �H;��H;�H;h�H;��H;��H;�H;�H;�H;��H;��H;��H;��H;��H;��H;)�H;��H;�H;��H;      ��H;��H;�H;��H;��H;��H;(�H;��H;�H;��H;�H;��H;��H;S�H;��H;��H;��H;��H;b�H;$�H;��H;�H;��H;��H;��H;.�H;<�H;B�H;S�H;I�H;T�H;Z�H;C�H;=�H;O�H;4�H;+�H;4�H;O�H;=�H;C�H;Z�H;T�H;I�H;S�H;B�H;<�H;.�H;��H;��H;��H;�H;��H;$�H;b�H;��H;��H;��H;��H;S�H;��H;��H;�H;��H;�H;��H;(�H;��H;��H;��H;�H;��H;      i�H;��H;=�H;I�H;��H;.�H;�H;��H;�H;N�H;v�H;��H;��H;|�H;B�H;��H;x�H;��H;��H;��H;��H;4�H;��H;(�H;��H;��H;��H;�H;6�H;J�H;a�H;T�H;E�H;E�H;c�H;U�H;6�H;U�H;c�H;E�H;E�H;T�H;a�H;J�H;6�H;�H;��H;��H;��H;(�H;��H;4�H;��H;��H;��H;��H;x�H;��H;B�H;|�H;��H;��H;v�H;N�H;�H;��H;�H;.�H;��H;I�H;=�H;��H;      ��H;ݶH;��H;8�H;*�H;��H;S�H;N�H;W�H;��H;��H;��H;��H;n�H;��H;�H;;�H;�H;��H;��H;��H;�H;��H;~�H;�H;R�H;��H;��H;�H;+�H;J�H;I�H;Y�H;h�H;P�H;b�H;{�H;b�H;P�H;h�H;Y�H;I�H;J�H;+�H;�H;��H;��H;R�H;�H;~�H;��H;�H;��H;��H;��H;�H;;�H;�H;��H;n�H;��H;��H;��H;��H;W�H;N�H;S�H;��H;*�H;8�H;��H;ݶH;      3�H;ϠH;[�H;ĤH;��H;��H;��H;�H;��H;H�H;��H;J�H;b�H;J�H;�H;2�H;��H;h�H;��H;��H;<�H;�H;��H;��H;8�H;��H;[�H;��H;��H;�H;6�H;S�H;j�H;l�H;j�H;u�H;u�H;u�H;j�H;l�H;j�H;S�H;6�H;�H;��H;��H;[�H;��H;8�H;��H;��H;�H;<�H;��H;��H;h�H;��H;2�H;�H;J�H;b�H;J�H;��H;H�H;��H;�H;��H;��H;��H;ĤH;[�H;ϠH;      �kH;[mH;�qH;�xH;r�H;ȊH;�H;ʜH;��H; �H;��H;�H;&�H;��H;��H;K�H;Y�H;��H;��H;w�H;��H;��H;�H;G�H;T�H;�H;��H;B�H;��H;��H;�H;B�H;k�H;l�H;��H;��H;��H;��H;��H;l�H;k�H;B�H;�H;��H;��H;B�H;��H;�H;T�H;G�H;�H;��H;��H;w�H;��H;��H;Y�H;K�H;��H;��H;&�H;�H;��H; �H;��H;ʜH;�H;ȊH;r�H;�xH;�qH;[mH;      =�G;��G;/�G;��G;�H;�/H;�KH;?eH;_{H;i�H;m�H;d�H;o�H;��H;žH;3�H;��H;��H;��H;i�H;d�H;��H;#�H;��H;�H;9�H;�H;��H;[�H;��H;��H;<�H;\�H;�H;��H;��H;��H;��H;��H;�H;\�H;<�H;��H;��H;[�H;��H;�H;9�H;�H;��H;#�H;��H;d�H;i�H;��H;��H;��H;3�H;žH;��H;o�H;d�H;m�H;i�H;_{H;?eH;�KH;�/H;�H;��G;/�G;��G;      UHF;3TF;RvF;G�F;��F;�7G;��G;��G;�H;�<H;/eH;p�H;ÖH;�H;��H;ϸH;��H;��H;T�H;Q�H;Y�H;��H;w�H;��H;��H;	�H;9�H;�H;��H;R�H;��H;.�H;C�H;}�H;��H;��H;��H;��H;��H;}�H;C�H;.�H;��H;R�H;��H;�H;9�H;	�H;��H;��H;w�H;��H;Y�H;Q�H;T�H;��H;��H;ϸH;��H;�H;ÖH;p�H;/eH;�<H;�H;��G;��G;�7G;��F;G�F;RvF;3TF;      �B;.�B;�C;ՏC;�/D;��D;1�E;�HF;��F;GiG;R�G;t#H;�[H;/�H;��H;�H;I�H;μH;��H;d�H;��H;��H;�H;5�H;��H;��H;�H;T�H;8�H;�H;��H;��H;=�H;��H;��H;��H;��H;��H;��H;��H;=�H;��H;��H;�H;8�H;T�H;�H;��H;��H;5�H;�H;��H;��H;d�H;��H;μH;I�H;�H;��H;/�H;�[H;t#H;R�G;GiG;��F;�HF;1�E;��D;�/D;ՏC;�C;.�B;      D�:;\�:;��;;'�<;3>;�?;FIA;��B;DED;6{E;WvF;�7G;��G;q&H; eH;s�H;_�H;m�H;��H;��H;�H;:�H;�H;��H;5�H;��H;��H;G�H;��H;~�H;(�H;��H;,�H;l�H;��H;��H;��H;��H;��H;l�H;,�H;��H;(�H;~�H;��H;G�H;��H;��H;5�H;��H;�H;:�H;�H;��H;��H;m�H;_�H;s�H; eH;q&H;��G;�7G;WvF;6{E;DED;��B;FIA;�?;3>;'�<;��;;\�:;      *;��*;�,;�c.;�X1;#�4;E+8;ӊ;;~�>;IA;jwC;�)E;kF;�MG;'�G;DH;"{H;A�H;��H;@�H;S�H;Y�H;��H;�H;�H;w�H;#�H;�H;��H;��H;��H;��H;��H;L�H;��H;��H;��H;��H;��H;L�H;��H;��H;��H;��H;��H;�H;#�H;w�H;�H;�H;��H;Y�H;S�H;@�H;��H;A�H;"{H;DH;'�G;�MG;kF;�)E;jwC;IA;~�>;ӊ;;E+8;#�4;�X1;�c.;�,;��*;      ��
;��;J�;[;��;7`;�C&;�-;�C3;t�8;?H=;��@;�C;c{E;��F;�G;k#H;,mH;��H;?�H;��H;��H;Y�H;:�H;��H;��H;��H;��H;�H;�H;4�H;�H;��H;1�H;r�H;��H;��H;��H;r�H;1�H;��H;�H;4�H;�H;�H;��H;��H;��H;��H;:�H;Y�H;��H;��H;?�H;��H;,mH;k#H;�G;��F;c{E;�C;��@;?H=;t�8;�C3;�-;�C&;7`;��;[;J�;��;      \�:���:��:Ҳ�:���:PO�:�z;i';4�;�}(;�X1;6t8;��=;Z�A;��D;&HF;�bG;�H;>cH;��H;m�H;��H;S�H;�H;��H;Y�H;d�H;��H;<�H;��H;��H;��H;m�H;��H;Y�H;��H;��H;��H;Y�H;��H;m�H;��H;��H;��H;<�H;��H;d�H;Y�H;��H;�H;S�H;��H;m�H;��H;>cH;�H;�bG;&HF;��D;Z�A;��=;6t8;�X1;�}(;4�;i';�z;PO�:���:Ҳ�:��:���:      �R�� ���7�<^9��:P�X:���:���:�O�:=�;7�;�);�C3;��:;� @;�C;k�E;8G;��G;�_H;��H;?�H;@�H;��H;d�H;Q�H;i�H;w�H;��H;��H;��H;$�H; �H;��H;@�H;{�H;{�H;{�H;@�H;��H; �H;$�H;��H;��H;��H;w�H;i�H;Q�H;d�H;��H;@�H;?�H;��H;�_H;��G;8G;k�E;�C;� @;��:;�C3;�);7�;=�;�O�:���:���:P�X:��:<^9��7�� �      ��)���$�����������=�\�
S���N�9�1j:a��:���:ڃ;�� ;%d.;+8;��>;qC;��E;�(G;��G;>cH;��H;��H;��H;��H;T�H;��H;��H;��H;��H;��H;b�H;��H;w�H;�H;I�H;c�H;I�H;�H;w�H;��H;b�H;��H;��H;��H;��H;��H;T�H;��H;��H;��H;��H;>cH;��G;�(G;��E;qC;��>;+8;%d.;�� ;ڃ;���:a��:�1j:�N�9
S��=�\�������������$�      q�ѻ�ͻP���mG�������d�*�$��Jɺ͇!��C^9��r:���:`0;y�;l�*;�Y6;>;n�B;��E;8G;�H;,mH;A�H;m�H;μH;��H;��H;��H;h�H;�H;��H;��H;�H;�H;��H;�H;<�H;�H;��H;�H;�H;��H;��H;�H;h�H;��H;��H;��H;μH;m�H;A�H;,mH;�H;8G;��E;n�B;>;�Y6;l�*;y�;`0;���:��r:�C^9͇!��Jɺ*�$���d����mG��P����ͻ      ��I�1�E��(;��O*�����<��?GĻ��t@�JҺ{��:�:�O�:O�; ~(;S�5;>;qC;k�E;�bG;k#H;"{H;_�H;I�H;��H;��H;Y�H;��H;;�H;x�H;��H;h�H;��H;Y�H;��H;�H;��H;Y�H;��H;h�H;��H;x�H;;�H;��H;Y�H;��H;��H;I�H;_�H;"{H;k#H;�bG;k�E;qC;>;S�5; ~(;O�;�O�:�:��:{��JҺt@���?GĻ�<������O*��(;�1�E�      &p��\x��ע��R��%��n�`��7�F��G�ѻ-��˃$��ǅ���09�:���:�; ~(;�Y6;��>;�C;&HF;�G;DH;s�H;�H;ϸH;3�H;K�H;2�H;�H;��H;��H;��H;,�H;�H;��H;��H;��H;�H;,�H;��H;��H;��H;�H;2�H;K�H;3�H;ϸH;�H;s�H;DH;�G;&HF;�C;��>;�Y6; ~(;�;���:�:��09�ǅ�˃$�-��G�ѻF���7�n�`�%���R��ע�\x��      &]� �%#�����u�ټ�ɺ������
v��(;�ר�c^��P6R�����	7����:���:O�;l�*;+8;� @;��D;��F;'�G; eH;��H;��H;žH;��H;�H;��H;B�H;��H;��H;��H;��H;B�H;u�H;B�H;��H;��H;��H;��H;B�H;��H;�H;��H;žH;��H;��H; eH;'�G;��F;��D;� @;+8;l�*;O�;���:���:�	7����P6R�c^��ר��(;��
v������ɺ�u�ټ����%#� �      ��_�\�<Q��f@�t +��5�����P�ļs�\�`����bͻfk��Iɺ�	7��:�O�:y�;%d.;��:;Z�A;c{E;�MG;q&H;/�H;�H;��H;��H;J�H;n�H;|�H;S�H;�H;��H;*�H;��H;�H;��H;*�H;��H;�H;S�H;|�H;n�H;J�H;��H;��H;�H;/�H;q&H;�MG;c{E;Z�A;��:;%d.;y�;�O�:�:�	7��Iɺfk�bͻ���\�`�s�P�ļ�����5�t +��f@�<Q�\�      �@���R��ڟ�绒�C����_�:�������$p���vz��O*�5ֻfk������09�:`0;�� ;�C3;��=;�C;kF;��G;�[H;ÖH;o�H;&�H;b�H;��H;��H;��H;�H;'�H;��H;o�H;��H;o�H;��H;'�H;�H;��H;��H;��H;b�H;&�H;o�H;ÖH;�[H;��G;kF;�C;��=;�C3;�� ;`0;�:��09���fk�5ֻ�O*��vz�$p����輙��:���_�C��绒�ڟ��R��      �` �j.��m��ڽ�b��gr��O��\�m +�� ��ɺ�<��O*�bͻP6R��ǅ���:���:ڃ;�);6t8;��@;�)E;�7G;t#H;p�H;d�H;�H;J�H;��H;��H;��H;�H;n�H;�H; �H;?�H; �H;�H;n�H;�H;��H;��H;��H;J�H;�H;d�H;p�H;t#H;�7G;�)E;��@;6t8;�);ڃ;���:��:�ǅ�P6R�bͻ�O*�<��ɺ�� �m +�\�O��gr���b����ڽm��j.��      �-=�1�9��k/�"�����i��y�Ľ�!��Tys�4�6�#��ɺ��vz����c^��˃$�{����r:���:7�;�X1;?H=;jwC;WvF;R�G;/eH;m�H;��H;��H;��H;v�H;�H;��H;��H;��H;��H;��H;��H;��H;��H;��H;�H;v�H;��H;��H;��H;m�H;/eH;R�G;WvF;jwC;?H=;�X1;7�;���:��r:{��˃$�c^������vz��ɺ�#�4�6�Tys��!��y�Ľi���"���k/�1�9�      �(��;l���.}�&ce�jPH���(�o
���ڽ�R����{�4�6�� �$p��\�`�ר�-��JҺ�C^9a��:=�;�}(;t�8;IA;6{E;GiG;�<H;i�H; �H;H�H;��H;N�H;��H;��H;��H;��H;�H;i�H;�H;��H;��H;��H;��H;N�H;��H;H�H; �H;i�H;�<H;GiG;6{E;IA;t�8;�}(;=�;a��:�C^9JҺ-��ר�\�`�$p��� �4�6���{��R����ڽo
���(�jPH�&ce��.}�;l��      �iþGD��)o���������� �i��-=�[t����R��Tys�m +����s񗼗(;�G�ѻt@�͇!��1j:�O�:4�;�C3;~�>;DED;��F;�H;_{H;��H;��H;W�H;�H;�H;��H;9�H;R�H;��H;�H;��H;R�H;9�H;��H;�H;�H;W�H;��H;��H;_{H;�H;��F;DED;~�>;�C3;4�;�O�:�1j:͇!�t@�G�ѻ�(;�s����m +�Tys��R����[t��-=� �i���������)o��GD��      ���
������޾HD���A���.}��D�[t���ڽ�!��\����P�ļ�
v�F�����Jɺ�N�9���:i';�-;ӊ;;��B;�HF;��G;?eH;ʜH;�H;N�H;��H;��H;��H;{�H;��H;�H;��H;�H;��H;{�H;��H;��H;��H;N�H;�H;ʜH;?eH;��G;�HF;��B;ӊ;;�-;i';���:�N�9�Jɺ��F���
v�P�ļ���\��!����ڽ[t��D��.}��A��HD���޾�����
�      ��7�Õ3��f'���\���о�����.}��-=�o
�y�ĽO��:����������7�?GĻ*�$�
S�����:�z;�C&;E+8;FIA;1�E;��G;�KH;�H;��H;S�H;�H;(�H;��H;��H;A�H;��H;5�H;��H;A�H;��H;��H;(�H;�H;S�H;��H;�H;�KH;��G;1�E;FIA;E+8;�C&;�z;���:
S��*�$�?GĻ�7���������:�O��y�Ľo
��-=��.}������о�\����f'�Õ3�      Io�PXi�s"Y���@�@�#��
��о�A�� �i���(�i��gr����_��5��ɺ�n�`��<����d�=�\�P�X:PO�:7`;#�4;�?;��D;�7G;�/H;ȊH;��H;��H;.�H;��H;��H;�H;��H;-�H;��H;-�H;��H;�H;��H;��H;.�H;��H;��H;ȊH;�/H;�7G;��D;�?;#�4;7`;PO�:P�X:=�\���d��<��n�`��ɺ��5���_�gr��i����(� �i��A���о�
�@�#���@�s"Y�PXi�      &����������Io��!J�@�#��\��HD������jPH�����b��C��t +�u�ټ%��������������:���:��;�X1;3>;�/D;��F;�H;r�H;��H;*�H;��H;��H;)�H;��H;p�H;��H;�H;��H;p�H;��H;)�H;��H;��H;*�H;��H;r�H;�H;��F;�/D;3>;�X1;��;���:��:����������%��u�ټt +�C���b�����jPH�����HD���\��@�#��!J�Io��������      2^������b���Io���@���޾����&ce�"����ڽ绒��f@������R���O*�mG�����<^9Ҳ�:[;�c.;'�<;ՏC;G�F;��G;�xH;ĤH;8�H;I�H;��H;��H;��H;�H;��H;7�H;��H;�H;��H;��H;��H;I�H;8�H;ĤH;�xH;��G;G�F;ՏC;'�<;�c.;[;Ҳ�:<^9���mG���O*��R�������f@�绒���ڽ"��&ce������޾���@�Io�b�������      �aǿ֊¿���������s"Y��f'�����)o���.}��k/�m��ڟ�<Q�%#�ע��(;�P��������7���:J�;�,;��;;�C;RvF;/�G;�qH;[�H;��H;=�H;�H;�H;��H;��H;j�H;��H;j�H;��H;��H;�H;�H;=�H;��H;[�H;�qH;/�G;RvF;�C;��;;�,;J�;��:��7����P����(;�ע�%#�<Q�ڟ�m���k/��.}�)o�������f'�s"Y����������֊¿      %�ֿ5pѿ֊¿������PXi�Õ3��
�GD��;l��1�9�j.���R��\� �\x��1�E��ͻ��$�� ����:��;��*;\�:;.�B;3TF;��G;[mH;ϠH;ݶH;��H;��H;��H;�H;��H;<�H;��H;<�H;��H;�H;��H;��H;��H;ݶH;ϠH;[mH;��G;3TF;.�B;\�:;��*;��;���:� ���$��ͻ1�E�\x�� �\��R��j.��1�9�;l��GD���
�Õ3�PXi�������֊¿5pѿ      �?��ph��2v��� ��$�X��O/�#y�-�;Ѱ��j+X�����ѽ����Gn;�>�＿����B(�嚩����/�e9��:^;Y.;��<;�VC;@ZF;�G;5/H;tiH;X�H;s�H;��H;E�H;��H;�H;��H;��H;��H;�H;��H;E�H;��H;s�H;X�H;tiH;5/H;�G;@ZF;�VC;��<;Y.;^;��:/�e9���嚩��B(�����>��Gn;�������ѽ��j+X�Ѱ��-�;#y��O/�$�X�� ��2v��ph��      ph��"���V�����y�EvS�aM+��v� 9ɾ�����T�]��[ν����`\8�����x���%�[��������9C,�:��;�.;N�<; nC;�cF;�G;�0H;!jH;ǋH;ңH;��H;��H;��H;��H;��H;��H;��H;��H;��H;��H;��H;ңH;ǋH;!jH;�0H;�G;�cF; nC;N�<;�.;��;C,�:��9���[����%��x�����`\8������[ν]��T����� 9ɾ�v�aM+�EvS���y�V���"���      2v��V���L ��M�h�%E�I��R���i㼾n���nH�È�a�ý�Ȅ��s/��o༼#�����4J���к��9$f�:Nl;�0;P\=; �C;6�F;��G;Q5H;^lH;H�H;ФH;��H;�H;b�H;��H;$�H;�H;$�H;��H;b�H;�H;��H;ФH;H�H;^lH;Q5H;��G;6�F; �C;P\=;�0;Nl;$f�:��9�к4J������#���o��s/��Ȅ�a�ýÈ��nH�n��i㼾R���I��%E�M�h�L ��V���      � ����y�M�h�ބN��O/����-�߾�A���*|�ؕ6�a}��㳽KSt�(�!�Wrμ(F{��_�
Y��f����:���:WZ;2;�N>;�D;��F;��G;J<H;�oH;��H;t�H;��H;��H;��H;��H;��H;�H;��H;��H;��H;��H;��H;t�H;��H;�oH;J<H;��G;��F;�D;�N>;2;WZ;���:�:f���
Y���_�(F{�Wrμ(�!�KSt��㳽a}�ؕ6��*|��A��-�߾����O/�ބN�M�h���y�      $�X�EvS�%E��O/��S�1W����������4S\�� �q�&�����Y�h��������]�|���S�b��Y���Y:�~�:�_;��4;�?;}�D;�F;/�G;5EH;tH;�H;��H;��H;3�H;��H;E�H;8�H;�H;8�H;E�H;��H;3�H;��H;��H;�H;tH;5EH;/�G;�F;}�D;�?;��4;�_;�~�:��Y:�Y�S�b�|�����]�����h����Y�&���q�� �4S\���������1W���S��O/�%E�EvS�      �O/�aM+�I�����1W�� 9ɾ0���Mw�� :�Y��_�ý�L��Dn;�>���bv���E<��˻(�-�����x�:^;%;�7;��@;V4E;�!G;,�G;iOH;1zH;�H;��H;��H;��H;�H;2�H;�H;��H;�H;2�H;�H;��H;��H;��H;�H;1zH;iOH;,�G;�!G;V4E;��@;�7;%;^;�x�:���(�-��˻�E<�bv��>���Dn;��L��_�ýY��� :��Mw�0�� 9ɾ1W�����I��aM+�      #y��v�R���-�߾����0��1����nH���(Ὁu��r�d�O�Prμ<"�����	��1���k89w:�:��;+;�{:;�6B;)�E;FaG;�H;ZH;��H;M�H;ĮH;�H;e�H;e�H;+�H;��H;��H;��H;+�H;e�H;e�H;�H;ĮH;M�H;��H;ZH;�H;FaG;)�E;�6B;�{:;+;��;w:�:�k891��	�����<"��PrμO�r�d��u��(����nH�1���0������-�߾R����v�      -�; 9ɾi㼾�A�������Mw��nH�����Z��㳽����Z\8�O#�������]N�J��-�b�VJx�z5:��:��;8�0;v\=;v�C;�ZF;�G;)H;eH;��H;G�H;g�H;��H;7�H;��H;P�H;��H;��H;��H;P�H;��H;7�H;��H;g�H;G�H;��H;eH;)H;�G;�ZF;v�C;v\=;8�0;��;��:z5:VJx�-�b�J���]N�����O#��Z\8������㳽�Z񽞯��nH��Mw������A��i㼾 9ɾ      Ѱ������n���*|�4S\�� :����Z�U$������K�c���Oļ����������x&�#��P.�:0^;��#;G6;��?;-�D;��F;��G;*?H;�oH;�H;��H;:�H;r�H;J�H;��H;��H;��H;��H;��H;��H;��H;J�H;r�H;:�H;��H;�H;�oH;*?H;��G;��F;-�D;��?;G6;��#;0^;P.�:#��x&������������Oļc���K����U$���Z���� :�4S\��*|�n������      j+X��T��nH�ؕ6�� �Y��(��㳽����mR����ټ�����E<��?ݻad\�a ��%:�c�:8�;z�,;��:;�6B;ͱE;�KG;jH;�RH;�zH;��H;
�H;9�H;`�H;n�H;+�H;��H;�H;��H;�H;��H;+�H;n�H;`�H;9�H;
�H;��H;�zH;�RH;jH;�KG;ͱE;�6B;��:;z�,;8�;�c�:%:a ��ad\��?ݻ�E<������ټ���mR�����㳽(�Y��� �ؕ6��nH��T�      ��]�È�a}�q�_�ý�u�������K����o�Wv���&R���e^���뺪@���:�A;�";��4;��>;�D;F;,�G;)H;�cH;��H;5�H;��H;N�H;M�H;��H;��H;<�H;(�H;��H;(�H;<�H;��H;��H;M�H;N�H;��H;5�H;��H;�cH;)H;,�G;F;�D;��>;��4;�";�A;��:�@���e^�����&R�Wv���o����K������u��_�ýq�a}�È�]�      ��ѽ�[νa�ý�㳽&����L��r�d�Z\8�c���ټWv����Y��_����y��]���Y:@��:�l; r-;R�:;��A;rnE;�!G;��G;�FH;�rH;�H;��H;�H;J�H;5�H;��H;��H;��H;B�H;�H;B�H;��H;��H;��H;5�H;J�H;�H;��H;�H;�rH;�FH;��G;�!G;rnE;��A;R�:; r-;�l;@��:��Y:]�y������_���Y�Wv���ټc��Z\8�r�d��L��&����㳽a�ý�[ν      ���������Ȅ�KSt���Y�Dn;�O�O#���Oļ�����&R��_������N3�,�Y�02:�:9�;A?&;)G6;�W?;�D;fwF;�G;c H;�]H;��H;�H;�H;a�H;$�H;�H;��H;(�H;��H;i�H;%�H;i�H;��H;(�H;��H;�H;$�H;a�H;�H;�H;��H;�]H;c H;�G;fwF;�D;�W?;)G6;A?&;9�;�:02:,�Y��N3������_��&R������OļO#��O�Dn;���Y�KSt��Ȅ�����      Gn;�`\8��s/�(�!�h��>���Prμ��������E<�������N3��Ix�f�9��:U^;� ;2;��<;.�B;�E;f4G;2�G;^EH;�pH;��H;h�H;гH;k�H;��H;��H;�H;��H;1�H;��H;�H;��H;1�H;��H;�H;��H;��H;k�H;гH;h�H;��H;�pH;^EH;2�G;f4G;�E;.�B;��<;2;� ;U^;��:f�9�Ix��N3�������E<��������Prμ>���h��(�!��s/�`\8�      >�Ｘ���o�Wrμ����bv��<"���]N�����?ݻe^��y��,�Y�f�9��:���:B�;��.;�{:;2>A;��D;`�F;�G;
)H;E`H;5�H;��H;�H;R�H;6�H;R�H;t�H;�H;/�H;k�H;��H;��H;��H;k�H;/�H;�H;t�H;R�H;6�H;R�H;�H;��H;5�H;E`H;
)H;�G;`�F;��D;2>A;�{:;��.;B�;���:��:f�9,�Y�y��e^���?ݻ����]N�<"��bv������Wrμ�o༸��      �����x���#��(F{���]��E<����J�뻱���ad\���]�02:��:���:�Z;��,;0�8;a @;0D;�ZF;QzG;
H;jOH;>uH;�H;\�H;�H;C�H;z�H;��H;��H;��H;��H;��H;��H;��H;��H;��H;��H;��H;��H;��H;z�H;C�H;�H;\�H;�H;>uH;jOH;
H;QzG;�ZF;0D;a @;0�8;��,;�Z;���:��:02:]���ad\�����J�뻛���E<���]�(F{��#���x��      �B(��%�����_�|����˻	��-�b�x&�a ���@���Y:�:U^;B�;��,;Z_8;��?;��C;�F;FG;u�G;?H;GjH;#�H; �H;
�H;k�H;��H;�H;��H;/�H;��H;��H;��H;��H;��H;��H;��H;��H;��H;/�H;��H;�H;��H;k�H;
�H; �H;#�H;GjH;?H;u�G;FG;�F;��C;��?;Z_8;��,;B�;U^;�:��Y:�@�a ��x&�-�b�	���˻|����_�����%�      嚩�[���4J��
Y��S�b�(�-�1��VJx�#��%:��:@��:9�;� ;��.;0�8;��?;2�C;�E;f"G;�G;1H;aH;gH;��H;��H;��H;��H;s�H;(�H;I�H;J�H;��H;(�H;��H;H�H;��H;H�H;��H;(�H;��H;J�H;I�H;(�H;s�H;��H;��H;��H;��H;gH;aH;1H;�G;f"G;�E;2�C;��?;0�8;��.;� ;9�;@��:��:%:#��VJx�1��(�-�S�b�
Y��4J��[���      �����뺶кf����Y�����k89z5:P.�:�c�:�A;�l;A?&;2;�{:;a @;��C;�E;�G;�G;}'H;ZH;�yH;X�H;��H;��H;{�H;��H;��H;l�H;��H;�H;[�H;<�H;W�H;
�H;��H;
�H;W�H;<�H;[�H;�H;��H;l�H;��H;��H;{�H;��H;��H;X�H;�yH;ZH;}'H;�G;�G;�E;��C;a @;�{:;2;A?&;�l;�A;�c�:P.�:z5:�k89����Y�f����к���      /�e9��9��9�:��Y:�x�:w:�:��:0^;8�;�"; r-;)G6;��<;2>A;0D;�F;f"G;�G;$H;VH;�uH;��H;Y�H;b�H;��H;!�H;��H;��H;E�H;��H;��H;��H;7�H;�H;��H;�H;��H;�H;7�H;��H;��H;��H;E�H;��H;��H;!�H;��H;b�H;Y�H;��H;�uH;VH;$H;�G;f"G;�F;0D;2>A;��<;)G6; r-;�";8�;0^;��:w:�:�x�:��Y:�:��9��9      ��:C,�:$f�:���:�~�:^;��;��;��#;z�,;��4;R�:;�W?;.�B;��D;�ZF;FG;�G;}'H;VH;�tH;��H;.�H;�H;<�H;
�H;��H;��H;��H;��H;��H;��H;��H;��H;��H;^�H;b�H;^�H;��H;��H;��H;��H;��H;��H;��H;��H;��H;
�H;<�H;�H;.�H;��H;�tH;VH;}'H;�G;FG;�ZF;��D;.�B;�W?;R�:;��4;z�,;��#;��;��;^;�~�:���:$f�:C,�:      ^;��;Nl;WZ;�_;%;+;8�0;G6;��:;��>;��A;�D;�E;`�F;QzG;u�G;1H;ZH;�uH;��H;g�H;ܫH;�H;��H;e�H;��H;��H;��H;��H;H�H;G�H;��H;��H;p�H;��H;��H;��H;p�H;��H;��H;G�H;H�H;��H;��H;��H;��H;e�H;��H;�H;ܫH;g�H;��H;�uH;ZH;1H;u�G;QzG;`�F;�E;�D;��A;��>;��:;G6;8�0;+;%;�_;WZ;Nl;��;      Y.;�.;�0;2;��4;�7;�{:;v\=;��?;�6B;�D;rnE;fwF;f4G;�G;
H;?H;aH;�yH;��H;.�H;ܫH;`�H;��H;�H;��H;��H;�H;)�H;��H;��H;h�H;c�H;O�H;��H;(�H;P�H;(�H;��H;O�H;c�H;h�H;��H;��H;)�H;�H;��H;��H;�H;��H;`�H;ܫH;.�H;��H;�yH;aH;?H;
H;�G;f4G;fwF;rnE;�D;�6B;��?;v\=;�{:;�7;��4;2;�0;�.;      ��<;N�<;P\=;�N>;�?;��@;�6B;v�C;-�D;ͱE;F;�!G;�G;2�G;
)H;jOH;GjH;gH;X�H;Y�H;�H;�H;��H;H�H;I�H;E�H;X�H;��H;,�H;B�H;�H;�H;�H;��H;I�H;��H;��H;��H;I�H;��H;�H;�H;�H;B�H;,�H;��H;X�H;E�H;I�H;H�H;��H;�H;�H;Y�H;X�H;gH;GjH;jOH;
)H;2�G;�G;�!G;F;ͱE;-�D;v�C;�6B;��@;�?;�N>;P\=;N�<;      �VC; nC; �C;�D;}�D;V4E;)�E;�ZF;��F;�KG;,�G;��G;c H;^EH;E`H;>uH;#�H;��H;��H;b�H;<�H;��H;�H;I�H;�H;�H;O�H;��H;��H;��H;��H;��H;��H;=�H;��H;��H;��H;��H;��H;=�H;��H;��H;��H;��H;��H;��H;O�H;�H;�H;I�H;�H;��H;<�H;b�H;��H;��H;#�H;>uH;E`H;^EH;c H;��G;,�G;�KG;��F;�ZF;)�E;V4E;}�D;�D; �C; nC;      @ZF;�cF;6�F;��F;�F;�!G;FaG;�G;��G;jH;)H;�FH;�]H;�pH;5�H;�H; �H;��H;��H;��H;
�H;e�H;��H;E�H;�H;6�H;��H;��H;u�H;��H;��H;��H;,�H;~�H;��H;�H;�H;�H;��H;~�H;,�H;��H;��H;��H;u�H;��H;��H;6�H;�H;E�H;��H;e�H;
�H;��H;��H;��H; �H;�H;5�H;�pH;�]H;�FH;)H;jH;��G;�G;FaG;�!G;�F;��F;6�F;�cF;      �G;�G;��G;��G;/�G;,�G;�H;)H;*?H;�RH;�cH;�rH;��H;��H;��H;\�H;
�H;��H;{�H;!�H;��H;��H;��H;X�H;O�H;��H;��H;J�H;��H;��H;j�H; �H;}�H;��H;�H;;�H;Y�H;;�H;�H;��H;}�H; �H;j�H;��H;��H;J�H;��H;��H;O�H;X�H;��H;��H;��H;!�H;{�H;��H;
�H;\�H;��H;��H;��H;�rH;�cH;�RH;*?H;)H;�H;,�G;/�G;��G;��G;�G;      5/H;�0H;Q5H;J<H;5EH;iOH;ZH;eH;�oH;�zH;��H;�H;�H;h�H;�H;�H;k�H;��H;��H;��H;��H;��H;�H;��H;��H;��H;J�H;��H;e�H;S�H;�H;j�H;��H;�H;E�H;[�H;M�H;[�H;E�H;�H;��H;j�H;�H;S�H;e�H;��H;J�H;��H;��H;��H;�H;��H;��H;��H;��H;��H;k�H;�H;�H;h�H;�H;�H;��H;�zH;�oH;eH;ZH;iOH;5EH;J<H;Q5H;�0H;      tiH;!jH;^lH;�oH;tH;1zH;��H;��H;�H;��H;5�H;��H;�H;гH;R�H;C�H;��H;s�H;��H;��H;��H;��H;)�H;,�H;��H;u�H;��H;e�H;[�H;��H;Z�H;��H;��H;5�H;e�H;o�H;b�H;o�H;e�H;5�H;��H;��H;Z�H;��H;[�H;e�H;��H;u�H;��H;,�H;)�H;��H;��H;��H;��H;s�H;��H;C�H;R�H;гH;�H;��H;5�H;��H;�H;��H;��H;1zH;tH;�oH;^lH;!jH;      X�H;ǋH;H�H;��H;�H;�H;M�H;G�H;��H;
�H;��H;�H;a�H;k�H;6�H;z�H;�H;(�H;l�H;E�H;��H;��H;��H;B�H;��H;��H;��H;S�H;��H;K�H;��H;��H;6�H;]�H;h�H;��H;��H;��H;h�H;]�H;6�H;��H;��H;K�H;��H;S�H;��H;��H;��H;B�H;��H;��H;��H;E�H;l�H;(�H;�H;z�H;6�H;k�H;a�H;�H;��H;
�H;��H;G�H;M�H;�H;�H;��H;H�H;ǋH;      s�H;ңH;ФH;t�H;��H;��H;ĮH;g�H;:�H;9�H;N�H;J�H;$�H;��H;R�H;��H;��H;I�H;��H;��H;��H;H�H;��H;�H;��H;��H;j�H;�H;Z�H;��H;��H;)�H;a�H;o�H;��H;��H;��H;��H;��H;o�H;a�H;)�H;��H;��H;Z�H;�H;j�H;��H;��H;�H;��H;H�H;��H;��H;��H;I�H;��H;��H;R�H;��H;$�H;J�H;N�H;9�H;:�H;g�H;ĮH;��H;��H;t�H;ФH;ңH;      ��H;��H;��H;��H;��H;��H;�H;��H;r�H;`�H;M�H;5�H;�H;��H;t�H;��H;/�H;J�H;�H;��H;��H;G�H;h�H;�H;��H;��H; �H;j�H;��H;��H;)�H;A�H;l�H;��H;��H;��H;��H;��H;��H;��H;l�H;A�H;)�H;��H;��H;j�H; �H;��H;��H;�H;h�H;G�H;��H;��H;�H;J�H;/�H;��H;t�H;��H;�H;5�H;M�H;`�H;r�H;��H;�H;��H;��H;��H;��H;��H;      E�H;��H;�H;��H;3�H;��H;e�H;7�H;J�H;n�H;��H;��H;��H;�H;�H;��H;��H;��H;[�H;��H;��H;��H;c�H;�H;��H;,�H;}�H;��H;��H;6�H;a�H;l�H;{�H;��H;��H;��H;��H;��H;��H;��H;{�H;l�H;a�H;6�H;��H;��H;}�H;,�H;��H;�H;c�H;��H;��H;��H;[�H;��H;��H;��H;�H;�H;��H;��H;��H;n�H;J�H;7�H;e�H;��H;3�H;��H;�H;��H;      ��H;��H;b�H;��H;��H;�H;e�H;��H;��H;+�H;��H;��H;(�H;��H;/�H;��H;��H;(�H;<�H;7�H;��H;��H;O�H;��H;=�H;~�H;��H;�H;5�H;]�H;o�H;��H;��H;��H;��H;��H;��H;��H;��H;��H;��H;��H;o�H;]�H;5�H;�H;��H;~�H;=�H;��H;O�H;��H;��H;7�H;<�H;(�H;��H;��H;/�H;��H;(�H;��H;��H;+�H;��H;��H;e�H;�H;��H;��H;b�H;��H;      �H;��H;��H;��H;E�H;2�H;+�H;P�H;��H;��H;<�H;��H;��H;1�H;k�H;��H;��H;��H;W�H;�H;��H;p�H;��H;I�H;��H;��H;�H;E�H;e�H;h�H;��H;��H;��H;��H;��H;��H;��H;��H;��H;��H;��H;��H;��H;h�H;e�H;E�H;�H;��H;��H;I�H;��H;p�H;��H;�H;W�H;��H;��H;��H;k�H;1�H;��H;��H;<�H;��H;��H;P�H;+�H;2�H;E�H;��H;��H;��H;      ��H;��H;$�H;��H;8�H;�H;��H;��H;��H;�H;(�H;B�H;i�H;��H;��H;��H;��H;H�H;
�H;��H;^�H;��H;(�H;��H;��H;�H;;�H;[�H;o�H;��H;��H;��H;��H;��H;��H;��H;��H;��H;��H;��H;��H;��H;��H;��H;o�H;[�H;;�H;�H;��H;��H;(�H;��H;^�H;��H;
�H;H�H;��H;��H;��H;��H;i�H;B�H;(�H;�H;��H;��H;��H;�H;8�H;��H;$�H;��H;      ��H;��H;�H;�H;�H;��H;��H;��H;��H;��H;��H;�H;%�H;�H;��H;��H;��H;��H;��H;�H;b�H;��H;P�H;��H;��H;�H;Y�H;M�H;b�H;��H;��H;��H;��H;��H;��H;��H;��H;��H;��H;��H;��H;��H;��H;��H;b�H;M�H;Y�H;�H;��H;��H;P�H;��H;b�H;�H;��H;��H;��H;��H;��H;�H;%�H;�H;��H;��H;��H;��H;��H;��H;�H;�H;�H;��H;      ��H;��H;$�H;��H;8�H;�H;��H;��H;��H;�H;(�H;B�H;i�H;��H;��H;��H;��H;H�H;
�H;��H;^�H;��H;(�H;��H;��H;�H;;�H;[�H;o�H;��H;��H;��H;��H;��H;��H;��H;��H;��H;��H;��H;��H;��H;��H;��H;o�H;[�H;;�H;�H;��H;��H;(�H;��H;^�H;��H;
�H;H�H;��H;��H;��H;��H;i�H;B�H;(�H;�H;��H;��H;��H;�H;8�H;��H;$�H;��H;      �H;��H;��H;��H;E�H;2�H;+�H;P�H;��H;��H;<�H;��H;��H;1�H;k�H;��H;��H;��H;W�H;�H;��H;p�H;��H;I�H;��H;��H;�H;E�H;e�H;h�H;��H;��H;��H;��H;��H;��H;��H;��H;��H;��H;��H;��H;��H;h�H;e�H;E�H;�H;��H;��H;I�H;��H;p�H;��H;�H;W�H;��H;��H;��H;k�H;1�H;��H;��H;<�H;��H;��H;P�H;+�H;2�H;E�H;��H;��H;��H;      ��H;��H;b�H;��H;��H;�H;e�H;��H;��H;+�H;��H;��H;(�H;��H;/�H;��H;��H;(�H;<�H;7�H;��H;��H;O�H;��H;=�H;~�H;��H;�H;5�H;]�H;o�H;��H;��H;��H;��H;��H;��H;��H;��H;��H;��H;��H;o�H;]�H;5�H;�H;��H;~�H;=�H;��H;O�H;��H;��H;7�H;<�H;(�H;��H;��H;/�H;��H;(�H;��H;��H;+�H;��H;��H;e�H;�H;��H;��H;b�H;��H;      E�H;��H;�H;��H;3�H;��H;e�H;7�H;J�H;n�H;��H;��H;��H;�H;�H;��H;��H;��H;[�H;��H;��H;��H;c�H;�H;��H;,�H;}�H;��H;��H;6�H;a�H;l�H;{�H;��H;��H;��H;��H;��H;��H;��H;{�H;l�H;a�H;6�H;��H;��H;}�H;,�H;��H;�H;c�H;��H;��H;��H;[�H;��H;��H;��H;�H;�H;��H;��H;��H;n�H;J�H;7�H;e�H;��H;3�H;��H;�H;��H;      ��H;��H;��H;��H;��H;��H;�H;��H;r�H;`�H;M�H;5�H;�H;��H;t�H;��H;/�H;J�H;�H;��H;��H;G�H;h�H;�H;��H;��H; �H;j�H;��H;��H;)�H;A�H;l�H;��H;��H;��H;��H;��H;��H;��H;l�H;A�H;)�H;��H;��H;j�H; �H;��H;��H;�H;h�H;G�H;��H;��H;�H;J�H;/�H;��H;t�H;��H;�H;5�H;M�H;`�H;r�H;��H;�H;��H;��H;��H;��H;��H;      s�H;ңH;ФH;t�H;��H;��H;ĮH;g�H;:�H;9�H;N�H;J�H;$�H;��H;R�H;��H;��H;I�H;��H;��H;��H;H�H;��H;�H;��H;��H;j�H;�H;Z�H;��H;��H;)�H;a�H;o�H;��H;��H;��H;��H;��H;o�H;a�H;)�H;��H;��H;Z�H;�H;j�H;��H;��H;�H;��H;H�H;��H;��H;��H;I�H;��H;��H;R�H;��H;$�H;J�H;N�H;9�H;:�H;g�H;ĮH;��H;��H;t�H;ФH;ңH;      X�H;ǋH;H�H;��H;�H;�H;M�H;G�H;��H;
�H;��H;�H;a�H;k�H;6�H;z�H;�H;(�H;l�H;E�H;��H;��H;��H;B�H;��H;��H;��H;S�H;��H;K�H;��H;��H;6�H;]�H;h�H;��H;��H;��H;h�H;]�H;6�H;��H;��H;K�H;��H;S�H;��H;��H;��H;B�H;��H;��H;��H;E�H;l�H;(�H;�H;z�H;6�H;k�H;a�H;�H;��H;
�H;��H;G�H;M�H;�H;�H;��H;H�H;ǋH;      tiH;!jH;^lH;�oH;tH;1zH;��H;��H;�H;��H;5�H;��H;�H;гH;R�H;C�H;��H;s�H;��H;��H;��H;��H;)�H;,�H;��H;u�H;��H;e�H;[�H;��H;Z�H;��H;��H;5�H;e�H;o�H;b�H;o�H;e�H;5�H;��H;��H;Z�H;��H;[�H;e�H;��H;u�H;��H;,�H;)�H;��H;��H;��H;��H;s�H;��H;C�H;R�H;гH;�H;��H;5�H;��H;�H;��H;��H;1zH;tH;�oH;^lH;!jH;      5/H;�0H;Q5H;J<H;5EH;iOH;ZH;eH;�oH;�zH;��H;�H;�H;h�H;�H;�H;k�H;��H;��H;��H;��H;��H;�H;��H;��H;��H;J�H;��H;e�H;S�H;�H;j�H;��H;�H;E�H;[�H;M�H;[�H;E�H;�H;��H;j�H;�H;S�H;e�H;��H;J�H;��H;��H;��H;�H;��H;��H;��H;��H;��H;k�H;�H;�H;h�H;�H;�H;��H;�zH;�oH;eH;ZH;iOH;5EH;J<H;Q5H;�0H;      �G;�G;��G;��G;/�G;,�G;�H;)H;*?H;�RH;�cH;�rH;��H;��H;��H;\�H;
�H;��H;{�H;!�H;��H;��H;��H;X�H;O�H;��H;��H;J�H;��H;��H;j�H; �H;}�H;��H;�H;;�H;Y�H;;�H;�H;��H;}�H; �H;j�H;��H;��H;J�H;��H;��H;O�H;X�H;��H;��H;��H;!�H;{�H;��H;
�H;\�H;��H;��H;��H;�rH;�cH;�RH;*?H;)H;�H;,�G;/�G;��G;��G;�G;      @ZF;�cF;6�F;��F;�F;�!G;FaG;�G;��G;jH;)H;�FH;�]H;�pH;5�H;�H; �H;��H;��H;��H;
�H;e�H;��H;E�H;�H;6�H;��H;��H;u�H;��H;��H;��H;,�H;~�H;��H;�H;�H;�H;��H;~�H;,�H;��H;��H;��H;u�H;��H;��H;6�H;�H;E�H;��H;e�H;
�H;��H;��H;��H; �H;�H;5�H;�pH;�]H;�FH;)H;jH;��G;�G;FaG;�!G;�F;��F;6�F;�cF;      �VC; nC; �C;�D;}�D;V4E;)�E;�ZF;��F;�KG;,�G;��G;c H;^EH;E`H;>uH;#�H;��H;��H;b�H;<�H;��H;�H;I�H;�H;�H;O�H;��H;��H;��H;��H;��H;��H;=�H;��H;��H;��H;��H;��H;=�H;��H;��H;��H;��H;��H;��H;O�H;�H;�H;I�H;�H;��H;<�H;b�H;��H;��H;#�H;>uH;E`H;^EH;c H;��G;,�G;�KG;��F;�ZF;)�E;V4E;}�D;�D; �C; nC;      ��<;N�<;P\=;�N>;�?;��@;�6B;v�C;-�D;ͱE;F;�!G;�G;2�G;
)H;jOH;GjH;gH;X�H;Y�H;�H;�H;��H;H�H;I�H;E�H;X�H;��H;,�H;B�H;�H;�H;�H;��H;I�H;��H;��H;��H;I�H;��H;�H;�H;�H;B�H;,�H;��H;X�H;E�H;I�H;H�H;��H;�H;�H;Y�H;X�H;gH;GjH;jOH;
)H;2�G;�G;�!G;F;ͱE;-�D;v�C;�6B;��@;�?;�N>;P\=;N�<;      Y.;�.;�0;2;��4;�7;�{:;v\=;��?;�6B;�D;rnE;fwF;f4G;�G;
H;?H;aH;�yH;��H;.�H;ܫH;`�H;��H;�H;��H;��H;�H;)�H;��H;��H;h�H;c�H;O�H;��H;(�H;P�H;(�H;��H;O�H;c�H;h�H;��H;��H;)�H;�H;��H;��H;�H;��H;`�H;ܫH;.�H;��H;�yH;aH;?H;
H;�G;f4G;fwF;rnE;�D;�6B;��?;v\=;�{:;�7;��4;2;�0;�.;      ^;��;Nl;WZ;�_;%;+;8�0;G6;��:;��>;��A;�D;�E;`�F;QzG;u�G;1H;ZH;�uH;��H;g�H;ܫH;�H;��H;e�H;��H;��H;��H;��H;H�H;G�H;��H;��H;p�H;��H;��H;��H;p�H;��H;��H;G�H;H�H;��H;��H;��H;��H;e�H;��H;�H;ܫH;g�H;��H;�uH;ZH;1H;u�G;QzG;`�F;�E;�D;��A;��>;��:;G6;8�0;+;%;�_;WZ;Nl;��;      ��:C,�:$f�:���:�~�:^;��;��;��#;z�,;��4;R�:;�W?;.�B;��D;�ZF;FG;�G;}'H;VH;�tH;��H;.�H;�H;<�H;
�H;��H;��H;��H;��H;��H;��H;��H;��H;��H;^�H;b�H;^�H;��H;��H;��H;��H;��H;��H;��H;��H;��H;
�H;<�H;�H;.�H;��H;�tH;VH;}'H;�G;FG;�ZF;��D;.�B;�W?;R�:;��4;z�,;��#;��;��;^;�~�:���:$f�:C,�:      /�e9��9��9�:��Y:�x�:w:�:��:0^;8�;�"; r-;)G6;��<;2>A;0D;�F;f"G;�G;$H;VH;�uH;��H;Y�H;b�H;��H;!�H;��H;��H;E�H;��H;��H;��H;7�H;�H;��H;�H;��H;�H;7�H;��H;��H;��H;E�H;��H;��H;!�H;��H;b�H;Y�H;��H;�uH;VH;$H;�G;f"G;�F;0D;2>A;��<;)G6; r-;�";8�;0^;��:w:�:�x�:��Y:�:��9��9      �����뺶кf����Y�����k89z5:P.�:�c�:�A;�l;A?&;2;�{:;a @;��C;�E;�G;�G;}'H;ZH;�yH;X�H;��H;��H;{�H;��H;��H;l�H;��H;�H;[�H;<�H;W�H;
�H;��H;
�H;W�H;<�H;[�H;�H;��H;l�H;��H;��H;{�H;��H;��H;X�H;�yH;ZH;}'H;�G;�G;�E;��C;a @;�{:;2;A?&;�l;�A;�c�:P.�:z5:�k89����Y�f����к���      嚩�[���4J��
Y��S�b�(�-�1��VJx�#��%:��:@��:9�;� ;��.;0�8;��?;2�C;�E;f"G;�G;1H;aH;gH;��H;��H;��H;��H;s�H;(�H;I�H;J�H;��H;(�H;��H;H�H;��H;H�H;��H;(�H;��H;J�H;I�H;(�H;s�H;��H;��H;��H;��H;gH;aH;1H;�G;f"G;�E;2�C;��?;0�8;��.;� ;9�;@��:��:%:#��VJx�1��(�-�S�b�
Y��4J��[���      �B(��%�����_�|����˻	��-�b�x&�a ���@���Y:�:U^;B�;��,;Z_8;��?;��C;�F;FG;u�G;?H;GjH;#�H; �H;
�H;k�H;��H;�H;��H;/�H;��H;��H;��H;��H;��H;��H;��H;��H;��H;/�H;��H;�H;��H;k�H;
�H; �H;#�H;GjH;?H;u�G;FG;�F;��C;��?;Z_8;��,;B�;U^;�:��Y:�@�a ��x&�-�b�	���˻|����_�����%�      �����x���#��(F{���]��E<����J�뻱���ad\���]�02:��:���:�Z;��,;0�8;a @;0D;�ZF;QzG;
H;jOH;>uH;�H;\�H;�H;C�H;z�H;��H;��H;��H;��H;��H;��H;��H;��H;��H;��H;��H;��H;��H;z�H;C�H;�H;\�H;�H;>uH;jOH;
H;QzG;�ZF;0D;a @;0�8;��,;�Z;���:��:02:]���ad\�����J�뻛���E<���]�(F{��#���x��      >�Ｘ���o�Wrμ����bv��<"���]N�����?ݻe^��y��,�Y�f�9��:���:B�;��.;�{:;2>A;��D;`�F;�G;
)H;E`H;5�H;��H;�H;R�H;6�H;R�H;t�H;�H;/�H;k�H;��H;��H;��H;k�H;/�H;�H;t�H;R�H;6�H;R�H;�H;��H;5�H;E`H;
)H;�G;`�F;��D;2>A;�{:;��.;B�;���:��:f�9,�Y�y��e^���?ݻ����]N�<"��bv������Wrμ�o༸��      Gn;�`\8��s/�(�!�h��>���Prμ��������E<�������N3��Ix�f�9��:U^;� ;2;��<;.�B;�E;f4G;2�G;^EH;�pH;��H;h�H;гH;k�H;��H;��H;�H;��H;1�H;��H;�H;��H;1�H;��H;�H;��H;��H;k�H;гH;h�H;��H;�pH;^EH;2�G;f4G;�E;.�B;��<;2;� ;U^;��:f�9�Ix��N3�������E<��������Prμ>���h��(�!��s/�`\8�      ���������Ȅ�KSt���Y�Dn;�O�O#���Oļ�����&R��_������N3�,�Y�02:�:9�;A?&;)G6;�W?;�D;fwF;�G;c H;�]H;��H;�H;�H;a�H;$�H;�H;��H;(�H;��H;i�H;%�H;i�H;��H;(�H;��H;�H;$�H;a�H;�H;�H;��H;�]H;c H;�G;fwF;�D;�W?;)G6;A?&;9�;�:02:,�Y��N3������_��&R������OļO#��O�Dn;���Y�KSt��Ȅ�����      ��ѽ�[νa�ý�㳽&����L��r�d�Z\8�c���ټWv����Y��_����y��]���Y:@��:�l; r-;R�:;��A;rnE;�!G;��G;�FH;�rH;�H;��H;�H;J�H;5�H;��H;��H;��H;B�H;�H;B�H;��H;��H;��H;5�H;J�H;�H;��H;�H;�rH;�FH;��G;�!G;rnE;��A;R�:; r-;�l;@��:��Y:]�y������_���Y�Wv���ټc��Z\8�r�d��L��&����㳽a�ý�[ν      ��]�È�a}�q�_�ý�u�������K����o�Wv���&R���e^���뺪@���:�A;�";��4;��>;�D;F;,�G;)H;�cH;��H;5�H;��H;N�H;M�H;��H;��H;<�H;(�H;��H;(�H;<�H;��H;��H;M�H;N�H;��H;5�H;��H;�cH;)H;,�G;F;�D;��>;��4;�";�A;��:�@���e^�����&R�Wv���o����K������u��_�ýq�a}�È�]�      j+X��T��nH�ؕ6�� �Y��(��㳽����mR����ټ�����E<��?ݻad\�a ��%:�c�:8�;z�,;��:;�6B;ͱE;�KG;jH;�RH;�zH;��H;
�H;9�H;`�H;n�H;+�H;��H;�H;��H;�H;��H;+�H;n�H;`�H;9�H;
�H;��H;�zH;�RH;jH;�KG;ͱE;�6B;��:;z�,;8�;�c�:%:a ��ad\��?ݻ�E<������ټ���mR�����㳽(�Y��� �ؕ6��nH��T�      Ѱ������n���*|�4S\�� :����Z�U$������K�c���Oļ����������x&�#��P.�:0^;��#;G6;��?;-�D;��F;��G;*?H;�oH;�H;��H;:�H;r�H;J�H;��H;��H;��H;��H;��H;��H;��H;J�H;r�H;:�H;��H;�H;�oH;*?H;��G;��F;-�D;��?;G6;��#;0^;P.�:#��x&������������Oļc���K����U$���Z���� :�4S\��*|�n������      -�; 9ɾi㼾�A�������Mw��nH�����Z��㳽����Z\8�O#�������]N�J��-�b�VJx�z5:��:��;8�0;v\=;v�C;�ZF;�G;)H;eH;��H;G�H;g�H;��H;7�H;��H;P�H;��H;��H;��H;P�H;��H;7�H;��H;g�H;G�H;��H;eH;)H;�G;�ZF;v�C;v\=;8�0;��;��:z5:VJx�-�b�J���]N�����O#��Z\8������㳽�Z񽞯��nH��Mw������A��i㼾 9ɾ      #y��v�R���-�߾����0��1����nH���(Ὁu��r�d�O�Prμ<"�����	��1���k89w:�:��;+;�{:;�6B;)�E;FaG;�H;ZH;��H;M�H;ĮH;�H;e�H;e�H;+�H;��H;��H;��H;+�H;e�H;e�H;�H;ĮH;M�H;��H;ZH;�H;FaG;)�E;�6B;�{:;+;��;w:�:�k891��	�����<"��PrμO�r�d��u��(����nH�1���0������-�߾R����v�      �O/�aM+�I�����1W�� 9ɾ0���Mw�� :�Y��_�ý�L��Dn;�>���bv���E<��˻(�-�����x�:^;%;�7;��@;V4E;�!G;,�G;iOH;1zH;�H;��H;��H;��H;�H;2�H;�H;��H;�H;2�H;�H;��H;��H;��H;�H;1zH;iOH;,�G;�!G;V4E;��@;�7;%;^;�x�:���(�-��˻�E<�bv��>���Dn;��L��_�ýY��� :��Mw�0�� 9ɾ1W�����I��aM+�      $�X�EvS�%E��O/��S�1W����������4S\�� �q�&�����Y�h��������]�|���S�b��Y���Y:�~�:�_;��4;�?;}�D;�F;/�G;5EH;tH;�H;��H;��H;3�H;��H;E�H;8�H;�H;8�H;E�H;��H;3�H;��H;��H;�H;tH;5EH;/�G;�F;}�D;�?;��4;�_;�~�:��Y:�Y�S�b�|�����]�����h����Y�&���q�� �4S\���������1W���S��O/�%E�EvS�      � ����y�M�h�ބN��O/����-�߾�A���*|�ؕ6�a}��㳽KSt�(�!�Wrμ(F{��_�
Y��f����:���:WZ;2;�N>;�D;��F;��G;J<H;�oH;��H;t�H;��H;��H;��H;��H;��H;�H;��H;��H;��H;��H;��H;t�H;��H;�oH;J<H;��G;��F;�D;�N>;2;WZ;���:�:f���
Y���_�(F{�Wrμ(�!�KSt��㳽a}�ؕ6��*|��A��-�߾����O/�ބN�M�h���y�      2v��V���L ��M�h�%E�I��R���i㼾n���nH�È�a�ý�Ȅ��s/��o༼#�����4J���к��9$f�:Nl;�0;P\=; �C;6�F;��G;Q5H;^lH;H�H;ФH;��H;�H;b�H;��H;$�H;�H;$�H;��H;b�H;�H;��H;ФH;H�H;^lH;Q5H;��G;6�F; �C;P\=;�0;Nl;$f�:��9�к4J������#���o��s/��Ȅ�a�ýÈ��nH�n��i㼾R���I��%E�M�h�L ��V���      ph��"���V�����y�EvS�aM+��v� 9ɾ�����T�]��[ν����`\8�����x���%�[��������9C,�:��;�.;N�<; nC;�cF;�G;�0H;!jH;ǋH;ңH;��H;��H;��H;��H;��H;��H;��H;��H;��H;��H;��H;ңH;ǋH;!jH;�0H;�G;�cF; nC;N�<;�.;��;C,�:��9���[����%��x�����`\8������[ν]��T����� 9ɾ�v�aM+�EvS���y�V���"���      .Eb�I]�tN�ߛ7����e� �{�˾��	�j��!,�J���0��m���,˼��x�E���1��`���T�:g�:3;��1;o+>;��C;�vF;�G;��G;>H;�gH;Z�H;w�H;9�H;�H;��H;(�H;��H;(�H;��H;�H;9�H;w�H;Z�H;�gH;>H;��G;�G;�vF;��C;o+>;��1;3;g�:T�:`����1��E����x�,˼��m�0��J����!,�	�j���{�˾e� ����ߛ7�tN�I]�      I]�N�W��TI�v3��D�������Ǿb���ȟf� )� ��W;���Fi��k�x�Ǽ�[t�8�	�(Ȅ�rX��џ:���:&�;�I2;�Y>;qD;�~F;\�G;+H;�>H;�hH;�H;�H;r�H;7�H;��H;S�H;��H;S�H;��H;7�H;r�H;�H;�H;�hH;�>H;+H;\�G;�~F;qD;�Y>;�I2;&�;���:џ:rX��(Ȅ�8�	��[t�x�Ǽ�k��Fi�W;�� �� )�ȟf�b�����Ǿ�����D�v3��TI�N�W�      tN��TI���;��'��k���i���f󐾖Z��K ��s�&����&^����"����g����Шu�Q!���1<:��:n
;�f3;-�>;�AD;֕F;�G;�H;UAH;jH;\�H;��H;(�H;ԻH;k�H;��H;B�H;��H;k�H;ԻH;(�H;��H;\�H;jH;UAH;�H;�G;֕F;�AD;-�>;�f3;n
;��:�1<:Q!��Шu������g��"�����&^�&����s潎K ��Z�f�i������k��'���;��TI�      ߛ7�v3��'����e� ��{Ծ
���6���]�F�����ӽ���;�L�1v�x뮼,T�Ƙ��PV�n�=�4(i:a��:!z ;�#5;�?;2�D;�F;�G;�H;�EH;�mH;��H;~�H;j�H;ۼH;4�H;P�H;��H;P�H;4�H;ۼH;j�H;~�H;��H;�mH;�EH;�H;�G;�F;2�D;�?;�#5;!z ;a��:4(i:n�=��PV�Ƙ�,T�x뮼1v�;�L�����ӽ���]�F�6���
����{Ծe� �����'�v3�      ����D��k�e� �<�ݾS���C͓�ȟf��>/�x��~'��n섽/�6�Rt��v��?�:�Tʻ�.�ݷ��s�:2;�$;�X7;��@;	E;;�F;Q�G;�H;EKH;�qH;��H;ɣH;�H;�H;.�H;E�H;��H;E�H;.�H;�H;�H;ɣH;��H;�qH;EKH;�H;Q�G;;�F;	E;��@;�X7;�$;2;�s�:ݷ��.�Tʻ?�:��v��Rt�/�6�n섽~'��x���>/�ȟf�C͓�S���<�ݾe� ��k��D�      e� ������쾻{ԾS���b���9�x�rSC��^�ͻ޽%���Q�e����ѼG������R�����դ8��:�X;��);6�9;.�A;��E;�G;3�G;t H;DRH;�vH;w�H;��H;:�H;��H;r�H;v�H;��H;v�H;r�H;��H;:�H;��H;w�H;�vH;DRH;t H;3�G;�G;��E;.�A;6�9;��);�X;��:դ8����R�����G���Ѽ��Q�e�%���ͻ޽�^�rSC�9�x�b���S����{Ծ�쾃���      {�˾��Ǿi���
���C͓�9�x�ؘJ��K �H��� �������?���t뮼�[�����3|��W��>�:w~�:	';�
/;�f<;�C;� F;�MG;��G;:,H;sZH;�|H;ȖH;éH;��H;��H;��H;��H;��H;��H;��H;��H;��H;éH;ȖH;�|H;sZH;:,H;��G;�MG;� F;�C;�f<;�
/;	';w~�:>�:�W��3|������[�t뮼����?���� ��H����K �ؘJ�9�x�C͓�
���i�����Ǿ      ��b���f�6���ȟf�rSC��K �Gn����Ž����Z��k��|ռX��Ey-����w.�s���O�:�*�:��;p4;t�>;)D;�vF;I�G;��G;�8H;\cH;x�H;��H;\�H;e�H;��H;��H;K�H;g�H;K�H;��H;��H;e�H;\�H;��H;x�H;\cH;�8H;��G;I�G;�vF;)D;t�>;p4;��;�*�:�O�:s��w.����Ey-�X���|ռ�k��Z������ŽGn���K �rSC�ȟf�6���f�b���      	�j�ȟf��Z�]�F��>/��^�H�����Ž- ���Fi�kQ+�Ot�PT��H�W�����1��hȺ�U�9�O�:	Y;��(;T�8;2A;�E;"�F;|�G;�H;�EH;�lH;��H;��H;8�H;d�H;��H;��H;��H;��H;��H;��H;��H;d�H;8�H;��H;��H;�lH;�EH;�H;|�G;"�F;�E;2A;T�8;��(;	Y;�O�:�U�9hȺ�1�����H�W�PT��Ot�kQ+��Fi�- ����ŽH����^��>/�]�F��Z�ȟf�      �!,� )��K ����x��ͻ޽ ������Fi���0�����跼z�x�����.��b�(�����)i:���:��;�0;��<;�C;��E;)<G;
�G;�#H;kSH;�vH;�H;�H;E�H;u�H;4�H;��H;��H;n�H;��H;��H;4�H;u�H;E�H;�H;�H;�vH;kSH;�#H;
�G;)<G;��E;�C;��<;�0;��;���:�)i:���b�(��.�����z�x��跼�����0��Fi���� ��ͻ޽x������K � )�      J��� ��s��ӽ~'��%�������Z�kQ+�����"��G����0���׻̕b��W���V�9�:�_;�)';0Y7;H#@;T�D;�F;+�G;��G;A7H;aH;��H;Z�H;��H;l�H;��H;��H;{�H;B�H;.�H;B�H;{�H;��H;��H;l�H;��H;Z�H;��H;aH;A7H;��G;+�G;�F;T�D;H#@;0Y7;�)';�_;�:�V�9�W��̕b���׻��0�G���"�����kQ+��Z����%���~'���ӽ�s� ��      0��W;��&������n섽Q�e���?��k�Ot��跼G��ee7�����Ǆ��0��t�_t�: +�:�
;�1;��<;��B;N�E;G;�G;iH;wIH;`nH;��H;��H;�H;��H;��H;�H;��H;�H;��H;�H;��H;�H;��H;��H;�H;��H;��H;`nH;wIH;iH;�G;G;N�E;��B;��<;�1;�
; +�:_t�:�t��0��Ǆ����ee7�G���跼Ot�k���?�Q�e�n섽���&���W;��      m��Fi��&^�;�L�/�6������|ռPT��z�x���0��������0���ڷ�{m`:��:��;��*;~�8;G�@;e�D;��F;}G;��G;�0H;�ZH;n{H;��H;֧H;�H;��H;��H;|�H;��H;��H;e�H;��H;��H;|�H;��H;��H;�H;֧H;��H;n{H;�ZH;�0H;��G;}G;��F;e�D;G�@;~�8;��*;��;��:{m`:�ڷ�0��������껢�0�z�x�PT���|ռ����/�6�;�L��&^��Fi�      ���k���1v�Rt��Ѽt뮼X��H�W������׻�Ǆ�0�����3<:w��:;Y;�s%;=$5;�Y>;.`C;��E;O)G;v�G;#H;GH;lkH;�H;��H;��H;ȻH;��H;��H;��H;g�H;_�H;�H;_�H;g�H;��H;��H;��H;ȻH;��H;��H;�H;lkH;GH;#H;v�G;O)G;��E;.`C;�Y>;=$5;�s%;;Y;w��:�3<:���0���Ǆ���׻���H�W�X��t뮼�ѼRt�1v����k�      ,˼x�Ǽ�"��x뮼�v��G���[�Ey-�����.��̕b��0㺄ڷ��3<:L�:_\;��!;2J2;�f<;/B;RBE;J�F;a�G; �G;�3H;�[H;{H;��H;��H;P�H;��H;6�H;��H;B�H;A�H;��H;��H;��H;A�H;B�H;��H;6�H;��H;P�H;��H;��H;{H;�[H;�3H; �G;a�G;J�F;RBE;/B;�f<;2J2;��!;_\;L�:�3<:�ڷ��0�̕b��.�����Ey-��[�G���v��x뮼�"��x�Ǽ      ��x��[t���g�,T�?�:������������1��b�(��W���t�{m`:w��:_\;pz ;�0;�;;9<A;?�D;�vF;�bG;e�G;� H;�LH;�nH;p�H;~�H;��H;��H;Z�H;��H;H�H;_�H;��H;��H;�H;��H;��H;_�H;H�H;��H;Z�H;��H;��H;~�H;p�H;�nH;�LH;� H;e�G;�bG;�vF;?�D;9<A;�;;�0;pz ;_\;w��:{m`:�t��W��b�(��1������������?�:�,T���g��[t�      E��8�	����Ƙ�Tʻ�R��3|�w.�hȺ����V�9_t�:��:;Y;��!;�0;.�:;�@;5BD;�1F;�7G;��G;�H;k?H;+cH;�H;n�H;;�H;<�H;>�H;��H;��H;��H;[�H;��H;��H;s�H;��H;��H;[�H;��H;��H;��H;>�H;<�H;;�H;n�H;�H;+cH;k?H;�H;��G;�7G;�1F;5BD;�@;.�:;�0;��!;;Y;��:_t�:�V�9���hȺw.�3|��R��TʻƘ����8�	�      �1��(Ȅ�Шu��PV��.�����W��s��U�9�)i:�: +�:��;�s%;2J2;�;;�@;�D;/F;?G;��G;�H;�4H;�YH;5wH;7�H;�H;	�H;�H;I�H;^�H;�H;�H;�H;*�H;E�H;��H;E�H;*�H;�H;�H;�H;^�H;I�H;�H;	�H;�H;7�H;5wH;�YH;�4H;�H;��G;?G;/F;�D;�@;�;;2J2;�s%;��; +�:�:�)i:�U�9s���W������.��PV�Шu�(Ȅ�      `���rX��Q!��n�=�ݷ�դ8>�:�O�:�O�:���:�_;�
;��*;=$5;�f<;9<A;5BD;/F;�G;��G;r�G;�,H;RH;UpH;�H;��H;r�H;�H;)�H;��H;��H;��H;?�H;��H;��H;|�H;��H;|�H;��H;��H;?�H;��H;��H;��H;)�H;�H;r�H;��H;�H;UpH;RH;�,H;r�G;��G;�G;/F;5BD;9<A;�f<;=$5;��*;�
;�_;���:�O�:�O�:>�:դ8ݷ�n�=�Q!��rX��      T�:џ:�1<:4(i:�s�:��:w~�:�*�:	Y;��;�)';�1;~�8;�Y>;/B;?�D;�1F;?G;��G;%�G;�(H;�MH;qkH;D�H;c�H;v�H;��H;�H;t�H;��H;$�H;�H;�H;D�H;��H;��H;��H;��H;��H;D�H;�H;�H;$�H;��H;t�H;�H;��H;v�H;c�H;D�H;qkH;�MH;�(H;%�G;��G;?G;�1F;?�D;/B;�Y>;~�8;�1;�)';��;	Y;�*�:w~�:��:�s�:4(i:�1<:џ:      g�:���:��:a��:2;�X;	';��;��(;�0;0Y7;��<;G�@;.`C;RBE;�vF;�7G;��G;r�G;�(H;�KH;�hH;.�H;O�H;��H;��H;��H;O�H;�H;��H;��H;A�H;��H;��H;��H;��H;��H;��H;��H;��H;��H;A�H;��H;��H;�H;O�H;��H;��H;��H;O�H;.�H;�hH;�KH;�(H;r�G;��G;�7G;�vF;RBE;.`C;G�@;��<;0Y7;�0;��(;��;	';�X;2;a��:��:���:      3;&�;n
;!z ;�$;��);�
/;p4;T�8;��<;H#@;��B;e�D;��E;J�F;�bG;��G;�H;�,H;�MH;�hH;B�H;��H;��H;ΰH;��H;��H;��H;2�H;��H;^�H;�H;1�H;��H;��H;P�H;��H;P�H;��H;��H;1�H;�H;^�H;��H;2�H;��H;��H;��H;ΰH;��H;��H;B�H;�hH;�MH;�,H;�H;��G;�bG;J�F;��E;e�D;��B;H#@;��<;T�8;p4;�
/;��);�$;!z ;n
;&�;      ��1;�I2;�f3;�#5;�X7;6�9;�f<;t�>;2A;�C;T�D;N�E;��F;O)G;a�G;e�G;�H;�4H;RH;qkH;.�H;��H;�H;ɯH;��H;V�H;L�H; �H;��H;��H;u�H;��H;o�H;��H;��H;�H;\�H;�H;��H;��H;o�H;��H;u�H;��H;��H; �H;L�H;V�H;��H;ɯH;�H;��H;.�H;qkH;RH;�4H;�H;e�G;a�G;O)G;��F;N�E;T�D;�C;2A;t�>;�f<;6�9;�X7;�#5;�f3;�I2;      o+>;�Y>;-�>;�?;��@;.�A;�C;)D;�E;��E;�F;G;}G;v�G; �G;� H;k?H;�YH;UpH;D�H;O�H;��H;ɯH;�H;��H;��H;6�H;��H;��H;��H;O�H; �H;��H;��H;H�H;��H;��H;��H;H�H;��H;��H; �H;O�H;��H;��H;��H;6�H;��H;��H;�H;ɯH;��H;O�H;D�H;UpH;�YH;k?H;� H; �G;v�G;}G;G;�F;��E;�E;)D;�C;.�A;��@;�?;-�>;�Y>;      ��C;qD;�AD;2�D;	E;��E;� F;�vF;"�F;)<G;+�G;�G;��G;#H;�3H;�LH;+cH;5wH;�H;c�H;��H;ΰH;��H;��H;=�H;��H;��H;^�H;c�H;��H;��H;g�H;��H;@�H;��H;D�H;L�H;D�H;��H;@�H;��H;g�H;��H;��H;c�H;^�H;��H;��H;=�H;��H;��H;ΰH;��H;c�H;�H;5wH;+cH;�LH;�3H;#H;��G;�G;+�G;)<G;"�F;�vF;� F;��E;	E;2�D;�AD;qD;      �vF;�~F;֕F;�F;;�F;�G;�MG;I�G;|�G;
�G;��G;iH;�0H;GH;�[H;�nH;�H;7�H;��H;v�H;��H;��H;V�H;��H;��H;W�H;$�H;�H;��H;��H;�H;S�H;6�H;��H;m�H;��H;��H;��H;m�H;��H;6�H;S�H;�H;��H;��H;�H;$�H;W�H;��H;��H;V�H;��H;��H;v�H;��H;7�H;�H;�nH;�[H;GH;�0H;iH;��G;
�G;|�G;I�G;�MG;�G;;�F;�F;֕F;�~F;      �G;\�G;�G;�G;Q�G;3�G;��G;��G;�H;�#H;A7H;wIH;�ZH;lkH;{H;p�H;n�H;�H;r�H;��H;��H;��H;L�H;6�H;��H;$�H;�H;h�H;J�H;��H;7�H;�H;��H;��H;��H;�H;�H;�H;��H;��H;��H;�H;7�H;��H;J�H;h�H;�H;$�H;��H;6�H;L�H;��H;��H;��H;r�H;�H;n�H;p�H;{H;lkH;�ZH;wIH;A7H;�#H;�H;��G;��G;3�G;Q�G;�G;�G;\�G;      ��G;+H;�H;�H;�H;t H;:,H;�8H;�EH;kSH;aH;`nH;n{H;�H;��H;~�H;;�H;	�H;�H;�H;O�H;��H; �H;��H;^�H;�H;h�H;]�H;��H;�H;�H;��H;z�H;��H;�H;^�H;g�H;^�H;�H;��H;z�H;��H;�H;�H;��H;]�H;h�H;�H;^�H;��H; �H;��H;O�H;�H;�H;	�H;;�H;~�H;��H;�H;n{H;`nH;aH;kSH;�EH;�8H;:,H;t H;�H;�H;�H;+H;      >H;�>H;UAH;�EH;EKH;DRH;sZH;\cH;�lH;�vH;��H;��H;��H;��H;��H;��H;<�H;�H;)�H;t�H;�H;2�H;��H;��H;c�H;��H;J�H;��H;$�H;��H;��H;k�H;��H;6�H;p�H;��H;��H;��H;p�H;6�H;��H;k�H;��H;��H;$�H;��H;J�H;��H;c�H;��H;��H;2�H;�H;t�H;)�H;�H;<�H;��H;��H;��H;��H;��H;��H;�vH;�lH;\cH;sZH;DRH;EKH;�EH;UAH;�>H;      �gH;�hH;jH;�mH;�qH;�vH;�|H;x�H;��H;�H;Z�H;��H;֧H;��H;P�H;��H;>�H;I�H;��H;��H;��H;��H;��H;��H;��H;��H;��H;�H;��H;��H;t�H;��H;%�H;z�H;��H;��H;��H;��H;��H;z�H;%�H;��H;t�H;��H;��H;�H;��H;��H;��H;��H;��H;��H;��H;��H;��H;I�H;>�H;��H;P�H;��H;֧H;��H;Z�H;�H;��H;x�H;�|H;�vH;�qH;�mH;jH;�hH;      Z�H;�H;\�H;��H;��H;w�H;ȖH;��H;��H;�H;��H;�H;�H;ȻH;��H;Z�H;��H;^�H;��H;$�H;��H;^�H;u�H;O�H;��H;�H;7�H;�H;��H;t�H;��H;.�H;��H;��H;��H;��H;��H;��H;��H;��H;��H;.�H;��H;t�H;��H;�H;7�H;�H;��H;O�H;u�H;^�H;��H;$�H;��H;^�H;��H;Z�H;��H;ȻH;�H;�H;��H;�H;��H;��H;ȖH;w�H;��H;��H;\�H;�H;      w�H;�H;��H;~�H;ɣH;��H;éH;\�H;8�H;E�H;l�H;��H;��H;��H;6�H;��H;��H;�H;��H;�H;A�H;�H;��H; �H;g�H;S�H;�H;��H;k�H;��H;.�H;{�H;��H;��H;��H;�H;�H;�H;��H;��H;��H;{�H;.�H;��H;k�H;��H;�H;S�H;g�H; �H;��H;�H;A�H;�H;��H;�H;��H;��H;6�H;��H;��H;��H;l�H;E�H;8�H;\�H;éH;��H;ɣH;~�H;��H;�H;      9�H;r�H;(�H;j�H;�H;:�H;��H;e�H;d�H;u�H;��H;��H;��H;��H;��H;H�H;��H;�H;?�H;�H;��H;1�H;o�H;��H;��H;6�H;��H;z�H;��H;%�H;��H;��H;��H;��H;�H;�H;�H;�H;�H;��H;��H;��H;��H;%�H;��H;z�H;��H;6�H;��H;��H;o�H;1�H;��H;�H;?�H;�H;��H;H�H;��H;��H;��H;��H;��H;u�H;d�H;e�H;��H;:�H;�H;j�H;(�H;r�H;      �H;7�H;ԻH;ۼH;�H;��H;��H;��H;��H;4�H;��H;�H;|�H;��H;B�H;_�H;[�H;�H;��H;D�H;��H;��H;��H;��H;@�H;��H;��H;��H;6�H;z�H;��H;��H;��H; �H;.�H;9�H;�H;9�H;.�H; �H;��H;��H;��H;z�H;6�H;��H;��H;��H;@�H;��H;��H;��H;��H;D�H;��H;�H;[�H;_�H;B�H;��H;|�H;�H;��H;4�H;��H;��H;��H;��H;�H;ۼH;ԻH;7�H;      ��H;��H;k�H;4�H;.�H;r�H;��H;��H;��H;��H;{�H;��H;��H;g�H;A�H;��H;��H;*�H;��H;��H;��H;��H;��H;H�H;��H;m�H;��H;�H;p�H;��H;��H;��H;�H;.�H;�H;.�H;J�H;.�H;�H;.�H;�H;��H;��H;��H;p�H;�H;��H;m�H;��H;H�H;��H;��H;��H;��H;��H;*�H;��H;��H;A�H;g�H;��H;��H;{�H;��H;��H;��H;��H;r�H;.�H;4�H;k�H;��H;      (�H;S�H;��H;P�H;E�H;v�H;��H;K�H;��H;��H;B�H;�H;��H;_�H;��H;��H;��H;E�H;|�H;��H;��H;P�H;�H;��H;D�H;��H;�H;^�H;��H;��H;��H;�H;�H;9�H;.�H;$�H;6�H;$�H;.�H;9�H;�H;�H;��H;��H;��H;^�H;�H;��H;D�H;��H;�H;P�H;��H;��H;|�H;E�H;��H;��H;��H;_�H;��H;�H;B�H;��H;��H;K�H;��H;v�H;E�H;P�H;��H;S�H;      ��H;��H;B�H;��H;��H;��H;��H;g�H;��H;n�H;.�H;��H;e�H;�H;��H;�H;s�H;��H;��H;��H;��H;��H;\�H;��H;L�H;��H;�H;g�H;��H;��H;��H;�H;�H;�H;J�H;6�H;#�H;6�H;J�H;�H;�H;�H;��H;��H;��H;g�H;�H;��H;L�H;��H;\�H;��H;��H;��H;��H;��H;s�H;�H;��H;�H;e�H;��H;.�H;n�H;��H;g�H;��H;��H;��H;��H;B�H;��H;      (�H;S�H;��H;P�H;E�H;v�H;��H;K�H;��H;��H;B�H;�H;��H;_�H;��H;��H;��H;E�H;|�H;��H;��H;P�H;�H;��H;D�H;��H;�H;^�H;��H;��H;��H;�H;�H;9�H;.�H;$�H;6�H;$�H;.�H;9�H;�H;�H;��H;��H;��H;^�H;�H;��H;D�H;��H;�H;P�H;��H;��H;|�H;E�H;��H;��H;��H;_�H;��H;�H;B�H;��H;��H;K�H;��H;v�H;E�H;P�H;��H;S�H;      ��H;��H;k�H;4�H;.�H;r�H;��H;��H;��H;��H;{�H;��H;��H;g�H;A�H;��H;��H;*�H;��H;��H;��H;��H;��H;H�H;��H;m�H;��H;�H;p�H;��H;��H;��H;�H;.�H;�H;.�H;J�H;.�H;�H;.�H;�H;��H;��H;��H;p�H;�H;��H;m�H;��H;H�H;��H;��H;��H;��H;��H;*�H;��H;��H;A�H;g�H;��H;��H;{�H;��H;��H;��H;��H;r�H;.�H;4�H;k�H;��H;      �H;7�H;ԻH;ۼH;�H;��H;��H;��H;��H;4�H;��H;�H;|�H;��H;B�H;_�H;[�H;�H;��H;D�H;��H;��H;��H;��H;@�H;��H;��H;��H;6�H;z�H;��H;��H;��H; �H;.�H;9�H;�H;9�H;.�H; �H;��H;��H;��H;z�H;6�H;��H;��H;��H;@�H;��H;��H;��H;��H;D�H;��H;�H;[�H;_�H;B�H;��H;|�H;�H;��H;4�H;��H;��H;��H;��H;�H;ۼH;ԻH;7�H;      9�H;r�H;(�H;j�H;�H;:�H;��H;e�H;d�H;u�H;��H;��H;��H;��H;��H;H�H;��H;�H;?�H;�H;��H;1�H;o�H;��H;��H;6�H;��H;z�H;��H;%�H;��H;��H;��H;��H;�H;�H;�H;�H;�H;��H;��H;��H;��H;%�H;��H;z�H;��H;6�H;��H;��H;o�H;1�H;��H;�H;?�H;�H;��H;H�H;��H;��H;��H;��H;��H;u�H;d�H;e�H;��H;:�H;�H;j�H;(�H;r�H;      w�H;�H;��H;~�H;ɣH;��H;éH;\�H;8�H;E�H;l�H;��H;��H;��H;6�H;��H;��H;�H;��H;�H;A�H;�H;��H; �H;g�H;S�H;�H;��H;k�H;��H;.�H;{�H;��H;��H;��H;�H;�H;�H;��H;��H;��H;{�H;.�H;��H;k�H;��H;�H;S�H;g�H; �H;��H;�H;A�H;�H;��H;�H;��H;��H;6�H;��H;��H;��H;l�H;E�H;8�H;\�H;éH;��H;ɣH;~�H;��H;�H;      Z�H;�H;\�H;��H;��H;w�H;ȖH;��H;��H;�H;��H;�H;�H;ȻH;��H;Z�H;��H;^�H;��H;$�H;��H;^�H;u�H;O�H;��H;�H;7�H;�H;��H;t�H;��H;.�H;��H;��H;��H;��H;��H;��H;��H;��H;��H;.�H;��H;t�H;��H;�H;7�H;�H;��H;O�H;u�H;^�H;��H;$�H;��H;^�H;��H;Z�H;��H;ȻH;�H;�H;��H;�H;��H;��H;ȖH;w�H;��H;��H;\�H;�H;      �gH;�hH;jH;�mH;�qH;�vH;�|H;x�H;��H;�H;Z�H;��H;֧H;��H;P�H;��H;>�H;I�H;��H;��H;��H;��H;��H;��H;��H;��H;��H;�H;��H;��H;t�H;��H;%�H;z�H;��H;��H;��H;��H;��H;z�H;%�H;��H;t�H;��H;��H;�H;��H;��H;��H;��H;��H;��H;��H;��H;��H;I�H;>�H;��H;P�H;��H;֧H;��H;Z�H;�H;��H;x�H;�|H;�vH;�qH;�mH;jH;�hH;      >H;�>H;UAH;�EH;EKH;DRH;sZH;\cH;�lH;�vH;��H;��H;��H;��H;��H;��H;<�H;�H;)�H;t�H;�H;2�H;��H;��H;c�H;��H;J�H;��H;$�H;��H;��H;k�H;��H;6�H;p�H;��H;��H;��H;p�H;6�H;��H;k�H;��H;��H;$�H;��H;J�H;��H;c�H;��H;��H;2�H;�H;t�H;)�H;�H;<�H;��H;��H;��H;��H;��H;��H;�vH;�lH;\cH;sZH;DRH;EKH;�EH;UAH;�>H;      ��G;+H;�H;�H;�H;t H;:,H;�8H;�EH;kSH;aH;`nH;n{H;�H;��H;~�H;;�H;	�H;�H;�H;O�H;��H; �H;��H;^�H;�H;h�H;]�H;��H;�H;�H;��H;z�H;��H;�H;^�H;g�H;^�H;�H;��H;z�H;��H;�H;�H;��H;]�H;h�H;�H;^�H;��H; �H;��H;O�H;�H;�H;	�H;;�H;~�H;��H;�H;n{H;`nH;aH;kSH;�EH;�8H;:,H;t H;�H;�H;�H;+H;      �G;\�G;�G;�G;Q�G;3�G;��G;��G;�H;�#H;A7H;wIH;�ZH;lkH;{H;p�H;n�H;�H;r�H;��H;��H;��H;L�H;6�H;��H;$�H;�H;h�H;J�H;��H;7�H;�H;��H;��H;��H;�H;�H;�H;��H;��H;��H;�H;7�H;��H;J�H;h�H;�H;$�H;��H;6�H;L�H;��H;��H;��H;r�H;�H;n�H;p�H;{H;lkH;�ZH;wIH;A7H;�#H;�H;��G;��G;3�G;Q�G;�G;�G;\�G;      �vF;�~F;֕F;�F;;�F;�G;�MG;I�G;|�G;
�G;��G;iH;�0H;GH;�[H;�nH;�H;7�H;��H;v�H;��H;��H;V�H;��H;��H;W�H;$�H;�H;��H;��H;�H;S�H;6�H;��H;m�H;��H;��H;��H;m�H;��H;6�H;S�H;�H;��H;��H;�H;$�H;W�H;��H;��H;V�H;��H;��H;v�H;��H;7�H;�H;�nH;�[H;GH;�0H;iH;��G;
�G;|�G;I�G;�MG;�G;;�F;�F;֕F;�~F;      ��C;qD;�AD;2�D;	E;��E;� F;�vF;"�F;)<G;+�G;�G;��G;#H;�3H;�LH;+cH;5wH;�H;c�H;��H;ΰH;��H;��H;=�H;��H;��H;^�H;c�H;��H;��H;g�H;��H;@�H;��H;D�H;L�H;D�H;��H;@�H;��H;g�H;��H;��H;c�H;^�H;��H;��H;=�H;��H;��H;ΰH;��H;c�H;�H;5wH;+cH;�LH;�3H;#H;��G;�G;+�G;)<G;"�F;�vF;� F;��E;	E;2�D;�AD;qD;      o+>;�Y>;-�>;�?;��@;.�A;�C;)D;�E;��E;�F;G;}G;v�G; �G;� H;k?H;�YH;UpH;D�H;O�H;��H;ɯH;�H;��H;��H;6�H;��H;��H;��H;O�H; �H;��H;��H;H�H;��H;��H;��H;H�H;��H;��H; �H;O�H;��H;��H;��H;6�H;��H;��H;�H;ɯH;��H;O�H;D�H;UpH;�YH;k?H;� H; �G;v�G;}G;G;�F;��E;�E;)D;�C;.�A;��@;�?;-�>;�Y>;      ��1;�I2;�f3;�#5;�X7;6�9;�f<;t�>;2A;�C;T�D;N�E;��F;O)G;a�G;e�G;�H;�4H;RH;qkH;.�H;��H;�H;ɯH;��H;V�H;L�H; �H;��H;��H;u�H;��H;o�H;��H;��H;�H;\�H;�H;��H;��H;o�H;��H;u�H;��H;��H; �H;L�H;V�H;��H;ɯH;�H;��H;.�H;qkH;RH;�4H;�H;e�G;a�G;O)G;��F;N�E;T�D;�C;2A;t�>;�f<;6�9;�X7;�#5;�f3;�I2;      3;&�;n
;!z ;�$;��);�
/;p4;T�8;��<;H#@;��B;e�D;��E;J�F;�bG;��G;�H;�,H;�MH;�hH;B�H;��H;��H;ΰH;��H;��H;��H;2�H;��H;^�H;�H;1�H;��H;��H;P�H;��H;P�H;��H;��H;1�H;�H;^�H;��H;2�H;��H;��H;��H;ΰH;��H;��H;B�H;�hH;�MH;�,H;�H;��G;�bG;J�F;��E;e�D;��B;H#@;��<;T�8;p4;�
/;��);�$;!z ;n
;&�;      g�:���:��:a��:2;�X;	';��;��(;�0;0Y7;��<;G�@;.`C;RBE;�vF;�7G;��G;r�G;�(H;�KH;�hH;.�H;O�H;��H;��H;��H;O�H;�H;��H;��H;A�H;��H;��H;��H;��H;��H;��H;��H;��H;��H;A�H;��H;��H;�H;O�H;��H;��H;��H;O�H;.�H;�hH;�KH;�(H;r�G;��G;�7G;�vF;RBE;.`C;G�@;��<;0Y7;�0;��(;��;	';�X;2;a��:��:���:      T�:џ:�1<:4(i:�s�:��:w~�:�*�:	Y;��;�)';�1;~�8;�Y>;/B;?�D;�1F;?G;��G;%�G;�(H;�MH;qkH;D�H;c�H;v�H;��H;�H;t�H;��H;$�H;�H;�H;D�H;��H;��H;��H;��H;��H;D�H;�H;�H;$�H;��H;t�H;�H;��H;v�H;c�H;D�H;qkH;�MH;�(H;%�G;��G;?G;�1F;?�D;/B;�Y>;~�8;�1;�)';��;	Y;�*�:w~�:��:�s�:4(i:�1<:џ:      `���rX��Q!��n�=�ݷ�դ8>�:�O�:�O�:���:�_;�
;��*;=$5;�f<;9<A;5BD;/F;�G;��G;r�G;�,H;RH;UpH;�H;��H;r�H;�H;)�H;��H;��H;��H;?�H;��H;��H;|�H;��H;|�H;��H;��H;?�H;��H;��H;��H;)�H;�H;r�H;��H;�H;UpH;RH;�,H;r�G;��G;�G;/F;5BD;9<A;�f<;=$5;��*;�
;�_;���:�O�:�O�:>�:դ8ݷ�n�=�Q!��rX��      �1��(Ȅ�Шu��PV��.�����W��s��U�9�)i:�: +�:��;�s%;2J2;�;;�@;�D;/F;?G;��G;�H;�4H;�YH;5wH;7�H;�H;	�H;�H;I�H;^�H;�H;�H;�H;*�H;E�H;��H;E�H;*�H;�H;�H;�H;^�H;I�H;�H;	�H;�H;7�H;5wH;�YH;�4H;�H;��G;?G;/F;�D;�@;�;;2J2;�s%;��; +�:�:�)i:�U�9s���W������.��PV�Шu�(Ȅ�      E��8�	����Ƙ�Tʻ�R��3|�w.�hȺ����V�9_t�:��:;Y;��!;�0;.�:;�@;5BD;�1F;�7G;��G;�H;k?H;+cH;�H;n�H;;�H;<�H;>�H;��H;��H;��H;[�H;��H;��H;s�H;��H;��H;[�H;��H;��H;��H;>�H;<�H;;�H;n�H;�H;+cH;k?H;�H;��G;�7G;�1F;5BD;�@;.�:;�0;��!;;Y;��:_t�:�V�9���hȺw.�3|��R��TʻƘ����8�	�      ��x��[t���g�,T�?�:������������1��b�(��W���t�{m`:w��:_\;pz ;�0;�;;9<A;?�D;�vF;�bG;e�G;� H;�LH;�nH;p�H;~�H;��H;��H;Z�H;��H;H�H;_�H;��H;��H;�H;��H;��H;_�H;H�H;��H;Z�H;��H;��H;~�H;p�H;�nH;�LH;� H;e�G;�bG;�vF;?�D;9<A;�;;�0;pz ;_\;w��:{m`:�t��W��b�(��1������������?�:�,T���g��[t�      ,˼x�Ǽ�"��x뮼�v��G���[�Ey-�����.��̕b��0㺄ڷ��3<:L�:_\;��!;2J2;�f<;/B;RBE;J�F;a�G; �G;�3H;�[H;{H;��H;��H;P�H;��H;6�H;��H;B�H;A�H;��H;��H;��H;A�H;B�H;��H;6�H;��H;P�H;��H;��H;{H;�[H;�3H; �G;a�G;J�F;RBE;/B;�f<;2J2;��!;_\;L�:�3<:�ڷ��0�̕b��.�����Ey-��[�G���v��x뮼�"��x�Ǽ      ���k���1v�Rt��Ѽt뮼X��H�W������׻�Ǆ�0�����3<:w��:;Y;�s%;=$5;�Y>;.`C;��E;O)G;v�G;#H;GH;lkH;�H;��H;��H;ȻH;��H;��H;��H;g�H;_�H;�H;_�H;g�H;��H;��H;��H;ȻH;��H;��H;�H;lkH;GH;#H;v�G;O)G;��E;.`C;�Y>;=$5;�s%;;Y;w��:�3<:���0���Ǆ���׻���H�W�X��t뮼�ѼRt�1v����k�      m��Fi��&^�;�L�/�6������|ռPT��z�x���0��������0���ڷ�{m`:��:��;��*;~�8;G�@;e�D;��F;}G;��G;�0H;�ZH;n{H;��H;֧H;�H;��H;��H;|�H;��H;��H;e�H;��H;��H;|�H;��H;��H;�H;֧H;��H;n{H;�ZH;�0H;��G;}G;��F;e�D;G�@;~�8;��*;��;��:{m`:�ڷ�0��������껢�0�z�x�PT���|ռ����/�6�;�L��&^��Fi�      0��W;��&������n섽Q�e���?��k�Ot��跼G��ee7�����Ǆ��0��t�_t�: +�:�
;�1;��<;��B;N�E;G;�G;iH;wIH;`nH;��H;��H;�H;��H;��H;�H;��H;�H;��H;�H;��H;�H;��H;��H;�H;��H;��H;`nH;wIH;iH;�G;G;N�E;��B;��<;�1;�
; +�:_t�:�t��0��Ǆ����ee7�G���跼Ot�k���?�Q�e�n섽���&���W;��      J��� ��s��ӽ~'��%�������Z�kQ+�����"��G����0���׻̕b��W���V�9�:�_;�)';0Y7;H#@;T�D;�F;+�G;��G;A7H;aH;��H;Z�H;��H;l�H;��H;��H;{�H;B�H;.�H;B�H;{�H;��H;��H;l�H;��H;Z�H;��H;aH;A7H;��G;+�G;�F;T�D;H#@;0Y7;�)';�_;�:�V�9�W��̕b���׻��0�G���"�����kQ+��Z����%���~'���ӽ�s� ��      �!,� )��K ����x��ͻ޽ ������Fi���0�����跼z�x�����.��b�(�����)i:���:��;�0;��<;�C;��E;)<G;
�G;�#H;kSH;�vH;�H;�H;E�H;u�H;4�H;��H;��H;n�H;��H;��H;4�H;u�H;E�H;�H;�H;�vH;kSH;�#H;
�G;)<G;��E;�C;��<;�0;��;���:�)i:���b�(��.�����z�x��跼�����0��Fi���� ��ͻ޽x������K � )�      	�j�ȟf��Z�]�F��>/��^�H�����Ž- ���Fi�kQ+�Ot�PT��H�W�����1��hȺ�U�9�O�:	Y;��(;T�8;2A;�E;"�F;|�G;�H;�EH;�lH;��H;��H;8�H;d�H;��H;��H;��H;��H;��H;��H;��H;d�H;8�H;��H;��H;�lH;�EH;�H;|�G;"�F;�E;2A;T�8;��(;	Y;�O�:�U�9hȺ�1�����H�W�PT��Ot�kQ+��Fi�- ����ŽH����^��>/�]�F��Z�ȟf�      ��b���f�6���ȟf�rSC��K �Gn����Ž����Z��k��|ռX��Ey-����w.�s���O�:�*�:��;p4;t�>;)D;�vF;I�G;��G;�8H;\cH;x�H;��H;\�H;e�H;��H;��H;K�H;g�H;K�H;��H;��H;e�H;\�H;��H;x�H;\cH;�8H;��G;I�G;�vF;)D;t�>;p4;��;�*�:�O�:s��w.����Ey-�X���|ռ�k��Z������ŽGn���K �rSC�ȟf�6���f�b���      {�˾��Ǿi���
���C͓�9�x�ؘJ��K �H��� �������?���t뮼�[�����3|��W��>�:w~�:	';�
/;�f<;�C;� F;�MG;��G;:,H;sZH;�|H;ȖH;éH;��H;��H;��H;��H;��H;��H;��H;��H;��H;éH;ȖH;�|H;sZH;:,H;��G;�MG;� F;�C;�f<;�
/;	';w~�:>�:�W��3|������[�t뮼����?���� ��H����K �ؘJ�9�x�C͓�
���i�����Ǿ      e� ������쾻{ԾS���b���9�x�rSC��^�ͻ޽%���Q�e����ѼG������R�����դ8��:�X;��);6�9;.�A;��E;�G;3�G;t H;DRH;�vH;w�H;��H;:�H;��H;r�H;v�H;��H;v�H;r�H;��H;:�H;��H;w�H;�vH;DRH;t H;3�G;�G;��E;.�A;6�9;��);�X;��:դ8����R�����G���Ѽ��Q�e�%���ͻ޽�^�rSC�9�x�b���S����{Ծ�쾃���      ����D��k�e� �<�ݾS���C͓�ȟf��>/�x��~'��n섽/�6�Rt��v��?�:�Tʻ�.�ݷ��s�:2;�$;�X7;��@;	E;;�F;Q�G;�H;EKH;�qH;��H;ɣH;�H;�H;.�H;E�H;��H;E�H;.�H;�H;�H;ɣH;��H;�qH;EKH;�H;Q�G;;�F;	E;��@;�X7;�$;2;�s�:ݷ��.�Tʻ?�:��v��Rt�/�6�n섽~'��x���>/�ȟf�C͓�S���<�ݾe� ��k��D�      ߛ7�v3��'����e� ��{Ծ
���6���]�F�����ӽ���;�L�1v�x뮼,T�Ƙ��PV�n�=�4(i:a��:!z ;�#5;�?;2�D;�F;�G;�H;�EH;�mH;��H;~�H;j�H;ۼH;4�H;P�H;��H;P�H;4�H;ۼH;j�H;~�H;��H;�mH;�EH;�H;�G;�F;2�D;�?;�#5;!z ;a��:4(i:n�=��PV�Ƙ�,T�x뮼1v�;�L�����ӽ���]�F�6���
����{Ծe� �����'�v3�      tN��TI���;��'��k���i���f󐾖Z��K ��s�&����&^����"����g����Шu�Q!���1<:��:n
;�f3;-�>;�AD;֕F;�G;�H;UAH;jH;\�H;��H;(�H;ԻH;k�H;��H;B�H;��H;k�H;ԻH;(�H;��H;\�H;jH;UAH;�H;�G;֕F;�AD;-�>;�f3;n
;��:�1<:Q!��Шu������g��"�����&^�&����s潎K ��Z�f�i������k��'���;��TI�      I]�N�W��TI�v3��D�������Ǿb���ȟf� )� ��W;���Fi��k�x�Ǽ�[t�8�	�(Ȅ�rX��џ:���:&�;�I2;�Y>;qD;�~F;\�G;+H;�>H;�hH;�H;�H;r�H;7�H;��H;S�H;��H;S�H;��H;7�H;r�H;�H;�H;�hH;�>H;+H;\�G;�~F;qD;�Y>;�I2;&�;���:џ:rX��(Ȅ�8�	��[t�x�Ǽ�k��Fi�W;�� �� )�ȟf�b�����Ǿ�����D�v3��TI�N�W�      �$��� ���������þ�*��
Dx�}�=����\Pν鰒��&K�xc����;�V�s���D^���S��v[:���:�d;��4;�_?;�lD;��F;puG;M�G;�H;�NH;�rH;�H;��H;��H;�H;q�H;E�H;q�H;�H;��H;��H;�H;�rH;�NH;�H;M�G;puG;��F;�lD;�_?;��4;�d;���:�v[:��S��D^�s��;�V����xc��&K�鰒�\Pν���}�=�
Dx��*���þ��������� �      �� �k��>��=���������0���s���:�N9���ʽZ����G��8��-��z5S�v���/X���D��Ad:�A�:� ;y�4;	�?;#~D;q�F;4xG;��G;�H;NOH;IsH;:�H;�H;�H;W�H;��H;U�H;��H;W�H;�H;�H;:�H;IsH;NOH;�H;��G;4xG;q�F;#~D;	�?;y�4;� ;�A�:�Ad:��D��/X�v��z5S��-���8���G�Z����ʽN9���:��s��0��������=��>��k��      ���>��&�
�����fYؾ���ȥ����f���0�C[�*8������ȟ>�|���#Ȥ�Y6H�,�ܻ�qF�-��7�}:���:�";��5;7�?;��D;��F;/�G;��G;s"H;�QH;�tH;z�H;�H;��H;�H;�H;��H;�H;�H;��H;�H;z�H;�tH;�QH;s"H;��G;/�G;��F;��D;7�?;��5;�";���:7�}:-���qF�,�ܻY6H�#Ȥ�|���ȟ>�����*8��C[���0���f�ȥ�����fYؾ����&�
�>��      ��=������I��þ�R��&���QS��Q"��s�����}��0���d���x�6��ƻ'}*����_�:�w;�%;Rl7;�@;�D;�F;��G;��G;3'H;UH;�wH;��H;f�H;ñH;ܺH;�H;��H;�H;ܺH;ñH;f�H;��H;�wH;UH;3'H;��G;��G;�F;�D;�@;Rl7;�%;�w;_�:���'}*��ƻx�6�d����켟0���}�����s��Q"�QS�&����R���þIᾁ���=��      ����fYؾ�þ�ê�f쏾jk���:�e�R�ؽ�����c�:y���Ҽݫ��� �B�'����'7��:�
;d�(;�^9;��A;�[E;��F;�G;��G;�-H;�YH;{H;�H;i�H;u�H;6�H;�H;��H;�H;6�H;u�H;i�H;�H;{H;�YH;�-H;��G;�G;��F;�[E;��A;�^9;d�(;�
;��:��'7'��B�� �ݫ����Ҽ:y��c�����R�ؽe���:�jk�f쏾�ê��þfYؾ��      �þ��������R��f쏾�s��H����������������D�vc�g����f�3,�����P����90��:6;�i-;��;;��B;,�E;�G;��G;��G;�5H;�_H;�H;{�H;��H;r�H;ɽH;r�H;��H;r�H;ɽH;r�H;��H;{�H;�H;�_H;�5H;��G;��G;�G;,�E;��B;��;;�i-;6;0��:��9�P�����3,��f�g���vc���D���������������H��s�f쏾�R���������      �*���0��ȥ��&���jk��H��#%�B[�ZPν�s��0�f�/%�d��`���G�=�n?ػfFL��D�d�R:D�:��;�2;�=;��C;�/F;�FG;�G;WH;?H;�fH;��H;V�H;ͫH;��H;��H;�H;��H;�H;��H;��H;ͫH;V�H;��H;�fH;?H;WH;�G;�FG;�/F;��C;�=;�2;��;D�:d�R:�D�fFL�n?ػG�=�`���d��/%�0�f��s��ZPνB[��#%��H�jk�&���ȥ���0��      
Dx��s���f�QS���:����B[��7ս�榽��}�u�;��8�)�����r����G������Ҭ����:��;}$;,�6;f�?;3�D;�F; pG;��G;H;XIH;dnH;i�H;��H;�H;[�H;��H;��H;G�H;��H;��H;[�H;�H;��H;i�H;dnH;XIH;H;��G; pG;�F;3�D;f�?;,�6;}$;��;���:�Ҭ����G�������r�)����8�u�;���}��榽�7սB[������:�QS���f��s�      }�=���:���0��Q"�e�����ZPν�榽%����G�����Ҽ���E:�	�ܻ�D^�͸��lh:���:P;�{,;�:;��A;~hE;��F;]�G;��G;�'H;eTH;�vH;��H;L�H;��H;�H;��H;��H;4�H;��H;��H;�H;��H;L�H;��H;�vH;eTH;�'H;��G;]�G;��F;~hE;��A;�:;�{,;P;���:lh:͸���D^�	�ܻE:������Ҽ����G�%���榽ZPν����e��Q"���0���:�      ���N9�C[��s�R�ؽ���s����}���G��K��	c��!�V�$,��*���������:@��:� ;ǂ3;0>;�C;#F;$8G;l�G;�H;7H;�_H;,H;�H; �H;g�H;�H;m�H;��H;3�H;��H;m�H;�H;g�H; �H;�H;,H;�_H;7H;�H;l�G;$8G;#F;�C;0>;ǂ3;� ;@��:��:������*��$,�!�V�	c��K�����G���}��s����R�ؽ�s�C[�N9�      \Pν��ʽ*8�������������0�f�u�;���K��Ȥ���f���#ߵ�>o5�1�D�O�-:���:Y>;H+;_9;�A;��D;\�F;�uG;�G;IH;�FH;�kH;�H;��H;�H;H�H;�H;��H;"�H;F�H;"�H;��H;�H;H�H;�H;��H;�H;�kH;�FH;IH;�G;�uG;\�F;��D;�A;_9;H+;Y>;���:O�-:1�D�>o5�#ߵ�����f�Ȥ�K����u�;�0�f������������*8����ʽ      鰒�Z��������}��c���D�/%��8���Ҽ	c����f�����ƻY/X�s������9h�:ȏ;G";�3;�>;�XC;��E;G;'�G;��G;�+H;/VH;9wH;��H;W�H;�H;.�H;�H;Q�H;a�H;O�H;a�H;Q�H;�H;.�H;�H;W�H;��H;9wH;/VH;�+H;��G;'�G;G;��E;�XC;�>;�3;G";ȏ;h�:���9s���Y/X��ƻ�����f�	c����Ҽ�8�/%���D��c���}�����Z��      �&K���G�ȟ>��0�:y�vc�d��)������!�V����ƻfod���ºQ(7�3�:���: �;^P.;:�:;ayA;y�D;�F;�mG;u�G;"H;�?H;MeH;��H;R�H;ժH;��H;�H;
�H;��H;��H;W�H;��H;��H;
�H;�H;��H;ժH;R�H;��H;MeH;�?H;"H;u�G;�mG;�F;y�D;ayA;:�:;^P.; �;���:�3�:Q(7��ºfod��ƻ��!�V����)���d��vc�:y��0�ȟ>���G�      xc��8�|����켔�Ҽg���`�����r�E:�$,�#ߵ�Y/X���º�ˬ�H�}:? �:w;��);�l7;j�?;�C;LF;�(G;F�G;��G;2)H;�RH;�sH;��H;��H;�H;μH;��H;��H;,�H;��H;l�H;��H;,�H;��H;��H;μH;�H;��H;��H;�sH;�RH;2)H;��G;F�G;�(G;LF;�C;j�?;�l7;��);w;? �:H�}:�ˬ���ºY/X�#ߵ�$,�E:���r�`���g�����Ҽ��|����8�      ����-��#Ȥ�d���ݫ���f�G�=����	�ܻ�*��>o5�s���Q(7H�}:�m�:��;>&;��4;C�=;�B;,�E;T�F;̀G;$�G;cH;�@H;�dH;d�H;��H;y�H;��H;��H;;�H;��H;��H;��H;l�H;��H;��H;��H;;�H;��H;��H;y�H;��H;d�H;�dH;�@H;cH;$�G;̀G;T�F;,�E;�B;C�=;��4;>&;��;�m�:H�}:Q(7s���>o5��*��	�ܻ���G�=��f�ݫ��d���#Ȥ��-��      ;�V�z5S�Y6H�x�6�� �3,�n?ػG���D^����1�D����9�3�:? �:��;^%;��3;p�<;�B;�
E;?�F;�WG;8�G;u�G;�/H;xVH;�uH;�H;��H;ܰH;��H;��H;��H;k�H;��H;��H;Q�H;��H;��H;k�H;��H;��H;��H;ܰH;��H;�H;�uH;xVH;�/H;u�G;8�G;�WG;?�F;�
E;�B;p�<;��3;^%;��;? �:�3�:���91�D�����D^�G��n?ػ3,�� �x�6�Y6H�z5S�      s��v��,�ܻ�ƻB󩻜��fFL����͸����O�-:h�:���:w;>&;��3;�8<;`�A;%�D;�YF;Z4G;3�G;�G;� H;aIH;VjH;ńH;ٙH;��H;��H;�H;��H;��H;��H;��H;v�H;�H;v�H;��H;��H;��H;��H;�H;��H;��H;ٙH;ńH;VjH;aIH;� H;�G;3�G;Z4G;�YF;%�D;`�A;�8<;��3;>&;w;���:h�:O�-:��͸�����fFL����B��ƻ,�ܻv��      �D^��/X��qF�'}*�'���P���D��Ҭ�lh:��:���:ȏ; �;��);��4;p�<;`�A;f�D;�8F;
G;��G;x�G;jH;C>H;�`H;6|H;��H;��H;��H;��H;��H;}�H;��H;4�H;��H;8�H;��H;8�H;��H;4�H;��H;}�H;��H;��H;��H;��H;��H;6|H;�`H;C>H;jH;x�G;��G;
G;�8F;f�D;`�A;p�<;��4;��); �;ȏ;���:��:lh:�Ҭ��D��P��'��'}*��qF��/X�      ��S���D�-�������'7��9d�R:���:���:@��:Y>;G";^P.;�l7;C�=;�B;%�D;�8F;YG;R�G;��G;�H;�5H;�XH;	uH;=�H;�H;�H;�H;��H;9�H;��H;-�H;M�H;r�H;��H;	�H;��H;r�H;M�H;-�H;��H;9�H;��H;�H;�H;�H;=�H;	uH;�XH;�5H;�H;��G;R�G;YG;�8F;%�D;�B;C�=;�l7;^P.;G";Y>;@��:���:���:d�R:��9��'7���-����D�      �v[:�Ad:7�}:_�:��:0��:D�:��;P;� ;H+;�3;:�:;j�?;�B;�
E;�YF;
G;R�G;��G;nH;�0H;�RH;�oH;�H;f�H;�H;��H;��H;��H;�H;��H;��H;5�H;�H;(�H;q�H;(�H;�H;5�H;��H;��H;�H;��H;��H;��H;�H;f�H;�H;�oH;�RH;�0H;nH;��G;R�G;
G;�YF;�
E;�B;j�?;:�:;�3;H+;� ;P;��;D�:0��:��:_�:7�}:�Ad:      ���:�A�:���:�w;�
;6;��;}$;�{,;ǂ3;_9;�>;ayA;�C;,�E;?�F;Z4G;��G;��G;nH;�.H;PH;'lH;i�H;��H;��H;��H;�H;��H;)�H;r�H;��H;��H;��H;z�H;W�H;��H;W�H;z�H;��H;��H;��H;r�H;)�H;��H;�H;��H;��H;��H;i�H;'lH;PH;�.H;nH;��G;��G;Z4G;?�F;,�E;�C;ayA;�>;_9;ǂ3;�{,;}$;��;6;�
;�w;���:�A�:      �d;� ;�";�%;d�(;�i-;�2;,�6;�:;0>;�A;�XC;y�D;LF;T�F;�WG;3�G;x�G;�H;�0H;PH;�jH;��H;��H;V�H;E�H;�H;��H;��H;�H;��H;��H;��H;�H;��H;j�H;��H;j�H;��H;�H;��H;��H;��H;�H;��H;��H;�H;E�H;V�H;��H;��H;�jH;PH;�0H;�H;x�G;3�G;�WG;T�F;LF;y�D;�XC;�A;0>;�:;,�6;�2;�i-;d�(;�%;�";� ;      ��4;y�4;��5;Rl7;�^9;��;;�=;f�?;��A;�C;��D;��E;�F;�(G;̀G;8�G;�G;jH;�5H;�RH;'lH;��H;̓H;$�H;گH;g�H;<�H;H�H;��H;��H;(�H;��H;C�H;��H;��H;m�H;��H;m�H;��H;��H;C�H;��H;(�H;��H;��H;H�H;<�H;g�H;گH;$�H;̓H;��H;'lH;�RH;�5H;jH;�G;8�G;̀G;�(G;�F;��E;��D;�C;��A;f�?;�=;��;;�^9;Rl7;��5;y�4;      �_?;	�?;7�?;�@;��A;��B;��C;3�D;~hE;#F;\�F;G;�mG;F�G;$�G;u�G;� H;C>H;�XH;�oH;i�H;��H;$�H;\�H;��H;<�H;Y�H;�H;��H;��H;g�H;��H;��H;��H;��H;E�H;^�H;E�H;��H;��H;��H;��H;g�H;��H;��H;�H;Y�H;<�H;��H;\�H;$�H;��H;i�H;�oH;�XH;C>H;� H;u�G;$�G;F�G;�mG;G;\�F;#F;~hE;3�D;��C;��B;��A;�@;7�?;	�?;      �lD;#~D;��D;�D;�[E;,�E;�/F;�F;��F;$8G;�uG;'�G;u�G;��G;cH;�/H;aIH;�`H;	uH;�H;��H;V�H;گH;��H;�H;��H;}�H;#�H;��H;�H;n�H;N�H;��H;��H;��H;��H;7�H;��H;��H;��H;��H;N�H;n�H;�H;��H;#�H;}�H;��H;�H;��H;گH;V�H;��H;�H;	uH;�`H;aIH;�/H;cH;��G;u�G;'�G;�uG;$8G;��F;�F;�/F;,�E;�[E;�D;��D;#~D;      ��F;q�F;��F;�F;��F;�G;�FG; pG;]�G;l�G;�G;��G;"H;2)H;�@H;xVH;VjH;6|H;=�H;f�H;��H;E�H;g�H;<�H;��H;E�H;��H;��H;��H;�H;�H;��H;��H;��H;C�H;��H;��H;��H;C�H;��H;��H;��H;�H;�H;��H;��H;��H;E�H;��H;<�H;g�H;E�H;��H;f�H;=�H;6|H;VjH;xVH;�@H;2)H;"H;��G;�G;l�G;]�G; pG;�FG;�G;��F;�F;��F;q�F;      puG;4xG;/�G;��G;�G;��G;�G;��G;��G;�H;IH;�+H;�?H;�RH;�dH;�uH;ńH;��H;�H;�H;��H;�H;<�H;Y�H;}�H;��H;t�H;m�H;��H;��H;n�H;��H;��H;L�H;��H;-�H;.�H;-�H;��H;L�H;��H;��H;n�H;��H;��H;m�H;t�H;��H;}�H;Y�H;<�H;�H;��H;�H;�H;��H;ńH;�uH;�dH;�RH;�?H;�+H;IH;�H;��G;��G;�G;��G;�G;��G;/�G;4xG;      M�G;��G;��G;��G;��G;��G;WH;H;�'H;7H;�FH;/VH;MeH;�sH;d�H;�H;ٙH;��H;�H;��H;�H;��H;H�H;�H;#�H;��H;m�H;��H;��H;p�H;��H;��H;c�H;��H;V�H;��H;��H;��H;V�H;��H;c�H;��H;��H;p�H;��H;��H;m�H;��H;#�H;�H;H�H;��H;�H;��H;�H;��H;ٙH;�H;d�H;�sH;MeH;/VH;�FH;7H;�'H;H;WH;��G;��G;��G;��G;��G;      �H;�H;s"H;3'H;�-H;�5H;?H;XIH;eTH;�_H;�kH;9wH;��H;��H;��H;��H;��H;��H;�H;��H;��H;��H;��H;��H;��H;��H;��H;��H;>�H;��H;��H;X�H;��H;y�H;��H;��H;��H;��H;��H;y�H;��H;X�H;��H;��H;>�H;��H;��H;��H;��H;��H;��H;��H;��H;��H;�H;��H;��H;��H;��H;��H;��H;9wH;�kH;�_H;eTH;XIH;?H;�5H;�-H;3'H;s"H;�H;      �NH;NOH;�QH;UH;�YH;�_H;�fH;dnH;�vH;,H;�H;��H;R�H;��H;y�H;ܰH;��H;��H;��H;��H;)�H;�H;��H;��H;�H;�H;��H;p�H;��H;��H;V�H;��H;q�H;��H;�H;%�H;?�H;%�H;�H;��H;q�H;��H;V�H;��H;��H;p�H;��H;�H;�H;��H;��H;�H;)�H;��H;��H;��H;��H;ܰH;y�H;��H;R�H;��H;�H;,H;�vH;dnH;�fH;�_H;�YH;UH;�QH;NOH;      �rH;IsH;�tH;�wH;{H;�H;��H;i�H;��H;�H;��H;W�H;ժH;�H;��H;��H;�H;��H;9�H;�H;r�H;��H;(�H;g�H;n�H;�H;n�H;��H;��H;V�H;��H;q�H;��H;�H;_�H;l�H;d�H;l�H;_�H;�H;��H;q�H;��H;V�H;��H;��H;n�H;�H;n�H;g�H;(�H;��H;r�H;�H;9�H;��H;�H;��H;��H;�H;ժH;W�H;��H;�H;��H;i�H;��H;�H;{H;�wH;�tH;IsH;      �H;:�H;z�H;��H;�H;{�H;V�H;��H;L�H; �H;�H;�H;��H;μH;��H;��H;��H;}�H;��H;��H;��H;��H;��H;��H;N�H;��H;��H;��H;X�H;��H;q�H;��H;�H;_�H;��H;��H;��H;��H;��H;_�H;�H;��H;q�H;��H;X�H;��H;��H;��H;N�H;��H;��H;��H;��H;��H;��H;}�H;��H;��H;��H;μH;��H;�H;�H; �H;L�H;��H;V�H;{�H;�H;��H;z�H;:�H;      ��H;�H;�H;f�H;i�H;��H;ͫH;�H;��H;g�H;H�H;.�H;�H;��H;;�H;��H;��H;��H;-�H;��H;��H;��H;C�H;��H;��H;��H;��H;c�H;��H;q�H;��H;�H;X�H;��H;��H;��H;��H;��H;��H;��H;X�H;�H;��H;q�H;��H;c�H;��H;��H;��H;��H;C�H;��H;��H;��H;-�H;��H;��H;��H;;�H;��H;�H;.�H;H�H;g�H;��H;�H;ͫH;��H;i�H;f�H;�H;�H;      ��H;�H;��H;ñH;u�H;r�H;��H;[�H;�H;�H;�H;�H;
�H;��H;��H;k�H;��H;4�H;M�H;5�H;��H;�H;��H;��H;��H;��H;L�H;��H;y�H;��H;�H;_�H;��H;��H;��H;��H;��H;��H;��H;��H;��H;_�H;�H;��H;y�H;��H;L�H;��H;��H;��H;��H;�H;��H;5�H;M�H;4�H;��H;k�H;��H;��H;
�H;�H;�H;�H;�H;[�H;��H;r�H;u�H;ñH;��H;�H;      �H;W�H;�H;ܺH;6�H;ɽH;��H;��H;��H;m�H;��H;Q�H;��H;,�H;��H;��H;��H;��H;r�H;�H;z�H;��H;��H;��H;��H;C�H;��H;V�H;��H;�H;_�H;��H;��H;��H;��H;��H;��H;��H;��H;��H;��H;��H;_�H;�H;��H;V�H;��H;C�H;��H;��H;��H;��H;z�H;�H;r�H;��H;��H;��H;��H;,�H;��H;Q�H;��H;m�H;��H;��H;��H;ɽH;6�H;ܺH;�H;W�H;      q�H;��H;�H;�H;�H;r�H;�H;��H;��H;��H;"�H;a�H;��H;��H;��H;��H;v�H;8�H;��H;(�H;W�H;j�H;m�H;E�H;��H;��H;-�H;��H;��H;%�H;l�H;��H;��H;��H;��H;��H;��H;��H;��H;��H;��H;��H;l�H;%�H;��H;��H;-�H;��H;��H;E�H;m�H;j�H;W�H;(�H;��H;8�H;v�H;��H;��H;��H;��H;a�H;"�H;��H;��H;��H;�H;r�H;�H;�H;�H;��H;      E�H;U�H;��H;��H;��H;��H;��H;G�H;4�H;3�H;F�H;O�H;W�H;l�H;l�H;Q�H;�H;��H;	�H;q�H;��H;��H;��H;^�H;7�H;��H;.�H;��H;��H;?�H;d�H;��H;��H;��H;��H;��H;��H;��H;��H;��H;��H;��H;d�H;?�H;��H;��H;.�H;��H;7�H;^�H;��H;��H;��H;q�H;	�H;��H;�H;Q�H;l�H;l�H;W�H;O�H;F�H;3�H;4�H;G�H;��H;��H;��H;��H;��H;U�H;      q�H;��H;�H;�H;�H;r�H;�H;��H;��H;��H;"�H;a�H;��H;��H;��H;��H;v�H;8�H;��H;(�H;W�H;j�H;m�H;E�H;��H;��H;-�H;��H;��H;%�H;l�H;��H;��H;��H;��H;��H;��H;��H;��H;��H;��H;��H;l�H;%�H;��H;��H;-�H;��H;��H;E�H;m�H;j�H;W�H;(�H;��H;8�H;v�H;��H;��H;��H;��H;a�H;"�H;��H;��H;��H;�H;r�H;�H;�H;�H;��H;      �H;W�H;�H;ܺH;6�H;ɽH;��H;��H;��H;m�H;��H;Q�H;��H;,�H;��H;��H;��H;��H;r�H;�H;z�H;��H;��H;��H;��H;C�H;��H;V�H;��H;�H;_�H;��H;��H;��H;��H;��H;��H;��H;��H;��H;��H;��H;_�H;�H;��H;V�H;��H;C�H;��H;��H;��H;��H;z�H;�H;r�H;��H;��H;��H;��H;,�H;��H;Q�H;��H;m�H;��H;��H;��H;ɽH;6�H;ܺH;�H;W�H;      ��H;�H;��H;ñH;u�H;r�H;��H;[�H;�H;�H;�H;�H;
�H;��H;��H;k�H;��H;4�H;M�H;5�H;��H;�H;��H;��H;��H;��H;L�H;��H;y�H;��H;�H;_�H;��H;��H;��H;��H;��H;��H;��H;��H;��H;_�H;�H;��H;y�H;��H;L�H;��H;��H;��H;��H;�H;��H;5�H;M�H;4�H;��H;k�H;��H;��H;
�H;�H;�H;�H;�H;[�H;��H;r�H;u�H;ñH;��H;�H;      ��H;�H;�H;f�H;i�H;��H;ͫH;�H;��H;g�H;H�H;.�H;�H;��H;;�H;��H;��H;��H;-�H;��H;��H;��H;C�H;��H;��H;��H;��H;c�H;��H;q�H;��H;�H;X�H;��H;��H;��H;��H;��H;��H;��H;X�H;�H;��H;q�H;��H;c�H;��H;��H;��H;��H;C�H;��H;��H;��H;-�H;��H;��H;��H;;�H;��H;�H;.�H;H�H;g�H;��H;�H;ͫH;��H;i�H;f�H;�H;�H;      �H;:�H;z�H;��H;�H;{�H;V�H;��H;L�H; �H;�H;�H;��H;μH;��H;��H;��H;}�H;��H;��H;��H;��H;��H;��H;N�H;��H;��H;��H;X�H;��H;q�H;��H;�H;_�H;��H;��H;��H;��H;��H;_�H;�H;��H;q�H;��H;X�H;��H;��H;��H;N�H;��H;��H;��H;��H;��H;��H;}�H;��H;��H;��H;μH;��H;�H;�H; �H;L�H;��H;V�H;{�H;�H;��H;z�H;:�H;      �rH;IsH;�tH;�wH;{H;�H;��H;i�H;��H;�H;��H;W�H;ժH;�H;��H;��H;�H;��H;9�H;�H;r�H;��H;(�H;g�H;n�H;�H;n�H;��H;��H;V�H;��H;q�H;��H;�H;_�H;l�H;d�H;l�H;_�H;�H;��H;q�H;��H;V�H;��H;��H;n�H;�H;n�H;g�H;(�H;��H;r�H;�H;9�H;��H;�H;��H;��H;�H;ժH;W�H;��H;�H;��H;i�H;��H;�H;{H;�wH;�tH;IsH;      �NH;NOH;�QH;UH;�YH;�_H;�fH;dnH;�vH;,H;�H;��H;R�H;��H;y�H;ܰH;��H;��H;��H;��H;)�H;�H;��H;��H;�H;�H;��H;p�H;��H;��H;V�H;��H;q�H;��H;�H;%�H;?�H;%�H;�H;��H;q�H;��H;V�H;��H;��H;p�H;��H;�H;�H;��H;��H;�H;)�H;��H;��H;��H;��H;ܰH;y�H;��H;R�H;��H;�H;,H;�vH;dnH;�fH;�_H;�YH;UH;�QH;NOH;      �H;�H;s"H;3'H;�-H;�5H;?H;XIH;eTH;�_H;�kH;9wH;��H;��H;��H;��H;��H;��H;�H;��H;��H;��H;��H;��H;��H;��H;��H;��H;>�H;��H;��H;X�H;��H;y�H;��H;��H;��H;��H;��H;y�H;��H;X�H;��H;��H;>�H;��H;��H;��H;��H;��H;��H;��H;��H;��H;�H;��H;��H;��H;��H;��H;��H;9wH;�kH;�_H;eTH;XIH;?H;�5H;�-H;3'H;s"H;�H;      M�G;��G;��G;��G;��G;��G;WH;H;�'H;7H;�FH;/VH;MeH;�sH;d�H;�H;ٙH;��H;�H;��H;�H;��H;H�H;�H;#�H;��H;m�H;��H;��H;p�H;��H;��H;c�H;��H;V�H;��H;��H;��H;V�H;��H;c�H;��H;��H;p�H;��H;��H;m�H;��H;#�H;�H;H�H;��H;�H;��H;�H;��H;ٙH;�H;d�H;�sH;MeH;/VH;�FH;7H;�'H;H;WH;��G;��G;��G;��G;��G;      puG;4xG;/�G;��G;�G;��G;�G;��G;��G;�H;IH;�+H;�?H;�RH;�dH;�uH;ńH;��H;�H;�H;��H;�H;<�H;Y�H;}�H;��H;t�H;m�H;��H;��H;n�H;��H;��H;L�H;��H;-�H;.�H;-�H;��H;L�H;��H;��H;n�H;��H;��H;m�H;t�H;��H;}�H;Y�H;<�H;�H;��H;�H;�H;��H;ńH;�uH;�dH;�RH;�?H;�+H;IH;�H;��G;��G;�G;��G;�G;��G;/�G;4xG;      ��F;q�F;��F;�F;��F;�G;�FG; pG;]�G;l�G;�G;��G;"H;2)H;�@H;xVH;VjH;6|H;=�H;f�H;��H;E�H;g�H;<�H;��H;E�H;��H;��H;��H;�H;�H;��H;��H;��H;C�H;��H;��H;��H;C�H;��H;��H;��H;�H;�H;��H;��H;��H;E�H;��H;<�H;g�H;E�H;��H;f�H;=�H;6|H;VjH;xVH;�@H;2)H;"H;��G;�G;l�G;]�G; pG;�FG;�G;��F;�F;��F;q�F;      �lD;#~D;��D;�D;�[E;,�E;�/F;�F;��F;$8G;�uG;'�G;u�G;��G;cH;�/H;aIH;�`H;	uH;�H;��H;V�H;گH;��H;�H;��H;}�H;#�H;��H;�H;n�H;N�H;��H;��H;��H;��H;7�H;��H;��H;��H;��H;N�H;n�H;�H;��H;#�H;}�H;��H;�H;��H;گH;V�H;��H;�H;	uH;�`H;aIH;�/H;cH;��G;u�G;'�G;�uG;$8G;��F;�F;�/F;,�E;�[E;�D;��D;#~D;      �_?;	�?;7�?;�@;��A;��B;��C;3�D;~hE;#F;\�F;G;�mG;F�G;$�G;u�G;� H;C>H;�XH;�oH;i�H;��H;$�H;\�H;��H;<�H;Y�H;�H;��H;��H;g�H;��H;��H;��H;��H;E�H;^�H;E�H;��H;��H;��H;��H;g�H;��H;��H;�H;Y�H;<�H;��H;\�H;$�H;��H;i�H;�oH;�XH;C>H;� H;u�G;$�G;F�G;�mG;G;\�F;#F;~hE;3�D;��C;��B;��A;�@;7�?;	�?;      ��4;y�4;��5;Rl7;�^9;��;;�=;f�?;��A;�C;��D;��E;�F;�(G;̀G;8�G;�G;jH;�5H;�RH;'lH;��H;̓H;$�H;گH;g�H;<�H;H�H;��H;��H;(�H;��H;C�H;��H;��H;m�H;��H;m�H;��H;��H;C�H;��H;(�H;��H;��H;H�H;<�H;g�H;گH;$�H;̓H;��H;'lH;�RH;�5H;jH;�G;8�G;̀G;�(G;�F;��E;��D;�C;��A;f�?;�=;��;;�^9;Rl7;��5;y�4;      �d;� ;�";�%;d�(;�i-;�2;,�6;�:;0>;�A;�XC;y�D;LF;T�F;�WG;3�G;x�G;�H;�0H;PH;�jH;��H;��H;V�H;E�H;�H;��H;��H;�H;��H;��H;��H;�H;��H;j�H;��H;j�H;��H;�H;��H;��H;��H;�H;��H;��H;�H;E�H;V�H;��H;��H;�jH;PH;�0H;�H;x�G;3�G;�WG;T�F;LF;y�D;�XC;�A;0>;�:;,�6;�2;�i-;d�(;�%;�";� ;      ���:�A�:���:�w;�
;6;��;}$;�{,;ǂ3;_9;�>;ayA;�C;,�E;?�F;Z4G;��G;��G;nH;�.H;PH;'lH;i�H;��H;��H;��H;�H;��H;)�H;r�H;��H;��H;��H;z�H;W�H;��H;W�H;z�H;��H;��H;��H;r�H;)�H;��H;�H;��H;��H;��H;i�H;'lH;PH;�.H;nH;��G;��G;Z4G;?�F;,�E;�C;ayA;�>;_9;ǂ3;�{,;}$;��;6;�
;�w;���:�A�:      �v[:�Ad:7�}:_�:��:0��:D�:��;P;� ;H+;�3;:�:;j�?;�B;�
E;�YF;
G;R�G;��G;nH;�0H;�RH;�oH;�H;f�H;�H;��H;��H;��H;�H;��H;��H;5�H;�H;(�H;q�H;(�H;�H;5�H;��H;��H;�H;��H;��H;��H;�H;f�H;�H;�oH;�RH;�0H;nH;��G;R�G;
G;�YF;�
E;�B;j�?;:�:;�3;H+;� ;P;��;D�:0��:��:_�:7�}:�Ad:      ��S���D�-�������'7��9d�R:���:���:@��:Y>;G";^P.;�l7;C�=;�B;%�D;�8F;YG;R�G;��G;�H;�5H;�XH;	uH;=�H;�H;�H;�H;��H;9�H;��H;-�H;M�H;r�H;��H;	�H;��H;r�H;M�H;-�H;��H;9�H;��H;�H;�H;�H;=�H;	uH;�XH;�5H;�H;��G;R�G;YG;�8F;%�D;�B;C�=;�l7;^P.;G";Y>;@��:���:���:d�R:��9��'7���-����D�      �D^��/X��qF�'}*�'���P���D��Ҭ�lh:��:���:ȏ; �;��);��4;p�<;`�A;f�D;�8F;
G;��G;x�G;jH;C>H;�`H;6|H;��H;��H;��H;��H;��H;}�H;��H;4�H;��H;8�H;��H;8�H;��H;4�H;��H;}�H;��H;��H;��H;��H;��H;6|H;�`H;C>H;jH;x�G;��G;
G;�8F;f�D;`�A;p�<;��4;��); �;ȏ;���:��:lh:�Ҭ��D��P��'��'}*��qF��/X�      s��v��,�ܻ�ƻB󩻜��fFL����͸����O�-:h�:���:w;>&;��3;�8<;`�A;%�D;�YF;Z4G;3�G;�G;� H;aIH;VjH;ńH;ٙH;��H;��H;�H;��H;��H;��H;��H;v�H;�H;v�H;��H;��H;��H;��H;�H;��H;��H;ٙH;ńH;VjH;aIH;� H;�G;3�G;Z4G;�YF;%�D;`�A;�8<;��3;>&;w;���:h�:O�-:��͸�����fFL����B��ƻ,�ܻv��      ;�V�z5S�Y6H�x�6�� �3,�n?ػG���D^����1�D����9�3�:? �:��;^%;��3;p�<;�B;�
E;?�F;�WG;8�G;u�G;�/H;xVH;�uH;�H;��H;ܰH;��H;��H;��H;k�H;��H;��H;Q�H;��H;��H;k�H;��H;��H;��H;ܰH;��H;�H;�uH;xVH;�/H;u�G;8�G;�WG;?�F;�
E;�B;p�<;��3;^%;��;? �:�3�:���91�D�����D^�G��n?ػ3,�� �x�6�Y6H�z5S�      ����-��#Ȥ�d���ݫ���f�G�=����	�ܻ�*��>o5�s���Q(7H�}:�m�:��;>&;��4;C�=;�B;,�E;T�F;̀G;$�G;cH;�@H;�dH;d�H;��H;y�H;��H;��H;;�H;��H;��H;��H;l�H;��H;��H;��H;;�H;��H;��H;y�H;��H;d�H;�dH;�@H;cH;$�G;̀G;T�F;,�E;�B;C�=;��4;>&;��;�m�:H�}:Q(7s���>o5��*��	�ܻ���G�=��f�ݫ��d���#Ȥ��-��      xc��8�|����켔�Ҽg���`�����r�E:�$,�#ߵ�Y/X���º�ˬ�H�}:? �:w;��);�l7;j�?;�C;LF;�(G;F�G;��G;2)H;�RH;�sH;��H;��H;�H;μH;��H;��H;,�H;��H;l�H;��H;,�H;��H;��H;μH;�H;��H;��H;�sH;�RH;2)H;��G;F�G;�(G;LF;�C;j�?;�l7;��);w;? �:H�}:�ˬ���ºY/X�#ߵ�$,�E:���r�`���g�����Ҽ��|����8�      �&K���G�ȟ>��0�:y�vc�d��)������!�V����ƻfod���ºQ(7�3�:���: �;^P.;:�:;ayA;y�D;�F;�mG;u�G;"H;�?H;MeH;��H;R�H;ժH;��H;�H;
�H;��H;��H;W�H;��H;��H;
�H;�H;��H;ժH;R�H;��H;MeH;�?H;"H;u�G;�mG;�F;y�D;ayA;:�:;^P.; �;���:�3�:Q(7��ºfod��ƻ��!�V����)���d��vc�:y��0�ȟ>���G�      鰒�Z��������}��c���D�/%��8���Ҽ	c����f�����ƻY/X�s������9h�:ȏ;G";�3;�>;�XC;��E;G;'�G;��G;�+H;/VH;9wH;��H;W�H;�H;.�H;�H;Q�H;a�H;O�H;a�H;Q�H;�H;.�H;�H;W�H;��H;9wH;/VH;�+H;��G;'�G;G;��E;�XC;�>;�3;G";ȏ;h�:���9s���Y/X��ƻ�����f�	c����Ҽ�8�/%���D��c���}�����Z��      \Pν��ʽ*8�������������0�f�u�;���K��Ȥ���f���#ߵ�>o5�1�D�O�-:���:Y>;H+;_9;�A;��D;\�F;�uG;�G;IH;�FH;�kH;�H;��H;�H;H�H;�H;��H;"�H;F�H;"�H;��H;�H;H�H;�H;��H;�H;�kH;�FH;IH;�G;�uG;\�F;��D;�A;_9;H+;Y>;���:O�-:1�D�>o5�#ߵ�����f�Ȥ�K����u�;�0�f������������*8����ʽ      ���N9�C[��s�R�ؽ���s����}���G��K��	c��!�V�$,��*���������:@��:� ;ǂ3;0>;�C;#F;$8G;l�G;�H;7H;�_H;,H;�H; �H;g�H;�H;m�H;��H;3�H;��H;m�H;�H;g�H; �H;�H;,H;�_H;7H;�H;l�G;$8G;#F;�C;0>;ǂ3;� ;@��:��:������*��$,�!�V�	c��K�����G���}��s����R�ؽ�s�C[�N9�      }�=���:���0��Q"�e�����ZPν�榽%����G�����Ҽ���E:�	�ܻ�D^�͸��lh:���:P;�{,;�:;��A;~hE;��F;]�G;��G;�'H;eTH;�vH;��H;L�H;��H;�H;��H;��H;4�H;��H;��H;�H;��H;L�H;��H;�vH;eTH;�'H;��G;]�G;��F;~hE;��A;�:;�{,;P;���:lh:͸���D^�	�ܻE:������Ҽ����G�%���榽ZPν����e��Q"���0���:�      
Dx��s���f�QS���:����B[��7ս�榽��}�u�;��8�)�����r����G������Ҭ����:��;}$;,�6;f�?;3�D;�F; pG;��G;H;XIH;dnH;i�H;��H;�H;[�H;��H;��H;G�H;��H;��H;[�H;�H;��H;i�H;dnH;XIH;H;��G; pG;�F;3�D;f�?;,�6;}$;��;���:�Ҭ����G�������r�)����8�u�;���}��榽�7սB[������:�QS���f��s�      �*���0��ȥ��&���jk��H��#%�B[�ZPν�s��0�f�/%�d��`���G�=�n?ػfFL��D�d�R:D�:��;�2;�=;��C;�/F;�FG;�G;WH;?H;�fH;��H;V�H;ͫH;��H;��H;�H;��H;�H;��H;��H;ͫH;V�H;��H;�fH;?H;WH;�G;�FG;�/F;��C;�=;�2;��;D�:d�R:�D�fFL�n?ػG�=�`���d��/%�0�f��s��ZPνB[��#%��H�jk�&���ȥ���0��      �þ��������R��f쏾�s��H����������������D�vc�g����f�3,�����P����90��:6;�i-;��;;��B;,�E;�G;��G;��G;�5H;�_H;�H;{�H;��H;r�H;ɽH;r�H;��H;r�H;ɽH;r�H;��H;{�H;�H;�_H;�5H;��G;��G;�G;,�E;��B;��;;�i-;6;0��:��9�P�����3,��f�g���vc���D���������������H��s�f쏾�R���������      ����fYؾ�þ�ê�f쏾jk���:�e�R�ؽ�����c�:y���Ҽݫ��� �B�'����'7��:�
;d�(;�^9;��A;�[E;��F;�G;��G;�-H;�YH;{H;�H;i�H;u�H;6�H;�H;��H;�H;6�H;u�H;i�H;�H;{H;�YH;�-H;��G;�G;��F;�[E;��A;�^9;d�(;�
;��:��'7'��B�� �ݫ����Ҽ:y��c�����R�ؽe���:�jk�f쏾�ê��þfYؾ��      ��=������I��þ�R��&���QS��Q"��s�����}��0���d���x�6��ƻ'}*����_�:�w;�%;Rl7;�@;�D;�F;��G;��G;3'H;UH;�wH;��H;f�H;ñH;ܺH;�H;��H;�H;ܺH;ñH;f�H;��H;�wH;UH;3'H;��G;��G;�F;�D;�@;Rl7;�%;�w;_�:���'}*��ƻx�6�d����켟0���}�����s��Q"�QS�&����R���þIᾁ���=��      ���>��&�
�����fYؾ���ȥ����f���0�C[�*8������ȟ>�|���#Ȥ�Y6H�,�ܻ�qF�-��7�}:���:�";��5;7�?;��D;��F;/�G;��G;s"H;�QH;�tH;z�H;�H;��H;�H;�H;��H;�H;�H;��H;�H;z�H;�tH;�QH;s"H;��G;/�G;��F;��D;7�?;��5;�";���:7�}:-���qF�,�ܻY6H�#Ȥ�|���ȟ>�����*8��C[���0���f�ȥ�����fYؾ����&�
�>��      �� �k��>��=���������0���s���:�N9���ʽZ����G��8��-��z5S�v���/X���D��Ad:�A�:� ;y�4;	�?;#~D;q�F;4xG;��G;�H;NOH;IsH;:�H;�H;�H;W�H;��H;U�H;��H;W�H;�H;�H;:�H;IsH;NOH;�H;��G;4xG;q�F;#~D;	�?;y�4;� ;�A�:�Ad:��D��/X�v��z5S��-���8���G�Z����ʽN9���:��s��0��������=��>��k��      3F�/h��ǰ�3Vھ�������~���S��#��o��S��Q₽�6�-���<y��FB��Eֻ^A?��	�Y�:���:�";�36;�@;��D;��F;�mG;&�G;>H;:?H;fH;w�H;P�H;��H;��H;�H;�H;�H;��H;��H;P�H;w�H;fH;:?H;>H;&�G;�mG;��F;��D;�@;�36;�";���:Y�:�	�^A?��EֻFB�<y��-����6�Q₽S���o���#��S��~��������3Vھǰ�/h��      /h���b���쾅*־�v������)�� �O�6� ��r�r���؀��3����ݜ��>��ѻ��9�����n�:�$ ;�L#;˃6;�@@;C�D;�F;<pG;��G;TH;@H;�fH;�H;��H;�H;>�H;�H;��H;�H;>�H;�H;��H;�H;�fH;@H;TH;��G;<pG;�F;C�D;�@@;˃6;�L#;�$ ;�n�:�����9��ѻ�>�ݜ�����3��؀��r���r�6� � �O��)������v���*־�쾼b��      ǰ�쾐�޾5ʾ/;���:����v��E�A'���L����u�X�+�aW缨A��r�4�m�Ļ�8)��j��W�:�;�%;kk7;g�@;B�D;4�F;wG;��G;vH;cBH;YhH;B�H;��H;ƩH;�H;��H;��H;��H;�H;ƩH;��H;B�H;YhH;cBH;vH;��G;wG;4�F;B�D;g�@;kk7;�%;�;W�:�j���8)�m�Ļr�4��A��aW�X�+���u�L����A'��E���v��:��/;��5ʾ��޾��      3Vھ�*־5ʾT��������M���9b��5���}�սn���Xc�ݟ���ռ�I��$�$�4T���Z�_����:��;��';��8;^QA;�8E;��F;�G;%�G;�H;-FH;@kH;u�H;[�H;�H;�H;��H;t�H;��H;�H;�H;[�H;u�H;@kH;-FH;�H;%�G;�G;��F;�8E;^QA;��8;��';��;��:_���Z�4T��$�$��I����ռݟ��Xc�n��}�ս���5��9b��M������T���5ʾ�*־      ���v��/;������:P���r�U�H�6� ��~��@������Q�K�<��վ���s�F��_�~ܺ3u9�%�:��;��+;��:;"B;��E;,�F;��G;�G;nH;[KH;(oH;k�H;��H;ƬH;_�H;��H;��H;��H;_�H;ƬH;��H;k�H;(oH;[KH;nH;�G;��G;,�F;��E;"B;��:;��+;��;�%�:3u9~ܺ_�F����s��վ�<�Q�K�����@���~��6� �U�H��r�:P������/;���v��      ��������:���M���r� �O��",�<�
��gٽKĥ�|�u�K1�(����Τ�m�P��Z�q.o�jp���:Դ�:|P;��/;��<;G
C;f�E;� G;^�G;6�G;�$H;�QH;�sH;%�H;f�H;��H;*�H;{�H;&�H;{�H;*�H;��H;f�H;%�H;�sH;�QH;�$H;6�G;^�G;� G;f�E;G
C;��<;��/;|P;Դ�:�:jp��q.o��Z�m�P��Τ�(���K1�|�u�Kĥ��gٽ<�
��",� �O��r��M���:�����      �~���)����v��9b�U�H��",�0Z���S��X^��e�N�{����μ�I���%+�ښ����.������i~:���:�l;@�3;��>;�C;�OF;�EG;|�G;"�G;�.H;'YH;�yH;q�H;��H;��H;F�H;K�H;��H;K�H;F�H;��H;��H;q�H;�yH;'YH;�.H;"�G;|�G;�EG;�OF;�C;��>;@�3;�l;���:�i~:������.�ښ���%+��I����μ{��e�N�X^��S����0Z��",�U�H��9b���v��)��      �S� �O��E��5�6� �<�
���|9��l���Xc���(����߈��Z�[����nݎ�ܺN99���:��	;�c';��7;��@;��D;/�F;biG;��G;�H;�9H;gaH;�H;0�H;P�H;g�H;��H;Y�H;��H;Y�H;��H;g�H;P�H;0�H;�H;gaH;�9H;�H;��G;biG;/�F;��D;��@;��7;�c';��	;���:N99ܺnݎ����Z�[�߈�������(��Xc�l��|9����<�
�6� ��5��E� �O�      �#�6� �A'����~���gٽS��l���j��3�ji��վ�T����(�P�Ļ+A?���B�8�@:[�:�P;w�.;Q�;;�sB;\�E;��F;l�G;'�G;H;�EH;KjH;��H;H�H;.�H;��H;0�H;��H;�H;��H;0�H;��H;.�H;H�H;��H;KjH;�EH;H;'�G;l�G;��F;\�E;�sB;Q�;;w�.;�P;[�:8�@:��B�+A?�P�Ļ�(�T����վ�ji��3��j�l��S���gٽ�~����A'�6� �      �o���r���}�ս@��Kĥ�X^���Xc��3���	���˼t]��FB��Z򻆜��CӺC��8�:{�;RM#;�<5;x?;��C;�?F;K9G;-�G;M�G;c&H;�QH;�sH;ۍH;��H;H�H;кH;��H;��H;a�H;��H;��H;кH;H�H;��H;ۍH;�sH;�QH;c&H;M�G;-�G;K9G;�?F;��C;x?;�<5;RM#;{�;�:C��8CӺ�����Z�FB�t]����˼��	��3��Xc�X^��Kĥ�@��}�ս���r�      S���r��L��n������|�u�e�N���(�ji���˼�A��b�P�=s��|������\:��:�;�m-;F�:;O�A;�+E;��F;mnG;,�G;�H;�6H;k^H;0}H;�H;&�H;��H;/�H;��H;Z�H;��H;Z�H;��H;/�H;��H;&�H;�H;0}H;k^H;�6H;�H;,�G;mnG;��F;�+E;O�A;F�:;�m-;�;��:�\:����|��=s�b�P��A����˼ji���(�e�N�|�u�����n��L���r��      Q₽�؀���u��Xc�Q�K�K1�{�����վ�t]��b�P�l��T��g�9� �o�n2�9�%�:��	;�%;��5;�>;��C;	F;� G;ޙG;�G;pH;�GH;�jH;ʆH;s�H;��H;̸H;��H;l�H;��H;��H;��H;l�H;��H;̸H;��H;s�H;ʆH;�jH;�GH;pH;�G;ޙG;� G;	F;��C;�>;��5;�%;��	;�%�:n2�9 �o�g�9�T��l��b�P�t]���վ����{��K1�Q�K��Xc���u��؀�      �6��3�X�+�ݟ�<�(�����μ߈��T���FB�=s�T����D��{���8u92q�:���:�X;at0;T�;;1B;D9E;/�F;:gG;�G;=�G;�/H;�WH;SwH;G�H;��H;$�H;�H; �H;2�H;I�H;S�H;I�H;2�H; �H;�H;$�H;��H;G�H;SwH;�WH;�/H;=�G;�G;:gG;/�F;D9E;1B;T�;;at0;�X;���:2q�:�8u9�{����D�T��=s�FB�T���߈����μ(���<�ݟ�X�+��3�      -������aW缐�ռ�վ��Τ��I��Z�[��(��Z�g�9��{���99�W�:�W�:�P;�,;�8;�@@;ZAD;�?F;�+G;ÛG;��G;�H;�CH;HgH;W�H;y�H;��H;�H;>�H;:�H;��H;��H;��H;��H;��H;:�H;>�H;�H;��H;y�H;W�H;HgH;�CH;�H;��G;ÛG;�+G;�?F;ZAD;�@@;�8;�,;�P;�W�:�W�:�99�{��g�9���Z��(�Z�[��I���Τ��վ���ռaW缧��      <y��ݜ��A���I����s�m�P��%+����P�Ļ����|� �o��8u9�W�::+�:�;^);8�6;ذ>;�OC;��E;:�F;�wG;a�G;� H;�0H;@WH;*vH;ԎH;9�H;$�H;��H;5�H;^�H;��H;�H;��H;�H;��H;^�H;5�H;��H;$�H;9�H;ԎH;*vH;@WH;�0H;� H;a�G;�wG;:�F;��E;�OC;ذ>;8�6;^);�;:+�:�W�:�8u9 �o�|�����P�Ļ����%+�m�P���s��I���A��ݜ�      FB��>�r�4�$�$�F���Z�ښ��nݎ�+A?�CӺ����n2�92q�:�W�:�;E�';�<5;֜=;[�B;jFE;��F;�TG;Z�G;�G;�H;�GH;9iH;�H;��H;g�H;T�H;f�H;��H;[�H;(�H;6�H;��H;6�H;(�H;[�H;��H;f�H;T�H;g�H;��H;�H;9iH;�GH;�H;�G;Z�G;�TG;��F;jFE;[�B;֜=;�<5;E�';�;�W�:2q�:n2�9����CӺ+A?�nݎ�ښ���Z�F��$�$�r�4��>�      �Eֻ�ѻm�Ļ4T��_�q.o���.�ܺ��B�C��8�\:�%�:���:�P;^);�<5;L:=;x"B;��D;!uF;,6G;��G;��G;�H;�9H;:]H;�yH;�H;��H;�H;'�H;��H;u�H;6�H;��H;B�H;��H;B�H;��H;6�H;u�H;��H;'�H;�H;��H;�H;�yH;:]H;�9H;�H;��G;��G;,6G;!uF;��D;x"B;L:=;�<5;^);�P;���:�%�:�\:C��8��B�ܺ��.�q.o�_�4T��m�Ļ�ѻ      ^A?���9��8)��Z�~ܺjp������N998�@:�:��:��	;�X;�,;8�6;֜=;x"B; �D;�WF;!G;��G;T�G;�H; .H;�RH;�pH;�H;ԜH;��H;׸H;��H;��H;��H;��H;��H;0�H;��H;0�H;��H;��H;��H;��H;��H;׸H;��H;ԜH;�H;�pH;�RH; .H;�H;T�G;��G;!G;�WF; �D;x"B;֜=;8�6;�,;�X;��	;��:�:8�@:N99����jp��~ܺ�Z��8)���9�      �	�����j��_��3u9�:�i~:���:[�:{�;�;�%;at0;�8;ذ>;[�B;��D;�WF;tG;��G;��G;��G;%H;.JH;�hH;�H;��H;T�H;��H;�H;x�H;��H;��H;H�H;��H;��H;i�H;��H;��H;H�H;��H;��H;x�H;�H;��H;T�H;��H;�H;�hH;.JH;%H;��G;��G;��G;tG;�WF;��D;[�B;ذ>;�8;at0;�%;�;{�;[�:���:�i~:�:3u9_���j�����      Y�:�n�:W�:��:�%�:Դ�:���:��	;�P;RM#;�m-;��5;T�;;�@@;�OC;jFE;!uF;!G;��G;�G;F�G;xH;7DH;�bH;e|H;��H;ԢH;��H;ۻH;��H;��H;B�H;j�H;e�H;^�H;��H;��H;��H;^�H;e�H;j�H;B�H;��H;��H;ۻH;��H;ԢH;��H;e|H;�bH;7DH;xH;F�G;�G;��G;!G;!uF;jFE;�OC;�@@;T�;;��5;�m-;RM#;�P;��	;���:Դ�:�%�:��:W�:�n�:      ���:�$ ;�;��;��;|P;�l;�c';w�.;�<5;F�:;�>;1B;ZAD;��E;��F;,6G;��G;��G;F�G;�H;AH;0_H;mxH;��H;<�H;m�H;��H;b�H;��H;��H;F�H;��H;S�H;�H;��H;[�H;��H;�H;S�H;��H;F�H;��H;��H;b�H;��H;m�H;<�H;��H;mxH;0_H;AH;�H;F�G;��G;��G;,6G;��F;��E;ZAD;1B;�>;F�:;�<5;w�.;�c';�l;|P;��;��;�;�$ ;      �";�L#;�%;��';��+;��/;@�3;��7;Q�;;x?;O�A;��C;D9E;�?F;:�F;�TG;��G;T�G;��G;xH;AH;�]H;hvH;9�H;��H;��H;��H;E�H;�H;7�H;1�H;��H;��H;��H;x�H;U�H;��H;U�H;x�H;��H;��H;��H;1�H;7�H;�H;E�H;��H;��H;��H;9�H;hvH;�]H;AH;xH;��G;T�G;��G;�TG;:�F;�?F;D9E;��C;O�A;x?;Q�;;��7;@�3;��/;��+;��';�%;�L#;      �36;˃6;kk7;��8;��:;��<;��>;��@;�sB;��C;�+E;	F;/�F;�+G;�wG;Z�G;��G;�H;%H;7DH;0_H;hvH;O�H;P�H;h�H;��H;��H;��H;��H;�H;=�H;Q�H;��H;m�H;��H;{�H;��H;{�H;��H;m�H;��H;Q�H;=�H;�H;��H;��H;��H;��H;h�H;P�H;O�H;hvH;0_H;7DH;%H;�H;��G;Z�G;�wG;�+G;/�F;	F;�+E;��C;�sB;��@;��>;��<;��:;��8;kk7;˃6;      �@;�@@;g�@;^QA;"B;G
C;�C;��D;\�E;�?F;��F;� G;:gG;ÛG;a�G;�G;�H; .H;.JH;�bH;mxH;9�H;P�H;ܨH;#�H;��H;��H;��H;"�H;\�H;��H;[�H;K�H;��H;��H;i�H;��H;i�H;��H;��H;K�H;[�H;��H;\�H;"�H;��H;��H;��H;#�H;ܨH;P�H;9�H;mxH;�bH;.JH; .H;�H;�G;a�G;ÛG;:gG;� G;��F;�?F;\�E;��D;�C;G
C;"B;^QA;g�@;�@@;      ��D;C�D;B�D;�8E;��E;f�E;�OF;/�F;��F;K9G;mnG;ޙG;�G;��G;� H;�H;�9H;�RH;�hH;e|H;��H;��H;h�H;#�H;U�H;��H;@�H;~�H;��H;9�H;��H;�H;��H;��H;��H;-�H;r�H;-�H;��H;��H;��H;�H;��H;9�H;��H;~�H;@�H;��H;U�H;#�H;h�H;��H;��H;e|H;�hH;�RH;�9H;�H;� H;��G;�G;ޙG;mnG;K9G;��F;/�F;�OF;f�E;��E;�8E;B�D;C�D;      ��F;�F;4�F;��F;,�F;� G;�EG;biG;l�G;-�G;,�G;�G;=�G;�H;�0H;�GH;:]H;�pH;�H;��H;<�H;��H;��H;��H;��H;�H;/�H;k�H;��H;��H;��H;��H;��H;��H;��H;��H;�H;��H;��H;��H;��H;��H;��H;��H;��H;k�H;/�H;�H;��H;��H;��H;��H;<�H;��H;�H;�pH;:]H;�GH;�0H;�H;=�G;�G;,�G;-�G;l�G;biG;�EG;� G;,�F;��F;4�F;�F;      �mG;<pG;wG;�G;��G;^�G;|�G;��G;'�G;M�G;�H;pH;�/H;�CH;@WH;9iH;�yH;�H;��H;ԢH;m�H;��H;��H;��H;@�H;/�H;N�H;��H;h�H;��H;X�H;��H;��H;��H;;�H;��H;��H;��H;;�H;��H;��H;��H;X�H;��H;h�H;��H;N�H;/�H;@�H;��H;��H;��H;m�H;ԢH;��H;�H;�yH;9iH;@WH;�CH;�/H;pH;�H;M�G;'�G;��G;|�G;^�G;��G;�G;wG;<pG;      &�G;��G;��G;%�G;�G;6�G;"�G;�H;H;c&H;�6H;�GH;�WH;HgH;*vH;�H;�H;ԜH;T�H;��H;��H;E�H;��H;��H;~�H;k�H;��H;G�H;��H;L�H;��H;��H;��H;k�H;��H;�H; �H;�H;��H;k�H;��H;��H;��H;L�H;��H;G�H;��H;k�H;~�H;��H;��H;E�H;��H;��H;T�H;ԜH;�H;�H;*vH;HgH;�WH;�GH;�6H;c&H;H;�H;"�G;6�G;�G;%�G;��G;��G;      >H;TH;vH;�H;nH;�$H;�.H;�9H;�EH;�QH;k^H;�jH;SwH;W�H;ԎH;��H;��H;��H;��H;ۻH;b�H;�H;��H;"�H;��H;��H;h�H;��H;-�H;��H;��H;��H;b�H;��H;L�H;�H;��H;�H;L�H;��H;b�H;��H;��H;��H;-�H;��H;h�H;��H;��H;"�H;��H;�H;b�H;ۻH;��H;��H;��H;��H;ԎH;W�H;SwH;�jH;k^H;�QH;�EH;�9H;�.H;�$H;nH;�H;vH;TH;      :?H;@H;cBH;-FH;[KH;�QH;'YH;gaH;KjH;�sH;0}H;ʆH;G�H;y�H;9�H;g�H;�H;׸H;�H;��H;��H;7�H;�H;\�H;9�H;��H;��H;L�H;��H;��H;��H;n�H;�H;T�H;��H;��H;��H;��H;��H;T�H;�H;n�H;��H;��H;��H;L�H;��H;��H;9�H;\�H;�H;7�H;��H;��H;�H;׸H;�H;g�H;9�H;y�H;G�H;ʆH;0}H;�sH;KjH;gaH;'YH;�QH;[KH;-FH;cBH;@H;      fH;�fH;YhH;@kH;(oH;�sH;�yH;�H;��H;ۍH;�H;s�H;��H;��H;$�H;T�H;'�H;��H;x�H;��H;��H;1�H;=�H;��H;��H;��H;X�H;��H;��H;��H;t�H;�H;h�H;��H;��H;�H;0�H;�H;��H;��H;h�H;�H;t�H;��H;��H;��H;X�H;��H;��H;��H;=�H;1�H;��H;��H;x�H;��H;'�H;T�H;$�H;��H;��H;s�H;�H;ۍH;��H;�H;�yH;�sH;(oH;@kH;YhH;�fH;      w�H;�H;B�H;u�H;k�H;%�H;q�H;0�H;H�H;��H;&�H;��H;$�H;�H;��H;f�H;��H;��H;��H;B�H;F�H;��H;Q�H;[�H;�H;��H;��H;��H;��H;n�H;�H;z�H;��H; �H;,�H;J�H;I�H;J�H;,�H; �H;��H;z�H;�H;n�H;��H;��H;��H;��H;�H;[�H;Q�H;��H;F�H;B�H;��H;��H;��H;f�H;��H;�H;$�H;��H;&�H;��H;H�H;0�H;q�H;%�H;k�H;u�H;B�H;�H;      P�H;��H;��H;[�H;��H;f�H;��H;P�H;.�H;H�H;��H;̸H;�H;>�H;5�H;��H;u�H;��H;��H;j�H;��H;��H;��H;K�H;��H;��H;��H;��H;b�H;�H;h�H;��H;	�H;:�H;X�H;��H;��H;��H;X�H;:�H;	�H;��H;h�H;�H;b�H;��H;��H;��H;��H;K�H;��H;��H;��H;j�H;��H;��H;u�H;��H;5�H;>�H;�H;̸H;��H;H�H;.�H;P�H;��H;f�H;��H;[�H;��H;��H;      ��H;�H;ƩH;�H;ƬH;��H;��H;g�H;��H;кH;/�H;��H; �H;:�H;^�H;[�H;6�H;��H;H�H;e�H;S�H;��H;m�H;��H;��H;��H;��H;k�H;��H;T�H;��H; �H;:�H;u�H;��H;��H;��H;��H;��H;u�H;:�H; �H;��H;T�H;��H;k�H;��H;��H;��H;��H;m�H;��H;S�H;e�H;H�H;��H;6�H;[�H;^�H;:�H; �H;��H;/�H;кH;��H;g�H;��H;��H;ƬH;�H;ƩH;�H;      ��H;>�H;�H;�H;_�H;*�H;F�H;��H;0�H;��H;��H;l�H;2�H;��H;��H;(�H;��H;��H;��H;^�H;�H;x�H;��H;��H;��H;��H;;�H;��H;L�H;��H;��H;,�H;X�H;��H;��H;��H;��H;��H;��H;��H;X�H;,�H;��H;��H;L�H;��H;;�H;��H;��H;��H;��H;x�H;�H;^�H;��H;��H;��H;(�H;��H;��H;2�H;l�H;��H;��H;0�H;��H;F�H;*�H;_�H;�H;�H;>�H;      �H;�H;��H;��H;��H;{�H;K�H;Y�H;��H;��H;Z�H;��H;I�H;��H;�H;6�H;B�H;0�H;��H;��H;��H;U�H;{�H;i�H;-�H;��H;��H;�H;�H;��H;�H;J�H;��H;��H;��H;��H;��H;��H;��H;��H;��H;J�H;�H;��H;�H;�H;��H;��H;-�H;i�H;{�H;U�H;��H;��H;��H;0�H;B�H;6�H;�H;��H;I�H;��H;Z�H;��H;��H;Y�H;K�H;{�H;��H;��H;��H;�H;      �H;��H;��H;t�H;��H;&�H;��H;��H;�H;a�H;��H;��H;S�H;��H;��H;��H;��H;��H;i�H;��H;[�H;��H;��H;��H;r�H;�H;��H; �H;��H;��H;0�H;I�H;��H;��H;��H;��H;��H;��H;��H;��H;��H;I�H;0�H;��H;��H; �H;��H;�H;r�H;��H;��H;��H;[�H;��H;i�H;��H;��H;��H;��H;��H;S�H;��H;��H;a�H;�H;��H;��H;&�H;��H;t�H;��H;��H;      �H;�H;��H;��H;��H;{�H;K�H;Y�H;��H;��H;Z�H;��H;I�H;��H;�H;6�H;B�H;0�H;��H;��H;��H;U�H;{�H;i�H;-�H;��H;��H;�H;�H;��H;�H;J�H;��H;��H;��H;��H;��H;��H;��H;��H;��H;J�H;�H;��H;�H;�H;��H;��H;-�H;i�H;{�H;U�H;��H;��H;��H;0�H;B�H;6�H;�H;��H;I�H;��H;Z�H;��H;��H;Y�H;K�H;{�H;��H;��H;��H;�H;      ��H;>�H;�H;�H;_�H;*�H;F�H;��H;0�H;��H;��H;l�H;2�H;��H;��H;(�H;��H;��H;��H;^�H;�H;x�H;��H;��H;��H;��H;;�H;��H;L�H;��H;��H;,�H;X�H;��H;��H;��H;��H;��H;��H;��H;X�H;,�H;��H;��H;L�H;��H;;�H;��H;��H;��H;��H;x�H;�H;^�H;��H;��H;��H;(�H;��H;��H;2�H;l�H;��H;��H;0�H;��H;F�H;*�H;_�H;�H;�H;>�H;      ��H;�H;ƩH;�H;ƬH;��H;��H;g�H;��H;кH;/�H;��H; �H;:�H;^�H;[�H;6�H;��H;H�H;e�H;S�H;��H;m�H;��H;��H;��H;��H;k�H;��H;T�H;��H; �H;:�H;u�H;��H;��H;��H;��H;��H;u�H;:�H; �H;��H;T�H;��H;k�H;��H;��H;��H;��H;m�H;��H;S�H;e�H;H�H;��H;6�H;[�H;^�H;:�H; �H;��H;/�H;кH;��H;g�H;��H;��H;ƬH;�H;ƩH;�H;      P�H;��H;��H;[�H;��H;f�H;��H;P�H;.�H;H�H;��H;̸H;�H;>�H;5�H;��H;u�H;��H;��H;j�H;��H;��H;��H;K�H;��H;��H;��H;��H;b�H;�H;h�H;��H;	�H;:�H;X�H;��H;��H;��H;X�H;:�H;	�H;��H;h�H;�H;b�H;��H;��H;��H;��H;K�H;��H;��H;��H;j�H;��H;��H;u�H;��H;5�H;>�H;�H;̸H;��H;H�H;.�H;P�H;��H;f�H;��H;[�H;��H;��H;      w�H;�H;B�H;u�H;k�H;%�H;q�H;0�H;H�H;��H;&�H;��H;$�H;�H;��H;f�H;��H;��H;��H;B�H;F�H;��H;Q�H;[�H;�H;��H;��H;��H;��H;n�H;�H;z�H;��H; �H;,�H;J�H;I�H;J�H;,�H; �H;��H;z�H;�H;n�H;��H;��H;��H;��H;�H;[�H;Q�H;��H;F�H;B�H;��H;��H;��H;f�H;��H;�H;$�H;��H;&�H;��H;H�H;0�H;q�H;%�H;k�H;u�H;B�H;�H;      fH;�fH;YhH;@kH;(oH;�sH;�yH;�H;��H;ۍH;�H;s�H;��H;��H;$�H;T�H;'�H;��H;x�H;��H;��H;1�H;=�H;��H;��H;��H;X�H;��H;��H;��H;t�H;�H;h�H;��H;��H;�H;0�H;�H;��H;��H;h�H;�H;t�H;��H;��H;��H;X�H;��H;��H;��H;=�H;1�H;��H;��H;x�H;��H;'�H;T�H;$�H;��H;��H;s�H;�H;ۍH;��H;�H;�yH;�sH;(oH;@kH;YhH;�fH;      :?H;@H;cBH;-FH;[KH;�QH;'YH;gaH;KjH;�sH;0}H;ʆH;G�H;y�H;9�H;g�H;�H;׸H;�H;��H;��H;7�H;�H;\�H;9�H;��H;��H;L�H;��H;��H;��H;n�H;�H;T�H;��H;��H;��H;��H;��H;T�H;�H;n�H;��H;��H;��H;L�H;��H;��H;9�H;\�H;�H;7�H;��H;��H;�H;׸H;�H;g�H;9�H;y�H;G�H;ʆH;0}H;�sH;KjH;gaH;'YH;�QH;[KH;-FH;cBH;@H;      >H;TH;vH;�H;nH;�$H;�.H;�9H;�EH;�QH;k^H;�jH;SwH;W�H;ԎH;��H;��H;��H;��H;ۻH;b�H;�H;��H;"�H;��H;��H;h�H;��H;-�H;��H;��H;��H;b�H;��H;L�H;�H;��H;�H;L�H;��H;b�H;��H;��H;��H;-�H;��H;h�H;��H;��H;"�H;��H;�H;b�H;ۻH;��H;��H;��H;��H;ԎH;W�H;SwH;�jH;k^H;�QH;�EH;�9H;�.H;�$H;nH;�H;vH;TH;      &�G;��G;��G;%�G;�G;6�G;"�G;�H;H;c&H;�6H;�GH;�WH;HgH;*vH;�H;�H;ԜH;T�H;��H;��H;E�H;��H;��H;~�H;k�H;��H;G�H;��H;L�H;��H;��H;��H;k�H;��H;�H; �H;�H;��H;k�H;��H;��H;��H;L�H;��H;G�H;��H;k�H;~�H;��H;��H;E�H;��H;��H;T�H;ԜH;�H;�H;*vH;HgH;�WH;�GH;�6H;c&H;H;�H;"�G;6�G;�G;%�G;��G;��G;      �mG;<pG;wG;�G;��G;^�G;|�G;��G;'�G;M�G;�H;pH;�/H;�CH;@WH;9iH;�yH;�H;��H;ԢH;m�H;��H;��H;��H;@�H;/�H;N�H;��H;h�H;��H;X�H;��H;��H;��H;;�H;��H;��H;��H;;�H;��H;��H;��H;X�H;��H;h�H;��H;N�H;/�H;@�H;��H;��H;��H;m�H;ԢH;��H;�H;�yH;9iH;@WH;�CH;�/H;pH;�H;M�G;'�G;��G;|�G;^�G;��G;�G;wG;<pG;      ��F;�F;4�F;��F;,�F;� G;�EG;biG;l�G;-�G;,�G;�G;=�G;�H;�0H;�GH;:]H;�pH;�H;��H;<�H;��H;��H;��H;��H;�H;/�H;k�H;��H;��H;��H;��H;��H;��H;��H;��H;�H;��H;��H;��H;��H;��H;��H;��H;��H;k�H;/�H;�H;��H;��H;��H;��H;<�H;��H;�H;�pH;:]H;�GH;�0H;�H;=�G;�G;,�G;-�G;l�G;biG;�EG;� G;,�F;��F;4�F;�F;      ��D;C�D;B�D;�8E;��E;f�E;�OF;/�F;��F;K9G;mnG;ޙG;�G;��G;� H;�H;�9H;�RH;�hH;e|H;��H;��H;h�H;#�H;U�H;��H;@�H;~�H;��H;9�H;��H;�H;��H;��H;��H;-�H;r�H;-�H;��H;��H;��H;�H;��H;9�H;��H;~�H;@�H;��H;U�H;#�H;h�H;��H;��H;e|H;�hH;�RH;�9H;�H;� H;��G;�G;ޙG;mnG;K9G;��F;/�F;�OF;f�E;��E;�8E;B�D;C�D;      �@;�@@;g�@;^QA;"B;G
C;�C;��D;\�E;�?F;��F;� G;:gG;ÛG;a�G;�G;�H; .H;.JH;�bH;mxH;9�H;P�H;ܨH;#�H;��H;��H;��H;"�H;\�H;��H;[�H;K�H;��H;��H;i�H;��H;i�H;��H;��H;K�H;[�H;��H;\�H;"�H;��H;��H;��H;#�H;ܨH;P�H;9�H;mxH;�bH;.JH; .H;�H;�G;a�G;ÛG;:gG;� G;��F;�?F;\�E;��D;�C;G
C;"B;^QA;g�@;�@@;      �36;˃6;kk7;��8;��:;��<;��>;��@;�sB;��C;�+E;	F;/�F;�+G;�wG;Z�G;��G;�H;%H;7DH;0_H;hvH;O�H;P�H;h�H;��H;��H;��H;��H;�H;=�H;Q�H;��H;m�H;��H;{�H;��H;{�H;��H;m�H;��H;Q�H;=�H;�H;��H;��H;��H;��H;h�H;P�H;O�H;hvH;0_H;7DH;%H;�H;��G;Z�G;�wG;�+G;/�F;	F;�+E;��C;�sB;��@;��>;��<;��:;��8;kk7;˃6;      �";�L#;�%;��';��+;��/;@�3;��7;Q�;;x?;O�A;��C;D9E;�?F;:�F;�TG;��G;T�G;��G;xH;AH;�]H;hvH;9�H;��H;��H;��H;E�H;�H;7�H;1�H;��H;��H;��H;x�H;U�H;��H;U�H;x�H;��H;��H;��H;1�H;7�H;�H;E�H;��H;��H;��H;9�H;hvH;�]H;AH;xH;��G;T�G;��G;�TG;:�F;�?F;D9E;��C;O�A;x?;Q�;;��7;@�3;��/;��+;��';�%;�L#;      ���:�$ ;�;��;��;|P;�l;�c';w�.;�<5;F�:;�>;1B;ZAD;��E;��F;,6G;��G;��G;F�G;�H;AH;0_H;mxH;��H;<�H;m�H;��H;b�H;��H;��H;F�H;��H;S�H;�H;��H;[�H;��H;�H;S�H;��H;F�H;��H;��H;b�H;��H;m�H;<�H;��H;mxH;0_H;AH;�H;F�G;��G;��G;,6G;��F;��E;ZAD;1B;�>;F�:;�<5;w�.;�c';�l;|P;��;��;�;�$ ;      Y�:�n�:W�:��:�%�:Դ�:���:��	;�P;RM#;�m-;��5;T�;;�@@;�OC;jFE;!uF;!G;��G;�G;F�G;xH;7DH;�bH;e|H;��H;ԢH;��H;ۻH;��H;��H;B�H;j�H;e�H;^�H;��H;��H;��H;^�H;e�H;j�H;B�H;��H;��H;ۻH;��H;ԢH;��H;e|H;�bH;7DH;xH;F�G;�G;��G;!G;!uF;jFE;�OC;�@@;T�;;��5;�m-;RM#;�P;��	;���:Դ�:�%�:��:W�:�n�:      �	�����j��_��3u9�:�i~:���:[�:{�;�;�%;at0;�8;ذ>;[�B;��D;�WF;tG;��G;��G;��G;%H;.JH;�hH;�H;��H;T�H;��H;�H;x�H;��H;��H;H�H;��H;��H;i�H;��H;��H;H�H;��H;��H;x�H;�H;��H;T�H;��H;�H;�hH;.JH;%H;��G;��G;��G;tG;�WF;��D;[�B;ذ>;�8;at0;�%;�;{�;[�:���:�i~:�:3u9_���j�����      ^A?���9��8)��Z�~ܺjp������N998�@:�:��:��	;�X;�,;8�6;֜=;x"B; �D;�WF;!G;��G;T�G;�H; .H;�RH;�pH;�H;ԜH;��H;׸H;��H;��H;��H;��H;��H;0�H;��H;0�H;��H;��H;��H;��H;��H;׸H;��H;ԜH;�H;�pH;�RH; .H;�H;T�G;��G;!G;�WF; �D;x"B;֜=;8�6;�,;�X;��	;��:�:8�@:N99����jp��~ܺ�Z��8)���9�      �Eֻ�ѻm�Ļ4T��_�q.o���.�ܺ��B�C��8�\:�%�:���:�P;^);�<5;L:=;x"B;��D;!uF;,6G;��G;��G;�H;�9H;:]H;�yH;�H;��H;�H;'�H;��H;u�H;6�H;��H;B�H;��H;B�H;��H;6�H;u�H;��H;'�H;�H;��H;�H;�yH;:]H;�9H;�H;��G;��G;,6G;!uF;��D;x"B;L:=;�<5;^);�P;���:�%�:�\:C��8��B�ܺ��.�q.o�_�4T��m�Ļ�ѻ      FB��>�r�4�$�$�F���Z�ښ��nݎ�+A?�CӺ����n2�92q�:�W�:�;E�';�<5;֜=;[�B;jFE;��F;�TG;Z�G;�G;�H;�GH;9iH;�H;��H;g�H;T�H;f�H;��H;[�H;(�H;6�H;��H;6�H;(�H;[�H;��H;f�H;T�H;g�H;��H;�H;9iH;�GH;�H;�G;Z�G;�TG;��F;jFE;[�B;֜=;�<5;E�';�;�W�:2q�:n2�9����CӺ+A?�nݎ�ښ���Z�F��$�$�r�4��>�      <y��ݜ��A���I����s�m�P��%+����P�Ļ����|� �o��8u9�W�::+�:�;^);8�6;ذ>;�OC;��E;:�F;�wG;a�G;� H;�0H;@WH;*vH;ԎH;9�H;$�H;��H;5�H;^�H;��H;�H;��H;�H;��H;^�H;5�H;��H;$�H;9�H;ԎH;*vH;@WH;�0H;� H;a�G;�wG;:�F;��E;�OC;ذ>;8�6;^);�;:+�:�W�:�8u9 �o�|�����P�Ļ����%+�m�P���s��I���A��ݜ�      -������aW缐�ռ�վ��Τ��I��Z�[��(��Z�g�9��{���99�W�:�W�:�P;�,;�8;�@@;ZAD;�?F;�+G;ÛG;��G;�H;�CH;HgH;W�H;y�H;��H;�H;>�H;:�H;��H;��H;��H;��H;��H;:�H;>�H;�H;��H;y�H;W�H;HgH;�CH;�H;��G;ÛG;�+G;�?F;ZAD;�@@;�8;�,;�P;�W�:�W�:�99�{��g�9���Z��(�Z�[��I���Τ��վ���ռaW缧��      �6��3�X�+�ݟ�<�(�����μ߈��T���FB�=s�T����D��{���8u92q�:���:�X;at0;T�;;1B;D9E;/�F;:gG;�G;=�G;�/H;�WH;SwH;G�H;��H;$�H;�H; �H;2�H;I�H;S�H;I�H;2�H; �H;�H;$�H;��H;G�H;SwH;�WH;�/H;=�G;�G;:gG;/�F;D9E;1B;T�;;at0;�X;���:2q�:�8u9�{����D�T��=s�FB�T���߈����μ(���<�ݟ�X�+��3�      Q₽�؀���u��Xc�Q�K�K1�{�����վ�t]��b�P�l��T��g�9� �o�n2�9�%�:��	;�%;��5;�>;��C;	F;� G;ޙG;�G;pH;�GH;�jH;ʆH;s�H;��H;̸H;��H;l�H;��H;��H;��H;l�H;��H;̸H;��H;s�H;ʆH;�jH;�GH;pH;�G;ޙG;� G;	F;��C;�>;��5;�%;��	;�%�:n2�9 �o�g�9�T��l��b�P�t]���վ����{��K1�Q�K��Xc���u��؀�      S���r��L��n������|�u�e�N���(�ji���˼�A��b�P�=s��|������\:��:�;�m-;F�:;O�A;�+E;��F;mnG;,�G;�H;�6H;k^H;0}H;�H;&�H;��H;/�H;��H;Z�H;��H;Z�H;��H;/�H;��H;&�H;�H;0}H;k^H;�6H;�H;,�G;mnG;��F;�+E;O�A;F�:;�m-;�;��:�\:����|��=s�b�P��A����˼ji���(�e�N�|�u�����n��L���r��      �o���r���}�ս@��Kĥ�X^���Xc��3���	���˼t]��FB��Z򻆜��CӺC��8�:{�;RM#;�<5;x?;��C;�?F;K9G;-�G;M�G;c&H;�QH;�sH;ۍH;��H;H�H;кH;��H;��H;a�H;��H;��H;кH;H�H;��H;ۍH;�sH;�QH;c&H;M�G;-�G;K9G;�?F;��C;x?;�<5;RM#;{�;�:C��8CӺ�����Z�FB�t]����˼��	��3��Xc�X^��Kĥ�@��}�ս���r�      �#�6� �A'����~���gٽS��l���j��3�ji��վ�T����(�P�Ļ+A?���B�8�@:[�:�P;w�.;Q�;;�sB;\�E;��F;l�G;'�G;H;�EH;KjH;��H;H�H;.�H;��H;0�H;��H;�H;��H;0�H;��H;.�H;H�H;��H;KjH;�EH;H;'�G;l�G;��F;\�E;�sB;Q�;;w�.;�P;[�:8�@:��B�+A?�P�Ļ�(�T����վ�ji��3��j�l��S���gٽ�~����A'�6� �      �S� �O��E��5�6� �<�
���|9��l���Xc���(����߈��Z�[����nݎ�ܺN99���:��	;�c';��7;��@;��D;/�F;biG;��G;�H;�9H;gaH;�H;0�H;P�H;g�H;��H;Y�H;��H;Y�H;��H;g�H;P�H;0�H;�H;gaH;�9H;�H;��G;biG;/�F;��D;��@;��7;�c';��	;���:N99ܺnݎ����Z�[�߈�������(��Xc�l��|9����<�
�6� ��5��E� �O�      �~���)����v��9b�U�H��",�0Z���S��X^��e�N�{����μ�I���%+�ښ����.������i~:���:�l;@�3;��>;�C;�OF;�EG;|�G;"�G;�.H;'YH;�yH;q�H;��H;��H;F�H;K�H;��H;K�H;F�H;��H;��H;q�H;�yH;'YH;�.H;"�G;|�G;�EG;�OF;�C;��>;@�3;�l;���:�i~:������.�ښ���%+��I����μ{��e�N�X^��S����0Z��",�U�H��9b���v��)��      ��������:���M���r� �O��",�<�
��gٽKĥ�|�u�K1�(����Τ�m�P��Z�q.o�jp���:Դ�:|P;��/;��<;G
C;f�E;� G;^�G;6�G;�$H;�QH;�sH;%�H;f�H;��H;*�H;{�H;&�H;{�H;*�H;��H;f�H;%�H;�sH;�QH;�$H;6�G;^�G;� G;f�E;G
C;��<;��/;|P;Դ�:�:jp��q.o��Z�m�P��Τ�(���K1�|�u�Kĥ��gٽ<�
��",� �O��r��M���:�����      ���v��/;������:P���r�U�H�6� ��~��@������Q�K�<��վ���s�F��_�~ܺ3u9�%�:��;��+;��:;"B;��E;,�F;��G;�G;nH;[KH;(oH;k�H;��H;ƬH;_�H;��H;��H;��H;_�H;ƬH;��H;k�H;(oH;[KH;nH;�G;��G;,�F;��E;"B;��:;��+;��;�%�:3u9~ܺ_�F����s��վ�<�Q�K�����@���~��6� �U�H��r�:P������/;���v��      3Vھ�*־5ʾT��������M���9b��5���}�սn���Xc�ݟ���ռ�I��$�$�4T���Z�_����:��;��';��8;^QA;�8E;��F;�G;%�G;�H;-FH;@kH;u�H;[�H;�H;�H;��H;t�H;��H;�H;�H;[�H;u�H;@kH;-FH;�H;%�G;�G;��F;�8E;^QA;��8;��';��;��:_���Z�4T��$�$��I����ռݟ��Xc�n��}�ս���5��9b��M������T���5ʾ�*־      ǰ�쾐�޾5ʾ/;���:����v��E�A'���L����u�X�+�aW缨A��r�4�m�Ļ�8)��j��W�:�;�%;kk7;g�@;B�D;4�F;wG;��G;vH;cBH;YhH;B�H;��H;ƩH;�H;��H;��H;��H;�H;ƩH;��H;B�H;YhH;cBH;vH;��G;wG;4�F;B�D;g�@;kk7;�%;�;W�:�j���8)�m�Ļr�4��A��aW�X�+���u�L����A'��E���v��:��/;��5ʾ��޾��      /h���b���쾅*־�v������)�� �O�6� ��r�r���؀��3����ݜ��>��ѻ��9�����n�:�$ ;�L#;˃6;�@@;C�D;�F;<pG;��G;TH;@H;�fH;�H;��H;�H;>�H;�H;��H;�H;>�H;�H;��H;�H;�fH;@H;TH;��G;<pG;�F;C�D;�@@;˃6;�L#;�$ ;�n�:�����9��ѻ�>�ݜ�����3��؀��r���r�6� � �O��)������v���*־�쾼b��      ����]�0_ݾ��ɾK*��Ы���zx��G�0,�U�뽘b�� @{�|�/�\���䙼�J;��ͻ��4�%Wṻ��:�;]�#;��6;VZ@;��D;��F;�kG;��G;{H;�9H;�aH;�H;M�H;V�H;�H;�H;��H;�H;�H;V�H;M�H;�H;�aH;�9H;{H;��G;�kG;��F;��D;VZ@;��6;]�#;�;���:%Wṫ�4��ͻ�J;��䙼\��|�/� @{��b��U��0,��G��zx�Ы��K*����ɾ0_ݾ�]�      �]����:پZ�žI�������8t�I�C�����罽���`w�-�l���_����7��Rɻ�K/� yƹd��:P/;f$;*7;~@;��D;��F;nG;-�G;hH;�:H;�bH;��H;��H;��H;5�H;M�H;B�H;M�H;5�H;��H;��H;��H;�bH;�:H;hH;-�G;nG;��F;��D;~@;*7;f$;P/;d��: yƹ�K/��Rɻ��7��_��l��-�`w����������I�C��8t����I���Z�ž�:پ��      0_ݾ�:پ�V;�*���Ƥ�3a����g�g$:��Z�?ݽkƣ�Al�:.%��߼=��m9.�����"V�2p��@�:�w;�'&;��7;�@;P
E;F�F;�tG;[�G;�
H;=H;|dH;��H;��H;t�H;ֱH;ݷH;عH;ݷH;ֱH;t�H;��H;��H;|dH;=H;�
H;[�G;�tG;F�F;P
E;�@;��7;�'&;�w;�@�:2p�"V�����m9.�=���߼:.%�Al�kƣ�?ݽ�Z�g$:���g�3a���Ƥ��*���V;�:پ      ��ɾZ�ž�*��Sת�Ы��	�����T��J+��a2̽ss���yZ����μ>y�����!Ϩ�+,�d��6���:��
;��(;�M9;D�A;�ME;��F;�~G;�G;�H;�@H;bgH;�H;`�H;��H;��H;ǸH;��H;ǸH;��H;��H;`�H;�H;bgH;�@H;�H;�G;�~G;��F;�ME;D�A;�M9;��(;��
;���:d��6+,�!Ϩ����>y��μ����yZ�ss��a2̽��J+���T�	���Ы��Sת��*��Z�ž      K*��I����Ƥ�Ы���/���c��G=����z�gж��ɇ� �C�����!��);k�z&�|-��E�˺SX�9
��:�8;hh,;9	;;@PB;��E; G;�G;�G;�H;2FH;}kH;/�H;��H;��H;e�H;'�H;��H;'�H;e�H;��H;��H;/�H;}kH;2FH;�H;�G;�G; G;��E;@PB;9	;;hh,;�8;
��:SX�9E�˺|-��z&�);k��!����� �C��ɇ�gж��z����G=��c��/��Ы���Ƥ�I���      Ы�����3a��	����c�J�C�Z#���$vϽ����Al�8g*�T��v
���I�W��p\c��쀺4t,:i��:v�;D_0;��<;�0C;2�E;�"G;}�G;B�G;GH;�LH;fpH;׊H;��H;�H;U�H;»H;��H;»H;U�H;�H;��H;׊H;fpH;�LH;GH;B�G;}�G;�"G;2�E;�0C;��<;D_0;v�;i��:4t,:�쀺p\c�W�軞I�v
��T��8g*�Al�����$vϽ��Z#�J�C��c�	���3a�����      �zx��8t���g���T��G=�Z#��5�?ݽ�b������G������Ǽ>y���$�&����$�vƹ裆:7&�:3� ;�~4;��>;�D;[F;�EG;��G;:�G;8)H;�TH;%vH;&�H;�H;��H;��H;��H;M�H;��H;��H;��H;�H;&�H;%vH;�TH;8)H;:�G;��G;�EG;[F;�D;��>;�~4;3� ;7&�:裆:vƹ�$�&����$�>y����Ǽ���G������b��?ݽ�5�Z#��G=���T���g��8t�      �G�I�C�g$:��J+�����?ݽ4���I���yZ�Ơ"�k�鼢���T�Y� ��L��h�˺�m9�ض:�;�_(;~8;��@;��D;'�F;�gG;��G;� H;e4H; ]H;�|H;�H;ۥH;z�H;�H;ʿH;X�H;ʿH;�H;z�H;ۥH;�H;�|H; ]H;e4H;� H;��G;�gG;'�F;��D;��@;~8;�_(;�;�ض:�m9h�˺�L��Y� �T�����k��Ơ"��yZ�I��4���?ݽ�����J+�g$:�I�C�      0,����Z���z�$vϽ�b��I��.]a�-�D� ��!��(�{��!�f���h�4�P(�?nQ:L�:��;I�/;:'<;B�B;=�E;)�F;φG;��G;hH;o@H;>fH;y�H;]�H;�H;��H;��H;�H;u�H;�H;��H;��H;�H;]�H;y�H;>fH;o@H;hH;��G;φG;)�F;=�E;B�B;:'<;I�/;��;L�:?nQ:P(�h�4�f����!�(�{��!��D� �-�.]a�I���b��$vϽ�z���Z���      U�뽱��?ݽa2̽gж����������yZ�-�����`ļ-O���J;�5��%�|�]�ºPM@9=��:�;Tf$;��5;)N?;�D;�KF;@:G;�G;$�G;� H;MH;�oH;��H;��H;K�H;�H;f�H;��H;��H;��H;f�H;�H;K�H;��H;��H;�oH;MH;� H;$�G;�G;@:G;�KF;�D;)N?;��5;Tf$;�;=��:PM@9]�º%�|�5�軃J;�-O���`ļ���-��yZ���������gж�a2̽?ݽ���      �b������kƣ�ss���ɇ�Al�G�Ơ"�D� ��`ļ6���I��C��ۙ��Ouƹ��k: ��:��;�=.;}	;;+�A;.AE;��F;OlG;��G;��G;�1H;ZH;�yH;�H;��H;��H;|�H;P�H;�H;3�H;�H;P�H;|�H;��H;��H;�H;�yH;ZH;�1H;��G;��G;OlG;��F;.AE;+�A;}	;;�=.;��; ��:��k:Ouƹ��ۙ��C��I�6���`ļD� �Ơ"�G�Al��ɇ�ss��kƣ�����       @{�`w�Al��yZ� �C�8g*����k���!��-O���I�|��Ψ�2K/�_$T��P:���:4�;6(&;^#6;%?;��C;�"F;:#G;^�G;��G;�H;XBH;gH;��H;��H;��H;�H;�H;@�H;��H;��H;��H;@�H;�H;�H;��H;��H;��H;gH;XBH;�H;��G;^�G;:#G;�"F;��C;%?;^#6;6(&;4�;���:�P:_$T�2K/��Ψ�|��I�-O���!��k�鼇��8g*� �C��yZ�Al�`w�      |�/�-�:.%�������T���Ǽ����(�{��J;��C��Ψ�	O:�����}Z�9N��:;�;�-1;l'<;%5B;%NE;Z�F;jeG;�G;h�G;"*H;
SH;�sH;F�H;�H;@�H;i�H;��H;�H;�H;=�H;�H;�H;��H;i�H;@�H;�H;F�H;�sH;
SH;"*H;h�G;�G;jeG;Z�F;%NE;%5B;l'<;�-1;�;;N��:}Z�9����	O:��Ψ��C��J;�(�{�������ǼT��������:.%�-�      \��l�鼟߼μ�!��v
��>y��T��!�5�軈ۙ�2K/�����wm9qA�:���:ƽ;��,;,N9;�~@;^D;
LF;�-G;�G;��G;�H;�>H;DcH;<�H;��H;+�H;��H;��H;��H;��H;��H;��H;��H;��H;��H;��H;��H;+�H;��H;<�H;DcH;�>H;�H;��G;�G;�-G;
LF;^D;�~@;,N9;��,;ƽ;���:qA�:wm9����2K/��ۙ�5���!�T�>y��v
���!��μ�߼l��      �䙼�_��=��>y��);k��I��$�Y� �f���%�|��_$T�}Z�9qA�:���:��;��);�7;=�>; tC;`�E;2�F;%uG;O�G;��G;/+H;�RH;�rH;��H;��H;0�H;�H;��H;S�H;��H;�H;��H;�H;��H;S�H;��H;�H;0�H;��H;��H;�rH;�RH;/+H;��G;O�G;%uG;2�F;`�E; tC;=�>;�7;��);��;���:qA�:}Z�9_$T��%�|�f���Y� ��$��I�);k�>y��=���_��      �J;���7�m9.����z&�W��&����L��h�4�]�ºOuƹ�P:N��:���:��;-�(;.�5;$�=;�B;�ZE;��F;TG;�G;��G;�H;�BH;:eH;�H;��H;�H;��H;�H;��H;p�H;�H;R�H;9�H;R�H;�H;p�H;��H;�H;��H;�H;��H;�H;:eH;�BH;�H;��G;�G;TG;��F;�ZE;�B;$�=;.�5;-�(;��;���:N��:�P:Ouƹ]�ºh�4��L��&���W��z&����m9.���7�      �ͻ�Rɻ����!Ϩ�|-��p\c��$�h�˺P(�PM@9��k:���:;ƽ;��);.�5;��=;vPB;�
E;6F;d7G;z�G;|�G;�H;�4H;�XH;gvH;��H;ѠH;�H;��H;��H;l�H;<�H;��H;��H;9�H;��H;��H;<�H;l�H;��H;��H;�H;ѠH;��H;gvH;�XH;�4H;�H;|�G;z�G;d7G;6F;�
E;vPB;��=;.�5;��);ƽ;;���:��k:PM@9P(�h�˺�$�p\c�|-��!Ϩ������Rɻ      ��4��K/�"V�+,�E�˺�쀺vƹ�m9?nQ:=��: ��:4�;�;��,;�7;$�=;vPB;�D;�bF;]#G;�G;�G;�G;�(H;�MH; mH;��H;�H;E�H;-�H;-�H;��H;��H;��H;��H;��H;'�H;��H;��H;��H;��H;��H;-�H;-�H;E�H;�H;��H; mH;�MH;�(H;�G;�G;�G;]#G;�bF;�D;vPB;$�=;�7;��,;�;4�; ��:=��:?nQ:�m9vƹ�쀺E�˺+,�"V��K/�      %W� yƹ2p�d��6SX�94t,:裆:�ض:L�:�;��;6(&;�-1;,N9;=�>;�B;�
E;�bF;,G;fG;�G;��G;�H;EH;�dH;�~H;ړH;�H;ҲH;��H;(�H;��H;��H;g�H;�H;Z�H;��H;Z�H;�H;g�H;��H;��H;(�H;��H;ҲH;�H;ړH;�~H;�dH;EH;�H;��G;�G;fG;,G;�bF;�
E;�B;=�>;,N9;�-1;6(&;��;�;L�:�ض:裆:4t,:SX�9d��62p� yƹ      ���:d��:�@�:���:
��:i��:7&�:�;��;Tf$;�=.;^#6;l'<;�~@; tC;�ZE;6F;]#G;fG;�G;L�G;�H;?H;�^H;yH;z�H;<�H;ҮH;J�H;��H;��H;d�H;��H;��H;��H;�H;|�H;�H;��H;��H;��H;d�H;��H;��H;J�H;ҮH;<�H;z�H;yH;�^H;?H;�H;L�G;�G;fG;]#G;6F;�ZE; tC;�~@;l'<;^#6;�=.;Tf$;��;�;7&�:i��:
��:���:�@�:d��:      �;P/;�w;��
;�8;v�;3� ;�_(;I�/;��5;}	;;%?;%5B;^D;`�E;��F;d7G;�G;�G;L�G;�H;�;H;�ZH;
uH;��H;q�H;U�H;U�H;��H;��H;��H;~�H;�H;��H;��H;��H;��H;��H;��H;��H;�H;~�H;��H;��H;��H;U�H;U�H;q�H;��H;
uH;�ZH;�;H;�H;L�G;�G;�G;d7G;��F;`�E;^D;%5B;%?;}	;;��5;I�/;�_(;3� ;v�;�8;��
;�w;P/;      ]�#;f$;�'&;��(;hh,;D_0;�~4;~8;:'<;)N?;+�A;��C;%NE;
LF;2�F;TG;z�G;�G;��G;�H;�;H;�YH;sH;�H;��H;��H;�H;�H;��H;)�H;Q�H;F�H;e�H;��H;��H;��H;%�H;��H;��H;��H;e�H;F�H;Q�H;)�H;��H;�H;�H;��H;��H;�H;sH;�YH;�;H;�H;��G;�G;z�G;TG;2�F;
LF;%NE;��C;+�A;)N?;:'<;~8;�~4;D_0;hh,;��(;�'&;f$;      ��6;*7;��7;�M9;9	;;��<;��>;��@;B�B;�D;.AE;�"F;Z�F;�-G;%uG;�G;|�G;�G;�H;?H;�ZH;sH;V�H;r�H;�H;?�H;�H;;�H;�H;4�H;d�H;��H;U�H;>�H;G�H;�H;@�H;�H;G�H;>�H;U�H;��H;d�H;4�H;�H;;�H;�H;?�H;�H;r�H;V�H;sH;�ZH;?H;�H;�G;|�G;�G;%uG;�-G;Z�F;�"F;.AE;�D;B�B;��@;��>;��<;9	;;�M9;��7;*7;      VZ@;~@;�@;D�A;@PB;�0C;�D;��D;=�E;�KF;��F;:#G;jeG;�G;O�G;��G;�H;�(H;EH;�^H;
uH;�H;r�H;}�H;W�H;/�H;@�H;��H;c�H;��H;�H;��H;��H;x�H;t�H;
�H;Q�H;
�H;t�H;x�H;��H;��H;�H;��H;c�H;��H;@�H;/�H;W�H;}�H;r�H;�H;
uH;�^H;EH;�(H;�H;��G;O�G;�G;jeG;:#G;��F;�KF;=�E;��D;�D;�0C;@PB;D�A;�@;~@;      ��D;��D;P
E;�ME;��E;2�E;[F;'�F;)�F;@:G;OlG;^�G;�G;��G;��G;�H;�4H;�MH;�dH;yH;��H;��H;�H;W�H;��H;��H;=�H;��H;�H;��H;c�H;��H;b�H;��H;��H;��H;�H;��H;��H;��H;b�H;��H;c�H;��H;�H;��H;=�H;��H;��H;W�H;�H;��H;��H;yH;�dH;�MH;�4H;�H;��G;��G;�G;^�G;OlG;@:G;)�F;'�F;[F;2�E;��E;�ME;P
E;��D;      ��F;��F;F�F;��F; G;�"G;�EG;�gG;φG;�G;��G;��G;h�G;�H;/+H;�BH;�XH; mH;�~H;z�H;q�H;��H;?�H;/�H;��H;�H;H�H;��H;$�H;)�H;k�H;�H;��H;��H;f�H;��H;��H;��H;f�H;��H;��H;�H;k�H;)�H;$�H;��H;H�H;�H;��H;/�H;?�H;��H;q�H;z�H;�~H; mH;�XH;�BH;/+H;�H;h�G;��G;��G;�G;φG;�gG;�EG;�"G; G;��F;F�F;��F;      �kG;nG;�tG;�~G;�G;}�G;��G;��G;��G;$�G;��G;�H;"*H;�>H;�RH;:eH;gvH;��H;ړH;<�H;U�H;�H;�H;@�H;=�H;H�H;e�H;��H;��H;5�H;*�H;t�H;��H;x�H;�H;d�H;��H;d�H;�H;x�H;��H;t�H;*�H;5�H;��H;��H;e�H;H�H;=�H;@�H;�H;�H;U�H;<�H;ړH;��H;gvH;:eH;�RH;�>H;"*H;�H;��G;$�G;��G;��G;��G;}�G;�G;�~G;�tG;nG;      ��G;-�G;[�G;�G;�G;B�G;:�G;� H;hH;� H;�1H;XBH;
SH;DcH;�rH;�H;��H;�H;�H;ҮH;U�H;�H;;�H;��H;��H;��H;��H;��H;�H;��H;q�H;��H;��H;B�H;��H;��H;#�H;��H;��H;B�H;��H;��H;q�H;��H;�H;��H;��H;��H;��H;��H;;�H;�H;U�H;ҮH;�H;�H;��H;�H;�rH;DcH;
SH;XBH;�1H;� H;hH;� H;:�G;B�G;�G;�G;[�G;-�G;      {H;hH;�
H;�H;�H;GH;8)H;e4H;o@H;MH;ZH;gH;�sH;<�H;��H;��H;ѠH;E�H;ҲH;J�H;��H;��H;�H;c�H;�H;$�H;��H;�H;��H;V�H;�H;��H;A�H;��H;�H;V�H;b�H;V�H;�H;��H;A�H;��H;�H;V�H;��H;�H;��H;$�H;�H;c�H;�H;��H;��H;J�H;ҲH;E�H;ѠH;��H;��H;<�H;�sH;gH;ZH;MH;o@H;e4H;8)H;GH;�H;�H;�
H;hH;      �9H;�:H;=H;�@H;2FH;�LH;�TH; ]H;>fH;�oH;�yH;��H;F�H;��H;��H;�H;�H;-�H;��H;��H;��H;)�H;4�H;��H;��H;)�H;5�H;��H;V�H;��H;w�H;1�H;��H;8�H;��H;��H;��H;��H;��H;8�H;��H;1�H;w�H;��H;V�H;��H;5�H;)�H;��H;��H;4�H;)�H;��H;��H;��H;-�H;�H;�H;��H;��H;F�H;��H;�yH;�oH;>fH; ]H;�TH;�LH;2FH;�@H;=H;�:H;      �aH;�bH;|dH;bgH;}kH;fpH;%vH;�|H;y�H;��H;�H;��H;�H;+�H;0�H;��H;��H;-�H;(�H;��H;��H;Q�H;d�H;�H;c�H;k�H;*�H;q�H;�H;w�H;I�H;��H;2�H;��H;��H;��H;�H;��H;��H;��H;2�H;��H;I�H;w�H;�H;q�H;*�H;k�H;c�H;�H;d�H;Q�H;��H;��H;(�H;-�H;��H;��H;0�H;+�H;�H;��H;�H;��H;y�H;�|H;%vH;fpH;}kH;bgH;|dH;�bH;      �H;��H;��H;�H;/�H;׊H;&�H;�H;]�H;��H;��H;��H;@�H;��H;�H;�H;��H;��H;��H;d�H;~�H;F�H;��H;��H;��H;�H;t�H;��H;��H;1�H;��H;C�H;��H;��H;�H;C�H;5�H;C�H;�H;��H;��H;C�H;��H;1�H;��H;��H;t�H;�H;��H;��H;��H;F�H;~�H;d�H;��H;��H;��H;�H;�H;��H;@�H;��H;��H;��H;]�H;�H;&�H;׊H;/�H;�H;��H;��H;      M�H;��H;��H;`�H;��H;��H;�H;ۥH;�H;K�H;��H;�H;i�H;��H;��H;��H;l�H;��H;��H;��H;�H;e�H;U�H;��H;b�H;��H;��H;��H;A�H;��H;2�H;��H;�H;�H;V�H;l�H;7�H;l�H;V�H;�H;�H;��H;2�H;��H;A�H;��H;��H;��H;b�H;��H;U�H;e�H;�H;��H;��H;��H;l�H;��H;��H;��H;i�H;�H;��H;K�H;�H;ۥH;�H;��H;��H;`�H;��H;��H;      V�H;��H;t�H;��H;��H;�H;��H;z�H;��H;�H;|�H;�H;��H;��H;S�H;p�H;<�H;��H;g�H;��H;��H;��H;>�H;x�H;��H;��H;x�H;B�H;��H;8�H;��H;��H;�H;M�H;m�H;y�H;��H;y�H;m�H;M�H;�H;��H;��H;8�H;��H;B�H;x�H;��H;��H;x�H;>�H;��H;��H;��H;g�H;��H;<�H;p�H;S�H;��H;��H;�H;|�H;�H;��H;z�H;��H;�H;��H;��H;t�H;��H;      �H;5�H;ֱH;��H;e�H;U�H;��H;�H;��H;f�H;P�H;@�H;�H;��H;��H;�H;��H;��H;�H;��H;��H;��H;G�H;t�H;��H;f�H;�H;��H;�H;��H;��H;�H;V�H;m�H;u�H;��H;��H;��H;u�H;m�H;V�H;�H;��H;��H;�H;��H;�H;f�H;��H;t�H;G�H;��H;��H;��H;�H;��H;��H;�H;��H;��H;�H;@�H;P�H;f�H;��H;�H;��H;U�H;e�H;��H;ֱH;5�H;      �H;M�H;ݷH;ǸH;'�H;»H;��H;ʿH;�H;��H;�H;��H;�H;��H;�H;R�H;��H;��H;Z�H;�H;��H;��H;�H;
�H;��H;��H;d�H;��H;V�H;��H;��H;C�H;l�H;y�H;��H;��H;��H;��H;��H;y�H;l�H;C�H;��H;��H;V�H;��H;d�H;��H;��H;
�H;�H;��H;��H;�H;Z�H;��H;��H;R�H;�H;��H;�H;��H;�H;��H;�H;ʿH;��H;»H;'�H;ǸH;ݷH;M�H;      ��H;B�H;عH;��H;��H;��H;M�H;X�H;u�H;��H;3�H;��H;=�H;��H;��H;9�H;9�H;'�H;��H;|�H;��H;%�H;@�H;Q�H;�H;��H;��H;#�H;b�H;��H;�H;5�H;7�H;��H;��H;��H;��H;��H;��H;��H;7�H;5�H;�H;��H;b�H;#�H;��H;��H;�H;Q�H;@�H;%�H;��H;|�H;��H;'�H;9�H;9�H;��H;��H;=�H;��H;3�H;��H;u�H;X�H;M�H;��H;��H;��H;عH;B�H;      �H;M�H;ݷH;ǸH;'�H;»H;��H;ʿH;�H;��H;�H;��H;�H;��H;�H;R�H;��H;��H;Z�H;�H;��H;��H;�H;
�H;��H;��H;d�H;��H;V�H;��H;��H;C�H;l�H;y�H;��H;��H;��H;��H;��H;y�H;l�H;C�H;��H;��H;V�H;��H;d�H;��H;��H;
�H;�H;��H;��H;�H;Z�H;��H;��H;R�H;�H;��H;�H;��H;�H;��H;�H;ʿH;��H;»H;'�H;ǸH;ݷH;M�H;      �H;5�H;ֱH;��H;e�H;U�H;��H;�H;��H;f�H;P�H;@�H;�H;��H;��H;�H;��H;��H;�H;��H;��H;��H;G�H;t�H;��H;f�H;�H;��H;�H;��H;��H;�H;V�H;m�H;u�H;��H;��H;��H;u�H;m�H;V�H;�H;��H;��H;�H;��H;�H;f�H;��H;t�H;G�H;��H;��H;��H;�H;��H;��H;�H;��H;��H;�H;@�H;P�H;f�H;��H;�H;��H;U�H;e�H;��H;ֱH;5�H;      V�H;��H;t�H;��H;��H;�H;��H;z�H;��H;�H;|�H;�H;��H;��H;S�H;p�H;<�H;��H;g�H;��H;��H;��H;>�H;x�H;��H;��H;x�H;B�H;��H;8�H;��H;��H;�H;M�H;m�H;y�H;��H;y�H;m�H;M�H;�H;��H;��H;8�H;��H;B�H;x�H;��H;��H;x�H;>�H;��H;��H;��H;g�H;��H;<�H;p�H;S�H;��H;��H;�H;|�H;�H;��H;z�H;��H;�H;��H;��H;t�H;��H;      M�H;��H;��H;`�H;��H;��H;�H;ۥH;�H;K�H;��H;�H;i�H;��H;��H;��H;l�H;��H;��H;��H;�H;e�H;U�H;��H;b�H;��H;��H;��H;A�H;��H;2�H;��H;�H;�H;V�H;l�H;7�H;l�H;V�H;�H;�H;��H;2�H;��H;A�H;��H;��H;��H;b�H;��H;U�H;e�H;�H;��H;��H;��H;l�H;��H;��H;��H;i�H;�H;��H;K�H;�H;ۥH;�H;��H;��H;`�H;��H;��H;      �H;��H;��H;�H;/�H;׊H;&�H;�H;]�H;��H;��H;��H;@�H;��H;�H;�H;��H;��H;��H;d�H;~�H;F�H;��H;��H;��H;�H;t�H;��H;��H;1�H;��H;C�H;��H;��H;�H;C�H;5�H;C�H;�H;��H;��H;C�H;��H;1�H;��H;��H;t�H;�H;��H;��H;��H;F�H;~�H;d�H;��H;��H;��H;�H;�H;��H;@�H;��H;��H;��H;]�H;�H;&�H;׊H;/�H;�H;��H;��H;      �aH;�bH;|dH;bgH;}kH;fpH;%vH;�|H;y�H;��H;�H;��H;�H;+�H;0�H;��H;��H;-�H;(�H;��H;��H;Q�H;d�H;�H;c�H;k�H;*�H;q�H;�H;w�H;I�H;��H;2�H;��H;��H;��H;�H;��H;��H;��H;2�H;��H;I�H;w�H;�H;q�H;*�H;k�H;c�H;�H;d�H;Q�H;��H;��H;(�H;-�H;��H;��H;0�H;+�H;�H;��H;�H;��H;y�H;�|H;%vH;fpH;}kH;bgH;|dH;�bH;      �9H;�:H;=H;�@H;2FH;�LH;�TH; ]H;>fH;�oH;�yH;��H;F�H;��H;��H;�H;�H;-�H;��H;��H;��H;)�H;4�H;��H;��H;)�H;5�H;��H;V�H;��H;w�H;1�H;��H;8�H;��H;��H;��H;��H;��H;8�H;��H;1�H;w�H;��H;V�H;��H;5�H;)�H;��H;��H;4�H;)�H;��H;��H;��H;-�H;�H;�H;��H;��H;F�H;��H;�yH;�oH;>fH; ]H;�TH;�LH;2FH;�@H;=H;�:H;      {H;hH;�
H;�H;�H;GH;8)H;e4H;o@H;MH;ZH;gH;�sH;<�H;��H;��H;ѠH;E�H;ҲH;J�H;��H;��H;�H;c�H;�H;$�H;��H;�H;��H;V�H;�H;��H;A�H;��H;�H;V�H;b�H;V�H;�H;��H;A�H;��H;�H;V�H;��H;�H;��H;$�H;�H;c�H;�H;��H;��H;J�H;ҲH;E�H;ѠH;��H;��H;<�H;�sH;gH;ZH;MH;o@H;e4H;8)H;GH;�H;�H;�
H;hH;      ��G;-�G;[�G;�G;�G;B�G;:�G;� H;hH;� H;�1H;XBH;
SH;DcH;�rH;�H;��H;�H;�H;ҮH;U�H;�H;;�H;��H;��H;��H;��H;��H;�H;��H;q�H;��H;��H;B�H;��H;��H;#�H;��H;��H;B�H;��H;��H;q�H;��H;�H;��H;��H;��H;��H;��H;;�H;�H;U�H;ҮH;�H;�H;��H;�H;�rH;DcH;
SH;XBH;�1H;� H;hH;� H;:�G;B�G;�G;�G;[�G;-�G;      �kG;nG;�tG;�~G;�G;}�G;��G;��G;��G;$�G;��G;�H;"*H;�>H;�RH;:eH;gvH;��H;ړH;<�H;U�H;�H;�H;@�H;=�H;H�H;e�H;��H;��H;5�H;*�H;t�H;��H;x�H;�H;d�H;��H;d�H;�H;x�H;��H;t�H;*�H;5�H;��H;��H;e�H;H�H;=�H;@�H;�H;�H;U�H;<�H;ړH;��H;gvH;:eH;�RH;�>H;"*H;�H;��G;$�G;��G;��G;��G;}�G;�G;�~G;�tG;nG;      ��F;��F;F�F;��F; G;�"G;�EG;�gG;φG;�G;��G;��G;h�G;�H;/+H;�BH;�XH; mH;�~H;z�H;q�H;��H;?�H;/�H;��H;�H;H�H;��H;$�H;)�H;k�H;�H;��H;��H;f�H;��H;��H;��H;f�H;��H;��H;�H;k�H;)�H;$�H;��H;H�H;�H;��H;/�H;?�H;��H;q�H;z�H;�~H; mH;�XH;�BH;/+H;�H;h�G;��G;��G;�G;φG;�gG;�EG;�"G; G;��F;F�F;��F;      ��D;��D;P
E;�ME;��E;2�E;[F;'�F;)�F;@:G;OlG;^�G;�G;��G;��G;�H;�4H;�MH;�dH;yH;��H;��H;�H;W�H;��H;��H;=�H;��H;�H;��H;c�H;��H;b�H;��H;��H;��H;�H;��H;��H;��H;b�H;��H;c�H;��H;�H;��H;=�H;��H;��H;W�H;�H;��H;��H;yH;�dH;�MH;�4H;�H;��G;��G;�G;^�G;OlG;@:G;)�F;'�F;[F;2�E;��E;�ME;P
E;��D;      VZ@;~@;�@;D�A;@PB;�0C;�D;��D;=�E;�KF;��F;:#G;jeG;�G;O�G;��G;�H;�(H;EH;�^H;
uH;�H;r�H;}�H;W�H;/�H;@�H;��H;c�H;��H;�H;��H;��H;x�H;t�H;
�H;Q�H;
�H;t�H;x�H;��H;��H;�H;��H;c�H;��H;@�H;/�H;W�H;}�H;r�H;�H;
uH;�^H;EH;�(H;�H;��G;O�G;�G;jeG;:#G;��F;�KF;=�E;��D;�D;�0C;@PB;D�A;�@;~@;      ��6;*7;��7;�M9;9	;;��<;��>;��@;B�B;�D;.AE;�"F;Z�F;�-G;%uG;�G;|�G;�G;�H;?H;�ZH;sH;V�H;r�H;�H;?�H;�H;;�H;�H;4�H;d�H;��H;U�H;>�H;G�H;�H;@�H;�H;G�H;>�H;U�H;��H;d�H;4�H;�H;;�H;�H;?�H;�H;r�H;V�H;sH;�ZH;?H;�H;�G;|�G;�G;%uG;�-G;Z�F;�"F;.AE;�D;B�B;��@;��>;��<;9	;;�M9;��7;*7;      ]�#;f$;�'&;��(;hh,;D_0;�~4;~8;:'<;)N?;+�A;��C;%NE;
LF;2�F;TG;z�G;�G;��G;�H;�;H;�YH;sH;�H;��H;��H;�H;�H;��H;)�H;Q�H;F�H;e�H;��H;��H;��H;%�H;��H;��H;��H;e�H;F�H;Q�H;)�H;��H;�H;�H;��H;��H;�H;sH;�YH;�;H;�H;��G;�G;z�G;TG;2�F;
LF;%NE;��C;+�A;)N?;:'<;~8;�~4;D_0;hh,;��(;�'&;f$;      �;P/;�w;��
;�8;v�;3� ;�_(;I�/;��5;}	;;%?;%5B;^D;`�E;��F;d7G;�G;�G;L�G;�H;�;H;�ZH;
uH;��H;q�H;U�H;U�H;��H;��H;��H;~�H;�H;��H;��H;��H;��H;��H;��H;��H;�H;~�H;��H;��H;��H;U�H;U�H;q�H;��H;
uH;�ZH;�;H;�H;L�G;�G;�G;d7G;��F;`�E;^D;%5B;%?;}	;;��5;I�/;�_(;3� ;v�;�8;��
;�w;P/;      ���:d��:�@�:���:
��:i��:7&�:�;��;Tf$;�=.;^#6;l'<;�~@; tC;�ZE;6F;]#G;fG;�G;L�G;�H;?H;�^H;yH;z�H;<�H;ҮH;J�H;��H;��H;d�H;��H;��H;��H;�H;|�H;�H;��H;��H;��H;d�H;��H;��H;J�H;ҮH;<�H;z�H;yH;�^H;?H;�H;L�G;�G;fG;]#G;6F;�ZE; tC;�~@;l'<;^#6;�=.;Tf$;��;�;7&�:i��:
��:���:�@�:d��:      %W� yƹ2p�d��6SX�94t,:裆:�ض:L�:�;��;6(&;�-1;,N9;=�>;�B;�
E;�bF;,G;fG;�G;��G;�H;EH;�dH;�~H;ړH;�H;ҲH;��H;(�H;��H;��H;g�H;�H;Z�H;��H;Z�H;�H;g�H;��H;��H;(�H;��H;ҲH;�H;ړH;�~H;�dH;EH;�H;��G;�G;fG;,G;�bF;�
E;�B;=�>;,N9;�-1;6(&;��;�;L�:�ض:裆:4t,:SX�9d��62p� yƹ      ��4��K/�"V�+,�E�˺�쀺vƹ�m9?nQ:=��: ��:4�;�;��,;�7;$�=;vPB;�D;�bF;]#G;�G;�G;�G;�(H;�MH; mH;��H;�H;E�H;-�H;-�H;��H;��H;��H;��H;��H;'�H;��H;��H;��H;��H;��H;-�H;-�H;E�H;�H;��H; mH;�MH;�(H;�G;�G;�G;]#G;�bF;�D;vPB;$�=;�7;��,;�;4�; ��:=��:?nQ:�m9vƹ�쀺E�˺+,�"V��K/�      �ͻ�Rɻ����!Ϩ�|-��p\c��$�h�˺P(�PM@9��k:���:;ƽ;��);.�5;��=;vPB;�
E;6F;d7G;z�G;|�G;�H;�4H;�XH;gvH;��H;ѠH;�H;��H;��H;l�H;<�H;��H;��H;9�H;��H;��H;<�H;l�H;��H;��H;�H;ѠH;��H;gvH;�XH;�4H;�H;|�G;z�G;d7G;6F;�
E;vPB;��=;.�5;��);ƽ;;���:��k:PM@9P(�h�˺�$�p\c�|-��!Ϩ������Rɻ      �J;���7�m9.����z&�W��&����L��h�4�]�ºOuƹ�P:N��:���:��;-�(;.�5;$�=;�B;�ZE;��F;TG;�G;��G;�H;�BH;:eH;�H;��H;�H;��H;�H;��H;p�H;�H;R�H;9�H;R�H;�H;p�H;��H;�H;��H;�H;��H;�H;:eH;�BH;�H;��G;�G;TG;��F;�ZE;�B;$�=;.�5;-�(;��;���:N��:�P:Ouƹ]�ºh�4��L��&���W��z&����m9.���7�      �䙼�_��=��>y��);k��I��$�Y� �f���%�|��_$T�}Z�9qA�:���:��;��);�7;=�>; tC;`�E;2�F;%uG;O�G;��G;/+H;�RH;�rH;��H;��H;0�H;�H;��H;S�H;��H;�H;��H;�H;��H;S�H;��H;�H;0�H;��H;��H;�rH;�RH;/+H;��G;O�G;%uG;2�F;`�E; tC;=�>;�7;��);��;���:qA�:}Z�9_$T��%�|�f���Y� ��$��I�);k�>y��=���_��      \��l�鼟߼μ�!��v
��>y��T��!�5�軈ۙ�2K/�����wm9qA�:���:ƽ;��,;,N9;�~@;^D;
LF;�-G;�G;��G;�H;�>H;DcH;<�H;��H;+�H;��H;��H;��H;��H;��H;��H;��H;��H;��H;��H;��H;+�H;��H;<�H;DcH;�>H;�H;��G;�G;�-G;
LF;^D;�~@;,N9;��,;ƽ;���:qA�:wm9����2K/��ۙ�5���!�T�>y��v
���!��μ�߼l��      |�/�-�:.%�������T���Ǽ����(�{��J;��C��Ψ�	O:�����}Z�9N��:;�;�-1;l'<;%5B;%NE;Z�F;jeG;�G;h�G;"*H;
SH;�sH;F�H;�H;@�H;i�H;��H;�H;�H;=�H;�H;�H;��H;i�H;@�H;�H;F�H;�sH;
SH;"*H;h�G;�G;jeG;Z�F;%NE;%5B;l'<;�-1;�;;N��:}Z�9����	O:��Ψ��C��J;�(�{�������ǼT��������:.%�-�       @{�`w�Al��yZ� �C�8g*����k���!��-O���I�|��Ψ�2K/�_$T��P:���:4�;6(&;^#6;%?;��C;�"F;:#G;^�G;��G;�H;XBH;gH;��H;��H;��H;�H;�H;@�H;��H;��H;��H;@�H;�H;�H;��H;��H;��H;gH;XBH;�H;��G;^�G;:#G;�"F;��C;%?;^#6;6(&;4�;���:�P:_$T�2K/��Ψ�|��I�-O���!��k�鼇��8g*� �C��yZ�Al�`w�      �b������kƣ�ss���ɇ�Al�G�Ơ"�D� ��`ļ6���I��C��ۙ��Ouƹ��k: ��:��;�=.;}	;;+�A;.AE;��F;OlG;��G;��G;�1H;ZH;�yH;�H;��H;��H;|�H;P�H;�H;3�H;�H;P�H;|�H;��H;��H;�H;�yH;ZH;�1H;��G;��G;OlG;��F;.AE;+�A;}	;;�=.;��; ��:��k:Ouƹ��ۙ��C��I�6���`ļD� �Ơ"�G�Al��ɇ�ss��kƣ�����      U�뽱��?ݽa2̽gж����������yZ�-�����`ļ-O���J;�5��%�|�]�ºPM@9=��:�;Tf$;��5;)N?;�D;�KF;@:G;�G;$�G;� H;MH;�oH;��H;��H;K�H;�H;f�H;��H;��H;��H;f�H;�H;K�H;��H;��H;�oH;MH;� H;$�G;�G;@:G;�KF;�D;)N?;��5;Tf$;�;=��:PM@9]�º%�|�5�軃J;�-O���`ļ���-��yZ���������gж�a2̽?ݽ���      0,����Z���z�$vϽ�b��I��.]a�-�D� ��!��(�{��!�f���h�4�P(�?nQ:L�:��;I�/;:'<;B�B;=�E;)�F;φG;��G;hH;o@H;>fH;y�H;]�H;�H;��H;��H;�H;u�H;�H;��H;��H;�H;]�H;y�H;>fH;o@H;hH;��G;φG;)�F;=�E;B�B;:'<;I�/;��;L�:?nQ:P(�h�4�f����!�(�{��!��D� �-�.]a�I���b��$vϽ�z���Z���      �G�I�C�g$:��J+�����?ݽ4���I���yZ�Ơ"�k�鼢���T�Y� ��L��h�˺�m9�ض:�;�_(;~8;��@;��D;'�F;�gG;��G;� H;e4H; ]H;�|H;�H;ۥH;z�H;�H;ʿH;X�H;ʿH;�H;z�H;ۥH;�H;�|H; ]H;e4H;� H;��G;�gG;'�F;��D;��@;~8;�_(;�;�ض:�m9h�˺�L��Y� �T�����k��Ơ"��yZ�I��4���?ݽ�����J+�g$:�I�C�      �zx��8t���g���T��G=�Z#��5�?ݽ�b������G������Ǽ>y���$�&����$�vƹ裆:7&�:3� ;�~4;��>;�D;[F;�EG;��G;:�G;8)H;�TH;%vH;&�H;�H;��H;��H;��H;M�H;��H;��H;��H;�H;&�H;%vH;�TH;8)H;:�G;��G;�EG;[F;�D;��>;�~4;3� ;7&�:裆:vƹ�$�&����$�>y����Ǽ���G������b��?ݽ�5�Z#��G=���T���g��8t�      Ы�����3a��	����c�J�C�Z#���$vϽ����Al�8g*�T��v
���I�W��p\c��쀺4t,:i��:v�;D_0;��<;�0C;2�E;�"G;}�G;B�G;GH;�LH;fpH;׊H;��H;�H;U�H;»H;��H;»H;U�H;�H;��H;׊H;fpH;�LH;GH;B�G;}�G;�"G;2�E;�0C;��<;D_0;v�;i��:4t,:�쀺p\c�W�軞I�v
��T��8g*�Al�����$vϽ��Z#�J�C��c�	���3a�����      K*��I����Ƥ�Ы���/���c��G=����z�gж��ɇ� �C�����!��);k�z&�|-��E�˺SX�9
��:�8;hh,;9	;;@PB;��E; G;�G;�G;�H;2FH;}kH;/�H;��H;��H;e�H;'�H;��H;'�H;e�H;��H;��H;/�H;}kH;2FH;�H;�G;�G; G;��E;@PB;9	;;hh,;�8;
��:SX�9E�˺|-��z&�);k��!����� �C��ɇ�gж��z����G=��c��/��Ы���Ƥ�I���      ��ɾZ�ž�*��Sת�Ы��	�����T��J+��a2̽ss���yZ����μ>y�����!Ϩ�+,�d��6���:��
;��(;�M9;D�A;�ME;��F;�~G;�G;�H;�@H;bgH;�H;`�H;��H;��H;ǸH;��H;ǸH;��H;��H;`�H;�H;bgH;�@H;�H;�G;�~G;��F;�ME;D�A;�M9;��(;��
;���:d��6+,�!Ϩ����>y��μ����yZ�ss��a2̽��J+���T�	���Ы��Sת��*��Z�ž      0_ݾ�:پ�V;�*���Ƥ�3a����g�g$:��Z�?ݽkƣ�Al�:.%��߼=��m9.�����"V�2p��@�:�w;�'&;��7;�@;P
E;F�F;�tG;[�G;�
H;=H;|dH;��H;��H;t�H;ֱH;ݷH;عH;ݷH;ֱH;t�H;��H;��H;|dH;=H;�
H;[�G;�tG;F�F;P
E;�@;��7;�'&;�w;�@�:2p�"V�����m9.�=���߼:.%�Al�kƣ�?ݽ�Z�g$:���g�3a���Ƥ��*���V;�:پ      �]����:پZ�žI�������8t�I�C�����罽���`w�-�l���_����7��Rɻ�K/� yƹd��:P/;f$;*7;~@;��D;��F;nG;-�G;hH;�:H;�bH;��H;��H;��H;5�H;M�H;B�H;M�H;5�H;��H;��H;��H;�bH;�:H;hH;-�G;nG;��F;��D;~@;*7;f$;P/;d��: yƹ�K/��Rɻ��7��_��l��-�`w����������I�C��8t����I���Z�ž�:پ��      3F�/h��ǰ�3Vھ�������~���S��#��o��S��Q₽�6�-���<y��FB��Eֻ^A?��	�Y�:���:�";�36;�@;��D;��F;�mG;&�G;>H;:?H;fH;w�H;P�H;��H;��H;�H;�H;�H;��H;��H;P�H;w�H;fH;:?H;>H;&�G;�mG;��F;��D;�@;�36;�";���:Y�:�	�^A?��EֻFB�<y��-����6�Q₽S���o���#��S��~��������3Vھǰ�/h��      /h���b���쾅*־�v������)�� �O�6� ��r�r���؀��3����ݜ��>��ѻ��9�����n�:�$ ;�L#;˃6;�@@;C�D;�F;<pG;��G;TH;@H;�fH;�H;��H;�H;>�H;�H;��H;�H;>�H;�H;��H;�H;�fH;@H;TH;��G;<pG;�F;C�D;�@@;˃6;�L#;�$ ;�n�:�����9��ѻ�>�ݜ�����3��؀��r���r�6� � �O��)������v���*־�쾼b��      ǰ�쾐�޾5ʾ/;���:����v��E�A'���L����u�X�+�aW缨A��r�4�m�Ļ�8)��j��W�:�;�%;kk7;g�@;B�D;4�F;wG;��G;vH;cBH;YhH;B�H;��H;ƩH;�H;��H;��H;��H;�H;ƩH;��H;B�H;YhH;cBH;vH;��G;wG;4�F;B�D;g�@;kk7;�%;�;W�:�j���8)�m�Ļr�4��A��aW�X�+���u�L����A'��E���v��:��/;��5ʾ��޾��      3Vھ�*־5ʾT��������M���9b��5���}�սn���Xc�ݟ���ռ�I��$�$�4T���Z�
_����:��;��';��8;^QA;�8E;��F;�G;%�G;�H;.FH;@kH;u�H;[�H;�H;�H;��H;t�H;��H;�H;�H;[�H;u�H;@kH;.FH;�H;%�G;�G;��F;�8E;^QA;��8;��';��;��:
_���Z�4T��$�$��I����ռݟ��Xc�n��}�ս���5��9b��M������T���5ʾ�*־      ���v��/;������:P���r�U�H�6� ��~��@������Q�K�<��վ���s�F��_�~ܺ3u9�%�:��;��+;��:;"B;��E;,�F;��G;�G;nH;[KH;(oH;k�H;��H;ƬH;_�H;��H;��H;��H;_�H;ƬH;��H;k�H;(oH;[KH;nH;�G;��G;,�F;��E;"B;��:;��+;��;�%�:3u9~ܺ_�F����s��վ�<�Q�K�����@���~��6� �U�H��r�:P������/;���v��      ��������:���M���r� �O��",�<�
��gٽKĥ�|�u�K1�(����Τ�m�P��Z�q.o�jp���:մ�:|P;��/;��<;G
C;f�E;� G;_�G;6�G;�$H;�QH;�sH;%�H;f�H;��H;+�H;{�H;&�H;{�H;+�H;��H;f�H;%�H;�sH;�QH;�$H;6�G;_�G;� G;f�E;G
C;��<;��/;|P;մ�:�:jp��q.o��Z�m�P��Τ�(���K1�|�u�Kĥ��gٽ<�
��",� �O��r��M���:�����      �~���)����v��9b�U�H��",�0Z���S��X^��e�N�{����μ�I���%+�ښ����.������i~:���:�l;A�3;��>;�C;�OF;�EG;|�G;"�G;�.H;'YH;�yH;q�H;��H;��H;F�H;K�H;��H;K�H;F�H;��H;��H;q�H;�yH;'YH;�.H;"�G;|�G;�EG;�OF;�C;��>;A�3;�l;���:�i~:������.�ښ���%+��I����μ{��e�N�X^��S����0Z��",�U�H��9b���v��)��      �S� �O��E��5�6� �<�
���|9��l���Xc���(����߈��Z�[����nݎ�ܺO99���:��	;�c';��7;��@;��D;/�F;biG;��G;�H;�9H;gaH;�H;0�H;P�H;g�H;��H;Y�H;��H;Y�H;��H;g�H;P�H;0�H;�H;gaH;�9H;�H;��G;biG;/�F;��D;��@;��7;�c';��	;���:O99ܺnݎ����Z�[�߈�������(��Xc�l��|9����<�
�6� ��5��E� �O�      �#�6� �A'����~���gٽS��l���j��3�ji��վ�T����(�P�Ļ+A?���B�8�@:[�:�P;w�.;Q�;;�sB;\�E;��F;l�G;'�G;H;�EH;KjH;��H;H�H;.�H;��H;0�H;��H;�H;��H;0�H;��H;.�H;H�H;��H;KjH;�EH;H;'�G;l�G;��F;\�E;�sB;Q�;;w�.;�P;[�:8�@:��B�+A?�P�Ļ�(�T����վ�ji��3��j�l��S���gٽ�~����A'�6� �      �o���r���}�ս@��Kĥ�X^���Xc��3���	���˼t]��FB��Z򻆜��CӺE��8�:{�;RM#;�<5;x?;��C;�?F;K9G;-�G;M�G;d&H;�QH;�sH;ۍH;��H;H�H;кH;��H;��H;a�H;��H;��H;кH;H�H;��H;ۍH;�sH;�QH;d&H;M�G;-�G;K9G;�?F;��C;x?;�<5;RM#;{�;�:E��8CӺ�����Z�FB�t]����˼��	��3��Xc�X^��Kĥ�@��}�ս���r�      S���r��L��n������|�u�e�N���(�ji���˼�A��b�P�=s��|������\:��:�;�m-;F�:;O�A;�+E;��F;mnG;,�G;�H;�6H;k^H;0}H;�H;&�H;��H;/�H;��H;Z�H;��H;Z�H;��H;/�H;��H;&�H;�H;0}H;k^H;�6H;�H;,�G;mnG;��F;�+E;O�A;F�:;�m-;�;��:�\:����|��=s�b�P��A����˼ji���(�e�N�|�u�����n��L���r��      Q₽�؀���u��Xc�Q�K�K1�{�����վ�t]��b�P�l��T��g�9���o�o2�9�%�:��	;�%;��5;�>;��C;	F;� G;ޙG;�G;pH;�GH;�jH;ʆH;s�H;��H;̸H;��H;l�H;��H;��H;��H;l�H;��H;̸H;��H;s�H;ʆH;�jH;�GH;pH;�G;ޙG;� G;	F;��C;�>;��5;�%;��	;�%�:o2�9��o�g�9�T��l��b�P�t]���վ����{��K1�Q�K��Xc���u��؀�      �6��3�X�+�ݟ�<�(�����μ߈��T���FB�=s�T����D��{���8u92q�:���:�X;at0;T�;;1B;D9E;/�F;:gG;�G;=�G;�/H;�WH;SwH;G�H;��H;$�H;�H; �H;2�H;I�H;S�H;I�H;2�H; �H;�H;$�H;��H;G�H;SwH;�WH;�/H;=�G;�G;:gG;/�F;D9E;1B;T�;;at0;�X;���:2q�:�8u9�{����D�T��=s�FB�T���߈����μ(���<�ݟ�X�+��3�      -������aW缐�ռ�վ��Τ��I��Z�[��(��Z�g�9��{���99�W�:�W�:�P;�,;�8;�@@;ZAD;�?F;�+G;ÛG;��G;�H;�CH;HgH;W�H;y�H;��H;�H;>�H;:�H;��H;��H;��H;��H;��H;:�H;>�H;�H;��H;y�H;W�H;HgH;�CH;�H;��G;ÛG;�+G;�?F;ZAD;�@@;�8;�,;�P;�W�:�W�:�99�{��g�9���Z��(�Z�[��I���Τ��վ���ռaW缧��      <y��ݜ��A���I����s�m�P��%+����P�Ļ����|���o��8u9�W�::+�:�;^);8�6;ذ>;�OC;��E;:�F;�wG;a�G;� H;�0H;@WH;*vH;ԎH;9�H;$�H;��H;5�H;^�H;��H;�H;��H;�H;��H;^�H;5�H;��H;$�H;9�H;ԎH;*vH;@WH;�0H;� H;a�G;�wG;:�F;��E;�OC;ذ>;8�6;^);�;:+�:�W�:�8u9��o�|�����P�Ļ����%+�m�P���s��I���A��ݜ�      FB��>�r�4�$�$�F���Z�ښ��nݎ�+A?�CӺ����o2�92q�:�W�:�;E�';�<5;֜=;[�B;jFE;��F;�TG;Z�G;�G;�H;�GH;9iH;�H;��H;g�H;T�H;f�H;��H;[�H;(�H;6�H;��H;6�H;(�H;[�H;��H;f�H;T�H;g�H;��H;�H;9iH;�GH;�H;�G;Z�G;�TG;��F;jFE;[�B;֜=;�<5;E�';�;�W�:2q�:o2�9����CӺ+A?�nݎ�ښ���Z�F��$�$�r�4��>�      �Eֻ�ѻm�Ļ4T��_�q.o���.�ܺ��B�E��8�\:�%�:���:�P;^);�<5;L:=;x"B;��D;!uF;,6G;��G;��G;�H;�9H;:]H;�yH;�H;��H;�H;'�H;��H;u�H;6�H;��H;B�H;��H;B�H;��H;6�H;u�H;��H;'�H;�H;��H;�H;�yH;:]H;�9H;�H;��G;��G;,6G;!uF;��D;x"B;L:=;�<5;^);�P;���:�%�:�\:E��8��B�ܺ��.�q.o�_�4T��m�Ļ�ѻ      ^A?���9��8)��Z�~ܺjp������O998�@:�:��:��	;�X;�,;8�6;֜=;x"B; �D;�WF;!G;��G;T�G;�H; .H;�RH;�pH;�H;ԜH;��H;׸H;��H;��H;��H;��H;��H;0�H;��H;0�H;��H;��H;��H;��H;��H;׸H;��H;ԜH;�H;�pH;�RH; .H;�H;T�G;��G;!G;�WF; �D;x"B;֜=;8�6;�,;�X;��	;��:�:8�@:O99����jp��~ܺ�Z��8)���9�      �	�����j��
_��3u9�:�i~:���:[�:{�;�;�%;at0;�8;ذ>;[�B;��D;�WF;tG;��G;��G;��G;%H;.JH;�hH;�H;��H;T�H;��H;�H;x�H;��H;��H;H�H;��H;��H;i�H;��H;��H;H�H;��H;��H;x�H;�H;��H;T�H;��H;�H;�hH;.JH;%H;��G;��G;��G;tG;�WF;��D;[�B;ذ>;�8;at0;�%;�;{�;[�:���:�i~:�:3u9
_���j�����      Y�:�n�:W�:��:�%�:մ�:���:��	;�P;RM#;�m-;��5;T�;;�@@;�OC;jFE;!uF;!G;��G;�G;F�G;xH;7DH;�bH;e|H;��H;ԢH;��H;ۻH;��H;��H;B�H;j�H;e�H;^�H;��H;��H;��H;^�H;e�H;j�H;B�H;��H;��H;ۻH;��H;ԢH;��H;e|H;�bH;7DH;xH;F�G;�G;��G;!G;!uF;jFE;�OC;�@@;T�;;��5;�m-;RM#;�P;��	;���:մ�:�%�:��:W�:�n�:      ���:�$ ;�;��;��;|P;�l;�c';w�.;�<5;F�:;�>;1B;ZAD;��E;��F;,6G;��G;��G;F�G;�H;AH;0_H;mxH;��H;<�H;m�H;��H;b�H;��H;��H;F�H;��H;S�H;�H;��H;[�H;��H;�H;S�H;��H;F�H;��H;��H;b�H;��H;m�H;<�H;��H;mxH;0_H;AH;�H;F�G;��G;��G;,6G;��F;��E;ZAD;1B;�>;F�:;�<5;w�.;�c';�l;|P;��;��;�;�$ ;      �";�L#;�%;��';��+;��/;A�3;��7;Q�;;x?;O�A;��C;D9E;�?F;:�F;�TG;��G;T�G;��G;xH;AH;�]H;hvH;9�H;��H;��H;��H;E�H;�H;7�H;1�H;��H;��H;��H;x�H;U�H;��H;U�H;x�H;��H;��H;��H;1�H;7�H;�H;E�H;��H;��H;��H;9�H;hvH;�]H;AH;xH;��G;T�G;��G;�TG;:�F;�?F;D9E;��C;O�A;x?;Q�;;��7;A�3;��/;��+;��';�%;�L#;      �36;˃6;kk7;��8;��:;��<;��>;��@;�sB;��C;�+E;	F;/�F;�+G;�wG;Z�G;��G;�H;%H;7DH;0_H;hvH;O�H;P�H;h�H;��H;��H;��H;��H;�H;=�H;Q�H;��H;m�H;��H;{�H;��H;{�H;��H;m�H;��H;Q�H;=�H;�H;��H;��H;��H;��H;h�H;P�H;O�H;hvH;0_H;7DH;%H;�H;��G;Z�G;�wG;�+G;/�F;	F;�+E;��C;�sB;��@;��>;��<;��:;��8;kk7;˃6;      �@;�@@;g�@;^QA;"B;G
C;�C;��D;\�E;�?F;��F;� G;:gG;ÛG;a�G;�G;�H; .H;.JH;�bH;mxH;9�H;P�H;ܨH;#�H;��H;��H;��H;"�H;\�H;��H;[�H;K�H;��H;��H;i�H;��H;i�H;��H;��H;K�H;[�H;��H;\�H;"�H;��H;��H;��H;#�H;ܨH;P�H;9�H;mxH;�bH;.JH; .H;�H;�G;a�G;ÛG;:gG;� G;��F;�?F;\�E;��D;�C;G
C;"B;^QA;g�@;�@@;      ��D;C�D;B�D;�8E;��E;f�E;�OF;/�F;��F;K9G;mnG;ޙG;�G;��G;� H;�H;�9H;�RH;�hH;e|H;��H;��H;h�H;#�H;U�H;��H;@�H;~�H;��H;9�H;��H;�H;��H;��H;��H;.�H;r�H;.�H;��H;��H;��H;�H;��H;9�H;��H;~�H;@�H;��H;U�H;#�H;h�H;��H;��H;e|H;�hH;�RH;�9H;�H;� H;��G;�G;ޙG;mnG;K9G;��F;/�F;�OF;f�E;��E;�8E;B�D;C�D;      ��F;�F;4�F;��F;,�F;� G;�EG;biG;l�G;-�G;,�G;�G;=�G;�H;�0H;�GH;:]H;�pH;�H;��H;<�H;��H;��H;��H;��H;�H;/�H;k�H;��H;��H;��H;��H;��H;��H;��H;��H;�H;��H;��H;��H;��H;��H;��H;��H;��H;k�H;/�H;�H;��H;��H;��H;��H;<�H;��H;�H;�pH;:]H;�GH;�0H;�H;=�G;�G;,�G;-�G;l�G;biG;�EG;� G;,�F;��F;4�F;�F;      �mG;<pG;wG;�G;��G;_�G;|�G;��G;'�G;M�G;�H;pH;�/H;�CH;@WH;9iH;�yH;�H;��H;ԢH;m�H;��H;��H;��H;@�H;/�H;N�H;��H;h�H;��H;X�H;��H;��H;��H;;�H;��H;��H;��H;;�H;��H;��H;��H;X�H;��H;h�H;��H;N�H;/�H;@�H;��H;��H;��H;m�H;ԢH;��H;�H;�yH;9iH;@WH;�CH;�/H;pH;�H;M�G;'�G;��G;|�G;_�G;��G;�G;wG;<pG;      &�G;��G;��G;%�G;�G;6�G;"�G;�H;H;d&H;�6H;�GH;�WH;HgH;*vH;�H;�H;ԜH;T�H;��H;��H;E�H;��H;��H;~�H;k�H;��H;G�H;��H;L�H;��H;��H;��H;k�H;��H;�H; �H;�H;��H;k�H;��H;��H;��H;L�H;��H;G�H;��H;k�H;~�H;��H;��H;E�H;��H;��H;T�H;ԜH;�H;�H;*vH;HgH;�WH;�GH;�6H;d&H;H;�H;"�G;6�G;�G;%�G;��G;��G;      >H;TH;vH;�H;nH;�$H;�.H;�9H;�EH;�QH;k^H;�jH;SwH;W�H;ԎH;��H;��H;��H;��H;ۻH;b�H;�H;��H;"�H;��H;��H;h�H;��H;-�H;��H;��H;��H;b�H;��H;L�H;�H;��H;�H;L�H;��H;b�H;��H;��H;��H;-�H;��H;h�H;��H;��H;"�H;��H;�H;b�H;ۻH;��H;��H;��H;��H;ԎH;W�H;SwH;�jH;k^H;�QH;�EH;�9H;�.H;�$H;nH;�H;vH;TH;      :?H;@H;cBH;.FH;[KH;�QH;'YH;gaH;KjH;�sH;0}H;ʆH;G�H;y�H;9�H;g�H;�H;׸H;�H;��H;��H;7�H;�H;\�H;9�H;��H;��H;L�H;��H;��H;��H;n�H;�H;T�H;��H;��H;��H;��H;��H;T�H;�H;n�H;��H;��H;��H;L�H;��H;��H;9�H;\�H;�H;7�H;��H;��H;�H;׸H;�H;g�H;9�H;y�H;G�H;ʆH;0}H;�sH;KjH;gaH;'YH;�QH;[KH;.FH;cBH;@H;      fH;�fH;YhH;@kH;(oH;�sH;�yH;�H;��H;ۍH;�H;s�H;��H;��H;$�H;T�H;'�H;��H;x�H;��H;��H;1�H;=�H;��H;��H;��H;X�H;��H;��H;��H;t�H;�H;h�H;��H;��H;�H;0�H;�H;��H;��H;h�H;�H;t�H;��H;��H;��H;X�H;��H;��H;��H;=�H;1�H;��H;��H;x�H;��H;'�H;T�H;$�H;��H;��H;s�H;�H;ۍH;��H;�H;�yH;�sH;(oH;@kH;YhH;�fH;      w�H;�H;B�H;u�H;k�H;%�H;q�H;0�H;H�H;��H;&�H;��H;$�H;�H;��H;f�H;��H;��H;��H;B�H;F�H;��H;Q�H;[�H;�H;��H;��H;��H;��H;n�H;�H;z�H;��H; �H;,�H;J�H;I�H;J�H;,�H; �H;��H;z�H;�H;n�H;��H;��H;��H;��H;�H;[�H;Q�H;��H;F�H;B�H;��H;��H;��H;f�H;��H;�H;$�H;��H;&�H;��H;H�H;0�H;q�H;%�H;k�H;u�H;B�H;�H;      P�H;��H;��H;[�H;��H;f�H;��H;P�H;.�H;H�H;��H;̸H;�H;>�H;5�H;��H;u�H;��H;��H;j�H;��H;��H;��H;K�H;��H;��H;��H;��H;b�H;�H;h�H;��H;	�H;:�H;X�H;��H;��H;��H;X�H;:�H;	�H;��H;h�H;�H;b�H;��H;��H;��H;��H;K�H;��H;��H;��H;j�H;��H;��H;u�H;��H;5�H;>�H;�H;̸H;��H;H�H;.�H;P�H;��H;f�H;��H;[�H;��H;��H;      ��H;�H;ƩH;�H;ƬH;��H;��H;g�H;��H;кH;/�H;��H; �H;:�H;^�H;[�H;6�H;��H;H�H;e�H;S�H;��H;m�H;��H;��H;��H;��H;k�H;��H;T�H;��H; �H;:�H;u�H;��H;��H;��H;��H;��H;u�H;:�H; �H;��H;T�H;��H;k�H;��H;��H;��H;��H;m�H;��H;S�H;e�H;H�H;��H;6�H;[�H;^�H;:�H; �H;��H;/�H;кH;��H;g�H;��H;��H;ƬH;�H;ƩH;�H;      ��H;>�H;�H;�H;_�H;+�H;F�H;��H;0�H;��H;��H;l�H;2�H;��H;��H;(�H;��H;��H;��H;^�H;�H;x�H;��H;��H;��H;��H;;�H;��H;L�H;��H;��H;,�H;X�H;��H;��H;��H;��H;��H;��H;��H;X�H;,�H;��H;��H;L�H;��H;;�H;��H;��H;��H;��H;x�H;�H;^�H;��H;��H;��H;(�H;��H;��H;2�H;l�H;��H;��H;0�H;��H;F�H;+�H;_�H;�H;�H;>�H;      �H;�H;��H;��H;��H;{�H;K�H;Y�H;��H;��H;Z�H;��H;I�H;��H;�H;6�H;B�H;0�H;��H;��H;��H;U�H;{�H;i�H;.�H;��H;��H;�H;�H;��H;�H;J�H;��H;��H;��H;��H;��H;��H;��H;��H;��H;J�H;�H;��H;�H;�H;��H;��H;.�H;i�H;{�H;U�H;��H;��H;��H;0�H;B�H;6�H;�H;��H;I�H;��H;Z�H;��H;��H;Y�H;K�H;{�H;��H;��H;��H;�H;      �H;��H;��H;t�H;��H;&�H;��H;��H;�H;a�H;��H;��H;S�H;��H;��H;��H;��H;��H;i�H;��H;[�H;��H;��H;��H;r�H;�H;��H; �H;��H;��H;0�H;I�H;��H;��H;��H;��H;��H;��H;��H;��H;��H;I�H;0�H;��H;��H; �H;��H;�H;r�H;��H;��H;��H;[�H;��H;i�H;��H;��H;��H;��H;��H;S�H;��H;��H;a�H;�H;��H;��H;&�H;��H;t�H;��H;��H;      �H;�H;��H;��H;��H;{�H;K�H;Y�H;��H;��H;Z�H;��H;I�H;��H;�H;6�H;B�H;0�H;��H;��H;��H;U�H;{�H;i�H;.�H;��H;��H;�H;�H;��H;�H;J�H;��H;��H;��H;��H;��H;��H;��H;��H;��H;J�H;�H;��H;�H;�H;��H;��H;.�H;i�H;{�H;U�H;��H;��H;��H;0�H;B�H;6�H;�H;��H;I�H;��H;Z�H;��H;��H;Y�H;K�H;{�H;��H;��H;��H;�H;      ��H;>�H;�H;�H;_�H;+�H;F�H;��H;0�H;��H;��H;l�H;2�H;��H;��H;(�H;��H;��H;��H;^�H;�H;x�H;��H;��H;��H;��H;;�H;��H;L�H;��H;��H;,�H;X�H;��H;��H;��H;��H;��H;��H;��H;X�H;,�H;��H;��H;L�H;��H;;�H;��H;��H;��H;��H;x�H;�H;^�H;��H;��H;��H;(�H;��H;��H;2�H;l�H;��H;��H;0�H;��H;F�H;+�H;_�H;�H;�H;>�H;      ��H;�H;ƩH;�H;ƬH;��H;��H;g�H;��H;кH;/�H;��H; �H;:�H;^�H;[�H;6�H;��H;H�H;e�H;S�H;��H;m�H;��H;��H;��H;��H;k�H;��H;T�H;��H; �H;:�H;u�H;��H;��H;��H;��H;��H;u�H;:�H; �H;��H;T�H;��H;k�H;��H;��H;��H;��H;m�H;��H;S�H;e�H;H�H;��H;6�H;[�H;^�H;:�H; �H;��H;/�H;кH;��H;g�H;��H;��H;ƬH;�H;ƩH;�H;      P�H;��H;��H;[�H;��H;f�H;��H;P�H;.�H;H�H;��H;̸H;�H;>�H;5�H;��H;u�H;��H;��H;j�H;��H;��H;��H;K�H;��H;��H;��H;��H;b�H;�H;h�H;��H;	�H;:�H;X�H;��H;��H;��H;X�H;:�H;	�H;��H;h�H;�H;b�H;��H;��H;��H;��H;K�H;��H;��H;��H;j�H;��H;��H;u�H;��H;5�H;>�H;�H;̸H;��H;H�H;.�H;P�H;��H;f�H;��H;[�H;��H;��H;      w�H;�H;B�H;u�H;k�H;%�H;q�H;0�H;H�H;��H;&�H;��H;$�H;�H;��H;f�H;��H;��H;��H;B�H;F�H;��H;Q�H;[�H;�H;��H;��H;��H;��H;n�H;�H;z�H;��H; �H;,�H;J�H;I�H;J�H;,�H; �H;��H;z�H;�H;n�H;��H;��H;��H;��H;�H;[�H;Q�H;��H;F�H;B�H;��H;��H;��H;f�H;��H;�H;$�H;��H;&�H;��H;H�H;0�H;q�H;%�H;k�H;u�H;B�H;�H;      fH;�fH;YhH;@kH;(oH;�sH;�yH;�H;��H;ۍH;�H;s�H;��H;��H;$�H;T�H;'�H;��H;x�H;��H;��H;1�H;=�H;��H;��H;��H;X�H;��H;��H;��H;t�H;�H;h�H;��H;��H;�H;0�H;�H;��H;��H;h�H;�H;t�H;��H;��H;��H;X�H;��H;��H;��H;=�H;1�H;��H;��H;x�H;��H;'�H;T�H;$�H;��H;��H;s�H;�H;ۍH;��H;�H;�yH;�sH;(oH;@kH;YhH;�fH;      :?H;@H;cBH;.FH;[KH;�QH;'YH;gaH;KjH;�sH;0}H;ʆH;G�H;y�H;9�H;g�H;�H;׸H;�H;��H;��H;7�H;�H;\�H;9�H;��H;��H;L�H;��H;��H;��H;n�H;�H;T�H;��H;��H;��H;��H;��H;T�H;�H;n�H;��H;��H;��H;L�H;��H;��H;9�H;\�H;�H;7�H;��H;��H;�H;׸H;�H;g�H;9�H;y�H;G�H;ʆH;0}H;�sH;KjH;gaH;'YH;�QH;[KH;.FH;cBH;@H;      >H;TH;vH;�H;nH;�$H;�.H;�9H;�EH;�QH;k^H;�jH;SwH;W�H;ԎH;��H;��H;��H;��H;ۻH;b�H;�H;��H;"�H;��H;��H;h�H;��H;-�H;��H;��H;��H;b�H;��H;L�H;�H;��H;�H;L�H;��H;b�H;��H;��H;��H;-�H;��H;h�H;��H;��H;"�H;��H;�H;b�H;ۻH;��H;��H;��H;��H;ԎH;W�H;SwH;�jH;k^H;�QH;�EH;�9H;�.H;�$H;nH;�H;vH;TH;      &�G;��G;��G;%�G;�G;6�G;"�G;�H;H;d&H;�6H;�GH;�WH;HgH;*vH;�H;�H;ԜH;T�H;��H;��H;E�H;��H;��H;~�H;k�H;��H;G�H;��H;L�H;��H;��H;��H;k�H;��H;�H; �H;�H;��H;k�H;��H;��H;��H;L�H;��H;G�H;��H;k�H;~�H;��H;��H;E�H;��H;��H;T�H;ԜH;�H;�H;*vH;HgH;�WH;�GH;�6H;d&H;H;�H;"�G;6�G;�G;%�G;��G;��G;      �mG;<pG;wG;�G;��G;_�G;|�G;��G;'�G;M�G;�H;pH;�/H;�CH;@WH;9iH;�yH;�H;��H;ԢH;m�H;��H;��H;��H;@�H;/�H;N�H;��H;h�H;��H;X�H;��H;��H;��H;;�H;��H;��H;��H;;�H;��H;��H;��H;X�H;��H;h�H;��H;N�H;/�H;@�H;��H;��H;��H;m�H;ԢH;��H;�H;�yH;9iH;@WH;�CH;�/H;pH;�H;M�G;'�G;��G;|�G;_�G;��G;�G;wG;<pG;      ��F;�F;4�F;��F;,�F;� G;�EG;biG;l�G;-�G;,�G;�G;=�G;�H;�0H;�GH;:]H;�pH;�H;��H;<�H;��H;��H;��H;��H;�H;/�H;k�H;��H;��H;��H;��H;��H;��H;��H;��H;�H;��H;��H;��H;��H;��H;��H;��H;��H;k�H;/�H;�H;��H;��H;��H;��H;<�H;��H;�H;�pH;:]H;�GH;�0H;�H;=�G;�G;,�G;-�G;l�G;biG;�EG;� G;,�F;��F;4�F;�F;      ��D;C�D;B�D;�8E;��E;f�E;�OF;/�F;��F;K9G;mnG;ޙG;�G;��G;� H;�H;�9H;�RH;�hH;e|H;��H;��H;h�H;#�H;U�H;��H;@�H;~�H;��H;9�H;��H;�H;��H;��H;��H;.�H;r�H;.�H;��H;��H;��H;�H;��H;9�H;��H;~�H;@�H;��H;U�H;#�H;h�H;��H;��H;e|H;�hH;�RH;�9H;�H;� H;��G;�G;ޙG;mnG;K9G;��F;/�F;�OF;f�E;��E;�8E;B�D;C�D;      �@;�@@;g�@;^QA;"B;G
C;�C;��D;\�E;�?F;��F;� G;:gG;ÛG;a�G;�G;�H; .H;.JH;�bH;mxH;9�H;P�H;ܨH;#�H;��H;��H;��H;"�H;\�H;��H;[�H;K�H;��H;��H;i�H;��H;i�H;��H;��H;K�H;[�H;��H;\�H;"�H;��H;��H;��H;#�H;ܨH;P�H;9�H;mxH;�bH;.JH; .H;�H;�G;a�G;ÛG;:gG;� G;��F;�?F;\�E;��D;�C;G
C;"B;^QA;g�@;�@@;      �36;˃6;kk7;��8;��:;��<;��>;��@;�sB;��C;�+E;	F;/�F;�+G;�wG;Z�G;��G;�H;%H;7DH;0_H;hvH;O�H;P�H;h�H;��H;��H;��H;��H;�H;=�H;Q�H;��H;m�H;��H;{�H;��H;{�H;��H;m�H;��H;Q�H;=�H;�H;��H;��H;��H;��H;h�H;P�H;O�H;hvH;0_H;7DH;%H;�H;��G;Z�G;�wG;�+G;/�F;	F;�+E;��C;�sB;��@;��>;��<;��:;��8;kk7;˃6;      �";�L#;�%;��';��+;��/;A�3;��7;Q�;;x?;O�A;��C;D9E;�?F;:�F;�TG;��G;T�G;��G;xH;AH;�]H;hvH;9�H;��H;��H;��H;E�H;�H;7�H;1�H;��H;��H;��H;x�H;U�H;��H;U�H;x�H;��H;��H;��H;1�H;7�H;�H;E�H;��H;��H;��H;9�H;hvH;�]H;AH;xH;��G;T�G;��G;�TG;:�F;�?F;D9E;��C;O�A;x?;Q�;;��7;A�3;��/;��+;��';�%;�L#;      ���:�$ ;�;��;��;|P;�l;�c';w�.;�<5;F�:;�>;1B;ZAD;��E;��F;,6G;��G;��G;F�G;�H;AH;0_H;mxH;��H;<�H;m�H;��H;b�H;��H;��H;F�H;��H;S�H;�H;��H;[�H;��H;�H;S�H;��H;F�H;��H;��H;b�H;��H;m�H;<�H;��H;mxH;0_H;AH;�H;F�G;��G;��G;,6G;��F;��E;ZAD;1B;�>;F�:;�<5;w�.;�c';�l;|P;��;��;�;�$ ;      Y�:�n�:W�:��:�%�:մ�:���:��	;�P;RM#;�m-;��5;T�;;�@@;�OC;jFE;!uF;!G;��G;�G;F�G;xH;7DH;�bH;e|H;��H;ԢH;��H;ۻH;��H;��H;B�H;j�H;e�H;^�H;��H;��H;��H;^�H;e�H;j�H;B�H;��H;��H;ۻH;��H;ԢH;��H;e|H;�bH;7DH;xH;F�G;�G;��G;!G;!uF;jFE;�OC;�@@;T�;;��5;�m-;RM#;�P;��	;���:մ�:�%�:��:W�:�n�:      �	�����j��
_��3u9�:�i~:���:[�:{�;�;�%;at0;�8;ذ>;[�B;��D;�WF;tG;��G;��G;��G;%H;.JH;�hH;�H;��H;T�H;��H;�H;x�H;��H;��H;H�H;��H;��H;i�H;��H;��H;H�H;��H;��H;x�H;�H;��H;T�H;��H;�H;�hH;.JH;%H;��G;��G;��G;tG;�WF;��D;[�B;ذ>;�8;at0;�%;�;{�;[�:���:�i~:�:3u9
_���j�����      ^A?���9��8)��Z�~ܺjp������O998�@:�:��:��	;�X;�,;8�6;֜=;x"B; �D;�WF;!G;��G;T�G;�H; .H;�RH;�pH;�H;ԜH;��H;׸H;��H;��H;��H;��H;��H;0�H;��H;0�H;��H;��H;��H;��H;��H;׸H;��H;ԜH;�H;�pH;�RH; .H;�H;T�G;��G;!G;�WF; �D;x"B;֜=;8�6;�,;�X;��	;��:�:8�@:O99����jp��~ܺ�Z��8)���9�      �Eֻ�ѻm�Ļ4T��_�q.o���.�ܺ��B�E��8�\:�%�:���:�P;^);�<5;L:=;x"B;��D;!uF;,6G;��G;��G;�H;�9H;:]H;�yH;�H;��H;�H;'�H;��H;u�H;6�H;��H;B�H;��H;B�H;��H;6�H;u�H;��H;'�H;�H;��H;�H;�yH;:]H;�9H;�H;��G;��G;,6G;!uF;��D;x"B;L:=;�<5;^);�P;���:�%�:�\:E��8��B�ܺ��.�q.o�_�4T��m�Ļ�ѻ      FB��>�r�4�$�$�F���Z�ښ��nݎ�+A?�CӺ����o2�92q�:�W�:�;E�';�<5;֜=;[�B;jFE;��F;�TG;Z�G;�G;�H;�GH;9iH;�H;��H;g�H;T�H;f�H;��H;[�H;(�H;6�H;��H;6�H;(�H;[�H;��H;f�H;T�H;g�H;��H;�H;9iH;�GH;�H;�G;Z�G;�TG;��F;jFE;[�B;֜=;�<5;E�';�;�W�:2q�:o2�9����CӺ+A?�nݎ�ښ���Z�F��$�$�r�4��>�      <y��ݜ��A���I����s�m�P��%+����P�Ļ����|���o��8u9�W�::+�:�;^);8�6;ذ>;�OC;��E;:�F;�wG;a�G;� H;�0H;@WH;*vH;ԎH;9�H;$�H;��H;5�H;^�H;��H;�H;��H;�H;��H;^�H;5�H;��H;$�H;9�H;ԎH;*vH;@WH;�0H;� H;a�G;�wG;:�F;��E;�OC;ذ>;8�6;^);�;:+�:�W�:�8u9��o�|�����P�Ļ����%+�m�P���s��I���A��ݜ�      -������aW缐�ռ�վ��Τ��I��Z�[��(��Z�g�9��{���99�W�:�W�:�P;�,;�8;�@@;ZAD;�?F;�+G;ÛG;��G;�H;�CH;HgH;W�H;y�H;��H;�H;>�H;:�H;��H;��H;��H;��H;��H;:�H;>�H;�H;��H;y�H;W�H;HgH;�CH;�H;��G;ÛG;�+G;�?F;ZAD;�@@;�8;�,;�P;�W�:�W�:�99�{��g�9���Z��(�Z�[��I���Τ��վ���ռaW缧��      �6��3�X�+�ݟ�<�(�����μ߈��T���FB�=s�T����D��{���8u92q�:���:�X;at0;T�;;1B;D9E;/�F;:gG;�G;=�G;�/H;�WH;SwH;G�H;��H;$�H;�H; �H;2�H;I�H;S�H;I�H;2�H; �H;�H;$�H;��H;G�H;SwH;�WH;�/H;=�G;�G;:gG;/�F;D9E;1B;T�;;at0;�X;���:2q�:�8u9�{����D�T��=s�FB�T���߈����μ(���<�ݟ�X�+��3�      Q₽�؀���u��Xc�Q�K�K1�{�����վ�t]��b�P�l��T��g�9���o�o2�9�%�:��	;�%;��5;�>;��C;	F;� G;ޙG;�G;pH;�GH;�jH;ʆH;s�H;��H;̸H;��H;l�H;��H;��H;��H;l�H;��H;̸H;��H;s�H;ʆH;�jH;�GH;pH;�G;ޙG;� G;	F;��C;�>;��5;�%;��	;�%�:o2�9��o�g�9�T��l��b�P�t]���վ����{��K1�Q�K��Xc���u��؀�      S���r��L��n������|�u�e�N���(�ji���˼�A��b�P�=s��|������\:��:�;�m-;F�:;O�A;�+E;��F;mnG;,�G;�H;�6H;k^H;0}H;�H;&�H;��H;/�H;��H;Z�H;��H;Z�H;��H;/�H;��H;&�H;�H;0}H;k^H;�6H;�H;,�G;mnG;��F;�+E;O�A;F�:;�m-;�;��:�\:����|��=s�b�P��A����˼ji���(�e�N�|�u�����n��L���r��      �o���r���}�ս@��Kĥ�X^���Xc��3���	���˼t]��FB��Z򻆜��CӺE��8�:{�;RM#;�<5;x?;��C;�?F;K9G;-�G;M�G;d&H;�QH;�sH;ۍH;��H;H�H;кH;��H;��H;a�H;��H;��H;кH;H�H;��H;ۍH;�sH;�QH;d&H;M�G;-�G;K9G;�?F;��C;x?;�<5;RM#;{�;�:E��8CӺ�����Z�FB�t]����˼��	��3��Xc�X^��Kĥ�@��}�ս���r�      �#�6� �A'����~���gٽS��l���j��3�ji��վ�T����(�P�Ļ+A?���B�8�@:[�:�P;w�.;Q�;;�sB;\�E;��F;l�G;'�G;H;�EH;KjH;��H;H�H;.�H;��H;0�H;��H;�H;��H;0�H;��H;.�H;H�H;��H;KjH;�EH;H;'�G;l�G;��F;\�E;�sB;Q�;;w�.;�P;[�:8�@:��B�+A?�P�Ļ�(�T����վ�ji��3��j�l��S���gٽ�~����A'�6� �      �S� �O��E��5�6� �<�
���|9��l���Xc���(����߈��Z�[����nݎ�ܺO99���:��	;�c';��7;��@;��D;/�F;biG;��G;�H;�9H;gaH;�H;0�H;P�H;g�H;��H;Y�H;��H;Y�H;��H;g�H;P�H;0�H;�H;gaH;�9H;�H;��G;biG;/�F;��D;��@;��7;�c';��	;���:O99ܺnݎ����Z�[�߈�������(��Xc�l��|9����<�
�6� ��5��E� �O�      �~���)����v��9b�U�H��",�0Z���S��X^��e�N�{����μ�I���%+�ښ����.������i~:���:�l;A�3;��>;�C;�OF;�EG;|�G;"�G;�.H;'YH;�yH;q�H;��H;��H;F�H;K�H;��H;K�H;F�H;��H;��H;q�H;�yH;'YH;�.H;"�G;|�G;�EG;�OF;�C;��>;A�3;�l;���:�i~:������.�ښ���%+��I����μ{��e�N�X^��S����0Z��",�U�H��9b���v��)��      ��������:���M���r� �O��",�<�
��gٽKĥ�|�u�K1�(����Τ�m�P��Z�q.o�jp���:մ�:|P;��/;��<;G
C;f�E;� G;_�G;6�G;�$H;�QH;�sH;%�H;f�H;��H;+�H;{�H;&�H;{�H;+�H;��H;f�H;%�H;�sH;�QH;�$H;6�G;_�G;� G;f�E;G
C;��<;��/;|P;մ�:�:jp��q.o��Z�m�P��Τ�(���K1�|�u�Kĥ��gٽ<�
��",� �O��r��M���:�����      ���v��/;������:P���r�U�H�6� ��~��@������Q�K�<��վ���s�F��_�~ܺ3u9�%�:��;��+;��:;"B;��E;,�F;��G;�G;nH;[KH;(oH;k�H;��H;ƬH;_�H;��H;��H;��H;_�H;ƬH;��H;k�H;(oH;[KH;nH;�G;��G;,�F;��E;"B;��:;��+;��;�%�:3u9~ܺ_�F����s��վ�<�Q�K�����@���~��6� �U�H��r�:P������/;���v��      3Vھ�*־5ʾT��������M���9b��5���}�սn���Xc�ݟ���ռ�I��$�$�4T���Z�
_����:��;��';��8;^QA;�8E;��F;�G;%�G;�H;.FH;@kH;u�H;[�H;�H;�H;��H;t�H;��H;�H;�H;[�H;u�H;@kH;.FH;�H;%�G;�G;��F;�8E;^QA;��8;��';��;��:
_���Z�4T��$�$��I����ռݟ��Xc�n��}�ս���5��9b��M������T���5ʾ�*־      ǰ�쾐�޾5ʾ/;���:����v��E�A'���L����u�X�+�aW缨A��r�4�m�Ļ�8)��j��W�:�;�%;kk7;g�@;B�D;4�F;wG;��G;vH;cBH;YhH;B�H;��H;ƩH;�H;��H;��H;��H;�H;ƩH;��H;B�H;YhH;cBH;vH;��G;wG;4�F;B�D;g�@;kk7;�%;�;W�:�j���8)�m�Ļr�4��A��aW�X�+���u�L����A'��E���v��:��/;��5ʾ��޾��      /h���b���쾅*־�v������)�� �O�6� ��r�r���؀��3����ݜ��>��ѻ��9�����n�:�$ ;�L#;˃6;�@@;C�D;�F;<pG;��G;TH;@H;�fH;�H;��H;�H;>�H;�H;��H;�H;>�H;�H;��H;�H;�fH;@H;TH;��G;<pG;�F;C�D;�@@;˃6;�L#;�$ ;�n�:�����9��ѻ�>�ݜ�����3��؀��r���r�6� � �O��)������v���*־�쾼b��      �$��� ���������þ�*��
Dx�}�=����\Pν鰒��&K�xc����;�V�s���D^���S��v[:���:�d;��4;�_?;�lD;��F;puG;M�G;�H;�NH;�rH;�H;��H;��H;�H;q�H;E�H;q�H;�H;��H;��H;�H;�rH;�NH;�H;M�G;puG;��F;�lD;�_?;��4;�d;���:�v[:��S��D^�s��;�V����xc��&K�鰒�\Pν���}�=�
Dx��*���þ��������� �      �� �k��>��=���������0���s���:�N9���ʽZ����G��8��-��z5S�v���/X���D��Ad:�A�:� ;y�4;	�?;#~D;q�F;4xG;��G;�H;NOH;IsH;:�H;�H;�H;W�H;��H;U�H;��H;W�H;�H;�H;:�H;IsH;NOH;�H;��G;4xG;q�F;#~D;	�?;y�4;� ;�A�:�Ad:��D��/X�v��z5S��-���8���G�Z����ʽN9���:��s��0��������=��>��k��      ���>��&�
�����fYؾ���ȥ����f���0�C[�*8������ȟ>�|���#Ȥ�X6H�,�ܻ�qF�,��7�}:���:�";��5;7�?;��D;��F;/�G;��G;t"H;�QH;�tH;z�H;�H;��H;�H;�H;��H;�H;�H;��H;�H;z�H;�tH;�QH;t"H;��G;/�G;��F;��D;7�?;��5;�";���:7�}:,���qF�,�ܻX6H�#Ȥ�|���ȟ>�����*8��C[���0���f�ȥ�����fYؾ����&�
�>��      ��=������I��þ�R��&���QS��Q"��s�����}��0���d���x�6��ƻ'}*����`�:�w;�%;Rl7;�@;�D;�F;��G;��G;3'H;UH;�wH;��H;f�H;ñH;ܺH;�H;��H;�H;ܺH;ñH;f�H;��H;�wH;UH;3'H;��G;��G;�F;�D;�@;Rl7;�%;�w;`�:���'}*��ƻx�6�d����켟0���}�����s��Q"�QS�&����R���þIᾁ���=��      ����fYؾ�þ�ê�f쏾jk���:�e�R�ؽ�����c�:y���Ҽݫ��� �B�'����'7��:�
;d�(;�^9;��A;�[E;��F;�G;��G;�-H;�YH;{H;�H;i�H;u�H;6�H;�H;��H;�H;6�H;u�H;i�H;�H;{H;�YH;�-H;��G;�G;��F;�[E;��A;�^9;d�(;�
;��:��'7'��B�� �ݫ����Ҽ:y��c�����R�ؽe���:�jk�f쏾�ê��þfYؾ��      �þ��������R��f쏾�s��H����������������D�vc�g����f�3,�����P����91��:6;�i-;��;;��B;,�E;�G;��G;��G;�5H;�_H;�H;{�H;��H;r�H;ɽH;r�H;��H;r�H;ɽH;r�H;��H;{�H;�H;�_H;�5H;��G;��G;�G;,�E;��B;��;;�i-;6;1��:��9�P�����3,��f�g���vc���D���������������H��s�f쏾�R���������      �*���0��ȥ��&���jk��H��#%�B[�ZPν�s��0�f�/%�d��`���G�=�n?ػfFL��D�d�R:D�:��;�2;�=;��C;�/F;�FG;�G;WH;?H;�fH;��H;W�H;ͫH;��H;��H;�H;��H;�H;��H;��H;ͫH;W�H;��H;�fH;?H;WH;�G;�FG;�/F;��C;�=;�2;��;D�:d�R:�D�fFL�n?ػG�=�`���d��/%�0�f��s��ZPνB[��#%��H�jk�&���ȥ���0��      
Dx��s���f�QS���:����B[��7ս�榽��}�u�;��8�)����r����G������Ҭ����:��;}$;,�6;f�?;4�D;�F; pG;��G;H;XIH;dnH;i�H;��H;�H;[�H;��H;��H;G�H;��H;��H;[�H;�H;��H;i�H;dnH;XIH;H;��G; pG;�F;4�D;f�?;,�6;}$;��;���:�Ҭ����G������r�)����8�u�;���}��榽�7սB[������:�QS���f��s�      }�=���:���0��Q"�e�����ZPν�榽%����G�����Ҽ���E:�	�ܻ�D^�͸��mh:���:P;�{,;�:;��A;~hE;��F;]�G;��G;�'H;eTH;�vH;��H;L�H;��H;�H;��H;��H;4�H;��H;��H;�H;��H;L�H;��H;�vH;eTH;�'H;��G;]�G;��F;~hE;��A;�:;�{,;P;���:mh:͸���D^�	�ܻE:������Ҽ����G�%���榽ZPν����e��Q"���0���:�      ���N9�C[��s�R�ؽ���s����}���G��K��	c��!�V�$,��*���������:A��:� ;ǂ3;0>;�C;#F;$8G;l�G;�H;7H;�_H;,H;�H; �H;h�H;�H;m�H;��H;3�H;��H;m�H;�H;h�H; �H;�H;,H;�_H;7H;�H;l�G;$8G;#F;�C;0>;ǂ3;� ;A��:��:������*��$,�!�V�	c��K�����G���}��s����R�ؽ�s�C[�N9�      \Pν��ʽ*8�������������0�f�u�;���K��Ȥ���f���#ߵ�>o5�1�D�P�-:���:Y>;H+;_9;�A;��D;\�F;�uG;�G;JH;�FH;�kH;�H;��H;�H;H�H;�H;��H;"�H;F�H;"�H;��H;�H;H�H;�H;��H;�H;�kH;�FH;JH;�G;�uG;\�F;��D;�A;_9;H+;Y>;���:P�-:1�D�>o5�#ߵ�����f�Ȥ�K����u�;�0�f������������*8����ʽ      鰒�Z��������}��c���D�/%��8���Ҽ	c����f�����ƻY/X�s������9h�:ɏ;G";�3;�>;�XC;��E;G;'�G;��G;�+H;/VH;9wH;��H;W�H;�H;.�H;�H;Q�H;a�H;O�H;a�H;Q�H;�H;.�H;�H;W�H;��H;9wH;/VH;�+H;��G;'�G;G;��E;�XC;�>;�3;G";ɏ;h�:���9s���Y/X��ƻ�����f�	c����Ҽ�8�/%���D��c���}�����Z��      �&K���G�ȟ>��0�:y�vc�d��)������!�V����ƻfod���º�Q(7�3�:���: �;^P.;:�:;ayA;z�D;�F;�mG;u�G;"H;�?H;MeH;��H;R�H;ժH;��H;�H;
�H;��H;��H;W�H;��H;��H;
�H;�H;��H;ժH;R�H;��H;MeH;�?H;"H;u�G;�mG;�F;z�D;ayA;:�:;^P.; �;���:�3�:�Q(7��ºfod��ƻ��!�V����)���d��vc�:y��0�ȟ>���G�      xc��8�|����켔�Ҽg���`����r�E:�$,�#ߵ�Y/X���º�ˬ�I�}:? �:w;��);�l7;j�?;�C;LF;�(G;F�G;��G;3)H;�RH;�sH;��H;��H;�H;μH;��H;��H;,�H;��H;l�H;��H;,�H;��H;��H;μH;�H;��H;��H;�sH;�RH;3)H;��G;F�G;�(G;LF;�C;j�?;�l7;��);w;? �:I�}:�ˬ���ºY/X�#ߵ�$,�E:��r�`���g�����Ҽ��|����8�      ����-��#Ȥ�d���ݫ���f�G�=����	�ܻ�*��>o5�s����Q(7I�}:�m�:��;>&;��4;C�=;�B;,�E;T�F;̀G;$�G;cH;�@H;�dH;d�H;��H;y�H;��H;��H;;�H;��H;��H;��H;l�H;��H;��H;��H;;�H;��H;��H;y�H;��H;d�H;�dH;�@H;cH;$�G;̀G;T�F;,�E;�B;C�=;��4;>&;��;�m�:I�}:�Q(7s���>o5��*��	�ܻ���G�=��f�ݫ��d���#Ȥ��-��      ;�V�z5S�X6H�x�6�� �3,�n?ػG���D^����1�D����9�3�:? �:��;^%;��3;p�<;�B;�
E;?�F;�WG;9�G;u�G;�/H;xVH;�uH;�H;��H;ܰH;��H;��H;��H;k�H;��H;��H;Q�H;��H;��H;k�H;��H;��H;��H;ܰH;��H;�H;�uH;xVH;�/H;u�G;9�G;�WG;?�F;�
E;�B;p�<;��3;^%;��;? �:�3�:���91�D�����D^�G��n?ػ3,�� �x�6�X6H�z5S�      s��v��,�ܻ�ƻB󩻜��fFL����͸����P�-:h�:���:w;>&;��3;�8<;`�A;%�D;�YF;Z4G;3�G;�G;� H;aIH;VjH;ńH;ٙH;��H;��H;�H;��H;��H;��H;��H;v�H;�H;v�H;��H;��H;��H;��H;�H;��H;��H;ٙH;ńH;VjH;aIH;� H;�G;3�G;Z4G;�YF;%�D;`�A;�8<;��3;>&;w;���:h�:P�-:��͸�����fFL����B��ƻ,�ܻv��      �D^��/X��qF�'}*�'���P���D��Ҭ�mh:��:���:ɏ; �;��);��4;p�<;`�A;f�D;�8F;
G;��G;x�G;jH;C>H;�`H;6|H;��H;��H;��H;��H;��H;}�H;��H;4�H;��H;8�H;��H;8�H;��H;4�H;��H;}�H;��H;��H;��H;��H;��H;6|H;�`H;C>H;jH;x�G;��G;
G;�8F;f�D;`�A;p�<;��4;��); �;ɏ;���:��:mh:�Ҭ��D��P��'��'}*��qF��/X�      ��S���D�,�������'7��9d�R:���:���:A��:Y>;G";^P.;�l7;C�=;�B;%�D;�8F;YG;R�G;��G;�H;�5H;�XH;	uH;=�H;�H;�H;�H;��H;9�H;��H;-�H;M�H;r�H;��H;	�H;��H;r�H;M�H;-�H;��H;9�H;��H;�H;�H;�H;=�H;	uH;�XH;�5H;�H;��G;R�G;YG;�8F;%�D;�B;C�=;�l7;^P.;G";Y>;A��:���:���:d�R:��9��'7���,����D�      �v[:�Ad:7�}:`�:��:1��:D�:��;P;� ;H+;�3;:�:;j�?;�B;�
E;�YF;
G;R�G;��G;oH;�0H;�RH;�oH;�H;f�H;�H;��H;��H;��H;�H;��H;��H;5�H;�H;(�H;r�H;(�H;�H;5�H;��H;��H;�H;��H;��H;��H;�H;f�H;�H;�oH;�RH;�0H;oH;��G;R�G;
G;�YF;�
E;�B;j�?;:�:;�3;H+;� ;P;��;D�:1��:��:`�:7�}:�Ad:      ���:�A�:���:�w;�
;6;��;}$;�{,;ǂ3;_9;�>;ayA;�C;,�E;?�F;Z4G;��G;��G;oH;�.H;PH;'lH;i�H;��H;��H;��H;�H;��H;)�H;r�H;��H;��H;��H;z�H;W�H;��H;W�H;z�H;��H;��H;��H;r�H;)�H;��H;�H;��H;��H;��H;i�H;'lH;PH;�.H;oH;��G;��G;Z4G;?�F;,�E;�C;ayA;�>;_9;ǂ3;�{,;}$;��;6;�
;�w;���:�A�:      �d;� ;�";�%;d�(;�i-;�2;,�6;�:;0>;�A;�XC;z�D;LF;T�F;�WG;3�G;x�G;�H;�0H;PH;�jH;��H;��H;V�H;E�H;�H;��H;��H;�H;��H;��H;��H;�H;��H;j�H;��H;j�H;��H;�H;��H;��H;��H;�H;��H;��H;�H;E�H;V�H;��H;��H;�jH;PH;�0H;�H;x�G;3�G;�WG;T�F;LF;z�D;�XC;�A;0>;�:;,�6;�2;�i-;d�(;�%;�";� ;      ��4;y�4;��5;Rl7;�^9;��;;�=;f�?;��A;�C;��D;��E;�F;�(G;̀G;9�G;�G;jH;�5H;�RH;'lH;��H;̓H;$�H;گH;g�H;=�H;H�H;��H;��H;(�H;��H;C�H;��H;��H;m�H;��H;m�H;��H;��H;C�H;��H;(�H;��H;��H;H�H;=�H;g�H;گH;$�H;̓H;��H;'lH;�RH;�5H;jH;�G;9�G;̀G;�(G;�F;��E;��D;�C;��A;f�?;�=;��;;�^9;Rl7;��5;y�4;      �_?;	�?;7�?;�@;��A;��B;��C;4�D;~hE;#F;\�F;G;�mG;F�G;$�G;u�G;� H;C>H;�XH;�oH;i�H;��H;$�H;\�H;��H;<�H;Y�H;�H;��H;��H;g�H;��H;��H;��H;��H;E�H;^�H;E�H;��H;��H;��H;��H;g�H;��H;��H;�H;Y�H;<�H;��H;\�H;$�H;��H;i�H;�oH;�XH;C>H;� H;u�G;$�G;F�G;�mG;G;\�F;#F;~hE;4�D;��C;��B;��A;�@;7�?;	�?;      �lD;#~D;��D;�D;�[E;,�E;�/F;�F;��F;$8G;�uG;'�G;u�G;��G;cH;�/H;aIH;�`H;	uH;�H;��H;V�H;گH;��H;�H;��H;}�H;#�H;��H;�H;n�H;N�H;��H;��H;��H;��H;7�H;��H;��H;��H;��H;N�H;n�H;�H;��H;#�H;}�H;��H;�H;��H;گH;V�H;��H;�H;	uH;�`H;aIH;�/H;cH;��G;u�G;'�G;�uG;$8G;��F;�F;�/F;,�E;�[E;�D;��D;#~D;      ��F;q�F;��F;�F;��F;�G;�FG; pG;]�G;l�G;�G;��G;"H;3)H;�@H;xVH;VjH;6|H;=�H;f�H;��H;E�H;g�H;<�H;��H;E�H;��H;��H;��H;�H;�H;��H;��H;��H;C�H;��H;��H;��H;C�H;��H;��H;��H;�H;�H;��H;��H;��H;E�H;��H;<�H;g�H;E�H;��H;f�H;=�H;6|H;VjH;xVH;�@H;3)H;"H;��G;�G;l�G;]�G; pG;�FG;�G;��F;�F;��F;q�F;      puG;4xG;/�G;��G;�G;��G;�G;��G;��G;�H;JH;�+H;�?H;�RH;�dH;�uH;ńH;��H;�H;�H;��H;�H;=�H;Y�H;}�H;��H;t�H;m�H;��H;��H;n�H;��H;��H;M�H;��H;-�H;.�H;-�H;��H;M�H;��H;��H;n�H;��H;��H;m�H;t�H;��H;}�H;Y�H;=�H;�H;��H;�H;�H;��H;ńH;�uH;�dH;�RH;�?H;�+H;JH;�H;��G;��G;�G;��G;�G;��G;/�G;4xG;      M�G;��G;��G;��G;��G;��G;WH;H;�'H;7H;�FH;/VH;MeH;�sH;d�H;�H;ٙH;��H;�H;��H;�H;��H;H�H;�H;#�H;��H;m�H;��H;��H;p�H;��H;��H;c�H;��H;V�H;��H;��H;��H;V�H;��H;c�H;��H;��H;p�H;��H;��H;m�H;��H;#�H;�H;H�H;��H;�H;��H;�H;��H;ٙH;�H;d�H;�sH;MeH;/VH;�FH;7H;�'H;H;WH;��G;��G;��G;��G;��G;      �H;�H;t"H;3'H;�-H;�5H;?H;XIH;eTH;�_H;�kH;9wH;��H;��H;��H;��H;��H;��H;�H;��H;��H;��H;��H;��H;��H;��H;��H;��H;>�H;��H;��H;X�H;��H;y�H;��H;��H;��H;��H;��H;y�H;��H;X�H;��H;��H;>�H;��H;��H;��H;��H;��H;��H;��H;��H;��H;�H;��H;��H;��H;��H;��H;��H;9wH;�kH;�_H;eTH;XIH;?H;�5H;�-H;3'H;t"H;�H;      �NH;NOH;�QH;UH;�YH;�_H;�fH;dnH;�vH;,H;�H;��H;R�H;��H;y�H;ܰH;��H;��H;��H;��H;)�H;�H;��H;��H;�H;�H;��H;p�H;��H;��H;V�H;��H;q�H;��H;�H;%�H;?�H;%�H;�H;��H;q�H;��H;V�H;��H;��H;p�H;��H;�H;�H;��H;��H;�H;)�H;��H;��H;��H;��H;ܰH;y�H;��H;R�H;��H;�H;,H;�vH;dnH;�fH;�_H;�YH;UH;�QH;NOH;      �rH;IsH;�tH;�wH;{H;�H;��H;i�H;��H;�H;��H;W�H;ժH;�H;��H;��H;�H;��H;9�H;�H;r�H;��H;(�H;g�H;n�H;�H;n�H;��H;��H;V�H;��H;q�H;��H;�H;_�H;l�H;d�H;l�H;_�H;�H;��H;q�H;��H;V�H;��H;��H;n�H;�H;n�H;g�H;(�H;��H;r�H;�H;9�H;��H;�H;��H;��H;�H;ժH;W�H;��H;�H;��H;i�H;��H;�H;{H;�wH;�tH;IsH;      �H;:�H;z�H;��H;�H;{�H;W�H;��H;L�H; �H;�H;�H;��H;μH;��H;��H;��H;}�H;��H;��H;��H;��H;��H;��H;N�H;��H;��H;��H;X�H;��H;q�H;��H;�H;_�H;��H;��H;��H;��H;��H;_�H;�H;��H;q�H;��H;X�H;��H;��H;��H;N�H;��H;��H;��H;��H;��H;��H;}�H;��H;��H;��H;μH;��H;�H;�H; �H;L�H;��H;W�H;{�H;�H;��H;z�H;:�H;      ��H;�H;�H;f�H;i�H;��H;ͫH;�H;��H;h�H;H�H;.�H;�H;��H;;�H;��H;��H;��H;-�H;��H;��H;��H;C�H;��H;��H;��H;��H;c�H;��H;q�H;��H;�H;X�H;��H;��H;��H;��H;��H;��H;��H;X�H;�H;��H;q�H;��H;c�H;��H;��H;��H;��H;C�H;��H;��H;��H;-�H;��H;��H;��H;;�H;��H;�H;.�H;H�H;h�H;��H;�H;ͫH;��H;i�H;f�H;�H;�H;      ��H;�H;��H;ñH;u�H;r�H;��H;[�H;�H;�H;�H;�H;
�H;��H;��H;k�H;��H;4�H;M�H;5�H;��H;�H;��H;��H;��H;��H;M�H;��H;y�H;��H;�H;_�H;��H;��H;��H;��H;��H;��H;��H;��H;��H;_�H;�H;��H;y�H;��H;M�H;��H;��H;��H;��H;�H;��H;5�H;M�H;4�H;��H;k�H;��H;��H;
�H;�H;�H;�H;�H;[�H;��H;r�H;u�H;ñH;��H;�H;      �H;W�H;�H;ܺH;6�H;ɽH;��H;��H;��H;m�H;��H;Q�H;��H;,�H;��H;��H;��H;��H;r�H;�H;z�H;��H;��H;��H;��H;C�H;��H;V�H;��H;�H;_�H;��H;��H;��H;��H;��H;��H;��H;��H;��H;��H;��H;_�H;�H;��H;V�H;��H;C�H;��H;��H;��H;��H;z�H;�H;r�H;��H;��H;��H;��H;,�H;��H;Q�H;��H;m�H;��H;��H;��H;ɽH;6�H;ܺH;�H;W�H;      q�H;��H;�H;�H;�H;r�H;�H;��H;��H;��H;"�H;a�H;��H;��H;��H;��H;v�H;8�H;��H;(�H;W�H;j�H;m�H;E�H;��H;��H;-�H;��H;��H;%�H;l�H;��H;��H;��H;��H;��H;��H;��H;��H;��H;��H;��H;l�H;%�H;��H;��H;-�H;��H;��H;E�H;m�H;j�H;W�H;(�H;��H;8�H;v�H;��H;��H;��H;��H;a�H;"�H;��H;��H;��H;�H;r�H;�H;�H;�H;��H;      E�H;U�H;��H;��H;��H;��H;��H;G�H;4�H;3�H;F�H;O�H;W�H;l�H;l�H;Q�H;�H;��H;	�H;r�H;��H;��H;��H;^�H;7�H;��H;.�H;��H;��H;?�H;d�H;��H;��H;��H;��H;��H;��H;��H;��H;��H;��H;��H;d�H;?�H;��H;��H;.�H;��H;7�H;^�H;��H;��H;��H;r�H;	�H;��H;�H;Q�H;l�H;l�H;W�H;O�H;F�H;3�H;4�H;G�H;��H;��H;��H;��H;��H;U�H;      q�H;��H;�H;�H;�H;r�H;�H;��H;��H;��H;"�H;a�H;��H;��H;��H;��H;v�H;8�H;��H;(�H;W�H;j�H;m�H;E�H;��H;��H;-�H;��H;��H;%�H;l�H;��H;��H;��H;��H;��H;��H;��H;��H;��H;��H;��H;l�H;%�H;��H;��H;-�H;��H;��H;E�H;m�H;j�H;W�H;(�H;��H;8�H;v�H;��H;��H;��H;��H;a�H;"�H;��H;��H;��H;�H;r�H;�H;�H;�H;��H;      �H;W�H;�H;ܺH;6�H;ɽH;��H;��H;��H;m�H;��H;Q�H;��H;,�H;��H;��H;��H;��H;r�H;�H;z�H;��H;��H;��H;��H;C�H;��H;V�H;��H;�H;_�H;��H;��H;��H;��H;��H;��H;��H;��H;��H;��H;��H;_�H;�H;��H;V�H;��H;C�H;��H;��H;��H;��H;z�H;�H;r�H;��H;��H;��H;��H;,�H;��H;Q�H;��H;m�H;��H;��H;��H;ɽH;6�H;ܺH;�H;W�H;      ��H;�H;��H;ñH;u�H;r�H;��H;[�H;�H;�H;�H;�H;
�H;��H;��H;k�H;��H;4�H;M�H;5�H;��H;�H;��H;��H;��H;��H;M�H;��H;y�H;��H;�H;_�H;��H;��H;��H;��H;��H;��H;��H;��H;��H;_�H;�H;��H;y�H;��H;M�H;��H;��H;��H;��H;�H;��H;5�H;M�H;4�H;��H;k�H;��H;��H;
�H;�H;�H;�H;�H;[�H;��H;r�H;u�H;ñH;��H;�H;      ��H;�H;�H;f�H;i�H;��H;ͫH;�H;��H;h�H;H�H;.�H;�H;��H;;�H;��H;��H;��H;-�H;��H;��H;��H;C�H;��H;��H;��H;��H;c�H;��H;q�H;��H;�H;X�H;��H;��H;��H;��H;��H;��H;��H;X�H;�H;��H;q�H;��H;c�H;��H;��H;��H;��H;C�H;��H;��H;��H;-�H;��H;��H;��H;;�H;��H;�H;.�H;H�H;h�H;��H;�H;ͫH;��H;i�H;f�H;�H;�H;      �H;:�H;z�H;��H;�H;{�H;W�H;��H;L�H; �H;�H;�H;��H;μH;��H;��H;��H;}�H;��H;��H;��H;��H;��H;��H;N�H;��H;��H;��H;X�H;��H;q�H;��H;�H;_�H;��H;��H;��H;��H;��H;_�H;�H;��H;q�H;��H;X�H;��H;��H;��H;N�H;��H;��H;��H;��H;��H;��H;}�H;��H;��H;��H;μH;��H;�H;�H; �H;L�H;��H;W�H;{�H;�H;��H;z�H;:�H;      �rH;IsH;�tH;�wH;{H;�H;��H;i�H;��H;�H;��H;W�H;ժH;�H;��H;��H;�H;��H;9�H;�H;r�H;��H;(�H;g�H;n�H;�H;n�H;��H;��H;V�H;��H;q�H;��H;�H;_�H;l�H;d�H;l�H;_�H;�H;��H;q�H;��H;V�H;��H;��H;n�H;�H;n�H;g�H;(�H;��H;r�H;�H;9�H;��H;�H;��H;��H;�H;ժH;W�H;��H;�H;��H;i�H;��H;�H;{H;�wH;�tH;IsH;      �NH;NOH;�QH;UH;�YH;�_H;�fH;dnH;�vH;,H;�H;��H;R�H;��H;y�H;ܰH;��H;��H;��H;��H;)�H;�H;��H;��H;�H;�H;��H;p�H;��H;��H;V�H;��H;q�H;��H;�H;%�H;?�H;%�H;�H;��H;q�H;��H;V�H;��H;��H;p�H;��H;�H;�H;��H;��H;�H;)�H;��H;��H;��H;��H;ܰH;y�H;��H;R�H;��H;�H;,H;�vH;dnH;�fH;�_H;�YH;UH;�QH;NOH;      �H;�H;t"H;3'H;�-H;�5H;?H;XIH;eTH;�_H;�kH;9wH;��H;��H;��H;��H;��H;��H;�H;��H;��H;��H;��H;��H;��H;��H;��H;��H;>�H;��H;��H;X�H;��H;y�H;��H;��H;��H;��H;��H;y�H;��H;X�H;��H;��H;>�H;��H;��H;��H;��H;��H;��H;��H;��H;��H;�H;��H;��H;��H;��H;��H;��H;9wH;�kH;�_H;eTH;XIH;?H;�5H;�-H;3'H;t"H;�H;      M�G;��G;��G;��G;��G;��G;WH;H;�'H;7H;�FH;/VH;MeH;�sH;d�H;�H;ٙH;��H;�H;��H;�H;��H;H�H;�H;#�H;��H;m�H;��H;��H;p�H;��H;��H;c�H;��H;V�H;��H;��H;��H;V�H;��H;c�H;��H;��H;p�H;��H;��H;m�H;��H;#�H;�H;H�H;��H;�H;��H;�H;��H;ٙH;�H;d�H;�sH;MeH;/VH;�FH;7H;�'H;H;WH;��G;��G;��G;��G;��G;      puG;4xG;/�G;��G;�G;��G;�G;��G;��G;�H;JH;�+H;�?H;�RH;�dH;�uH;ńH;��H;�H;�H;��H;�H;=�H;Y�H;}�H;��H;t�H;m�H;��H;��H;n�H;��H;��H;M�H;��H;-�H;.�H;-�H;��H;M�H;��H;��H;n�H;��H;��H;m�H;t�H;��H;}�H;Y�H;=�H;�H;��H;�H;�H;��H;ńH;�uH;�dH;�RH;�?H;�+H;JH;�H;��G;��G;�G;��G;�G;��G;/�G;4xG;      ��F;q�F;��F;�F;��F;�G;�FG; pG;]�G;l�G;�G;��G;"H;3)H;�@H;xVH;VjH;6|H;=�H;f�H;��H;E�H;g�H;<�H;��H;E�H;��H;��H;��H;�H;�H;��H;��H;��H;C�H;��H;��H;��H;C�H;��H;��H;��H;�H;�H;��H;��H;��H;E�H;��H;<�H;g�H;E�H;��H;f�H;=�H;6|H;VjH;xVH;�@H;3)H;"H;��G;�G;l�G;]�G; pG;�FG;�G;��F;�F;��F;q�F;      �lD;#~D;��D;�D;�[E;,�E;�/F;�F;��F;$8G;�uG;'�G;u�G;��G;cH;�/H;aIH;�`H;	uH;�H;��H;V�H;گH;��H;�H;��H;}�H;#�H;��H;�H;n�H;N�H;��H;��H;��H;��H;7�H;��H;��H;��H;��H;N�H;n�H;�H;��H;#�H;}�H;��H;�H;��H;گH;V�H;��H;�H;	uH;�`H;aIH;�/H;cH;��G;u�G;'�G;�uG;$8G;��F;�F;�/F;,�E;�[E;�D;��D;#~D;      �_?;	�?;7�?;�@;��A;��B;��C;4�D;~hE;#F;\�F;G;�mG;F�G;$�G;u�G;� H;C>H;�XH;�oH;i�H;��H;$�H;\�H;��H;<�H;Y�H;�H;��H;��H;g�H;��H;��H;��H;��H;E�H;^�H;E�H;��H;��H;��H;��H;g�H;��H;��H;�H;Y�H;<�H;��H;\�H;$�H;��H;i�H;�oH;�XH;C>H;� H;u�G;$�G;F�G;�mG;G;\�F;#F;~hE;4�D;��C;��B;��A;�@;7�?;	�?;      ��4;y�4;��5;Rl7;�^9;��;;�=;f�?;��A;�C;��D;��E;�F;�(G;̀G;9�G;�G;jH;�5H;�RH;'lH;��H;̓H;$�H;گH;g�H;=�H;H�H;��H;��H;(�H;��H;C�H;��H;��H;m�H;��H;m�H;��H;��H;C�H;��H;(�H;��H;��H;H�H;=�H;g�H;گH;$�H;̓H;��H;'lH;�RH;�5H;jH;�G;9�G;̀G;�(G;�F;��E;��D;�C;��A;f�?;�=;��;;�^9;Rl7;��5;y�4;      �d;� ;�";�%;d�(;�i-;�2;,�6;�:;0>;�A;�XC;z�D;LF;T�F;�WG;3�G;x�G;�H;�0H;PH;�jH;��H;��H;V�H;E�H;�H;��H;��H;�H;��H;��H;��H;�H;��H;j�H;��H;j�H;��H;�H;��H;��H;��H;�H;��H;��H;�H;E�H;V�H;��H;��H;�jH;PH;�0H;�H;x�G;3�G;�WG;T�F;LF;z�D;�XC;�A;0>;�:;,�6;�2;�i-;d�(;�%;�";� ;      ���:�A�:���:�w;�
;6;��;}$;�{,;ǂ3;_9;�>;ayA;�C;,�E;?�F;Z4G;��G;��G;oH;�.H;PH;'lH;i�H;��H;��H;��H;�H;��H;)�H;r�H;��H;��H;��H;z�H;W�H;��H;W�H;z�H;��H;��H;��H;r�H;)�H;��H;�H;��H;��H;��H;i�H;'lH;PH;�.H;oH;��G;��G;Z4G;?�F;,�E;�C;ayA;�>;_9;ǂ3;�{,;}$;��;6;�
;�w;���:�A�:      �v[:�Ad:7�}:`�:��:1��:D�:��;P;� ;H+;�3;:�:;j�?;�B;�
E;�YF;
G;R�G;��G;oH;�0H;�RH;�oH;�H;f�H;�H;��H;��H;��H;�H;��H;��H;5�H;�H;(�H;r�H;(�H;�H;5�H;��H;��H;�H;��H;��H;��H;�H;f�H;�H;�oH;�RH;�0H;oH;��G;R�G;
G;�YF;�
E;�B;j�?;:�:;�3;H+;� ;P;��;D�:1��:��:`�:7�}:�Ad:      ��S���D�,�������'7��9d�R:���:���:A��:Y>;G";^P.;�l7;C�=;�B;%�D;�8F;YG;R�G;��G;�H;�5H;�XH;	uH;=�H;�H;�H;�H;��H;9�H;��H;-�H;M�H;r�H;��H;	�H;��H;r�H;M�H;-�H;��H;9�H;��H;�H;�H;�H;=�H;	uH;�XH;�5H;�H;��G;R�G;YG;�8F;%�D;�B;C�=;�l7;^P.;G";Y>;A��:���:���:d�R:��9��'7���,����D�      �D^��/X��qF�'}*�'���P���D��Ҭ�mh:��:���:ɏ; �;��);��4;p�<;`�A;f�D;�8F;
G;��G;x�G;jH;C>H;�`H;6|H;��H;��H;��H;��H;��H;}�H;��H;4�H;��H;8�H;��H;8�H;��H;4�H;��H;}�H;��H;��H;��H;��H;��H;6|H;�`H;C>H;jH;x�G;��G;
G;�8F;f�D;`�A;p�<;��4;��); �;ɏ;���:��:mh:�Ҭ��D��P��'��'}*��qF��/X�      s��v��,�ܻ�ƻB󩻜��fFL����͸����P�-:h�:���:w;>&;��3;�8<;`�A;%�D;�YF;Z4G;3�G;�G;� H;aIH;VjH;ńH;ٙH;��H;��H;�H;��H;��H;��H;��H;v�H;�H;v�H;��H;��H;��H;��H;�H;��H;��H;ٙH;ńH;VjH;aIH;� H;�G;3�G;Z4G;�YF;%�D;`�A;�8<;��3;>&;w;���:h�:P�-:��͸�����fFL����B��ƻ,�ܻv��      ;�V�z5S�X6H�x�6�� �3,�n?ػG���D^����1�D����9�3�:? �:��;^%;��3;p�<;�B;�
E;?�F;�WG;9�G;u�G;�/H;xVH;�uH;�H;��H;ܰH;��H;��H;��H;k�H;��H;��H;Q�H;��H;��H;k�H;��H;��H;��H;ܰH;��H;�H;�uH;xVH;�/H;u�G;9�G;�WG;?�F;�
E;�B;p�<;��3;^%;��;? �:�3�:���91�D�����D^�G��n?ػ3,�� �x�6�X6H�z5S�      ����-��#Ȥ�d���ݫ���f�G�=����	�ܻ�*��>o5�s����Q(7I�}:�m�:��;>&;��4;C�=;�B;,�E;T�F;̀G;$�G;cH;�@H;�dH;d�H;��H;y�H;��H;��H;;�H;��H;��H;��H;l�H;��H;��H;��H;;�H;��H;��H;y�H;��H;d�H;�dH;�@H;cH;$�G;̀G;T�F;,�E;�B;C�=;��4;>&;��;�m�:I�}:�Q(7s���>o5��*��	�ܻ���G�=��f�ݫ��d���#Ȥ��-��      xc��8�|����켔�Ҽg���`����r�E:�$,�#ߵ�Y/X���º�ˬ�I�}:? �:w;��);�l7;j�?;�C;LF;�(G;F�G;��G;3)H;�RH;�sH;��H;��H;�H;μH;��H;��H;,�H;��H;l�H;��H;,�H;��H;��H;μH;�H;��H;��H;�sH;�RH;3)H;��G;F�G;�(G;LF;�C;j�?;�l7;��);w;? �:I�}:�ˬ���ºY/X�#ߵ�$,�E:��r�`���g�����Ҽ��|����8�      �&K���G�ȟ>��0�:y�vc�d��)������!�V����ƻfod���º�Q(7�3�:���: �;^P.;:�:;ayA;z�D;�F;�mG;u�G;"H;�?H;MeH;��H;R�H;ժH;��H;�H;
�H;��H;��H;W�H;��H;��H;
�H;�H;��H;ժH;R�H;��H;MeH;�?H;"H;u�G;�mG;�F;z�D;ayA;:�:;^P.; �;���:�3�:�Q(7��ºfod��ƻ��!�V����)���d��vc�:y��0�ȟ>���G�      鰒�Z��������}��c���D�/%��8���Ҽ	c����f�����ƻY/X�s������9h�:ɏ;G";�3;�>;�XC;��E;G;'�G;��G;�+H;/VH;9wH;��H;W�H;�H;.�H;�H;Q�H;a�H;O�H;a�H;Q�H;�H;.�H;�H;W�H;��H;9wH;/VH;�+H;��G;'�G;G;��E;�XC;�>;�3;G";ɏ;h�:���9s���Y/X��ƻ�����f�	c����Ҽ�8�/%���D��c���}�����Z��      \Pν��ʽ*8�������������0�f�u�;���K��Ȥ���f���#ߵ�>o5�1�D�P�-:���:Y>;H+;_9;�A;��D;\�F;�uG;�G;JH;�FH;�kH;�H;��H;�H;H�H;�H;��H;"�H;F�H;"�H;��H;�H;H�H;�H;��H;�H;�kH;�FH;JH;�G;�uG;\�F;��D;�A;_9;H+;Y>;���:P�-:1�D�>o5�#ߵ�����f�Ȥ�K����u�;�0�f������������*8����ʽ      ���N9�C[��s�R�ؽ���s����}���G��K��	c��!�V�$,��*���������:A��:� ;ǂ3;0>;�C;#F;$8G;l�G;�H;7H;�_H;,H;�H; �H;h�H;�H;m�H;��H;3�H;��H;m�H;�H;h�H; �H;�H;,H;�_H;7H;�H;l�G;$8G;#F;�C;0>;ǂ3;� ;A��:��:������*��$,�!�V�	c��K�����G���}��s����R�ؽ�s�C[�N9�      }�=���:���0��Q"�e�����ZPν�榽%����G�����Ҽ���E:�	�ܻ�D^�͸��mh:���:P;�{,;�:;��A;~hE;��F;]�G;��G;�'H;eTH;�vH;��H;L�H;��H;�H;��H;��H;4�H;��H;��H;�H;��H;L�H;��H;�vH;eTH;�'H;��G;]�G;��F;~hE;��A;�:;�{,;P;���:mh:͸���D^�	�ܻE:������Ҽ����G�%���榽ZPν����e��Q"���0���:�      
Dx��s���f�QS���:����B[��7ս�榽��}�u�;��8�)����r����G������Ҭ����:��;}$;,�6;f�?;4�D;�F; pG;��G;H;XIH;dnH;i�H;��H;�H;[�H;��H;��H;G�H;��H;��H;[�H;�H;��H;i�H;dnH;XIH;H;��G; pG;�F;4�D;f�?;,�6;}$;��;���:�Ҭ����G������r�)����8�u�;���}��榽�7սB[������:�QS���f��s�      �*���0��ȥ��&���jk��H��#%�B[�ZPν�s��0�f�/%�d��`���G�=�n?ػfFL��D�d�R:D�:��;�2;�=;��C;�/F;�FG;�G;WH;?H;�fH;��H;W�H;ͫH;��H;��H;�H;��H;�H;��H;��H;ͫH;W�H;��H;�fH;?H;WH;�G;�FG;�/F;��C;�=;�2;��;D�:d�R:�D�fFL�n?ػG�=�`���d��/%�0�f��s��ZPνB[��#%��H�jk�&���ȥ���0��      �þ��������R��f쏾�s��H����������������D�vc�g����f�3,�����P����91��:6;�i-;��;;��B;,�E;�G;��G;��G;�5H;�_H;�H;{�H;��H;r�H;ɽH;r�H;��H;r�H;ɽH;r�H;��H;{�H;�H;�_H;�5H;��G;��G;�G;,�E;��B;��;;�i-;6;1��:��9�P�����3,��f�g���vc���D���������������H��s�f쏾�R���������      ����fYؾ�þ�ê�f쏾jk���:�e�R�ؽ�����c�:y���Ҽݫ��� �B�'����'7��:�
;d�(;�^9;��A;�[E;��F;�G;��G;�-H;�YH;{H;�H;i�H;u�H;6�H;�H;��H;�H;6�H;u�H;i�H;�H;{H;�YH;�-H;��G;�G;��F;�[E;��A;�^9;d�(;�
;��:��'7'��B�� �ݫ����Ҽ:y��c�����R�ؽe���:�jk�f쏾�ê��þfYؾ��      ��=������I��þ�R��&���QS��Q"��s�����}��0���d���x�6��ƻ'}*����`�:�w;�%;Rl7;�@;�D;�F;��G;��G;3'H;UH;�wH;��H;f�H;ñH;ܺH;�H;��H;�H;ܺH;ñH;f�H;��H;�wH;UH;3'H;��G;��G;�F;�D;�@;Rl7;�%;�w;`�:���'}*��ƻx�6�d����켟0���}�����s��Q"�QS�&����R���þIᾁ���=��      ���>��&�
�����fYؾ���ȥ����f���0�C[�*8������ȟ>�|���#Ȥ�X6H�,�ܻ�qF�,��7�}:���:�";��5;7�?;��D;��F;/�G;��G;t"H;�QH;�tH;z�H;�H;��H;�H;�H;��H;�H;�H;��H;�H;z�H;�tH;�QH;t"H;��G;/�G;��F;��D;7�?;��5;�";���:7�}:,���qF�,�ܻX6H�#Ȥ�|���ȟ>�����*8��C[���0���f�ȥ�����fYؾ����&�
�>��      �� �k��>��=���������0���s���:�N9���ʽZ����G��8��-��z5S�v���/X���D��Ad:�A�:� ;y�4;	�?;#~D;q�F;4xG;��G;�H;NOH;IsH;:�H;�H;�H;W�H;��H;U�H;��H;W�H;�H;�H;:�H;IsH;NOH;�H;��G;4xG;q�F;#~D;	�?;y�4;� ;�A�:�Ad:��D��/X�v��z5S��-���8���G�Z����ʽN9���:��s��0��������=��>��k��      .Eb�I]�tN�ߛ7����e� �{�˾��	�j��!,�J���0��m���,˼��x�E���1��_���U�:g�:3;��1;o+>;��C;�vF;�G;��G;>H;�gH;Z�H;w�H;9�H;�H;��H;(�H;��H;(�H;��H;�H;9�H;w�H;Z�H;�gH;>H;��G;�G;�vF;��C;o+>;��1;3;g�:U�:_����1��E����x�,˼��m�0��J����!,�	�j���{�˾e� ����ߛ7�tN�I]�      I]�N�W��TI�v3��D�������Ǿb���ȟf� )� ��W;���Fi��k�x�Ǽ�[t�8�	�(Ȅ�rX��ҟ:���:&�;�I2;�Y>;qD;�~F;\�G;,H;�>H;�hH;�H;�H;r�H;7�H;��H;S�H;��H;S�H;��H;7�H;r�H;�H;�H;�hH;�>H;,H;\�G;�~F;qD;�Y>;�I2;&�;���:ҟ:rX��(Ȅ�8�	��[t�x�Ǽ�k��Fi�W;�� �� )�ȟf�b�����Ǿ�����D�v3��TI�N�W�      tN��TI���;��'��k���i���f󐾖Z��K ��s�&����&^����"����g����Шu�Q!���1<:��:n
;�f3;-�>;�AD;֕F;�G;�H;UAH;jH;]�H;��H;(�H;ԻH;k�H;��H;B�H;��H;k�H;ԻH;(�H;��H;]�H;jH;UAH;�H;�G;֕F;�AD;-�>;�f3;n
;��:�1<:Q!��Шu������g��"�����&^�&����s潎K ��Z�f�i������k��'���;��TI�      ߛ7�v3��'����e� ��{Ծ
���6���]�F�����ӽ���;�L�1v�x뮼,T�Ƙ��PV�m�=�5(i:a��:"z ;�#5;�?;2�D;�F;�G;�H;�EH;�mH;��H;~�H;j�H;ۼH;4�H;P�H;��H;P�H;4�H;ۼH;j�H;~�H;��H;�mH;�EH;�H;�G;�F;2�D;�?;�#5;"z ;a��:5(i:m�=��PV�Ƙ�,T�x뮼1v�;�L�����ӽ���]�F�6���
����{Ծe� �����'�v3�      ����D��k�e� �<�ݾS���C͓�ȟf��>/�x��~'��n섽/�6�Rt��v��?�:�Tʻ�.�ݷ��s�:2;�$;�X7;��@;	E;;�F;Q�G;�H;EKH;�qH;��H;ʣH;�H;�H;/�H;E�H;��H;E�H;/�H;�H;�H;ʣH;��H;�qH;EKH;�H;Q�G;;�F;	E;��@;�X7;�$;2;�s�:ݷ��.�Tʻ?�:��v��Rt�/�6�n섽~'��x���>/�ȟf�C͓�S���<�ݾe� ��k��D�      e� ������쾻{ԾS���b���9�x�rSC��^�ͻ޽%���Q�e����ѼG������R�����դ8��:�X;��);6�9;.�A;��E;�G;3�G;t H;ERH;�vH;w�H;��H;:�H;��H;r�H;v�H;��H;v�H;r�H;��H;:�H;��H;w�H;�vH;ERH;t H;3�G;�G;��E;.�A;6�9;��);�X;��:դ8����R�����G���Ѽ��Q�e�%���ͻ޽�^�rSC�9�x�b���S����{Ծ�쾃���      {�˾��Ǿi���
���C͓�9�x�ؘJ��K �H��� �������?���t뮼�[�����3|��W��?�:w~�:	';�
/;�f<;�C;� F;�MG;��G;:,H;sZH;�|H;ȖH;éH;��H;��H;��H;��H;��H;��H;��H;��H;��H;éH;ȖH;�|H;sZH;:,H;��G;�MG;� F;�C;�f<;�
/;	';w~�:?�:�W��3|������[�t뮼����?���� ��H����K �ؘJ�9�x�C͓�
���i�����Ǿ      ��b���f�6���ȟf�rSC��K �Gn����Ž����Z��k��|ռX��Ey-����w.�q���O�:�*�:��;p4;t�>;*D;�vF;I�G;��G;�8H;\cH;x�H;��H;\�H;e�H;��H;��H;K�H;g�H;K�H;��H;��H;e�H;\�H;��H;x�H;\cH;�8H;��G;I�G;�vF;*D;t�>;p4;��;�*�:�O�:q��w.����Ey-�X���|ռ�k��Z������ŽGn���K �rSC�ȟf�6���f�b���      	�j�ȟf��Z�]�F��>/��^�H�����Ž- ���Fi�kQ+�Nt�PT��G�W�����1��hȺ�U�9�O�:
Y;��(;T�8;2A;�E;"�F;|�G;�H;�EH;�lH;��H;��H;8�H;d�H;��H;��H;��H;��H;��H;��H;��H;d�H;8�H;��H;��H;�lH;�EH;�H;|�G;"�F;�E;2A;T�8;��(;
Y;�O�:�U�9hȺ�1�����G�W�PT��Nt�kQ+��Fi�- ����ŽH����^��>/�]�F��Z�ȟf�      �!,� )��K ����x��ͻ޽ ������Fi���0�����跼z�x�����.��a�(�����)i:���:��;�0;��<;�C;��E;*<G;�G;�#H;kSH;�vH;�H;�H;F�H;u�H;4�H;��H;��H;n�H;��H;��H;4�H;u�H;F�H;�H;�H;�vH;kSH;�#H;�G;*<G;��E;�C;��<;�0;��;���:�)i:���a�(��.�����z�x��跼�����0��Fi���� ��ͻ޽x������K � )�      J��� ��s��ӽ~'��%�������Z�kQ+�����"��G����0���׻̕b��W���V�9���:�_;�)';0Y7;H#@;T�D;�F;+�G;��G;A7H;aH;��H;Z�H;��H;l�H;��H;��H;{�H;B�H;.�H;B�H;{�H;��H;��H;l�H;��H;Z�H;��H;aH;A7H;��G;+�G;�F;T�D;H#@;0Y7;�)';�_;���:�V�9�W��̕b���׻��0�G���"�����kQ+��Z����%���~'���ӽ�s� ��      0��W;��&������n섽Q�e���?��k�Nt��跼G��ee7�����Ǆ��0��t�`t�: +�:�
;�1;��<;��B;N�E;G;�G;jH;wIH;`nH;��H;��H;�H;��H;��H;�H;��H;�H;��H;�H;��H;�H;��H;��H;�H;��H;��H;`nH;wIH;jH;�G;G;N�E;��B;��<;�1;�
; +�:`t�:�t��0��Ǆ����ee7�G���跼Nt�k���?�Q�e�n섽���&���W;��      m��Fi��&^�;�L�/�6������|ռPT��z�x���0��������0���ڷ�{m`:��:��;��*;~�8;G�@;e�D;��F;}G;��G;�0H;�ZH;n{H;��H;קH;�H;��H;��H;|�H;��H;��H;e�H;��H;��H;|�H;��H;��H;�H;קH;��H;n{H;�ZH;�0H;��G;}G;��F;e�D;G�@;~�8;��*;��;��:{m`:�ڷ�0��������껢�0�z�x�PT���|ռ����/�6�;�L��&^��Fi�      ���k���1v�Rt��Ѽt뮼X��G�W������׻�Ǆ�0�����3<:x��:;Y;�s%;=$5;�Y>;.`C;��E;O)G;v�G;#H;GH;lkH;�H;��H;��H;ȻH;��H;��H;��H;g�H;_�H;�H;_�H;g�H;��H;��H;��H;ȻH;��H;��H;�H;lkH;GH;#H;v�G;O)G;��E;.`C;�Y>;=$5;�s%;;Y;x��:�3<:���0���Ǆ���׻���G�W�X��t뮼�ѼRt�1v����k�      ,˼x�Ǽ�"��x뮼�v��G���[�Ey-�����.��̕b��0㺂ڷ��3<:L�:_\;��!;2J2;�f<;�/B;RBE;K�F;a�G; �G;�3H;�[H;{H;��H;��H;P�H;��H;6�H;��H;B�H;A�H;��H;��H;��H;A�H;B�H;��H;6�H;��H;P�H;��H;��H;{H;�[H;�3H; �G;a�G;K�F;RBE;�/B;�f<;2J2;��!;_\;L�:�3<:�ڷ��0�̕b��.�����Ey-��[�G���v��x뮼�"��x�Ǽ      ��x��[t���g�,T�?�:������������1��a�(��W���t�{m`:x��:_\;qz ;�0;�;;:<A;?�D;�vF;�bG;e�G;� H;�LH;�nH;p�H;~�H;��H;��H;Z�H;��H;I�H;_�H;��H;��H;�H;��H;��H;_�H;I�H;��H;Z�H;��H;��H;~�H;p�H;�nH;�LH;� H;e�G;�bG;�vF;?�D;:<A;�;;�0;qz ;_\;x��:{m`:�t��W��a�(��1������������?�:�,T���g��[t�      E��8�	����Ƙ�Tʻ�R��3|�w.�hȺ����V�9`t�:��:;Y;��!;�0;.�:;�@;5BD;�1F;�7G;��G;�H;k?H;+cH;�H;n�H;;�H;<�H;>�H;��H;��H;��H;[�H;��H;��H;s�H;��H;��H;[�H;��H;��H;��H;>�H;<�H;;�H;n�H;�H;+cH;k?H;�H;��G;�7G;�1F;5BD;�@;.�:;�0;��!;;Y;��:`t�:�V�9���hȺw.�3|��R��TʻƘ����8�	�      �1��(Ȅ�Шu��PV��.�����W��q��U�9�)i:���: +�:��;�s%;2J2;�;;�@;�D;/F;?G;��G;�H;�4H;�YH;5wH;7�H;�H;	�H;�H;I�H;^�H;�H;�H;�H;*�H;E�H;��H;E�H;*�H;�H;�H;�H;^�H;I�H;�H;	�H;�H;7�H;5wH;�YH;�4H;�H;��G;?G;/F;�D;�@;�;;2J2;�s%;��; +�:���:�)i:�U�9q���W������.��PV�Шu�(Ȅ�      _���rX��Q!��m�=�ݷ�դ8?�:�O�:�O�:���:�_;�
;��*;=$5;�f<;:<A;5BD;/F;�G;��G;r�G;�,H;RH;UpH;�H;��H;r�H;�H;)�H;��H;��H;��H;?�H;��H;��H;|�H;��H;|�H;��H;��H;?�H;��H;��H;��H;)�H;�H;r�H;��H;�H;UpH;RH;�,H;r�G;��G;�G;/F;5BD;:<A;�f<;=$5;��*;�
;�_;���:�O�:�O�:?�:դ8ݷ�m�=�Q!��rX��      U�:ҟ:�1<:5(i:�s�:��:w~�:�*�:
Y;��;�)';�1;~�8;�Y>;�/B;?�D;�1F;?G;��G;&�G;�(H;�MH;qkH;D�H;c�H;v�H;��H;�H;t�H;��H;$�H;�H;�H;D�H;��H;��H;��H;��H;��H;D�H;�H;�H;$�H;��H;t�H;�H;��H;v�H;c�H;D�H;qkH;�MH;�(H;&�G;��G;?G;�1F;?�D;�/B;�Y>;~�8;�1;�)';��;
Y;�*�:w~�:��:�s�:5(i:�1<:ҟ:      g�:���:��:a��:2;�X;	';��;��(;�0;0Y7;��<;G�@;.`C;RBE;�vF;�7G;��G;r�G;�(H;�KH;�hH;.�H;O�H;��H;��H;��H;O�H;�H;��H;��H;A�H;��H;��H;��H;��H;��H;��H;��H;��H;��H;A�H;��H;��H;�H;O�H;��H;��H;��H;O�H;.�H;�hH;�KH;�(H;r�G;��G;�7G;�vF;RBE;.`C;G�@;��<;0Y7;�0;��(;��;	';�X;2;a��:��:���:      3;&�;n
;"z ;�$;��);�
/;p4;T�8;��<;H#@;��B;e�D;��E;K�F;�bG;��G;�H;�,H;�MH;�hH;B�H;��H;��H;ΰH;��H;��H;��H;2�H;��H;^�H;�H;1�H;��H;��H;P�H;��H;P�H;��H;��H;1�H;�H;^�H;��H;2�H;��H;��H;��H;ΰH;��H;��H;B�H;�hH;�MH;�,H;�H;��G;�bG;K�F;��E;e�D;��B;H#@;��<;T�8;p4;�
/;��);�$;"z ;n
;&�;      ��1;�I2;�f3;�#5;�X7;6�9;�f<;t�>;2A;�C;T�D;N�E;��F;O)G;a�G;e�G;�H;�4H;RH;qkH;.�H;��H;�H;ɯH;��H;V�H;L�H; �H;��H;��H;u�H;��H;o�H;��H;��H;�H;\�H;�H;��H;��H;o�H;��H;u�H;��H;��H; �H;L�H;V�H;��H;ɯH;�H;��H;.�H;qkH;RH;�4H;�H;e�G;a�G;O)G;��F;N�E;T�D;�C;2A;t�>;�f<;6�9;�X7;�#5;�f3;�I2;      o+>;�Y>;-�>;�?;��@;.�A;�C;*D;�E;��E;�F;G;}G;v�G; �G;� H;k?H;�YH;UpH;D�H;O�H;��H;ɯH;�H;��H;��H;6�H;��H;��H;��H;P�H; �H;��H;��H;H�H;��H;��H;��H;H�H;��H;��H; �H;P�H;��H;��H;��H;6�H;��H;��H;�H;ɯH;��H;O�H;D�H;UpH;�YH;k?H;� H; �G;v�G;}G;G;�F;��E;�E;*D;�C;.�A;��@;�?;-�>;�Y>;      ��C;qD;�AD;2�D;	E;��E;� F;�vF;"�F;*<G;+�G;�G;��G;#H;�3H;�LH;+cH;5wH;�H;c�H;��H;ΰH;��H;��H;=�H;��H;��H;^�H;c�H;��H;��H;g�H;��H;@�H;��H;D�H;L�H;D�H;��H;@�H;��H;g�H;��H;��H;c�H;^�H;��H;��H;=�H;��H;��H;ΰH;��H;c�H;�H;5wH;+cH;�LH;�3H;#H;��G;�G;+�G;*<G;"�F;�vF;� F;��E;	E;2�D;�AD;qD;      �vF;�~F;֕F;�F;;�F;�G;�MG;I�G;|�G;�G;��G;jH;�0H;GH;�[H;�nH;�H;7�H;��H;v�H;��H;��H;V�H;��H;��H;W�H;$�H;�H;��H;��H;�H;T�H;6�H;��H;m�H;��H;��H;��H;m�H;��H;6�H;T�H;�H;��H;��H;�H;$�H;W�H;��H;��H;V�H;��H;��H;v�H;��H;7�H;�H;�nH;�[H;GH;�0H;jH;��G;�G;|�G;I�G;�MG;�G;;�F;�F;֕F;�~F;      �G;\�G;�G;�G;Q�G;3�G;��G;��G;�H;�#H;A7H;wIH;�ZH;lkH;{H;p�H;n�H;�H;r�H;��H;��H;��H;L�H;6�H;��H;$�H;�H;h�H;J�H;��H;7�H;�H;��H;��H;��H;�H;�H;�H;��H;��H;��H;�H;7�H;��H;J�H;h�H;�H;$�H;��H;6�H;L�H;��H;��H;��H;r�H;�H;n�H;p�H;{H;lkH;�ZH;wIH;A7H;�#H;�H;��G;��G;3�G;Q�G;�G;�G;\�G;      ��G;,H;�H;�H;�H;t H;:,H;�8H;�EH;kSH;aH;`nH;n{H;�H;��H;~�H;;�H;	�H;�H;�H;O�H;��H; �H;��H;^�H;�H;h�H;]�H;��H;�H;�H;��H;z�H;��H;�H;^�H;g�H;^�H;�H;��H;z�H;��H;�H;�H;��H;]�H;h�H;�H;^�H;��H; �H;��H;O�H;�H;�H;	�H;;�H;~�H;��H;�H;n{H;`nH;aH;kSH;�EH;�8H;:,H;t H;�H;�H;�H;,H;      >H;�>H;UAH;�EH;EKH;ERH;sZH;\cH;�lH;�vH;��H;��H;��H;��H;��H;��H;<�H;�H;)�H;t�H;�H;2�H;��H;��H;c�H;��H;J�H;��H;$�H;��H;��H;k�H;��H;6�H;p�H;��H;��H;��H;p�H;6�H;��H;k�H;��H;��H;$�H;��H;J�H;��H;c�H;��H;��H;2�H;�H;t�H;)�H;�H;<�H;��H;��H;��H;��H;��H;��H;�vH;�lH;\cH;sZH;ERH;EKH;�EH;UAH;�>H;      �gH;�hH;jH;�mH;�qH;�vH;�|H;x�H;��H;�H;Z�H;��H;קH;��H;P�H;��H;>�H;I�H;��H;��H;��H;��H;��H;��H;��H;��H;��H;�H;��H;��H;t�H;��H;%�H;z�H;��H;��H;��H;��H;��H;z�H;%�H;��H;t�H;��H;��H;�H;��H;��H;��H;��H;��H;��H;��H;��H;��H;I�H;>�H;��H;P�H;��H;קH;��H;Z�H;�H;��H;x�H;�|H;�vH;�qH;�mH;jH;�hH;      Z�H;�H;]�H;��H;��H;w�H;ȖH;��H;��H;�H;��H;�H;�H;ȻH;��H;Z�H;��H;^�H;��H;$�H;��H;^�H;u�H;P�H;��H;�H;7�H;�H;��H;t�H;��H;.�H;��H;��H;��H;��H;��H;��H;��H;��H;��H;.�H;��H;t�H;��H;�H;7�H;�H;��H;P�H;u�H;^�H;��H;$�H;��H;^�H;��H;Z�H;��H;ȻH;�H;�H;��H;�H;��H;��H;ȖH;w�H;��H;��H;]�H;�H;      w�H;�H;��H;~�H;ʣH;��H;éH;\�H;8�H;F�H;l�H;��H;��H;��H;6�H;��H;��H;�H;��H;�H;A�H;�H;��H; �H;g�H;T�H;�H;��H;k�H;��H;.�H;{�H;��H;��H;��H;�H;�H;�H;��H;��H;��H;{�H;.�H;��H;k�H;��H;�H;T�H;g�H; �H;��H;�H;A�H;�H;��H;�H;��H;��H;6�H;��H;��H;��H;l�H;F�H;8�H;\�H;éH;��H;ʣH;~�H;��H;�H;      9�H;r�H;(�H;j�H;�H;:�H;��H;e�H;d�H;u�H;��H;��H;��H;��H;��H;I�H;��H;�H;?�H;�H;��H;1�H;o�H;��H;��H;6�H;��H;z�H;��H;%�H;��H;��H;��H;��H;�H;�H;�H;�H;�H;��H;��H;��H;��H;%�H;��H;z�H;��H;6�H;��H;��H;o�H;1�H;��H;�H;?�H;�H;��H;I�H;��H;��H;��H;��H;��H;u�H;d�H;e�H;��H;:�H;�H;j�H;(�H;r�H;      �H;7�H;ԻH;ۼH;�H;��H;��H;��H;��H;4�H;��H;�H;|�H;��H;B�H;_�H;[�H;�H;��H;D�H;��H;��H;��H;��H;@�H;��H;��H;��H;6�H;z�H;��H;��H;��H; �H;.�H;9�H;�H;9�H;.�H; �H;��H;��H;��H;z�H;6�H;��H;��H;��H;@�H;��H;��H;��H;��H;D�H;��H;�H;[�H;_�H;B�H;��H;|�H;�H;��H;4�H;��H;��H;��H;��H;�H;ۼH;ԻH;7�H;      ��H;��H;k�H;4�H;/�H;r�H;��H;��H;��H;��H;{�H;��H;��H;g�H;A�H;��H;��H;*�H;��H;��H;��H;��H;��H;H�H;��H;m�H;��H;�H;p�H;��H;��H;��H;�H;.�H;�H;.�H;J�H;.�H;�H;.�H;�H;��H;��H;��H;p�H;�H;��H;m�H;��H;H�H;��H;��H;��H;��H;��H;*�H;��H;��H;A�H;g�H;��H;��H;{�H;��H;��H;��H;��H;r�H;/�H;4�H;k�H;��H;      (�H;S�H;��H;P�H;E�H;v�H;��H;K�H;��H;��H;B�H;�H;��H;_�H;��H;��H;��H;E�H;|�H;��H;��H;P�H;�H;��H;D�H;��H;�H;^�H;��H;��H;��H;�H;�H;9�H;.�H;$�H;6�H;$�H;.�H;9�H;�H;�H;��H;��H;��H;^�H;�H;��H;D�H;��H;�H;P�H;��H;��H;|�H;E�H;��H;��H;��H;_�H;��H;�H;B�H;��H;��H;K�H;��H;v�H;E�H;P�H;��H;S�H;      ��H;��H;B�H;��H;��H;��H;��H;g�H;��H;n�H;.�H;��H;e�H;�H;��H;�H;s�H;��H;��H;��H;��H;��H;\�H;��H;L�H;��H;�H;g�H;��H;��H;��H;�H;�H;�H;J�H;6�H;#�H;6�H;J�H;�H;�H;�H;��H;��H;��H;g�H;�H;��H;L�H;��H;\�H;��H;��H;��H;��H;��H;s�H;�H;��H;�H;e�H;��H;.�H;n�H;��H;g�H;��H;��H;��H;��H;B�H;��H;      (�H;S�H;��H;P�H;E�H;v�H;��H;K�H;��H;��H;B�H;�H;��H;_�H;��H;��H;��H;E�H;|�H;��H;��H;P�H;�H;��H;D�H;��H;�H;^�H;��H;��H;��H;�H;�H;9�H;.�H;$�H;6�H;$�H;.�H;9�H;�H;�H;��H;��H;��H;^�H;�H;��H;D�H;��H;�H;P�H;��H;��H;|�H;E�H;��H;��H;��H;_�H;��H;�H;B�H;��H;��H;K�H;��H;v�H;E�H;P�H;��H;S�H;      ��H;��H;k�H;4�H;/�H;r�H;��H;��H;��H;��H;{�H;��H;��H;g�H;A�H;��H;��H;*�H;��H;��H;��H;��H;��H;H�H;��H;m�H;��H;�H;p�H;��H;��H;��H;�H;.�H;�H;.�H;J�H;.�H;�H;.�H;�H;��H;��H;��H;p�H;�H;��H;m�H;��H;H�H;��H;��H;��H;��H;��H;*�H;��H;��H;A�H;g�H;��H;��H;{�H;��H;��H;��H;��H;r�H;/�H;4�H;k�H;��H;      �H;7�H;ԻH;ۼH;�H;��H;��H;��H;��H;4�H;��H;�H;|�H;��H;B�H;_�H;[�H;�H;��H;D�H;��H;��H;��H;��H;@�H;��H;��H;��H;6�H;z�H;��H;��H;��H; �H;.�H;9�H;�H;9�H;.�H; �H;��H;��H;��H;z�H;6�H;��H;��H;��H;@�H;��H;��H;��H;��H;D�H;��H;�H;[�H;_�H;B�H;��H;|�H;�H;��H;4�H;��H;��H;��H;��H;�H;ۼH;ԻH;7�H;      9�H;r�H;(�H;j�H;�H;:�H;��H;e�H;d�H;u�H;��H;��H;��H;��H;��H;I�H;��H;�H;?�H;�H;��H;1�H;o�H;��H;��H;6�H;��H;z�H;��H;%�H;��H;��H;��H;��H;�H;�H;�H;�H;�H;��H;��H;��H;��H;%�H;��H;z�H;��H;6�H;��H;��H;o�H;1�H;��H;�H;?�H;�H;��H;I�H;��H;��H;��H;��H;��H;u�H;d�H;e�H;��H;:�H;�H;j�H;(�H;r�H;      w�H;�H;��H;~�H;ʣH;��H;éH;\�H;8�H;F�H;l�H;��H;��H;��H;6�H;��H;��H;�H;��H;�H;A�H;�H;��H; �H;g�H;T�H;�H;��H;k�H;��H;.�H;{�H;��H;��H;��H;�H;�H;�H;��H;��H;��H;{�H;.�H;��H;k�H;��H;�H;T�H;g�H; �H;��H;�H;A�H;�H;��H;�H;��H;��H;6�H;��H;��H;��H;l�H;F�H;8�H;\�H;éH;��H;ʣH;~�H;��H;�H;      Z�H;�H;]�H;��H;��H;w�H;ȖH;��H;��H;�H;��H;�H;�H;ȻH;��H;Z�H;��H;^�H;��H;$�H;��H;^�H;u�H;P�H;��H;�H;7�H;�H;��H;t�H;��H;.�H;��H;��H;��H;��H;��H;��H;��H;��H;��H;.�H;��H;t�H;��H;�H;7�H;�H;��H;P�H;u�H;^�H;��H;$�H;��H;^�H;��H;Z�H;��H;ȻH;�H;�H;��H;�H;��H;��H;ȖH;w�H;��H;��H;]�H;�H;      �gH;�hH;jH;�mH;�qH;�vH;�|H;x�H;��H;�H;Z�H;��H;קH;��H;P�H;��H;>�H;I�H;��H;��H;��H;��H;��H;��H;��H;��H;��H;�H;��H;��H;t�H;��H;%�H;z�H;��H;��H;��H;��H;��H;z�H;%�H;��H;t�H;��H;��H;�H;��H;��H;��H;��H;��H;��H;��H;��H;��H;I�H;>�H;��H;P�H;��H;קH;��H;Z�H;�H;��H;x�H;�|H;�vH;�qH;�mH;jH;�hH;      >H;�>H;UAH;�EH;EKH;ERH;sZH;\cH;�lH;�vH;��H;��H;��H;��H;��H;��H;<�H;�H;)�H;t�H;�H;2�H;��H;��H;c�H;��H;J�H;��H;$�H;��H;��H;k�H;��H;6�H;p�H;��H;��H;��H;p�H;6�H;��H;k�H;��H;��H;$�H;��H;J�H;��H;c�H;��H;��H;2�H;�H;t�H;)�H;�H;<�H;��H;��H;��H;��H;��H;��H;�vH;�lH;\cH;sZH;ERH;EKH;�EH;UAH;�>H;      ��G;,H;�H;�H;�H;t H;:,H;�8H;�EH;kSH;aH;`nH;n{H;�H;��H;~�H;;�H;	�H;�H;�H;O�H;��H; �H;��H;^�H;�H;h�H;]�H;��H;�H;�H;��H;z�H;��H;�H;^�H;g�H;^�H;�H;��H;z�H;��H;�H;�H;��H;]�H;h�H;�H;^�H;��H; �H;��H;O�H;�H;�H;	�H;;�H;~�H;��H;�H;n{H;`nH;aH;kSH;�EH;�8H;:,H;t H;�H;�H;�H;,H;      �G;\�G;�G;�G;Q�G;3�G;��G;��G;�H;�#H;A7H;wIH;�ZH;lkH;{H;p�H;n�H;�H;r�H;��H;��H;��H;L�H;6�H;��H;$�H;�H;h�H;J�H;��H;7�H;�H;��H;��H;��H;�H;�H;�H;��H;��H;��H;�H;7�H;��H;J�H;h�H;�H;$�H;��H;6�H;L�H;��H;��H;��H;r�H;�H;n�H;p�H;{H;lkH;�ZH;wIH;A7H;�#H;�H;��G;��G;3�G;Q�G;�G;�G;\�G;      �vF;�~F;֕F;�F;;�F;�G;�MG;I�G;|�G;�G;��G;jH;�0H;GH;�[H;�nH;�H;7�H;��H;v�H;��H;��H;V�H;��H;��H;W�H;$�H;�H;��H;��H;�H;T�H;6�H;��H;m�H;��H;��H;��H;m�H;��H;6�H;T�H;�H;��H;��H;�H;$�H;W�H;��H;��H;V�H;��H;��H;v�H;��H;7�H;�H;�nH;�[H;GH;�0H;jH;��G;�G;|�G;I�G;�MG;�G;;�F;�F;֕F;�~F;      ��C;qD;�AD;2�D;	E;��E;� F;�vF;"�F;*<G;+�G;�G;��G;#H;�3H;�LH;+cH;5wH;�H;c�H;��H;ΰH;��H;��H;=�H;��H;��H;^�H;c�H;��H;��H;g�H;��H;@�H;��H;D�H;L�H;D�H;��H;@�H;��H;g�H;��H;��H;c�H;^�H;��H;��H;=�H;��H;��H;ΰH;��H;c�H;�H;5wH;+cH;�LH;�3H;#H;��G;�G;+�G;*<G;"�F;�vF;� F;��E;	E;2�D;�AD;qD;      o+>;�Y>;-�>;�?;��@;.�A;�C;*D;�E;��E;�F;G;}G;v�G; �G;� H;k?H;�YH;UpH;D�H;O�H;��H;ɯH;�H;��H;��H;6�H;��H;��H;��H;P�H; �H;��H;��H;H�H;��H;��H;��H;H�H;��H;��H; �H;P�H;��H;��H;��H;6�H;��H;��H;�H;ɯH;��H;O�H;D�H;UpH;�YH;k?H;� H; �G;v�G;}G;G;�F;��E;�E;*D;�C;.�A;��@;�?;-�>;�Y>;      ��1;�I2;�f3;�#5;�X7;6�9;�f<;t�>;2A;�C;T�D;N�E;��F;O)G;a�G;e�G;�H;�4H;RH;qkH;.�H;��H;�H;ɯH;��H;V�H;L�H; �H;��H;��H;u�H;��H;o�H;��H;��H;�H;\�H;�H;��H;��H;o�H;��H;u�H;��H;��H; �H;L�H;V�H;��H;ɯH;�H;��H;.�H;qkH;RH;�4H;�H;e�G;a�G;O)G;��F;N�E;T�D;�C;2A;t�>;�f<;6�9;�X7;�#5;�f3;�I2;      3;&�;n
;"z ;�$;��);�
/;p4;T�8;��<;H#@;��B;e�D;��E;K�F;�bG;��G;�H;�,H;�MH;�hH;B�H;��H;��H;ΰH;��H;��H;��H;2�H;��H;^�H;�H;1�H;��H;��H;P�H;��H;P�H;��H;��H;1�H;�H;^�H;��H;2�H;��H;��H;��H;ΰH;��H;��H;B�H;�hH;�MH;�,H;�H;��G;�bG;K�F;��E;e�D;��B;H#@;��<;T�8;p4;�
/;��);�$;"z ;n
;&�;      g�:���:��:a��:2;�X;	';��;��(;�0;0Y7;��<;G�@;.`C;RBE;�vF;�7G;��G;r�G;�(H;�KH;�hH;.�H;O�H;��H;��H;��H;O�H;�H;��H;��H;A�H;��H;��H;��H;��H;��H;��H;��H;��H;��H;A�H;��H;��H;�H;O�H;��H;��H;��H;O�H;.�H;�hH;�KH;�(H;r�G;��G;�7G;�vF;RBE;.`C;G�@;��<;0Y7;�0;��(;��;	';�X;2;a��:��:���:      U�:ҟ:�1<:5(i:�s�:��:w~�:�*�:
Y;��;�)';�1;~�8;�Y>;�/B;?�D;�1F;?G;��G;&�G;�(H;�MH;qkH;D�H;c�H;v�H;��H;�H;t�H;��H;$�H;�H;�H;D�H;��H;��H;��H;��H;��H;D�H;�H;�H;$�H;��H;t�H;�H;��H;v�H;c�H;D�H;qkH;�MH;�(H;&�G;��G;?G;�1F;?�D;�/B;�Y>;~�8;�1;�)';��;
Y;�*�:w~�:��:�s�:5(i:�1<:ҟ:      _���rX��Q!��m�=�ݷ�դ8?�:�O�:�O�:���:�_;�
;��*;=$5;�f<;:<A;5BD;/F;�G;��G;r�G;�,H;RH;UpH;�H;��H;r�H;�H;)�H;��H;��H;��H;?�H;��H;��H;|�H;��H;|�H;��H;��H;?�H;��H;��H;��H;)�H;�H;r�H;��H;�H;UpH;RH;�,H;r�G;��G;�G;/F;5BD;:<A;�f<;=$5;��*;�
;�_;���:�O�:�O�:?�:դ8ݷ�m�=�Q!��rX��      �1��(Ȅ�Шu��PV��.�����W��q��U�9�)i:���: +�:��;�s%;2J2;�;;�@;�D;/F;?G;��G;�H;�4H;�YH;5wH;7�H;�H;	�H;�H;I�H;^�H;�H;�H;�H;*�H;E�H;��H;E�H;*�H;�H;�H;�H;^�H;I�H;�H;	�H;�H;7�H;5wH;�YH;�4H;�H;��G;?G;/F;�D;�@;�;;2J2;�s%;��; +�:���:�)i:�U�9q���W������.��PV�Шu�(Ȅ�      E��8�	����Ƙ�Tʻ�R��3|�w.�hȺ����V�9`t�:��:;Y;��!;�0;.�:;�@;5BD;�1F;�7G;��G;�H;k?H;+cH;�H;n�H;;�H;<�H;>�H;��H;��H;��H;[�H;��H;��H;s�H;��H;��H;[�H;��H;��H;��H;>�H;<�H;;�H;n�H;�H;+cH;k?H;�H;��G;�7G;�1F;5BD;�@;.�:;�0;��!;;Y;��:`t�:�V�9���hȺw.�3|��R��TʻƘ����8�	�      ��x��[t���g�,T�?�:������������1��a�(��W���t�{m`:x��:_\;qz ;�0;�;;:<A;?�D;�vF;�bG;e�G;� H;�LH;�nH;p�H;~�H;��H;��H;Z�H;��H;I�H;_�H;��H;��H;�H;��H;��H;_�H;I�H;��H;Z�H;��H;��H;~�H;p�H;�nH;�LH;� H;e�G;�bG;�vF;?�D;:<A;�;;�0;qz ;_\;x��:{m`:�t��W��a�(��1������������?�:�,T���g��[t�      ,˼x�Ǽ�"��x뮼�v��G���[�Ey-�����.��̕b��0㺂ڷ��3<:L�:_\;��!;2J2;�f<;�/B;RBE;K�F;a�G; �G;�3H;�[H;{H;��H;��H;P�H;��H;6�H;��H;B�H;A�H;��H;��H;��H;A�H;B�H;��H;6�H;��H;P�H;��H;��H;{H;�[H;�3H; �G;a�G;K�F;RBE;�/B;�f<;2J2;��!;_\;L�:�3<:�ڷ��0�̕b��.�����Ey-��[�G���v��x뮼�"��x�Ǽ      ���k���1v�Rt��Ѽt뮼X��G�W������׻�Ǆ�0�����3<:x��:;Y;�s%;=$5;�Y>;.`C;��E;O)G;v�G;#H;GH;lkH;�H;��H;��H;ȻH;��H;��H;��H;g�H;_�H;�H;_�H;g�H;��H;��H;��H;ȻH;��H;��H;�H;lkH;GH;#H;v�G;O)G;��E;.`C;�Y>;=$5;�s%;;Y;x��:�3<:���0���Ǆ���׻���G�W�X��t뮼�ѼRt�1v����k�      m��Fi��&^�;�L�/�6������|ռPT��z�x���0��������0���ڷ�{m`:��:��;��*;~�8;G�@;e�D;��F;}G;��G;�0H;�ZH;n{H;��H;קH;�H;��H;��H;|�H;��H;��H;e�H;��H;��H;|�H;��H;��H;�H;קH;��H;n{H;�ZH;�0H;��G;}G;��F;e�D;G�@;~�8;��*;��;��:{m`:�ڷ�0��������껢�0�z�x�PT���|ռ����/�6�;�L��&^��Fi�      0��W;��&������n섽Q�e���?��k�Nt��跼G��ee7�����Ǆ��0��t�`t�: +�:�
;�1;��<;��B;N�E;G;�G;jH;wIH;`nH;��H;��H;�H;��H;��H;�H;��H;�H;��H;�H;��H;�H;��H;��H;�H;��H;��H;`nH;wIH;jH;�G;G;N�E;��B;��<;�1;�
; +�:`t�:�t��0��Ǆ����ee7�G���跼Nt�k���?�Q�e�n섽���&���W;��      J��� ��s��ӽ~'��%�������Z�kQ+�����"��G����0���׻̕b��W���V�9���:�_;�)';0Y7;H#@;T�D;�F;+�G;��G;A7H;aH;��H;Z�H;��H;l�H;��H;��H;{�H;B�H;.�H;B�H;{�H;��H;��H;l�H;��H;Z�H;��H;aH;A7H;��G;+�G;�F;T�D;H#@;0Y7;�)';�_;���:�V�9�W��̕b���׻��0�G���"�����kQ+��Z����%���~'���ӽ�s� ��      �!,� )��K ����x��ͻ޽ ������Fi���0�����跼z�x�����.��a�(�����)i:���:��;�0;��<;�C;��E;*<G;�G;�#H;kSH;�vH;�H;�H;F�H;u�H;4�H;��H;��H;n�H;��H;��H;4�H;u�H;F�H;�H;�H;�vH;kSH;�#H;�G;*<G;��E;�C;��<;�0;��;���:�)i:���a�(��.�����z�x��跼�����0��Fi���� ��ͻ޽x������K � )�      	�j�ȟf��Z�]�F��>/��^�H�����Ž- ���Fi�kQ+�Nt�PT��G�W�����1��hȺ�U�9�O�:
Y;��(;T�8;2A;�E;"�F;|�G;�H;�EH;�lH;��H;��H;8�H;d�H;��H;��H;��H;��H;��H;��H;��H;d�H;8�H;��H;��H;�lH;�EH;�H;|�G;"�F;�E;2A;T�8;��(;
Y;�O�:�U�9hȺ�1�����G�W�PT��Nt�kQ+��Fi�- ����ŽH����^��>/�]�F��Z�ȟf�      ��b���f�6���ȟf�rSC��K �Gn����Ž����Z��k��|ռX��Ey-����w.�q���O�:�*�:��;p4;t�>;*D;�vF;I�G;��G;�8H;\cH;x�H;��H;\�H;e�H;��H;��H;K�H;g�H;K�H;��H;��H;e�H;\�H;��H;x�H;\cH;�8H;��G;I�G;�vF;*D;t�>;p4;��;�*�:�O�:q��w.����Ey-�X���|ռ�k��Z������ŽGn���K �rSC�ȟf�6���f�b���      {�˾��Ǿi���
���C͓�9�x�ؘJ��K �H��� �������?���t뮼�[�����3|��W��?�:w~�:	';�
/;�f<;�C;� F;�MG;��G;:,H;sZH;�|H;ȖH;éH;��H;��H;��H;��H;��H;��H;��H;��H;��H;éH;ȖH;�|H;sZH;:,H;��G;�MG;� F;�C;�f<;�
/;	';w~�:?�:�W��3|������[�t뮼����?���� ��H����K �ؘJ�9�x�C͓�
���i�����Ǿ      e� ������쾻{ԾS���b���9�x�rSC��^�ͻ޽%���Q�e����ѼG������R�����դ8��:�X;��);6�9;.�A;��E;�G;3�G;t H;ERH;�vH;w�H;��H;:�H;��H;r�H;v�H;��H;v�H;r�H;��H;:�H;��H;w�H;�vH;ERH;t H;3�G;�G;��E;.�A;6�9;��);�X;��:դ8����R�����G���Ѽ��Q�e�%���ͻ޽�^�rSC�9�x�b���S����{Ծ�쾃���      ����D��k�e� �<�ݾS���C͓�ȟf��>/�x��~'��n섽/�6�Rt��v��?�:�Tʻ�.�ݷ��s�:2;�$;�X7;��@;	E;;�F;Q�G;�H;EKH;�qH;��H;ʣH;�H;�H;/�H;E�H;��H;E�H;/�H;�H;�H;ʣH;��H;�qH;EKH;�H;Q�G;;�F;	E;��@;�X7;�$;2;�s�:ݷ��.�Tʻ?�:��v��Rt�/�6�n섽~'��x���>/�ȟf�C͓�S���<�ݾe� ��k��D�      ߛ7�v3��'����e� ��{Ծ
���6���]�F�����ӽ���;�L�1v�x뮼,T�Ƙ��PV�m�=�5(i:a��:"z ;�#5;�?;2�D;�F;�G;�H;�EH;�mH;��H;~�H;j�H;ۼH;4�H;P�H;��H;P�H;4�H;ۼH;j�H;~�H;��H;�mH;�EH;�H;�G;�F;2�D;�?;�#5;"z ;a��:5(i:m�=��PV�Ƙ�,T�x뮼1v�;�L�����ӽ���]�F�6���
����{Ծe� �����'�v3�      tN��TI���;��'��k���i���f󐾖Z��K ��s�&����&^����"����g����Шu�Q!���1<:��:n
;�f3;-�>;�AD;֕F;�G;�H;UAH;jH;]�H;��H;(�H;ԻH;k�H;��H;B�H;��H;k�H;ԻH;(�H;��H;]�H;jH;UAH;�H;�G;֕F;�AD;-�>;�f3;n
;��:�1<:Q!��Шu������g��"�����&^�&����s潎K ��Z�f�i������k��'���;��TI�      I]�N�W��TI�v3��D�������Ǿb���ȟf� )� ��W;���Fi��k�x�Ǽ�[t�8�	�(Ȅ�rX��ҟ:���:&�;�I2;�Y>;qD;�~F;\�G;,H;�>H;�hH;�H;�H;r�H;7�H;��H;S�H;��H;S�H;��H;7�H;r�H;�H;�H;�hH;�>H;,H;\�G;�~F;qD;�Y>;�I2;&�;���:ҟ:rX��(Ȅ�8�	��[t�x�Ǽ�k��Fi�W;�� �� )�ȟf�b�����Ǿ�����D�v3��TI�N�W�      �?��ph��2v��� ��$�X��O/�#y�-�;Ѱ��j+X�����ѽ����Gn;�>�＿����B(�嚩����2�e9��:^;Y.;��<;�VC;@ZF;�G;5/H;tiH;X�H;s�H;��H;F�H;��H;�H;��H;��H;��H;�H;��H;F�H;��H;s�H;X�H;tiH;5/H;�G;@ZF;�VC;��<;Y.;^;��:2�e9���嚩��B(�����>��Gn;�������ѽ��j+X�Ѱ��-�;#y��O/�$�X�� ��2v��ph��      ph��"���V�����y�EvS�aM+��v� 9ɾ�����T�]��[ν����`\8�����x���%�[��������9C,�:��;�.;N�<;!nC;�cF;�G;�0H;"jH;ȋH;ңH;��H;��H;��H;��H;��H;��H;��H;��H;��H;��H;��H;ңH;ȋH;"jH;�0H;�G;�cF;!nC;N�<;�.;��;C,�:��9���[����%��x�����`\8������[ν]��T����� 9ɾ�v�aM+�EvS���y�V���"���      2v��V���L ��M�h�%E�I��R���i㼾n���nH�È�a�ý�Ȅ��s/��o༼#�����3J���к��9$f�:Nl;�0;Q\=; �C;6�F;��G;Q5H;^lH;H�H;ФH;��H;�H;b�H;��H;$�H;�H;$�H;��H;b�H;�H;��H;ФH;H�H;^lH;Q5H;��G;6�F; �C;Q\=;�0;Nl;$f�:��9�к3J������#���o��s/��Ȅ�a�ýÈ��nH�n��i㼾R���I��%E�M�h�L ��V���      � ����y�M�h�ބN��O/����-�߾�A���*|�ؕ6�a}��㳽JSt�(�!�Wrμ(F{��_�
Y��f����:���:WZ;2;�N>;�D;��F;��G;J<H;�oH;��H;t�H;��H;��H;��H;��H;��H;�H;��H;��H;��H;��H;��H;t�H;��H;�oH;J<H;��G;��F;�D;�N>;2;WZ;���:�:f���
Y���_�(F{�Wrμ(�!�JSt��㳽a}�ؕ6��*|��A��-�߾����O/�ބN�M�h���y�      $�X�EvS�%E��O/��S�1W����������4S\�� �q�&�����Y�h��������]�|���S�b��Y���Y:�~�:�_;��4; �?;}�D;�F;/�G;6EH;tH;�H;��H;��H;3�H;��H;E�H;8�H;�H;8�H;E�H;��H;3�H;��H;��H;�H;tH;6EH;/�G;�F;}�D; �?;��4;�_;�~�:��Y:�Y�S�b�|�����]�����h����Y�&���q�� �4S\���������1W���S��O/�%E�EvS�      �O/�aM+�I�����1W�� 9ɾ0���Mw�� :�Y��_�ý�L��Dn;�>���bv���E<��˻(�-�����x�:^;%;�7;��@;V4E;�!G;,�G;iOH;1zH;�H;��H;��H;��H;�H;2�H;�H;��H;�H;2�H;�H;��H;��H;��H;�H;1zH;iOH;,�G;�!G;V4E;��@;�7;%;^;�x�:���(�-��˻�E<�bv��>���Dn;��L��_�ýY��� :��Mw�0�� 9ɾ1W�����I��aM+�      #y��v�R���-�߾����0��1����nH���(Ὁu��r�d�O�Prμ<"�����	��1���k89w:�:��;+;�{:;�6B;)�E;FaG;�H;ZH;��H;M�H;ĮH;�H;f�H;e�H;+�H;��H;��H;��H;+�H;e�H;f�H;�H;ĮH;M�H;��H;ZH;�H;FaG;)�E;�6B;�{:;+;��;w:�:�k891��	�����<"��PrμO�r�d��u��(����nH�1���0������-�߾R����v�      -�; 9ɾi㼾�A�������Mw��nH�����Z��㳽����Z\8�O#�������]N�J��-�b�UJx�{5:��:��;8�0;v\=;v�C;�ZF;�G;)H;eH;��H;G�H;g�H;��H;7�H;��H;P�H;��H;��H;��H;P�H;��H;7�H;��H;g�H;G�H;��H;eH;)H;�G;�ZF;v�C;v\=;8�0;��;��:{5:UJx�-�b�J���]N�����O#��Z\8������㳽�Z񽞯��nH��Mw������A��i㼾 9ɾ      Ѱ������n���*|�4S\�� :����Z�U$������K�c���Oļ����������x&���P.�:0^;��#;G6;��?;-�D;��F;��G;*?H;�oH;�H;��H;:�H;r�H;J�H;��H;��H;��H;��H;��H;��H;��H;J�H;r�H;:�H;��H;�H;�oH;*?H;��G;��F;-�D;��?;G6;��#;0^;P.�:��x&������������Oļc���K����U$���Z���� :�4S\��*|�n������      j+X��T��nH�ؕ6�� �Y��(��㳽����mR����ټ�����E<��?ݻad\�a ��&:�c�:8�;z�,;��:;�6B;ͱE;�KG;jH;�RH;�zH;��H;
�H;9�H;`�H;n�H;+�H;��H;�H;��H;�H;��H;+�H;n�H;`�H;9�H;
�H;��H;�zH;�RH;jH;�KG;ͱE;�6B;��:;z�,;8�;�c�:&:a ��ad\��?ݻ�E<������ټ���mR�����㳽(�Y��� �ؕ6��nH��T�      ��]�È�a}�q�_�ý�u�������K����o�Wv���&R���e^���뺾@���:�A;�";��4;��>;�D;F;-�G;)H;�cH;��H;5�H;��H;N�H;N�H;��H;��H;<�H;(�H;��H;(�H;<�H;��H;��H;N�H;N�H;��H;5�H;��H;�cH;)H;-�G;F;�D;��>;��4;�";�A;��:�@���e^�����&R�Wv���o����K������u��_�ýq�a}�È�]�      ��ѽ�[νa�ý�㳽&����L��r�d�Z\8�c���ټWv����Y��_����y��]���Y:A��:�l; r-;R�:;��A;rnE;�!G;��G;�FH;�rH;�H;��H;�H;J�H;5�H;��H;��H;��H;B�H;�H;B�H;��H;��H;��H;5�H;J�H;�H;��H;�H;�rH;�FH;��G;�!G;rnE;��A;R�:; r-;�l;A��:��Y:]�y������_���Y�Wv���ټc��Z\8�r�d��L��&����㳽a�ý�[ν      ���������Ȅ�JSt���Y�Dn;�O�O#���Oļ�����&R��_������N3�+�Y�12:�:9�;A?&;)G6;�W?;�D;gwF;�G;c H;�]H;��H;�H;�H;a�H;$�H;�H;��H;(�H;��H;j�H;%�H;j�H;��H;(�H;��H;�H;$�H;a�H;�H;�H;��H;�]H;c H;�G;gwF;�D;�W?;)G6;A?&;9�;�:12:+�Y��N3������_��&R������OļO#��O�Dn;���Y�JSt��Ȅ�����      Gn;�`\8��s/�(�!�h��>���Prμ��������E<�������N3��Ix�h�9��:U^;� ;2;��<;/�B;�E;f4G;2�G;^EH;�pH;��H;h�H;гH;k�H;��H;��H;�H;��H;1�H;��H;�H;��H;1�H;��H;�H;��H;��H;k�H;гH;h�H;��H;�pH;^EH;2�G;f4G;�E;/�B;��<;2;� ;U^;��:h�9�Ix��N3�������E<��������Prμ>���h��(�!��s/�`\8�      >�Ｘ���o�Wrμ����bv��<"���]N�����?ݻe^��y��+�Y�h�9��:���:B�;��.;�{:;3>A;��D;`�F;�G;
)H;E`H;5�H;��H;�H;S�H;6�H;R�H;t�H;�H;/�H;k�H;��H;��H;��H;k�H;/�H;�H;t�H;R�H;6�H;S�H;�H;��H;5�H;E`H;
)H;�G;`�F;��D;3>A;�{:;��.;B�;���:��:h�9+�Y�y��e^���?ݻ����]N�<"��bv������Wrμ�o༸��      �����x���#��(F{���]��E<����J�뻱���ad\���]�12:��:���:�Z;��,;0�8;a @;0D;�ZF;QzG;
H;jOH;>uH;�H;\�H;�H;C�H;z�H;��H;��H;��H;��H;��H;��H;��H;��H;��H;��H;��H;��H;��H;z�H;C�H;�H;\�H;�H;>uH;jOH;
H;QzG;�ZF;0D;a @;0�8;��,;�Z;���:��:12:]���ad\�����J�뻛���E<���]�(F{��#���x��      �B(��%�����_�|����˻	��-�b�x&�a ���@���Y:�:U^;B�;��,;[_8;��?;��C;�F;FG;u�G;?H;GjH;#�H; �H;
�H;k�H;��H;�H;��H;/�H;��H;��H;��H;��H;��H;��H;��H;��H;��H;/�H;��H;�H;��H;k�H;
�H; �H;#�H;GjH;?H;u�G;FG;�F;��C;��?;[_8;��,;B�;U^;�:��Y:�@�a ��x&�-�b�	���˻|����_�����%�      嚩�[���3J��
Y��S�b�(�-�1��UJx���&:��:A��:9�;� ;��.;0�8;��?;2�C;�E;f"G;�G;1H;aH;gH;��H;��H;��H;��H;s�H;(�H;I�H;J�H;��H;(�H;��H;H�H;��H;H�H;��H;(�H;��H;J�H;I�H;(�H;s�H;��H;��H;��H;��H;gH;aH;1H;�G;f"G;�E;2�C;��?;0�8;��.;� ;9�;A��:��:&:��UJx�1��(�-�S�b�
Y��3J��[���      �����뺶кf����Y�����k89{5:P.�:�c�:�A;�l;A?&;2;�{:;a @;��C;�E;�G;�G;}'H;ZH;�yH;X�H;��H;��H;{�H;��H;��H;l�H;��H;�H;[�H;<�H;W�H;
�H;��H;
�H;W�H;<�H;[�H;�H;��H;l�H;��H;��H;{�H;��H;��H;X�H;�yH;ZH;}'H;�G;�G;�E;��C;a @;�{:;2;A?&;�l;�A;�c�:P.�:{5:�k89����Y�f����к���      2�e9��9��9�:��Y:�x�:w:�:��:0^;8�;�"; r-;)G6;��<;3>A;0D;�F;f"G;�G;$H;VH;�uH;��H;Y�H;b�H;��H;!�H;��H;��H;E�H;��H;��H;��H;7�H;�H;��H;�H;��H;�H;7�H;��H;��H;��H;E�H;��H;��H;!�H;��H;b�H;Y�H;��H;�uH;VH;$H;�G;f"G;�F;0D;3>A;��<;)G6; r-;�";8�;0^;��:w:�:�x�:��Y:�:��9��9      ��:C,�:$f�:���:�~�:^;��;��;��#;z�,;��4;R�:;�W?;/�B;��D;�ZF;FG;�G;}'H;VH;�tH;��H;.�H;�H;<�H;
�H;��H;��H;��H;��H;��H;��H;��H;��H;��H;^�H;b�H;^�H;��H;��H;��H;��H;��H;��H;��H;��H;��H;
�H;<�H;�H;.�H;��H;�tH;VH;}'H;�G;FG;�ZF;��D;/�B;�W?;R�:;��4;z�,;��#;��;��;^;�~�:���:$f�:C,�:      ^;��;Nl;WZ;�_;%;+;8�0;G6;��:;��>;��A;�D;�E;`�F;QzG;u�G;1H;ZH;�uH;��H;g�H;ܫH;�H;��H;f�H;��H;��H;��H;��H;H�H;G�H;��H;��H;p�H;��H;��H;��H;p�H;��H;��H;G�H;H�H;��H;��H;��H;��H;f�H;��H;�H;ܫH;g�H;��H;�uH;ZH;1H;u�G;QzG;`�F;�E;�D;��A;��>;��:;G6;8�0;+;%;�_;WZ;Nl;��;      Y.;�.;�0;2;��4;�7;�{:;v\=;��?;�6B;�D;rnE;gwF;f4G;�G;
H;?H;aH;�yH;��H;.�H;ܫH;`�H;��H;��H;��H;��H;�H;)�H;��H;��H;h�H;c�H;O�H;��H;(�H;P�H;(�H;��H;O�H;c�H;h�H;��H;��H;)�H;�H;��H;��H;��H;��H;`�H;ܫH;.�H;��H;�yH;aH;?H;
H;�G;f4G;gwF;rnE;�D;�6B;��?;v\=;�{:;�7;��4;2;�0;�.;      ��<;N�<;Q\=;�N>; �?;��@;�6B;v�C;-�D;ͱE;F;�!G;�G;2�G;
)H;jOH;GjH;gH;X�H;Y�H;�H;�H;��H;H�H;I�H;E�H;X�H;��H;,�H;B�H;�H;�H;�H;��H;I�H;��H;��H;��H;I�H;��H;�H;�H;�H;B�H;,�H;��H;X�H;E�H;I�H;H�H;��H;�H;�H;Y�H;X�H;gH;GjH;jOH;
)H;2�G;�G;�!G;F;ͱE;-�D;v�C;�6B;��@; �?;�N>;Q\=;N�<;      �VC;!nC; �C;�D;}�D;V4E;)�E;�ZF;��F;�KG;-�G;��G;c H;^EH;E`H;>uH;#�H;��H;��H;b�H;<�H;��H;��H;I�H;�H;�H;O�H;��H;��H;��H;��H;��H;��H;=�H;��H;��H;��H;��H;��H;=�H;��H;��H;��H;��H;��H;��H;O�H;�H;�H;I�H;��H;��H;<�H;b�H;��H;��H;#�H;>uH;E`H;^EH;c H;��G;-�G;�KG;��F;�ZF;)�E;V4E;}�D;�D; �C;!nC;      @ZF;�cF;6�F;��F;�F;�!G;FaG;�G;��G;jH;)H;�FH;�]H;�pH;5�H;�H; �H;��H;��H;��H;
�H;f�H;��H;E�H;�H;6�H;��H;��H;u�H;��H;��H;��H;,�H;�H;��H;�H;�H;�H;��H;�H;,�H;��H;��H;��H;u�H;��H;��H;6�H;�H;E�H;��H;f�H;
�H;��H;��H;��H; �H;�H;5�H;�pH;�]H;�FH;)H;jH;��G;�G;FaG;�!G;�F;��F;6�F;�cF;      �G;�G;��G;��G;/�G;,�G;�H;)H;*?H;�RH;�cH;�rH;��H;��H;��H;\�H;
�H;��H;{�H;!�H;��H;��H;��H;X�H;O�H;��H;��H;J�H;��H;��H;j�H; �H;}�H;��H;�H;;�H;Y�H;;�H;�H;��H;}�H; �H;j�H;��H;��H;J�H;��H;��H;O�H;X�H;��H;��H;��H;!�H;{�H;��H;
�H;\�H;��H;��H;��H;�rH;�cH;�RH;*?H;)H;�H;,�G;/�G;��G;��G;�G;      5/H;�0H;Q5H;J<H;6EH;iOH;ZH;eH;�oH;�zH;��H;�H;�H;h�H;�H;�H;k�H;��H;��H;��H;��H;��H;�H;��H;��H;��H;J�H;��H;e�H;T�H;�H;j�H;��H;�H;E�H;[�H;M�H;[�H;E�H;�H;��H;j�H;�H;T�H;e�H;��H;J�H;��H;��H;��H;�H;��H;��H;��H;��H;��H;k�H;�H;�H;h�H;�H;�H;��H;�zH;�oH;eH;ZH;iOH;6EH;J<H;Q5H;�0H;      tiH;"jH;^lH;�oH;tH;1zH;��H;��H;�H;��H;5�H;��H;�H;гH;S�H;C�H;��H;s�H;��H;��H;��H;��H;)�H;,�H;��H;u�H;��H;e�H;[�H;��H;Z�H;��H;��H;5�H;e�H;o�H;b�H;o�H;e�H;5�H;��H;��H;Z�H;��H;[�H;e�H;��H;u�H;��H;,�H;)�H;��H;��H;��H;��H;s�H;��H;C�H;S�H;гH;�H;��H;5�H;��H;�H;��H;��H;1zH;tH;�oH;^lH;"jH;      X�H;ȋH;H�H;��H;�H;�H;M�H;G�H;��H;
�H;��H;�H;a�H;k�H;6�H;z�H;�H;(�H;l�H;E�H;��H;��H;��H;B�H;��H;��H;��H;T�H;��H;K�H;��H;��H;6�H;]�H;h�H;��H;��H;��H;h�H;]�H;6�H;��H;��H;K�H;��H;T�H;��H;��H;��H;B�H;��H;��H;��H;E�H;l�H;(�H;�H;z�H;6�H;k�H;a�H;�H;��H;
�H;��H;G�H;M�H;�H;�H;��H;H�H;ȋH;      s�H;ңH;ФH;t�H;��H;��H;ĮH;g�H;:�H;9�H;N�H;J�H;$�H;��H;R�H;��H;��H;I�H;��H;��H;��H;H�H;��H;�H;��H;��H;j�H;�H;Z�H;��H;��H;)�H;a�H;o�H;��H;��H;��H;��H;��H;o�H;a�H;)�H;��H;��H;Z�H;�H;j�H;��H;��H;�H;��H;H�H;��H;��H;��H;I�H;��H;��H;R�H;��H;$�H;J�H;N�H;9�H;:�H;g�H;ĮH;��H;��H;t�H;ФH;ңH;      ��H;��H;��H;��H;��H;��H;�H;��H;r�H;`�H;N�H;5�H;�H;��H;t�H;��H;/�H;J�H;�H;��H;��H;G�H;h�H;�H;��H;��H; �H;j�H;��H;��H;)�H;A�H;l�H;��H;��H;��H;��H;��H;��H;��H;l�H;A�H;)�H;��H;��H;j�H; �H;��H;��H;�H;h�H;G�H;��H;��H;�H;J�H;/�H;��H;t�H;��H;�H;5�H;N�H;`�H;r�H;��H;�H;��H;��H;��H;��H;��H;      F�H;��H;�H;��H;3�H;��H;f�H;7�H;J�H;n�H;��H;��H;��H;�H;�H;��H;��H;��H;[�H;��H;��H;��H;c�H;�H;��H;,�H;}�H;��H;��H;6�H;a�H;l�H;{�H;��H;��H;��H;��H;��H;��H;��H;{�H;l�H;a�H;6�H;��H;��H;}�H;,�H;��H;�H;c�H;��H;��H;��H;[�H;��H;��H;��H;�H;�H;��H;��H;��H;n�H;J�H;7�H;f�H;��H;3�H;��H;�H;��H;      ��H;��H;b�H;��H;��H;�H;e�H;��H;��H;+�H;��H;��H;(�H;��H;/�H;��H;��H;(�H;<�H;7�H;��H;��H;O�H;��H;=�H;�H;��H;�H;5�H;]�H;o�H;��H;��H;��H;��H;��H;��H;��H;��H;��H;��H;��H;o�H;]�H;5�H;�H;��H;�H;=�H;��H;O�H;��H;��H;7�H;<�H;(�H;��H;��H;/�H;��H;(�H;��H;��H;+�H;��H;��H;e�H;�H;��H;��H;b�H;��H;      �H;��H;��H;��H;E�H;2�H;+�H;P�H;��H;��H;<�H;��H;��H;1�H;k�H;��H;��H;��H;W�H;�H;��H;p�H;��H;I�H;��H;��H;�H;E�H;e�H;h�H;��H;��H;��H;��H;��H;��H;��H;��H;��H;��H;��H;��H;��H;h�H;e�H;E�H;�H;��H;��H;I�H;��H;p�H;��H;�H;W�H;��H;��H;��H;k�H;1�H;��H;��H;<�H;��H;��H;P�H;+�H;2�H;E�H;��H;��H;��H;      ��H;��H;$�H;��H;8�H;�H;��H;��H;��H;�H;(�H;B�H;j�H;��H;��H;��H;��H;H�H;
�H;��H;^�H;��H;(�H;��H;��H;�H;;�H;[�H;o�H;��H;��H;��H;��H;��H;��H;��H;��H;��H;��H;��H;��H;��H;��H;��H;o�H;[�H;;�H;�H;��H;��H;(�H;��H;^�H;��H;
�H;H�H;��H;��H;��H;��H;j�H;B�H;(�H;�H;��H;��H;��H;�H;8�H;��H;$�H;��H;      ��H;��H;�H;�H;�H;��H;��H;��H;��H;��H;��H;�H;%�H;�H;��H;��H;��H;��H;��H;�H;b�H;��H;P�H;��H;��H;�H;Y�H;M�H;b�H;��H;��H;��H;��H;��H;��H;��H;��H;��H;��H;��H;��H;��H;��H;��H;b�H;M�H;Y�H;�H;��H;��H;P�H;��H;b�H;�H;��H;��H;��H;��H;��H;�H;%�H;�H;��H;��H;��H;��H;��H;��H;�H;�H;�H;��H;      ��H;��H;$�H;��H;8�H;�H;��H;��H;��H;�H;(�H;B�H;j�H;��H;��H;��H;��H;H�H;
�H;��H;^�H;��H;(�H;��H;��H;�H;;�H;[�H;o�H;��H;��H;��H;��H;��H;��H;��H;��H;��H;��H;��H;��H;��H;��H;��H;o�H;[�H;;�H;�H;��H;��H;(�H;��H;^�H;��H;
�H;H�H;��H;��H;��H;��H;j�H;B�H;(�H;�H;��H;��H;��H;�H;8�H;��H;$�H;��H;      �H;��H;��H;��H;E�H;2�H;+�H;P�H;��H;��H;<�H;��H;��H;1�H;k�H;��H;��H;��H;W�H;�H;��H;p�H;��H;I�H;��H;��H;�H;E�H;e�H;h�H;��H;��H;��H;��H;��H;��H;��H;��H;��H;��H;��H;��H;��H;h�H;e�H;E�H;�H;��H;��H;I�H;��H;p�H;��H;�H;W�H;��H;��H;��H;k�H;1�H;��H;��H;<�H;��H;��H;P�H;+�H;2�H;E�H;��H;��H;��H;      ��H;��H;b�H;��H;��H;�H;e�H;��H;��H;+�H;��H;��H;(�H;��H;/�H;��H;��H;(�H;<�H;7�H;��H;��H;O�H;��H;=�H;�H;��H;�H;5�H;]�H;o�H;��H;��H;��H;��H;��H;��H;��H;��H;��H;��H;��H;o�H;]�H;5�H;�H;��H;�H;=�H;��H;O�H;��H;��H;7�H;<�H;(�H;��H;��H;/�H;��H;(�H;��H;��H;+�H;��H;��H;e�H;�H;��H;��H;b�H;��H;      F�H;��H;�H;��H;3�H;��H;f�H;7�H;J�H;n�H;��H;��H;��H;�H;�H;��H;��H;��H;[�H;��H;��H;��H;c�H;�H;��H;,�H;}�H;��H;��H;6�H;a�H;l�H;{�H;��H;��H;��H;��H;��H;��H;��H;{�H;l�H;a�H;6�H;��H;��H;}�H;,�H;��H;�H;c�H;��H;��H;��H;[�H;��H;��H;��H;�H;�H;��H;��H;��H;n�H;J�H;7�H;f�H;��H;3�H;��H;�H;��H;      ��H;��H;��H;��H;��H;��H;�H;��H;r�H;`�H;N�H;5�H;�H;��H;t�H;��H;/�H;J�H;�H;��H;��H;G�H;h�H;�H;��H;��H; �H;j�H;��H;��H;)�H;A�H;l�H;��H;��H;��H;��H;��H;��H;��H;l�H;A�H;)�H;��H;��H;j�H; �H;��H;��H;�H;h�H;G�H;��H;��H;�H;J�H;/�H;��H;t�H;��H;�H;5�H;N�H;`�H;r�H;��H;�H;��H;��H;��H;��H;��H;      s�H;ңH;ФH;t�H;��H;��H;ĮH;g�H;:�H;9�H;N�H;J�H;$�H;��H;R�H;��H;��H;I�H;��H;��H;��H;H�H;��H;�H;��H;��H;j�H;�H;Z�H;��H;��H;)�H;a�H;o�H;��H;��H;��H;��H;��H;o�H;a�H;)�H;��H;��H;Z�H;�H;j�H;��H;��H;�H;��H;H�H;��H;��H;��H;I�H;��H;��H;R�H;��H;$�H;J�H;N�H;9�H;:�H;g�H;ĮH;��H;��H;t�H;ФH;ңH;      X�H;ȋH;H�H;��H;�H;�H;M�H;G�H;��H;
�H;��H;�H;a�H;k�H;6�H;z�H;�H;(�H;l�H;E�H;��H;��H;��H;B�H;��H;��H;��H;T�H;��H;K�H;��H;��H;6�H;]�H;h�H;��H;��H;��H;h�H;]�H;6�H;��H;��H;K�H;��H;T�H;��H;��H;��H;B�H;��H;��H;��H;E�H;l�H;(�H;�H;z�H;6�H;k�H;a�H;�H;��H;
�H;��H;G�H;M�H;�H;�H;��H;H�H;ȋH;      tiH;"jH;^lH;�oH;tH;1zH;��H;��H;�H;��H;5�H;��H;�H;гH;S�H;C�H;��H;s�H;��H;��H;��H;��H;)�H;,�H;��H;u�H;��H;e�H;[�H;��H;Z�H;��H;��H;5�H;e�H;o�H;b�H;o�H;e�H;5�H;��H;��H;Z�H;��H;[�H;e�H;��H;u�H;��H;,�H;)�H;��H;��H;��H;��H;s�H;��H;C�H;S�H;гH;�H;��H;5�H;��H;�H;��H;��H;1zH;tH;�oH;^lH;"jH;      5/H;�0H;Q5H;J<H;6EH;iOH;ZH;eH;�oH;�zH;��H;�H;�H;h�H;�H;�H;k�H;��H;��H;��H;��H;��H;�H;��H;��H;��H;J�H;��H;e�H;T�H;�H;j�H;��H;�H;E�H;[�H;M�H;[�H;E�H;�H;��H;j�H;�H;T�H;e�H;��H;J�H;��H;��H;��H;�H;��H;��H;��H;��H;��H;k�H;�H;�H;h�H;�H;�H;��H;�zH;�oH;eH;ZH;iOH;6EH;J<H;Q5H;�0H;      �G;�G;��G;��G;/�G;,�G;�H;)H;*?H;�RH;�cH;�rH;��H;��H;��H;\�H;
�H;��H;{�H;!�H;��H;��H;��H;X�H;O�H;��H;��H;J�H;��H;��H;j�H; �H;}�H;��H;�H;;�H;Y�H;;�H;�H;��H;}�H; �H;j�H;��H;��H;J�H;��H;��H;O�H;X�H;��H;��H;��H;!�H;{�H;��H;
�H;\�H;��H;��H;��H;�rH;�cH;�RH;*?H;)H;�H;,�G;/�G;��G;��G;�G;      @ZF;�cF;6�F;��F;�F;�!G;FaG;�G;��G;jH;)H;�FH;�]H;�pH;5�H;�H; �H;��H;��H;��H;
�H;f�H;��H;E�H;�H;6�H;��H;��H;u�H;��H;��H;��H;,�H;�H;��H;�H;�H;�H;��H;�H;,�H;��H;��H;��H;u�H;��H;��H;6�H;�H;E�H;��H;f�H;
�H;��H;��H;��H; �H;�H;5�H;�pH;�]H;�FH;)H;jH;��G;�G;FaG;�!G;�F;��F;6�F;�cF;      �VC;!nC; �C;�D;}�D;V4E;)�E;�ZF;��F;�KG;-�G;��G;c H;^EH;E`H;>uH;#�H;��H;��H;b�H;<�H;��H;��H;I�H;�H;�H;O�H;��H;��H;��H;��H;��H;��H;=�H;��H;��H;��H;��H;��H;=�H;��H;��H;��H;��H;��H;��H;O�H;�H;�H;I�H;��H;��H;<�H;b�H;��H;��H;#�H;>uH;E`H;^EH;c H;��G;-�G;�KG;��F;�ZF;)�E;V4E;}�D;�D; �C;!nC;      ��<;N�<;Q\=;�N>; �?;��@;�6B;v�C;-�D;ͱE;F;�!G;�G;2�G;
)H;jOH;GjH;gH;X�H;Y�H;�H;�H;��H;H�H;I�H;E�H;X�H;��H;,�H;B�H;�H;�H;�H;��H;I�H;��H;��H;��H;I�H;��H;�H;�H;�H;B�H;,�H;��H;X�H;E�H;I�H;H�H;��H;�H;�H;Y�H;X�H;gH;GjH;jOH;
)H;2�G;�G;�!G;F;ͱE;-�D;v�C;�6B;��@; �?;�N>;Q\=;N�<;      Y.;�.;�0;2;��4;�7;�{:;v\=;��?;�6B;�D;rnE;gwF;f4G;�G;
H;?H;aH;�yH;��H;.�H;ܫH;`�H;��H;��H;��H;��H;�H;)�H;��H;��H;h�H;c�H;O�H;��H;(�H;P�H;(�H;��H;O�H;c�H;h�H;��H;��H;)�H;�H;��H;��H;��H;��H;`�H;ܫH;.�H;��H;�yH;aH;?H;
H;�G;f4G;gwF;rnE;�D;�6B;��?;v\=;�{:;�7;��4;2;�0;�.;      ^;��;Nl;WZ;�_;%;+;8�0;G6;��:;��>;��A;�D;�E;`�F;QzG;u�G;1H;ZH;�uH;��H;g�H;ܫH;�H;��H;f�H;��H;��H;��H;��H;H�H;G�H;��H;��H;p�H;��H;��H;��H;p�H;��H;��H;G�H;H�H;��H;��H;��H;��H;f�H;��H;�H;ܫH;g�H;��H;�uH;ZH;1H;u�G;QzG;`�F;�E;�D;��A;��>;��:;G6;8�0;+;%;�_;WZ;Nl;��;      ��:C,�:$f�:���:�~�:^;��;��;��#;z�,;��4;R�:;�W?;/�B;��D;�ZF;FG;�G;}'H;VH;�tH;��H;.�H;�H;<�H;
�H;��H;��H;��H;��H;��H;��H;��H;��H;��H;^�H;b�H;^�H;��H;��H;��H;��H;��H;��H;��H;��H;��H;
�H;<�H;�H;.�H;��H;�tH;VH;}'H;�G;FG;�ZF;��D;/�B;�W?;R�:;��4;z�,;��#;��;��;^;�~�:���:$f�:C,�:      2�e9��9��9�:��Y:�x�:w:�:��:0^;8�;�"; r-;)G6;��<;3>A;0D;�F;f"G;�G;$H;VH;�uH;��H;Y�H;b�H;��H;!�H;��H;��H;E�H;��H;��H;��H;7�H;�H;��H;�H;��H;�H;7�H;��H;��H;��H;E�H;��H;��H;!�H;��H;b�H;Y�H;��H;�uH;VH;$H;�G;f"G;�F;0D;3>A;��<;)G6; r-;�";8�;0^;��:w:�:�x�:��Y:�:��9��9      �����뺶кf����Y�����k89{5:P.�:�c�:�A;�l;A?&;2;�{:;a @;��C;�E;�G;�G;}'H;ZH;�yH;X�H;��H;��H;{�H;��H;��H;l�H;��H;�H;[�H;<�H;W�H;
�H;��H;
�H;W�H;<�H;[�H;�H;��H;l�H;��H;��H;{�H;��H;��H;X�H;�yH;ZH;}'H;�G;�G;�E;��C;a @;�{:;2;A?&;�l;�A;�c�:P.�:{5:�k89����Y�f����к���      嚩�[���3J��
Y��S�b�(�-�1��UJx���&:��:A��:9�;� ;��.;0�8;��?;2�C;�E;f"G;�G;1H;aH;gH;��H;��H;��H;��H;s�H;(�H;I�H;J�H;��H;(�H;��H;H�H;��H;H�H;��H;(�H;��H;J�H;I�H;(�H;s�H;��H;��H;��H;��H;gH;aH;1H;�G;f"G;�E;2�C;��?;0�8;��.;� ;9�;A��:��:&:��UJx�1��(�-�S�b�
Y��3J��[���      �B(��%�����_�|����˻	��-�b�x&�a ���@���Y:�:U^;B�;��,;[_8;��?;��C;�F;FG;u�G;?H;GjH;#�H; �H;
�H;k�H;��H;�H;��H;/�H;��H;��H;��H;��H;��H;��H;��H;��H;��H;/�H;��H;�H;��H;k�H;
�H; �H;#�H;GjH;?H;u�G;FG;�F;��C;��?;[_8;��,;B�;U^;�:��Y:�@�a ��x&�-�b�	���˻|����_�����%�      �����x���#��(F{���]��E<����J�뻱���ad\���]�12:��:���:�Z;��,;0�8;a @;0D;�ZF;QzG;
H;jOH;>uH;�H;\�H;�H;C�H;z�H;��H;��H;��H;��H;��H;��H;��H;��H;��H;��H;��H;��H;��H;z�H;C�H;�H;\�H;�H;>uH;jOH;
H;QzG;�ZF;0D;a @;0�8;��,;�Z;���:��:12:]���ad\�����J�뻛���E<���]�(F{��#���x��      >�Ｘ���o�Wrμ����bv��<"���]N�����?ݻe^��y��+�Y�h�9��:���:B�;��.;�{:;3>A;��D;`�F;�G;
)H;E`H;5�H;��H;�H;S�H;6�H;R�H;t�H;�H;/�H;k�H;��H;��H;��H;k�H;/�H;�H;t�H;R�H;6�H;S�H;�H;��H;5�H;E`H;
)H;�G;`�F;��D;3>A;�{:;��.;B�;���:��:h�9+�Y�y��e^���?ݻ����]N�<"��bv������Wrμ�o༸��      Gn;�`\8��s/�(�!�h��>���Prμ��������E<�������N3��Ix�h�9��:U^;� ;2;��<;/�B;�E;f4G;2�G;^EH;�pH;��H;h�H;гH;k�H;��H;��H;�H;��H;1�H;��H;�H;��H;1�H;��H;�H;��H;��H;k�H;гH;h�H;��H;�pH;^EH;2�G;f4G;�E;/�B;��<;2;� ;U^;��:h�9�Ix��N3�������E<��������Prμ>���h��(�!��s/�`\8�      ���������Ȅ�JSt���Y�Dn;�O�O#���Oļ�����&R��_������N3�+�Y�12:�:9�;A?&;)G6;�W?;�D;gwF;�G;c H;�]H;��H;�H;�H;a�H;$�H;�H;��H;(�H;��H;j�H;%�H;j�H;��H;(�H;��H;�H;$�H;a�H;�H;�H;��H;�]H;c H;�G;gwF;�D;�W?;)G6;A?&;9�;�:12:+�Y��N3������_��&R������OļO#��O�Dn;���Y�JSt��Ȅ�����      ��ѽ�[νa�ý�㳽&����L��r�d�Z\8�c���ټWv����Y��_����y��]���Y:A��:�l; r-;R�:;��A;rnE;�!G;��G;�FH;�rH;�H;��H;�H;J�H;5�H;��H;��H;��H;B�H;�H;B�H;��H;��H;��H;5�H;J�H;�H;��H;�H;�rH;�FH;��G;�!G;rnE;��A;R�:; r-;�l;A��:��Y:]�y������_���Y�Wv���ټc��Z\8�r�d��L��&����㳽a�ý�[ν      ��]�È�a}�q�_�ý�u�������K����o�Wv���&R���e^���뺾@���:�A;�";��4;��>;�D;F;-�G;)H;�cH;��H;5�H;��H;N�H;N�H;��H;��H;<�H;(�H;��H;(�H;<�H;��H;��H;N�H;N�H;��H;5�H;��H;�cH;)H;-�G;F;�D;��>;��4;�";�A;��:�@���e^�����&R�Wv���o����K������u��_�ýq�a}�È�]�      j+X��T��nH�ؕ6�� �Y��(��㳽����mR����ټ�����E<��?ݻad\�a ��&:�c�:8�;z�,;��:;�6B;ͱE;�KG;jH;�RH;�zH;��H;
�H;9�H;`�H;n�H;+�H;��H;�H;��H;�H;��H;+�H;n�H;`�H;9�H;
�H;��H;�zH;�RH;jH;�KG;ͱE;�6B;��:;z�,;8�;�c�:&:a ��ad\��?ݻ�E<������ټ���mR�����㳽(�Y��� �ؕ6��nH��T�      Ѱ������n���*|�4S\�� :����Z�U$������K�c���Oļ����������x&���P.�:0^;��#;G6;��?;-�D;��F;��G;*?H;�oH;�H;��H;:�H;r�H;J�H;��H;��H;��H;��H;��H;��H;��H;J�H;r�H;:�H;��H;�H;�oH;*?H;��G;��F;-�D;��?;G6;��#;0^;P.�:��x&������������Oļc���K����U$���Z���� :�4S\��*|�n������      -�; 9ɾi㼾�A�������Mw��nH�����Z��㳽����Z\8�O#�������]N�J��-�b�UJx�{5:��:��;8�0;v\=;v�C;�ZF;�G;)H;eH;��H;G�H;g�H;��H;7�H;��H;P�H;��H;��H;��H;P�H;��H;7�H;��H;g�H;G�H;��H;eH;)H;�G;�ZF;v�C;v\=;8�0;��;��:{5:UJx�-�b�J���]N�����O#��Z\8������㳽�Z񽞯��nH��Mw������A��i㼾 9ɾ      #y��v�R���-�߾����0��1����nH���(Ὁu��r�d�O�Prμ<"�����	��1���k89w:�:��;+;�{:;�6B;)�E;FaG;�H;ZH;��H;M�H;ĮH;�H;f�H;e�H;+�H;��H;��H;��H;+�H;e�H;f�H;�H;ĮH;M�H;��H;ZH;�H;FaG;)�E;�6B;�{:;+;��;w:�:�k891��	�����<"��PrμO�r�d��u��(����nH�1���0������-�߾R����v�      �O/�aM+�I�����1W�� 9ɾ0���Mw�� :�Y��_�ý�L��Dn;�>���bv���E<��˻(�-�����x�:^;%;�7;��@;V4E;�!G;,�G;iOH;1zH;�H;��H;��H;��H;�H;2�H;�H;��H;�H;2�H;�H;��H;��H;��H;�H;1zH;iOH;,�G;�!G;V4E;��@;�7;%;^;�x�:���(�-��˻�E<�bv��>���Dn;��L��_�ýY��� :��Mw�0�� 9ɾ1W�����I��aM+�      $�X�EvS�%E��O/��S�1W����������4S\�� �q�&�����Y�h��������]�|���S�b��Y���Y:�~�:�_;��4; �?;}�D;�F;/�G;6EH;tH;�H;��H;��H;3�H;��H;E�H;8�H;�H;8�H;E�H;��H;3�H;��H;��H;�H;tH;6EH;/�G;�F;}�D; �?;��4;�_;�~�:��Y:�Y�S�b�|�����]�����h����Y�&���q�� �4S\���������1W���S��O/�%E�EvS�      � ����y�M�h�ބN��O/����-�߾�A���*|�ؕ6�a}��㳽JSt�(�!�Wrμ(F{��_�
Y��f����:���:WZ;2;�N>;�D;��F;��G;J<H;�oH;��H;t�H;��H;��H;��H;��H;��H;�H;��H;��H;��H;��H;��H;t�H;��H;�oH;J<H;��G;��F;�D;�N>;2;WZ;���:�:f���
Y���_�(F{�Wrμ(�!�JSt��㳽a}�ؕ6��*|��A��-�߾����O/�ބN�M�h���y�      2v��V���L ��M�h�%E�I��R���i㼾n���nH�È�a�ý�Ȅ��s/��o༼#�����3J���к��9$f�:Nl;�0;Q\=; �C;6�F;��G;Q5H;^lH;H�H;ФH;��H;�H;b�H;��H;$�H;�H;$�H;��H;b�H;�H;��H;ФH;H�H;^lH;Q5H;��G;6�F; �C;Q\=;�0;Nl;$f�:��9�к3J������#���o��s/��Ȅ�a�ýÈ��nH�n��i㼾R���I��%E�M�h�L ��V���      ph��"���V�����y�EvS�aM+��v� 9ɾ�����T�]��[ν����`\8�����x���%�[��������9C,�:��;�.;N�<;!nC;�cF;�G;�0H;"jH;ȋH;ңH;��H;��H;��H;��H;��H;��H;��H;��H;��H;��H;��H;ңH;ȋH;"jH;�0H;�G;�cF;!nC;N�<;�.;��;C,�:��9���[����%��x�����`\8������[ν]��T����� 9ɾ�v�aM+�EvS���y�V���"���      Vܿ%�ֿ�aǿ2^��&���Io���7����iþ�(���-=��` ��@����_�&]�&p����I�q�ѻ��)��R�]�:��
;*;D�:;�B;VHF;=�G;�kH;4�H;��H;i�H;��H;��H;p�H;��H;)�H;��H;)�H;��H;p�H;��H;��H;i�H;��H;4�H;�kH;=�G;VHF;�B;D�:;*;��
;]�:�R���)�q�ѻ��I�&p��&]���_��@���` ��-=��(���iþ����7�Io�&���2^���aǿ%�ֿ      %�ֿ5pѿ֊¿������PXi�Õ3��
�GD��;l��1�9�j.���R��\� �\x��1�E��ͻ��$�� ����:��;��*;\�:;.�B;4TF;��G;[mH;ϠH;ݶH;��H;��H;��H;�H;��H;<�H;��H;<�H;��H;�H;��H;��H;��H;ݶH;ϠH;[mH;��G;4TF;.�B;\�:;��*;��;���:� ���$��ͻ1�E�\x�� �\��R��j.��1�9�;l��GD���
�Õ3�PXi�������֊¿5pѿ      �aǿ֊¿���������s"Y��f'�����)o���.}��k/�m��ڟ�<Q�$#�ע��(;�P������B�7���:J�;�,;��;;�C;SvF;0�G;�qH;[�H;��H;=�H;�H;�H;��H;��H;j�H;��H;j�H;��H;��H;�H;�H;=�H;��H;[�H;�qH;0�G;SvF;�C;��;;�,;J�;��:B�7����P����(;�ע�$#�<Q�ڟ�m���k/��.}�)o�������f'�s"Y����������֊¿      2^������b���Io���@���޾����&ce�"����ڽ绒��f@������R���O*�mG������<^9Ӳ�:\;�c.;'�<;ՏC;G�F;��G;�xH;ĤH;8�H;J�H;��H;��H;��H;�H;��H;7�H;��H;�H;��H;��H;��H;J�H;8�H;ĤH;�xH;��G;G�F;ՏC;'�<;�c.;\;Ӳ�:�<^9���mG���O*��R�������f@�绒���ڽ"��&ce������޾���@�Io�b�������      &����������Io��!J�@�#��\��HD������jPH�����b��C��t +�u�ټ%��������������:���:��;�X1;3>;�/D;��F;�H;s�H;��H;*�H;��H;��H;)�H;��H;p�H;��H;�H;��H;p�H;��H;)�H;��H;��H;*�H;��H;s�H;�H;��F;�/D;3>;�X1;��;���:��:����������%��u�ټt +�C���b�����jPH�����HD���\��@�#��!J�Io��������      Io�PXi�s"Y���@�@�#��
��о�A�� �i���(�i��gr����_��5��ɺ�n�`��<����d�<�\�Q�X:PO�:7`;$�4;�?;��D;�7G;�/H;ȊH;��H;��H;.�H;��H;��H;�H;��H;-�H;��H;-�H;��H;�H;��H;��H;.�H;��H;��H;ȊH;�/H;�7G;��D;�?;$�4;7`;PO�:Q�X:<�\���d��<��n�`��ɺ��5���_�gr��i����(� �i��A���о�
�@�#���@�s"Y�PXi�      ��7�Õ3��f'���\���о�����.}��-=�o
�y�ĽO��:����������7�?GĻ*�$�S�����:�z;�C&;E+8;FIA;1�E;��G;�KH;�H;��H;S�H;�H;(�H;��H;��H;A�H;��H;5�H;��H;A�H;��H;��H;(�H;�H;S�H;��H;�H;�KH;��G;1�E;FIA;E+8;�C&;�z;���:S��*�$�?GĻ�7���������:�O��y�Ľo
��-=��.}������о�\����f'�Õ3�      ���
������޾HD���A���.}��D�[t���ڽ�!��\����P�ļ�
v�F�����Jɺ�N�9���:i';�-;ӊ;;��B;�HF;��G;?eH;ʜH;�H;N�H;��H;��H;��H;{�H;��H;�H;��H;�H;��H;{�H;��H;��H;��H;N�H;�H;ʜH;?eH;��G;�HF;��B;ӊ;;�-;i';���:�N�9�Jɺ��F���
v�P�ļ���\��!����ڽ[t��D��.}��A��HD���޾�����
�      �iþGD��)o���������� �i��-=�[t����R��Tys�m +����s񗼗(;�G�ѻt@�̇!��1j:�O�:4�;�C3;~�>;DED;��F;�H;`{H;��H;��H;W�H;�H;�H;��H;9�H;S�H;��H;�H;��H;S�H;9�H;��H;�H;�H;W�H;��H;��H;`{H;�H;��F;DED;~�>;�C3;4�;�O�:�1j:̇!�t@�G�ѻ�(;�s����m +�Tys��R����[t��-=� �i���������)o��GD��      �(��;l���.}�&ce�jPH���(�o
���ڽ�R����{�4�6�� �$p��\�`�ר�-��JҺ�C^9a��:>�;�}(;t�8;IA;6{E;GiG;�<H;i�H; �H;H�H;��H;N�H;��H;��H;��H;��H;�H;i�H;�H;��H;��H;��H;��H;N�H;��H;H�H; �H;i�H;�<H;GiG;6{E;IA;t�8;�}(;>�;a��:�C^9JҺ-��ר�\�`�$p��� �4�6���{��R����ڽo
���(�jPH�&ce��.}�;l��      �-=�1�9��k/�"�����i��y�Ľ�!��Tys�4�6�#��ɺ��vz����c^��˃$�y����r:���:7�;�X1;?H=;jwC;WvF;S�G;/eH;m�H;��H;��H;��H;v�H;�H;��H;��H;��H;��H;��H;��H;��H;��H;��H;�H;v�H;��H;��H;��H;m�H;/eH;S�G;WvF;jwC;?H=;�X1;7�;���:��r:y��˃$�c^������vz��ɺ�#�4�6�Tys��!��y�Ľi���"���k/�1�9�      �` �j.��m��ڽ�b��gr��O��\�m +�� ��ɺ�<��O*�bͻP6R��ǅ���:���:ۃ;�);6t8;��@;�)E;�7G;t#H;p�H;d�H;�H;J�H;��H;��H;��H;�H;n�H;�H; �H;?�H; �H;�H;n�H;�H;��H;��H;��H;J�H;�H;d�H;p�H;t#H;�7G;�)E;��@;6t8;�);ۃ;���:��:�ǅ�P6R�bͻ�O*�<��ɺ�� �m +�\�O��gr���b����ڽm��j.��      �@���R��ڟ�绒�C����_�:�������$p���vz��O*�5ֻek������09�:`0;�� ;�C3;��=;�C;kF;��G;�[H;ÖH;o�H;&�H;b�H;��H;��H;��H;�H;'�H;��H;o�H;��H;o�H;��H;'�H;�H;��H;��H;��H;b�H;&�H;o�H;ÖH;�[H;��G;kF;�C;��=;�C3;�� ;`0;�:��09���ek�5ֻ�O*��vz�$p����輙��:���_�C��绒�ڟ��R��      ��_�\�<Q��f@�t +��5�����P�ļs�\�`����bͻek��IɺW	7��:�O�:y�;%d.;��:;Z�A;d{E;�MG;q&H;/�H;�H;��H;��H;J�H;n�H;|�H;S�H;�H;��H;*�H;��H;�H;��H;*�H;��H;�H;S�H;|�H;n�H;J�H;��H;��H;�H;/�H;q&H;�MG;d{E;Z�A;��:;%d.;y�;�O�:�:W	7��Iɺek�bͻ���\�`�s�P�ļ�����5�t +��f@�<Q�\�      &]� �$#�����u�ټ�ɺ������
v��(;�ר�c^��P6R����W	7����:���:O�;l�*;+8;� @;��D;��F;'�G;eH;��H;��H;žH;��H;�H;��H;B�H;��H;��H;��H;��H;B�H;u�H;B�H;��H;��H;��H;��H;B�H;��H;�H;��H;žH;��H;��H;eH;'�G;��F;��D;� @;+8;l�*;O�;���:���:W	7����P6R�c^��ר��(;��
v������ɺ�u�ټ����$#� �      &p��\x��ע��R��%��n�`��7�F��G�ѻ-��˃$��ǅ���09�:���:�;!~(;�Y6;��>;�C;&HF;�G;DH;s�H;�H;ϸH;3�H;K�H;2�H;�H;��H;��H;��H;,�H;�H;��H;��H;��H;�H;,�H;��H;��H;��H;�H;2�H;K�H;3�H;ϸH;�H;s�H;DH;�G;&HF;�C;��>;�Y6;!~(;�;���:�:��09�ǅ�˃$�-��G�ѻF���7�n�`�%���R��ע�\x��      ��I�1�E��(;��O*�����<��?GĻ��t@�JҺy��:�:�O�:O�;!~(;S�5;>;qC;k�E;�bG;k#H;"{H;_�H;I�H;��H;��H;Y�H;��H;;�H;x�H;��H;i�H;��H;Y�H;��H;�H;��H;Y�H;��H;i�H;��H;x�H;;�H;��H;Y�H;��H;��H;I�H;_�H;"{H;k#H;�bG;k�E;qC;>;S�5;!~(;O�;�O�:�:��:y��JҺt@���?GĻ�<������O*��(;�1�E�      q�ѻ�ͻP���mG�������d�*�$��Jɺ̇!��C^9��r:���:`0;y�;l�*;�Y6;>;o�B;��E;8G;�H;,mH;A�H;m�H;μH;��H;��H;��H;h�H;�H;��H;��H;�H;�H;��H;�H;<�H;�H;��H;�H;�H;��H;��H;�H;h�H;��H;��H;��H;μH;m�H;A�H;,mH;�H;8G;��E;o�B;>;�Y6;l�*;y�;`0;���:��r:�C^9̇!��Jɺ*�$���d����mG��P����ͻ      ��)���$�����������<�\�S���N�9�1j:a��:���:ۃ;�� ;%d.;+8;��>;qC;��E;�(G;��G;>cH;��H;��H;��H;��H;U�H;��H;��H;��H;��H;��H;b�H;��H;w�H;�H;I�H;c�H;I�H;�H;w�H;��H;b�H;��H;��H;��H;��H;��H;U�H;��H;��H;��H;��H;>cH;��G;�(G;��E;qC;��>;+8;%d.;�� ;ۃ;���:a��:�1j:�N�9S��<�\�������������$�      �R�� �B�7��<^9��:Q�X:���:���:�O�:>�;7�;�);�C3;��:;� @;�C;k�E;8G;��G;�_H;��H;?�H;@�H;��H;e�H;Q�H;i�H;x�H;��H;��H;��H;$�H; �H;��H;@�H;{�H;{�H;{�H;@�H;��H; �H;$�H;��H;��H;��H;x�H;i�H;Q�H;e�H;��H;@�H;?�H;��H;�_H;��G;8G;k�E;�C;� @;��:;�C3;�);7�;>�;�O�:���:���:Q�X:��:�<^9B�7�� �      ]�:���:��:Ӳ�:���:PO�:�z;i';4�;�}(;�X1;6t8;��=;Z�A;��D;&HF;�bG;�H;>cH;��H;n�H;��H;S�H;�H;��H;Y�H;d�H;��H;<�H;��H;��H;��H;m�H;��H;Y�H;��H;��H;��H;Y�H;��H;m�H;��H;��H;��H;<�H;��H;d�H;Y�H;��H;�H;S�H;��H;n�H;��H;>cH;�H;�bG;&HF;��D;Z�A;��=;6t8;�X1;�}(;4�;i';�z;PO�:���:Ӳ�:��:���:      ��
;��;J�;\;��;7`;�C&;�-;�C3;t�8;?H=;��@;�C;d{E;��F;�G;k#H;,mH;��H;?�H;��H;��H;Y�H;:�H;��H;��H;��H;��H;�H;�H;4�H;�H;��H;1�H;r�H;��H;��H;��H;r�H;1�H;��H;�H;4�H;�H;�H;��H;��H;��H;��H;:�H;Y�H;��H;��H;?�H;��H;,mH;k#H;�G;��F;d{E;�C;��@;?H=;t�8;�C3;�-;�C&;7`;��;\;J�;��;      *;��*;�,;�c.;�X1;$�4;E+8;ӊ;;~�>;IA;jwC;�)E;kF;�MG;'�G;DH;"{H;A�H;��H;@�H;S�H;Y�H;��H;�H;�H;w�H;#�H;�H;��H;��H;��H;��H;��H;L�H;��H;��H;��H;��H;��H;L�H;��H;��H;��H;��H;��H;�H;#�H;w�H;�H;�H;��H;Y�H;S�H;@�H;��H;A�H;"{H;DH;'�G;�MG;kF;�)E;jwC;IA;~�>;ӊ;;E+8;$�4;�X1;�c.;�,;��*;      D�:;\�:;��;;'�<;3>;�?;FIA;��B;DED;6{E;WvF;�7G;��G;q&H;eH;s�H;_�H;m�H;��H;��H;�H;:�H;�H;��H;5�H;��H;��H;G�H;��H;~�H;(�H;��H;,�H;l�H;��H;��H;��H;��H;��H;l�H;,�H;��H;(�H;~�H;��H;G�H;��H;��H;5�H;��H;�H;:�H;�H;��H;��H;m�H;_�H;s�H;eH;q&H;��G;�7G;WvF;6{E;DED;��B;FIA;�?;3>;'�<;��;;\�:;      �B;.�B;�C;ՏC;�/D;��D;1�E;�HF;��F;GiG;S�G;t#H;�[H;/�H;��H;�H;I�H;μH;��H;e�H;��H;��H;�H;5�H;��H;��H;�H;T�H;8�H;�H;��H;��H;=�H;��H;��H;��H;��H;��H;��H;��H;=�H;��H;��H;�H;8�H;T�H;�H;��H;��H;5�H;�H;��H;��H;e�H;��H;μH;I�H;�H;��H;/�H;�[H;t#H;S�G;GiG;��F;�HF;1�E;��D;�/D;ՏC;�C;.�B;      VHF;4TF;SvF;G�F;��F;�7G;��G;��G;�H;�<H;/eH;p�H;ÖH;�H;��H;ϸH;��H;��H;U�H;Q�H;Y�H;��H;w�H;��H;��H;	�H;9�H;�H;��H;R�H;��H;.�H;C�H;}�H;��H;��H;��H;��H;��H;}�H;C�H;.�H;��H;R�H;��H;�H;9�H;	�H;��H;��H;w�H;��H;Y�H;Q�H;U�H;��H;��H;ϸH;��H;�H;ÖH;p�H;/eH;�<H;�H;��G;��G;�7G;��F;G�F;SvF;4TF;      =�G;��G;0�G;��G;�H;�/H;�KH;?eH;`{H;i�H;m�H;d�H;o�H;��H;žH;3�H;��H;��H;��H;i�H;d�H;��H;#�H;��H;�H;9�H;�H;��H;[�H;��H;��H;<�H;\�H;�H;��H;��H;��H;��H;��H;�H;\�H;<�H;��H;��H;[�H;��H;�H;9�H;�H;��H;#�H;��H;d�H;i�H;��H;��H;��H;3�H;žH;��H;o�H;d�H;m�H;i�H;`{H;?eH;�KH;�/H;�H;��G;0�G;��G;      �kH;[mH;�qH;�xH;s�H;ȊH;�H;ʜH;��H; �H;��H;�H;&�H;��H;��H;K�H;Y�H;��H;��H;x�H;��H;��H;�H;G�H;T�H;�H;��H;B�H;��H;��H;�H;B�H;k�H;l�H;��H;��H;��H;��H;��H;l�H;k�H;B�H;�H;��H;��H;B�H;��H;�H;T�H;G�H;�H;��H;��H;x�H;��H;��H;Y�H;K�H;��H;��H;&�H;�H;��H; �H;��H;ʜH;�H;ȊH;s�H;�xH;�qH;[mH;      4�H;ϠH;[�H;ĤH;��H;��H;��H;�H;��H;H�H;��H;J�H;b�H;J�H;�H;2�H;��H;h�H;��H;��H;<�H;�H;��H;��H;8�H;��H;[�H;��H;��H;�H;6�H;S�H;j�H;l�H;j�H;u�H;v�H;u�H;j�H;l�H;j�H;S�H;6�H;�H;��H;��H;[�H;��H;8�H;��H;��H;�H;<�H;��H;��H;h�H;��H;2�H;�H;J�H;b�H;J�H;��H;H�H;��H;�H;��H;��H;��H;ĤH;[�H;ϠH;      ��H;ݶH;��H;8�H;*�H;��H;S�H;N�H;W�H;��H;��H;��H;��H;n�H;��H;�H;;�H;�H;��H;��H;��H;�H;��H;~�H;�H;R�H;��H;��H;�H;+�H;J�H;I�H;Y�H;h�H;P�H;b�H;{�H;b�H;P�H;h�H;Y�H;I�H;J�H;+�H;�H;��H;��H;R�H;�H;~�H;��H;�H;��H;��H;��H;�H;;�H;�H;��H;n�H;��H;��H;��H;��H;W�H;N�H;S�H;��H;*�H;8�H;��H;ݶH;      i�H;��H;=�H;J�H;��H;.�H;�H;��H;�H;N�H;v�H;��H;��H;|�H;B�H;��H;x�H;��H;��H;��H;��H;4�H;��H;(�H;��H;��H;��H;�H;6�H;J�H;a�H;T�H;E�H;E�H;c�H;U�H;6�H;U�H;c�H;E�H;E�H;T�H;a�H;J�H;6�H;�H;��H;��H;��H;(�H;��H;4�H;��H;��H;��H;��H;x�H;��H;B�H;|�H;��H;��H;v�H;N�H;�H;��H;�H;.�H;��H;J�H;=�H;��H;      ��H;��H;�H;��H;��H;��H;(�H;��H;�H;��H;�H;��H;��H;S�H;��H;��H;��H;��H;b�H;$�H;��H;�H;��H;��H;��H;.�H;<�H;B�H;S�H;I�H;T�H;Z�H;D�H;=�H;O�H;4�H;+�H;4�H;O�H;=�H;D�H;Z�H;T�H;I�H;S�H;B�H;<�H;.�H;��H;��H;��H;�H;��H;$�H;b�H;��H;��H;��H;��H;S�H;��H;��H;�H;��H;�H;��H;(�H;��H;��H;��H;�H;��H;      ��H;��H;�H;��H;)�H;��H;��H;��H;��H;��H;��H;�H;�H;�H;��H;��H;i�H;�H;��H; �H;m�H;��H;��H;,�H;=�H;C�H;\�H;k�H;j�H;Y�H;E�H;D�H;H�H;C�H;#�H;#�H;S�H;#�H;#�H;C�H;H�H;D�H;E�H;Y�H;j�H;k�H;\�H;C�H;=�H;,�H;��H;��H;m�H; �H;��H;�H;i�H;��H;��H;�H;�H;�H;��H;��H;��H;��H;��H;��H;)�H;��H;�H;��H;      p�H;�H;��H;��H;��H;�H;��H;{�H;9�H;��H;��H;n�H;'�H;��H;��H;,�H;��H;�H;w�H;��H;��H;1�H;L�H;l�H;��H;}�H;�H;l�H;l�H;h�H;E�H;=�H;C�H;-�H;�H;$�H;)�H;$�H;�H;-�H;C�H;=�H;E�H;h�H;l�H;l�H;�H;}�H;��H;l�H;L�H;1�H;��H;��H;w�H;�H;��H;,�H;��H;��H;'�H;n�H;��H;��H;9�H;{�H;��H;�H;��H;��H;��H;�H;      ��H;��H;��H;�H;p�H;��H;A�H;��H;S�H;��H;��H;�H;��H;*�H;��H;�H;Y�H;��H;�H;@�H;Y�H;r�H;��H;��H;��H;��H;��H;��H;j�H;P�H;c�H;O�H;#�H;�H;'�H;�H;�H;�H;'�H;�H;#�H;O�H;c�H;P�H;j�H;��H;��H;��H;��H;��H;��H;r�H;Y�H;@�H;�H;��H;Y�H;�H;��H;*�H;��H;�H;��H;��H;S�H;��H;A�H;��H;p�H;�H;��H;��H;      )�H;<�H;j�H;��H;��H;-�H;��H;�H;��H;�H;��H; �H;o�H;��H;B�H;��H;��H;�H;I�H;{�H;��H;��H;��H;��H;��H;��H;��H;��H;u�H;b�H;U�H;4�H;#�H;$�H;�H;�H;�H;�H;�H;$�H;#�H;4�H;U�H;b�H;u�H;��H;��H;��H;��H;��H;��H;��H;��H;{�H;I�H;�H;��H;��H;B�H;��H;o�H; �H;��H;�H;��H;�H;��H;-�H;��H;��H;j�H;<�H;      ��H;��H;��H;7�H;�H;��H;5�H;��H;�H;i�H;��H;?�H;��H;�H;u�H;��H;�H;<�H;c�H;{�H;��H;��H;��H;��H;��H;��H;��H;��H;v�H;{�H;6�H;+�H;S�H;)�H;�H;�H;�H;�H;�H;)�H;S�H;+�H;6�H;{�H;v�H;��H;��H;��H;��H;��H;��H;��H;��H;{�H;c�H;<�H;�H;��H;u�H;�H;��H;?�H;��H;i�H;�H;��H;5�H;��H;�H;7�H;��H;��H;      )�H;<�H;j�H;��H;��H;-�H;��H;�H;��H;�H;��H; �H;o�H;��H;B�H;��H;��H;�H;I�H;{�H;��H;��H;��H;��H;��H;��H;��H;��H;u�H;b�H;U�H;4�H;#�H;$�H;�H;�H;�H;�H;�H;$�H;#�H;4�H;U�H;b�H;u�H;��H;��H;��H;��H;��H;��H;��H;��H;{�H;I�H;�H;��H;��H;B�H;��H;o�H; �H;��H;�H;��H;�H;��H;-�H;��H;��H;j�H;<�H;      ��H;��H;��H;�H;p�H;��H;A�H;��H;S�H;��H;��H;�H;��H;*�H;��H;�H;Y�H;��H;�H;@�H;Y�H;r�H;��H;��H;��H;��H;��H;��H;j�H;P�H;c�H;O�H;#�H;�H;'�H;�H;�H;�H;'�H;�H;#�H;O�H;c�H;P�H;j�H;��H;��H;��H;��H;��H;��H;r�H;Y�H;@�H;�H;��H;Y�H;�H;��H;*�H;��H;�H;��H;��H;S�H;��H;A�H;��H;p�H;�H;��H;��H;      p�H;�H;��H;��H;��H;�H;��H;{�H;9�H;��H;��H;n�H;'�H;��H;��H;,�H;��H;�H;w�H;��H;��H;1�H;L�H;l�H;��H;}�H;�H;l�H;l�H;h�H;E�H;=�H;C�H;-�H;�H;$�H;)�H;$�H;�H;-�H;C�H;=�H;E�H;h�H;l�H;l�H;�H;}�H;��H;l�H;L�H;1�H;��H;��H;w�H;�H;��H;,�H;��H;��H;'�H;n�H;��H;��H;9�H;{�H;��H;�H;��H;��H;��H;�H;      ��H;��H;�H;��H;)�H;��H;��H;��H;��H;��H;��H;�H;�H;�H;��H;��H;i�H;�H;��H; �H;m�H;��H;��H;,�H;=�H;C�H;\�H;k�H;j�H;Y�H;E�H;D�H;H�H;C�H;#�H;#�H;S�H;#�H;#�H;C�H;H�H;D�H;E�H;Y�H;j�H;k�H;\�H;C�H;=�H;,�H;��H;��H;m�H; �H;��H;�H;i�H;��H;��H;�H;�H;�H;��H;��H;��H;��H;��H;��H;)�H;��H;�H;��H;      ��H;��H;�H;��H;��H;��H;(�H;��H;�H;��H;�H;��H;��H;S�H;��H;��H;��H;��H;b�H;$�H;��H;�H;��H;��H;��H;.�H;<�H;B�H;S�H;I�H;T�H;Z�H;D�H;=�H;O�H;4�H;+�H;4�H;O�H;=�H;D�H;Z�H;T�H;I�H;S�H;B�H;<�H;.�H;��H;��H;��H;�H;��H;$�H;b�H;��H;��H;��H;��H;S�H;��H;��H;�H;��H;�H;��H;(�H;��H;��H;��H;�H;��H;      i�H;��H;=�H;J�H;��H;.�H;�H;��H;�H;N�H;v�H;��H;��H;|�H;B�H;��H;x�H;��H;��H;��H;��H;4�H;��H;(�H;��H;��H;��H;�H;6�H;J�H;a�H;T�H;E�H;E�H;c�H;U�H;6�H;U�H;c�H;E�H;E�H;T�H;a�H;J�H;6�H;�H;��H;��H;��H;(�H;��H;4�H;��H;��H;��H;��H;x�H;��H;B�H;|�H;��H;��H;v�H;N�H;�H;��H;�H;.�H;��H;J�H;=�H;��H;      ��H;ݶH;��H;8�H;*�H;��H;S�H;N�H;W�H;��H;��H;��H;��H;n�H;��H;�H;;�H;�H;��H;��H;��H;�H;��H;~�H;�H;R�H;��H;��H;�H;+�H;J�H;I�H;Y�H;h�H;P�H;b�H;{�H;b�H;P�H;h�H;Y�H;I�H;J�H;+�H;�H;��H;��H;R�H;�H;~�H;��H;�H;��H;��H;��H;�H;;�H;�H;��H;n�H;��H;��H;��H;��H;W�H;N�H;S�H;��H;*�H;8�H;��H;ݶH;      4�H;ϠH;[�H;ĤH;��H;��H;��H;�H;��H;H�H;��H;J�H;b�H;J�H;�H;2�H;��H;h�H;��H;��H;<�H;�H;��H;��H;8�H;��H;[�H;��H;��H;�H;6�H;S�H;j�H;l�H;j�H;u�H;v�H;u�H;j�H;l�H;j�H;S�H;6�H;�H;��H;��H;[�H;��H;8�H;��H;��H;�H;<�H;��H;��H;h�H;��H;2�H;�H;J�H;b�H;J�H;��H;H�H;��H;�H;��H;��H;��H;ĤH;[�H;ϠH;      �kH;[mH;�qH;�xH;s�H;ȊH;�H;ʜH;��H; �H;��H;�H;&�H;��H;��H;K�H;Y�H;��H;��H;x�H;��H;��H;�H;G�H;T�H;�H;��H;B�H;��H;��H;�H;B�H;k�H;l�H;��H;��H;��H;��H;��H;l�H;k�H;B�H;�H;��H;��H;B�H;��H;�H;T�H;G�H;�H;��H;��H;x�H;��H;��H;Y�H;K�H;��H;��H;&�H;�H;��H; �H;��H;ʜH;�H;ȊH;s�H;�xH;�qH;[mH;      =�G;��G;0�G;��G;�H;�/H;�KH;?eH;`{H;i�H;m�H;d�H;o�H;��H;žH;3�H;��H;��H;��H;i�H;d�H;��H;#�H;��H;�H;9�H;�H;��H;[�H;��H;��H;<�H;\�H;�H;��H;��H;��H;��H;��H;�H;\�H;<�H;��H;��H;[�H;��H;�H;9�H;�H;��H;#�H;��H;d�H;i�H;��H;��H;��H;3�H;žH;��H;o�H;d�H;m�H;i�H;`{H;?eH;�KH;�/H;�H;��G;0�G;��G;      VHF;4TF;SvF;G�F;��F;�7G;��G;��G;�H;�<H;/eH;p�H;ÖH;�H;��H;ϸH;��H;��H;U�H;Q�H;Y�H;��H;w�H;��H;��H;	�H;9�H;�H;��H;R�H;��H;.�H;C�H;}�H;��H;��H;��H;��H;��H;}�H;C�H;.�H;��H;R�H;��H;�H;9�H;	�H;��H;��H;w�H;��H;Y�H;Q�H;U�H;��H;��H;ϸH;��H;�H;ÖH;p�H;/eH;�<H;�H;��G;��G;�7G;��F;G�F;SvF;4TF;      �B;.�B;�C;ՏC;�/D;��D;1�E;�HF;��F;GiG;S�G;t#H;�[H;/�H;��H;�H;I�H;μH;��H;e�H;��H;��H;�H;5�H;��H;��H;�H;T�H;8�H;�H;��H;��H;=�H;��H;��H;��H;��H;��H;��H;��H;=�H;��H;��H;�H;8�H;T�H;�H;��H;��H;5�H;�H;��H;��H;e�H;��H;μH;I�H;�H;��H;/�H;�[H;t#H;S�G;GiG;��F;�HF;1�E;��D;�/D;ՏC;�C;.�B;      D�:;\�:;��;;'�<;3>;�?;FIA;��B;DED;6{E;WvF;�7G;��G;q&H;eH;s�H;_�H;m�H;��H;��H;�H;:�H;�H;��H;5�H;��H;��H;G�H;��H;~�H;(�H;��H;,�H;l�H;��H;��H;��H;��H;��H;l�H;,�H;��H;(�H;~�H;��H;G�H;��H;��H;5�H;��H;�H;:�H;�H;��H;��H;m�H;_�H;s�H;eH;q&H;��G;�7G;WvF;6{E;DED;��B;FIA;�?;3>;'�<;��;;\�:;      *;��*;�,;�c.;�X1;$�4;E+8;ӊ;;~�>;IA;jwC;�)E;kF;�MG;'�G;DH;"{H;A�H;��H;@�H;S�H;Y�H;��H;�H;�H;w�H;#�H;�H;��H;��H;��H;��H;��H;L�H;��H;��H;��H;��H;��H;L�H;��H;��H;��H;��H;��H;�H;#�H;w�H;�H;�H;��H;Y�H;S�H;@�H;��H;A�H;"{H;DH;'�G;�MG;kF;�)E;jwC;IA;~�>;ӊ;;E+8;$�4;�X1;�c.;�,;��*;      ��
;��;J�;\;��;7`;�C&;�-;�C3;t�8;?H=;��@;�C;d{E;��F;�G;k#H;,mH;��H;?�H;��H;��H;Y�H;:�H;��H;��H;��H;��H;�H;�H;4�H;�H;��H;1�H;r�H;��H;��H;��H;r�H;1�H;��H;�H;4�H;�H;�H;��H;��H;��H;��H;:�H;Y�H;��H;��H;?�H;��H;,mH;k#H;�G;��F;d{E;�C;��@;?H=;t�8;�C3;�-;�C&;7`;��;\;J�;��;      ]�:���:��:Ӳ�:���:PO�:�z;i';4�;�}(;�X1;6t8;��=;Z�A;��D;&HF;�bG;�H;>cH;��H;n�H;��H;S�H;�H;��H;Y�H;d�H;��H;<�H;��H;��H;��H;m�H;��H;Y�H;��H;��H;��H;Y�H;��H;m�H;��H;��H;��H;<�H;��H;d�H;Y�H;��H;�H;S�H;��H;n�H;��H;>cH;�H;�bG;&HF;��D;Z�A;��=;6t8;�X1;�}(;4�;i';�z;PO�:���:Ӳ�:��:���:      �R�� �B�7��<^9��:Q�X:���:���:�O�:>�;7�;�);�C3;��:;� @;�C;k�E;8G;��G;�_H;��H;?�H;@�H;��H;e�H;Q�H;i�H;x�H;��H;��H;��H;$�H; �H;��H;@�H;{�H;{�H;{�H;@�H;��H; �H;$�H;��H;��H;��H;x�H;i�H;Q�H;e�H;��H;@�H;?�H;��H;�_H;��G;8G;k�E;�C;� @;��:;�C3;�);7�;>�;�O�:���:���:Q�X:��:�<^9B�7�� �      ��)���$�����������<�\�S���N�9�1j:a��:���:ۃ;�� ;%d.;+8;��>;qC;��E;�(G;��G;>cH;��H;��H;��H;��H;U�H;��H;��H;��H;��H;��H;b�H;��H;w�H;�H;I�H;c�H;I�H;�H;w�H;��H;b�H;��H;��H;��H;��H;��H;U�H;��H;��H;��H;��H;>cH;��G;�(G;��E;qC;��>;+8;%d.;�� ;ۃ;���:a��:�1j:�N�9S��<�\�������������$�      q�ѻ�ͻP���mG�������d�*�$��Jɺ̇!��C^9��r:���:`0;y�;l�*;�Y6;>;o�B;��E;8G;�H;,mH;A�H;m�H;μH;��H;��H;��H;h�H;�H;��H;��H;�H;�H;��H;�H;<�H;�H;��H;�H;�H;��H;��H;�H;h�H;��H;��H;��H;μH;m�H;A�H;,mH;�H;8G;��E;o�B;>;�Y6;l�*;y�;`0;���:��r:�C^9̇!��Jɺ*�$���d����mG��P����ͻ      ��I�1�E��(;��O*�����<��?GĻ��t@�JҺy��:�:�O�:O�;!~(;S�5;>;qC;k�E;�bG;k#H;"{H;_�H;I�H;��H;��H;Y�H;��H;;�H;x�H;��H;i�H;��H;Y�H;��H;�H;��H;Y�H;��H;i�H;��H;x�H;;�H;��H;Y�H;��H;��H;I�H;_�H;"{H;k#H;�bG;k�E;qC;>;S�5;!~(;O�;�O�:�:��:y��JҺt@���?GĻ�<������O*��(;�1�E�      &p��\x��ע��R��%��n�`��7�F��G�ѻ-��˃$��ǅ���09�:���:�;!~(;�Y6;��>;�C;&HF;�G;DH;s�H;�H;ϸH;3�H;K�H;2�H;�H;��H;��H;��H;,�H;�H;��H;��H;��H;�H;,�H;��H;��H;��H;�H;2�H;K�H;3�H;ϸH;�H;s�H;DH;�G;&HF;�C;��>;�Y6;!~(;�;���:�:��09�ǅ�˃$�-��G�ѻF���7�n�`�%���R��ע�\x��      &]� �$#�����u�ټ�ɺ������
v��(;�ר�c^��P6R����W	7����:���:O�;l�*;+8;� @;��D;��F;'�G;eH;��H;��H;žH;��H;�H;��H;B�H;��H;��H;��H;��H;B�H;u�H;B�H;��H;��H;��H;��H;B�H;��H;�H;��H;žH;��H;��H;eH;'�G;��F;��D;� @;+8;l�*;O�;���:���:W	7����P6R�c^��ר��(;��
v������ɺ�u�ټ����$#� �      ��_�\�<Q��f@�t +��5�����P�ļs�\�`����bͻek��IɺW	7��:�O�:y�;%d.;��:;Z�A;d{E;�MG;q&H;/�H;�H;��H;��H;J�H;n�H;|�H;S�H;�H;��H;*�H;��H;�H;��H;*�H;��H;�H;S�H;|�H;n�H;J�H;��H;��H;�H;/�H;q&H;�MG;d{E;Z�A;��:;%d.;y�;�O�:�:W	7��Iɺek�bͻ���\�`�s�P�ļ�����5�t +��f@�<Q�\�      �@���R��ڟ�绒�C����_�:�������$p���vz��O*�5ֻek������09�:`0;�� ;�C3;��=;�C;kF;��G;�[H;ÖH;o�H;&�H;b�H;��H;��H;��H;�H;'�H;��H;o�H;��H;o�H;��H;'�H;�H;��H;��H;��H;b�H;&�H;o�H;ÖH;�[H;��G;kF;�C;��=;�C3;�� ;`0;�:��09���ek�5ֻ�O*��vz�$p����輙��:���_�C��绒�ڟ��R��      �` �j.��m��ڽ�b��gr��O��\�m +�� ��ɺ�<��O*�bͻP6R��ǅ���:���:ۃ;�);6t8;��@;�)E;�7G;t#H;p�H;d�H;�H;J�H;��H;��H;��H;�H;n�H;�H; �H;?�H; �H;�H;n�H;�H;��H;��H;��H;J�H;�H;d�H;p�H;t#H;�7G;�)E;��@;6t8;�);ۃ;���:��:�ǅ�P6R�bͻ�O*�<��ɺ�� �m +�\�O��gr���b����ڽm��j.��      �-=�1�9��k/�"�����i��y�Ľ�!��Tys�4�6�#��ɺ��vz����c^��˃$�y����r:���:7�;�X1;?H=;jwC;WvF;S�G;/eH;m�H;��H;��H;��H;v�H;�H;��H;��H;��H;��H;��H;��H;��H;��H;��H;�H;v�H;��H;��H;��H;m�H;/eH;S�G;WvF;jwC;?H=;�X1;7�;���:��r:y��˃$�c^������vz��ɺ�#�4�6�Tys��!��y�Ľi���"���k/�1�9�      �(��;l���.}�&ce�jPH���(�o
���ڽ�R����{�4�6�� �$p��\�`�ר�-��JҺ�C^9a��:>�;�}(;t�8;IA;6{E;GiG;�<H;i�H; �H;H�H;��H;N�H;��H;��H;��H;��H;�H;i�H;�H;��H;��H;��H;��H;N�H;��H;H�H; �H;i�H;�<H;GiG;6{E;IA;t�8;�}(;>�;a��:�C^9JҺ-��ר�\�`�$p��� �4�6���{��R����ڽo
���(�jPH�&ce��.}�;l��      �iþGD��)o���������� �i��-=�[t����R��Tys�m +����s񗼗(;�G�ѻt@�̇!��1j:�O�:4�;�C3;~�>;DED;��F;�H;`{H;��H;��H;W�H;�H;�H;��H;9�H;S�H;��H;�H;��H;S�H;9�H;��H;�H;�H;W�H;��H;��H;`{H;�H;��F;DED;~�>;�C3;4�;�O�:�1j:̇!�t@�G�ѻ�(;�s����m +�Tys��R����[t��-=� �i���������)o��GD��      ���
������޾HD���A���.}��D�[t���ڽ�!��\����P�ļ�
v�F�����Jɺ�N�9���:i';�-;ӊ;;��B;�HF;��G;?eH;ʜH;�H;N�H;��H;��H;��H;{�H;��H;�H;��H;�H;��H;{�H;��H;��H;��H;N�H;�H;ʜH;?eH;��G;�HF;��B;ӊ;;�-;i';���:�N�9�Jɺ��F���
v�P�ļ���\��!����ڽ[t��D��.}��A��HD���޾�����
�      ��7�Õ3��f'���\���о�����.}��-=�o
�y�ĽO��:����������7�?GĻ*�$�S�����:�z;�C&;E+8;FIA;1�E;��G;�KH;�H;��H;S�H;�H;(�H;��H;��H;A�H;��H;5�H;��H;A�H;��H;��H;(�H;�H;S�H;��H;�H;�KH;��G;1�E;FIA;E+8;�C&;�z;���:S��*�$�?GĻ�7���������:�O��y�Ľo
��-=��.}������о�\����f'�Õ3�      Io�PXi�s"Y���@�@�#��
��о�A�� �i���(�i��gr����_��5��ɺ�n�`��<����d�<�\�Q�X:PO�:7`;$�4;�?;��D;�7G;�/H;ȊH;��H;��H;.�H;��H;��H;�H;��H;-�H;��H;-�H;��H;�H;��H;��H;.�H;��H;��H;ȊH;�/H;�7G;��D;�?;$�4;7`;PO�:Q�X:<�\���d��<��n�`��ɺ��5���_�gr��i����(� �i��A���о�
�@�#���@�s"Y�PXi�      &����������Io��!J�@�#��\��HD������jPH�����b��C��t +�u�ټ%��������������:���:��;�X1;3>;�/D;��F;�H;s�H;��H;*�H;��H;��H;)�H;��H;p�H;��H;�H;��H;p�H;��H;)�H;��H;��H;*�H;��H;s�H;�H;��F;�/D;3>;�X1;��;���:��:����������%��u�ټt +�C���b�����jPH�����HD���\��@�#��!J�Io��������      2^������b���Io���@���޾����&ce�"����ڽ绒��f@������R���O*�mG������<^9Ӳ�:\;�c.;'�<;ՏC;G�F;��G;�xH;ĤH;8�H;J�H;��H;��H;��H;�H;��H;7�H;��H;�H;��H;��H;��H;J�H;8�H;ĤH;�xH;��G;G�F;ՏC;'�<;�c.;\;Ӳ�:�<^9���mG���O*��R�������f@�绒���ڽ"��&ce������޾���@�Io�b�������      �aǿ֊¿���������s"Y��f'�����)o���.}��k/�m��ڟ�<Q�$#�ע��(;�P������B�7���:J�;�,;��;;�C;SvF;0�G;�qH;[�H;��H;=�H;�H;�H;��H;��H;j�H;��H;j�H;��H;��H;�H;�H;=�H;��H;[�H;�qH;0�G;SvF;�C;��;;�,;J�;��:B�7����P����(;�ע�$#�<Q�ڟ�m���k/��.}�)o�������f'�s"Y����������֊¿      %�ֿ5pѿ֊¿������PXi�Õ3��
�GD��;l��1�9�j.���R��\� �\x��1�E��ͻ��$�� ����:��;��*;\�:;.�B;4TF;��G;[mH;ϠH;ݶH;��H;��H;��H;�H;��H;<�H;��H;<�H;��H;�H;��H;��H;��H;ݶH;ϠH;[mH;��G;4TF;.�B;\�:;��*;��;���:� ���$��ͻ1�E�\x�� �\��R��j.��1�9�;l��GD���
�Õ3�PXi�������֊¿5pѿ      ���$������꿥�ſ�ޞ�3s��2�/����� j���nHͽ������'�B<ͼ��n������Q^�0.��:�V;�R%;n8;��A;nCF;�H;��H;��H;��H;L�H;>�H;C�H;��H;��H;��H;+�H;��H;��H;��H;C�H;>�H;L�H;��H;��H;��H;�H;nCF;��A;n8;�R%;�V;�:0.��Q^�������n�B<ͼ��'�����nHͽ�� j���/����2�3s��ޞ���ſ������$�      $��������~�����cm�L�-�����Fh��Ide�-�̪ɽ�v��#�$���ɼ�mj�o����X�4��oĆ:�w;j�%;M�8;B;{QF;H;5�H;U�H;	�H;q�H;B�H;6�H;��H;��H;��H;$�H;��H;��H;��H;6�H;B�H;q�H;	�H;U�H;5�H;H;{QF;B;M�8;j�%;�w;oĆ:4���X�o����mj���ɼ#�$��v��̪ɽ-�Ide�Fh������L�-�cm����~���忖����      ������{���ԿBw�����/�\��"����b��M0X�}���;����w����������]�W��UF�*��pȒ:1�;_�';؎9;2oB;�yF;� H;��H;8�H;�H;��H;F�H;:�H;��H;��H;��H;�H;��H;��H;��H;:�H;F�H;��H;�H;8�H;��H;� H;�yF;2oB;؎9;_�';1�;pȒ:*��UF�W�黼�]����������w��;��}��M0X�b������"�/�\����Bw���Կ{�𿖏�      ������Կp���ޞ�RF�]�C�$E��;�I��sD�|�"��]�c�y��֯���J�O�ѻ\�)���K����:Q�
;M*;��:;�C;�F;�7H;Z�H;��H;w�H;��H;?�H;:�H;��H;��H;��H;��H;��H;��H;��H;:�H;?�H;��H;w�H;��H;Z�H;�7H;�F;�C;��:;M*;Q�
;���:��K�\�)�O�ѻ��J��֯�y�]�c�"��|�sD��I���;$E�]�C�RF��ޞ�p���Կ��      ��ſ~��Bw���ޞ�|���3�W�,�%�����^ɰ��|x�\{+�ű����J��  �Ҷ��n�1�f����+�
9s�:�;5�-;��<;��C;�G;�SH;R�H;��H;��H;��H;V�H;3�H;��H;��H;��H;��H;��H;��H;��H;3�H;V�H;��H;��H;��H;R�H;�SH;�G;��C;��<;5�-;�;s�:
9�+�f���n�1�Ҷ���  ��J���ű�\{+��|x�^ɰ�����,�%�3�W�|����ޞ�Bw��~��      �ޞ�������RF�3�W�M�-���4Kɾ�G����O�z��ƽ����Ȅ-���ۼㄼK4�[ǐ�+ж��Z:o��:�;˕1;c>;|�D;�[G;KrH;��H;j�H;f�H;'�H;u�H;)�H;i�H;��H;|�H;��H;|�H;��H;i�H;)�H;u�H;'�H;f�H;j�H;��H;KrH;�[G;|�D;c>;˕1;�;o��:�Z:+ж�[ǐ�K4�ㄼ��ۼȄ-�����ƽz����O��G��4Kɾ��M�-�3�W�RF�������      3s�cm�/�\�]�C�,�%����TҾa����i��C(����UP����[�x������Y�k���X���<���k:���:*� ;�5;[Q@;ptE;�G;9�H;M�H;��H;�H;J�H;l�H;$�H;c�H;s�H;X�H;��H;X�H;s�H;c�H;$�H;l�H;J�H;�H;��H;M�H;9�H;�G;ptE;[Q@;�5;*� ;���:��k:��<��X�k����Y����x���[�UP����콡C(���i�a���TҾ��,�%�]�C�/�\�cm�      �2�L�-��"�$E�����4Kɾa��w�s�.�5�y�k㻽�v��z0��;��+��-�*�R����6�jS�L�:��	;��(;6�9;�.B;�CF;YH;ժH;��H;��H;��H;w�H;��H;�H;0�H;C�H;<�H;Y�H;<�H;C�H;0�H;�H;��H;w�H;��H;��H;��H;ժH;YH;�CF;�.B;6�9;��(;��	;L�:jS��6�R���-�*��+���;�z0��v��k㻽y�.�5�w�s�a��4Kɾ����$E��"�L�-�      /�����������;^ɰ��G����i�.�5��	�ĪɽR����J�p���沼��]�I���U
x��
���k:6��:v;��/;�,=;��C;N�F;#HH;��H;(�H;��H;$�H;��H;��H;��H;�H;�H;�H;$�H;�H;�H;�H;��H;��H;��H;$�H;��H;(�H;��H;#HH;N�F;��C;�,=;��/;v;6��:�k:�
��U
x�I�����]��沼p���J�R���Īɽ�	�.�5���i��G��^ɰ��;��徨���      ��Fh��b���I���|x���O��C(�y�Īɽ����IDX�D��'<ͼㄼ�X!�t��gX��K����:�x;8�#;$H6;IQ@;�OE;��G;��H;��H;2�H;��H;��H;��H;v�H;��H;��H;��H;��H;��H;��H;��H;��H;��H;v�H;��H;��H;��H;2�H;��H;��H;��G;�OE;IQ@;$H6;8�#;�x;���:�K�gX�t���X!�ㄼ'<ͼD��IDX�����Īɽy��C(���O��|x��I��b��Fh��       j�Ide�M0X�sD�\{+�z�����k㻽R���IDX������ۼо����;�>ۻ�X���y�?<":K��:��;��-;��;;�B;�yF;�H;��H;|�H;&�H;��H;��H;��H;n�H;��H;��H;��H;��H;z�H;��H;��H;��H;��H;n�H;��H;��H;��H;&�H;|�H;��H;�H;�yF;�B;��;;��-;��;K��:?<":��y��X�>ۻ��;�о����ۼ���IDX�R���k㻽���z��\{+�sD�M0X�Ide�      ��-�}��|�ű�ƽUP���v���J�D����ۼ��u�J������+���sѺ3
9gL�: �;�$;#�5;�?;��D;j[G;eH;��H;��H;��H;��H;!�H;��H;T�H;n�H;Z�H;T�H;a�H;7�H;a�H;T�H;Z�H;n�H;T�H;��H;!�H;��H;��H;��H;��H;eH;j[G;��D;�?;#�5;�$; �;gL�:3
9�sѺ�+������u�J�����ۼD���J��v��UP��ƽű�|�}��-�      nHͽ̪ɽ�;��"����������[�z0�p��'<ͼо��u�J���k��+��(����:�`�:}�;�/;�K<;!C;:lF;��G;�H;�H;�H;�H;A�H;T�H;��H;%�H;/�H;�H;�H;�H;��H;�H;�H;�H;/�H;%�H;��H;T�H;A�H;�H;�H;�H;�H;��G;:lF;!C;�K<;�/;}�;�`�:���:�(�+�k����u�J�о��'<ͼp��z0���[�������"���;��̪ɽ      �����v����w�]�c��J�Ȅ-�x��;缈沼ㄼ��;�����k��56�a��N<Q:ף�:�h;M*;��8;��@;�OE;�tG;DhH;��H;��H;�H;#�H;��H;z�H;��H;��H;��H;��H;��H;��H;��H;��H;��H;��H;��H;��H;��H;z�H;��H;#�H;�H;��H;��H;DhH;�tG;�OE;��@;��8;M*;�h;ף�:N<Q:a��56�k��������;�ㄼ�沼�;�x�Ȅ-��J�]�c���w��v��      ��'�#�$����y��  ���ۼ����+����]��X!�>ۻ�+��+�a���>:]��:@�;[�%;	�5;��>;�'D;�F;� H;8�H;[�H;��H;��H;��H;��H;k�H;��H;��H;��H;��H;h�H;K�H;m�H;K�H;h�H;��H;��H;��H;��H;k�H;��H;��H;��H;��H;[�H;8�H;� H;�F;�'D;��>;	�5;[�%;@�;]��:�>:a��+��+��>ۻ�X!���]��+�������ۼ�  �y����#�$�      B<ͼ��ɼ�����֯�Ҷ��ㄼ��Y�-�*�I���t���X��sѺ�(�N<Q:]��:��
;v�#;��3;�b=;#C;3CF;�G;�H;��H;�H;9�H;��H;X�H;!�H;d�H;��H;b�H;5�H;O�H;	�H;��H;�H;��H;	�H;O�H;5�H;b�H;��H;d�H;!�H;X�H;��H;9�H;�H;��H;�H;�G;3CF;#C;�b=;��3;v�#;��
;]��:N<Q:�(��sѺ�X�t��I���-�*���Y�ㄼҶ���֯�������ɼ      ��n��mj���]���J�n�1�K4�k��R���U
x�gX���y�3
9���:ף�:@�;v�#;w�2;�<;�oB;7�E;��G;�dH;��H;8�H;��H;��H;��H;��H;9�H;F�H;8�H;�H;��H;��H;��H;��H;��H;��H;��H;��H;��H;�H;8�H;F�H;9�H;��H;��H;��H;��H;8�H;��H;�dH;��G;7�E;�oB;�<;w�2;v�#;@�;ף�:���:3
9��y�gX�U
x�R���k��K4�n�1���J���]��mj�      ����o���W��O�ѻf���[ǐ��X��6��
���K�?<":gL�:�`�:�h;[�%;��3;�<;Y/B;��E;�[G;�GH;N�H;��H;b�H;�H;7�H;=�H;��H;�H;�H;��H;��H;��H;]�H;O�H;K�H;'�H;K�H;O�H;]�H;��H;��H;��H;�H;�H;��H;=�H;7�H;�H;b�H;��H;N�H;�GH;�[G;��E;Y/B;�<;��3;[�%;�h;�`�:gL�:?<":�K��
���6��X�[ǐ�f���O�ѻW��o���      �Q^��X�UF�\�)��+�+ж���<�jS��k:���:K��: �;}�;M*;	�5;�b=;�oB;��E;�IG;]7H;s�H;��H;�H;-�H;��H;��H;��H;��H;��H;��H;��H;u�H;P�H;��H;��H;��H;��H;��H;��H;��H;P�H;u�H;��H;��H;��H;��H;��H;��H;��H;-�H;�H;��H;s�H;]7H;�IG;��E;�oB;�b=;	�5;M*;}�; �;K��:���:�k:jS���<�+ж��+�\�)�UF��X�      0.�4��*�깖�K�
9�Z:��k:L�:6��:�x;��;�$;�/;��8;��>;#C;7�E;�[G;]7H;ͤH;�H;&�H;��H;5�H;��H;P�H;��H;��H;��H;z�H;6�H;�H;��H;��H;��H;��H;u�H;��H;��H;��H;��H;�H;6�H;z�H;��H;��H;��H;P�H;��H;5�H;��H;&�H;�H;ͤH;]7H;�[G;7�E;#C;��>;��8;�/;�$;��;�x;6��:L�:��k:�Z:
9��K�*��4��      �:oĆ:pȒ:���:s�:o��:���:��	;v;8�#;��-;#�5;�K<;��@;�'D;3CF;��G;�GH;s�H;�H;��H;P�H;��H;]�H;#�H;��H;��H;��H;[�H;�H;��H;��H;m�H;[�H;*�H;�H;�H;�H;*�H;[�H;m�H;��H;��H;�H;[�H;��H;��H;��H;#�H;]�H;��H;P�H;��H;�H;s�H;�GH;��G;3CF;�'D;��@;�K<;#�5;��-;8�#;v;��	;���:o��:s�:���:pȒ:oĆ:      �V;�w;1�;Q�
;�;�;*� ;��(;��/;$H6;��;;�?;!C;�OE;�F;�G;�dH;N�H;��H;&�H;P�H;��H;1�H;��H;f�H;�H;��H;b�H;��H;��H;��H;B�H;�H;�H;��H;��H;��H;��H;��H;�H;�H;B�H;��H;��H;��H;b�H;��H;�H;f�H;��H;1�H;��H;P�H;&�H;��H;N�H;�dH;�G;�F;�OE;!C;�?;��;;$H6;��/;��(;*� ;�;�;Q�
;1�;�w;      �R%;j�%;_�';M*;5�-;˕1;�5;6�9;�,=;IQ@;�B;��D;:lF;�tG;� H;�H;��H;��H;�H;��H;��H;1�H;�H;b�H;��H;r�H;5�H;��H;��H;��H;�H;��H;��H;��H;}�H;e�H;L�H;e�H;}�H;��H;��H;��H;�H;��H;��H;��H;5�H;r�H;��H;b�H;�H;1�H;��H;��H;�H;��H;��H;�H;� H;�tG;:lF;��D;�B;IQ@;�,=;6�9;�5;˕1;5�-;M*;_�';j�%;      n8;M�8;؎9;��:;��<;c>;[Q@;�.B;��C;�OE;�yF;j[G;��G;DhH;8�H;��H;8�H;b�H;-�H;5�H;]�H;��H;b�H;k�H;j�H;D�H;��H;��H;e�H;	�H;��H;��H;Y�H;(�H;"�H;�H;��H;�H;"�H;(�H;Y�H;��H;��H;	�H;e�H;��H;��H;D�H;j�H;k�H;b�H;��H;]�H;5�H;-�H;b�H;8�H;��H;8�H;DhH;��G;j[G;�yF;�OE;��C;�.B;[Q@;c>;��<;��:;؎9;M�8;      ��A;B;2oB;�C;��C;|�D;ptE;�CF;N�F;��G;�H;eH;�H;��H;[�H;�H;��H;�H;��H;��H;#�H;f�H;��H;j�H;-�H;��H;��H;i�H; �H;��H;r�H;@�H;�H;��H;��H;��H;��H;��H;��H;��H;�H;@�H;r�H;��H; �H;i�H;��H;��H;-�H;j�H;��H;f�H;#�H;��H;��H;�H;��H;�H;[�H;��H;�H;eH;�H;��G;N�F;�CF;ptE;|�D;��C;�C;2oB;B;      nCF;{QF;�yF;�F;�G;�[G;�G;YH;#HH;��H;��H;��H;�H;��H;��H;9�H;��H;7�H;��H;P�H;��H;�H;r�H;D�H;��H;��H;_�H;��H;��H;a�H;�H;��H;��H;��H;p�H;\�H;n�H;\�H;p�H;��H;��H;��H;�H;a�H;��H;��H;_�H;��H;��H;D�H;r�H;�H;��H;P�H;��H;7�H;��H;9�H;��H;��H;�H;��H;��H;��H;#HH;YH;�G;�[G;�G;�F;�yF;{QF;      �H;H;� H;�7H;�SH;KrH;9�H;ժH;��H;��H;|�H;��H;�H;�H;��H;��H;��H;=�H;��H;��H;��H;��H;5�H;��H;��H;_�H;��H;��H;H�H;�H;��H;��H;b�H;D�H;(�H;�H;�H;�H;(�H;D�H;b�H;��H;��H;�H;H�H;��H;��H;_�H;��H;��H;5�H;��H;��H;��H;��H;=�H;��H;��H;��H;�H;�H;��H;|�H;��H;��H;ժH;9�H;KrH;�SH;�7H;� H;H;      ��H;5�H;��H;Z�H;R�H;��H;M�H;��H;(�H;2�H;&�H;��H;�H;#�H;��H;X�H;��H;��H;��H;��H;��H;b�H;��H;��H;i�H;��H;��H;W�H;�H;��H;u�H;F�H;!�H;��H;��H;��H;��H;��H;��H;��H;!�H;F�H;u�H;��H;�H;W�H;��H;��H;i�H;��H;��H;b�H;��H;��H;��H;��H;��H;X�H;��H;#�H;�H;��H;&�H;2�H;(�H;��H;M�H;��H;R�H;Z�H;��H;5�H;      ��H;U�H;8�H;��H;��H;j�H;��H;��H;��H;��H;��H;��H;A�H;��H;��H;!�H;9�H;�H;��H;��H;[�H;��H;��H;e�H; �H;��H;H�H;�H;��H;k�H;7�H;��H;��H;��H;��H;��H;�H;��H;��H;��H;��H;��H;7�H;k�H;��H;�H;H�H;��H; �H;e�H;��H;��H;[�H;��H;��H;�H;9�H;!�H;��H;��H;A�H;��H;��H;��H;��H;��H;��H;j�H;��H;��H;8�H;U�H;      ��H;	�H;�H;w�H;��H;f�H;�H;��H;$�H;��H;��H;!�H;T�H;z�H;k�H;d�H;F�H;�H;��H;z�H;�H;��H;��H;	�H;��H;a�H;�H;��H;k�H;-�H;��H;��H;��H;��H;d�H;K�H;B�H;K�H;d�H;��H;��H;��H;��H;-�H;k�H;��H;�H;a�H;��H;	�H;��H;��H;�H;z�H;��H;�H;F�H;d�H;k�H;z�H;T�H;!�H;��H;��H;$�H;��H;�H;f�H;��H;w�H;�H;	�H;      L�H;q�H;��H;��H;��H;'�H;J�H;w�H;��H;��H;��H;��H;��H;��H;��H;��H;8�H;��H;��H;6�H;��H;��H;�H;��H;r�H;�H;��H;u�H;7�H;��H;��H;��H;w�H;@�H;�H;'�H;(�H;'�H;�H;@�H;w�H;��H;��H;��H;7�H;u�H;��H;�H;r�H;��H;�H;��H;��H;6�H;��H;��H;8�H;��H;��H;��H;��H;��H;��H;��H;��H;w�H;J�H;'�H;��H;��H;��H;q�H;      >�H;B�H;F�H;?�H;V�H;u�H;l�H;��H;��H;v�H;n�H;T�H;%�H;��H;��H;b�H;�H;��H;u�H;�H;��H;B�H;��H;��H;@�H;��H;��H;F�H;��H;��H;��H;_�H;A�H;�H;��H;��H;��H;��H;��H;�H;A�H;_�H;��H;��H;��H;F�H;��H;��H;@�H;��H;��H;B�H;��H;�H;u�H;��H;�H;b�H;��H;��H;%�H;T�H;n�H;v�H;��H;��H;l�H;u�H;V�H;?�H;F�H;B�H;      C�H;6�H;:�H;:�H;3�H;)�H;$�H;�H;��H;��H;��H;n�H;/�H;��H;��H;5�H;��H;��H;P�H;��H;m�H;�H;��H;Y�H;�H;��H;b�H;!�H;��H;��H;w�H;A�H;��H;��H;��H;��H;��H;��H;��H;��H;��H;A�H;w�H;��H;��H;!�H;b�H;��H;�H;Y�H;��H;�H;m�H;��H;P�H;��H;��H;5�H;��H;��H;/�H;n�H;��H;��H;��H;�H;$�H;)�H;3�H;:�H;:�H;6�H;      ��H;��H;��H;��H;��H;i�H;c�H;0�H;�H;��H;��H;Z�H;�H;��H;��H;O�H;��H;]�H;��H;��H;[�H;�H;��H;(�H;��H;��H;D�H;��H;��H;��H;@�H;�H;��H;��H;��H;��H;��H;��H;��H;��H;��H;�H;@�H;��H;��H;��H;D�H;��H;��H;(�H;��H;�H;[�H;��H;��H;]�H;��H;O�H;��H;��H;�H;Z�H;��H;��H;�H;0�H;c�H;i�H;��H;��H;��H;��H;      ��H;��H;��H;��H;��H;��H;s�H;C�H;�H;��H;��H;T�H;�H;��H;h�H;	�H;��H;O�H;��H;��H;*�H;��H;}�H;"�H;��H;p�H;(�H;��H;��H;d�H;�H;��H;��H;��H;��H;��H;��H;��H;��H;��H;��H;��H;�H;d�H;��H;��H;(�H;p�H;��H;"�H;}�H;��H;*�H;��H;��H;O�H;��H;	�H;h�H;��H;�H;T�H;��H;��H;�H;C�H;s�H;��H;��H;��H;��H;��H;      ��H;��H;��H;��H;��H;|�H;X�H;<�H;�H;��H;��H;a�H;�H;��H;K�H;��H;��H;K�H;��H;��H;�H;��H;e�H;�H;��H;\�H;�H;��H;��H;K�H;'�H;��H;��H;��H;��H;��H;��H;��H;��H;��H;��H;��H;'�H;K�H;��H;��H;�H;\�H;��H;�H;e�H;��H;�H;��H;��H;K�H;��H;��H;K�H;��H;�H;a�H;��H;��H;�H;<�H;X�H;|�H;��H;��H;��H;��H;      +�H;$�H;�H;��H;��H;��H;��H;Y�H;$�H;��H;z�H;7�H;��H;��H;m�H;�H;��H;'�H;��H;u�H;�H;��H;L�H;��H;��H;n�H;�H;��H;�H;B�H;(�H;��H;��H;��H;��H;��H;~�H;��H;��H;��H;��H;��H;(�H;B�H;�H;��H;�H;n�H;��H;��H;L�H;��H;�H;u�H;��H;'�H;��H;�H;m�H;��H;��H;7�H;z�H;��H;$�H;Y�H;��H;��H;��H;��H;�H;$�H;      ��H;��H;��H;��H;��H;|�H;X�H;<�H;�H;��H;��H;a�H;�H;��H;K�H;��H;��H;K�H;��H;��H;�H;��H;e�H;�H;��H;\�H;�H;��H;��H;K�H;'�H;��H;��H;��H;��H;��H;��H;��H;��H;��H;��H;��H;'�H;K�H;��H;��H;�H;\�H;��H;�H;e�H;��H;�H;��H;��H;K�H;��H;��H;K�H;��H;�H;a�H;��H;��H;�H;<�H;X�H;|�H;��H;��H;��H;��H;      ��H;��H;��H;��H;��H;��H;s�H;C�H;�H;��H;��H;T�H;�H;��H;h�H;	�H;��H;O�H;��H;��H;*�H;��H;}�H;"�H;��H;p�H;(�H;��H;��H;d�H;�H;��H;��H;��H;��H;��H;��H;��H;��H;��H;��H;��H;�H;d�H;��H;��H;(�H;p�H;��H;"�H;}�H;��H;*�H;��H;��H;O�H;��H;	�H;h�H;��H;�H;T�H;��H;��H;�H;C�H;s�H;��H;��H;��H;��H;��H;      ��H;��H;��H;��H;��H;i�H;c�H;0�H;�H;��H;��H;Z�H;�H;��H;��H;O�H;��H;]�H;��H;��H;[�H;�H;��H;(�H;��H;��H;D�H;��H;��H;��H;@�H;�H;��H;��H;��H;��H;��H;��H;��H;��H;��H;�H;@�H;��H;��H;��H;D�H;��H;��H;(�H;��H;�H;[�H;��H;��H;]�H;��H;O�H;��H;��H;�H;Z�H;��H;��H;�H;0�H;c�H;i�H;��H;��H;��H;��H;      C�H;6�H;:�H;:�H;3�H;)�H;$�H;�H;��H;��H;��H;n�H;/�H;��H;��H;5�H;��H;��H;P�H;��H;m�H;�H;��H;Y�H;�H;��H;b�H;!�H;��H;��H;w�H;A�H;��H;��H;��H;��H;��H;��H;��H;��H;��H;A�H;w�H;��H;��H;!�H;b�H;��H;�H;Y�H;��H;�H;m�H;��H;P�H;��H;��H;5�H;��H;��H;/�H;n�H;��H;��H;��H;�H;$�H;)�H;3�H;:�H;:�H;6�H;      >�H;B�H;F�H;?�H;V�H;u�H;l�H;��H;��H;v�H;n�H;T�H;%�H;��H;��H;b�H;�H;��H;u�H;�H;��H;B�H;��H;��H;@�H;��H;��H;F�H;��H;��H;��H;_�H;A�H;�H;��H;��H;��H;��H;��H;�H;A�H;_�H;��H;��H;��H;F�H;��H;��H;@�H;��H;��H;B�H;��H;�H;u�H;��H;�H;b�H;��H;��H;%�H;T�H;n�H;v�H;��H;��H;l�H;u�H;V�H;?�H;F�H;B�H;      L�H;q�H;��H;��H;��H;'�H;J�H;w�H;��H;��H;��H;��H;��H;��H;��H;��H;8�H;��H;��H;6�H;��H;��H;�H;��H;r�H;�H;��H;u�H;7�H;��H;��H;��H;w�H;@�H;�H;'�H;(�H;'�H;�H;@�H;w�H;��H;��H;��H;7�H;u�H;��H;�H;r�H;��H;�H;��H;��H;6�H;��H;��H;8�H;��H;��H;��H;��H;��H;��H;��H;��H;w�H;J�H;'�H;��H;��H;��H;q�H;      ��H;	�H;�H;w�H;��H;f�H;�H;��H;$�H;��H;��H;!�H;T�H;z�H;k�H;d�H;F�H;�H;��H;z�H;�H;��H;��H;	�H;��H;a�H;�H;��H;k�H;-�H;��H;��H;��H;��H;d�H;K�H;B�H;K�H;d�H;��H;��H;��H;��H;-�H;k�H;��H;�H;a�H;��H;	�H;��H;��H;�H;z�H;��H;�H;F�H;d�H;k�H;z�H;T�H;!�H;��H;��H;$�H;��H;�H;f�H;��H;w�H;�H;	�H;      ��H;U�H;8�H;��H;��H;j�H;��H;��H;��H;��H;��H;��H;A�H;��H;��H;!�H;9�H;�H;��H;��H;[�H;��H;��H;e�H; �H;��H;H�H;�H;��H;k�H;7�H;��H;��H;��H;��H;��H;�H;��H;��H;��H;��H;��H;7�H;k�H;��H;�H;H�H;��H; �H;e�H;��H;��H;[�H;��H;��H;�H;9�H;!�H;��H;��H;A�H;��H;��H;��H;��H;��H;��H;j�H;��H;��H;8�H;U�H;      ��H;5�H;��H;Z�H;R�H;��H;M�H;��H;(�H;2�H;&�H;��H;�H;#�H;��H;X�H;��H;��H;��H;��H;��H;b�H;��H;��H;i�H;��H;��H;W�H;�H;��H;u�H;F�H;!�H;��H;��H;��H;��H;��H;��H;��H;!�H;F�H;u�H;��H;�H;W�H;��H;��H;i�H;��H;��H;b�H;��H;��H;��H;��H;��H;X�H;��H;#�H;�H;��H;&�H;2�H;(�H;��H;M�H;��H;R�H;Z�H;��H;5�H;      �H;H;� H;�7H;�SH;KrH;9�H;ժH;��H;��H;|�H;��H;�H;�H;��H;��H;��H;=�H;��H;��H;��H;��H;5�H;��H;��H;_�H;��H;��H;H�H;�H;��H;��H;b�H;D�H;(�H;�H;�H;�H;(�H;D�H;b�H;��H;��H;�H;H�H;��H;��H;_�H;��H;��H;5�H;��H;��H;��H;��H;=�H;��H;��H;��H;�H;�H;��H;|�H;��H;��H;ժH;9�H;KrH;�SH;�7H;� H;H;      nCF;{QF;�yF;�F;�G;�[G;�G;YH;#HH;��H;��H;��H;�H;��H;��H;9�H;��H;7�H;��H;P�H;��H;�H;r�H;D�H;��H;��H;_�H;��H;��H;a�H;�H;��H;��H;��H;p�H;\�H;n�H;\�H;p�H;��H;��H;��H;�H;a�H;��H;��H;_�H;��H;��H;D�H;r�H;�H;��H;P�H;��H;7�H;��H;9�H;��H;��H;�H;��H;��H;��H;#HH;YH;�G;�[G;�G;�F;�yF;{QF;      ��A;B;2oB;�C;��C;|�D;ptE;�CF;N�F;��G;�H;eH;�H;��H;[�H;�H;��H;�H;��H;��H;#�H;f�H;��H;j�H;-�H;��H;��H;i�H; �H;��H;r�H;@�H;�H;��H;��H;��H;��H;��H;��H;��H;�H;@�H;r�H;��H; �H;i�H;��H;��H;-�H;j�H;��H;f�H;#�H;��H;��H;�H;��H;�H;[�H;��H;�H;eH;�H;��G;N�F;�CF;ptE;|�D;��C;�C;2oB;B;      n8;M�8;؎9;��:;��<;c>;[Q@;�.B;��C;�OE;�yF;j[G;��G;DhH;8�H;��H;8�H;b�H;-�H;5�H;]�H;��H;b�H;k�H;j�H;D�H;��H;��H;e�H;	�H;��H;��H;Y�H;(�H;"�H;�H;��H;�H;"�H;(�H;Y�H;��H;��H;	�H;e�H;��H;��H;D�H;j�H;k�H;b�H;��H;]�H;5�H;-�H;b�H;8�H;��H;8�H;DhH;��G;j[G;�yF;�OE;��C;�.B;[Q@;c>;��<;��:;؎9;M�8;      �R%;j�%;_�';M*;5�-;˕1;�5;6�9;�,=;IQ@;�B;��D;:lF;�tG;� H;�H;��H;��H;�H;��H;��H;1�H;�H;b�H;��H;r�H;5�H;��H;��H;��H;�H;��H;��H;��H;}�H;e�H;L�H;e�H;}�H;��H;��H;��H;�H;��H;��H;��H;5�H;r�H;��H;b�H;�H;1�H;��H;��H;�H;��H;��H;�H;� H;�tG;:lF;��D;�B;IQ@;�,=;6�9;�5;˕1;5�-;M*;_�';j�%;      �V;�w;1�;Q�
;�;�;*� ;��(;��/;$H6;��;;�?;!C;�OE;�F;�G;�dH;N�H;��H;&�H;P�H;��H;1�H;��H;f�H;�H;��H;b�H;��H;��H;��H;B�H;�H;�H;��H;��H;��H;��H;��H;�H;�H;B�H;��H;��H;��H;b�H;��H;�H;f�H;��H;1�H;��H;P�H;&�H;��H;N�H;�dH;�G;�F;�OE;!C;�?;��;;$H6;��/;��(;*� ;�;�;Q�
;1�;�w;      �:oĆ:pȒ:���:s�:o��:���:��	;v;8�#;��-;#�5;�K<;��@;�'D;3CF;��G;�GH;s�H;�H;��H;P�H;��H;]�H;#�H;��H;��H;��H;[�H;�H;��H;��H;m�H;[�H;*�H;�H;�H;�H;*�H;[�H;m�H;��H;��H;�H;[�H;��H;��H;��H;#�H;]�H;��H;P�H;��H;�H;s�H;�GH;��G;3CF;�'D;��@;�K<;#�5;��-;8�#;v;��	;���:o��:s�:���:pȒ:oĆ:      0.�4��*�깖�K�
9�Z:��k:L�:6��:�x;��;�$;�/;��8;��>;#C;7�E;�[G;]7H;ͤH;�H;&�H;��H;5�H;��H;P�H;��H;��H;��H;z�H;6�H;�H;��H;��H;��H;��H;u�H;��H;��H;��H;��H;�H;6�H;z�H;��H;��H;��H;P�H;��H;5�H;��H;&�H;�H;ͤH;]7H;�[G;7�E;#C;��>;��8;�/;�$;��;�x;6��:L�:��k:�Z:
9��K�*��4��      �Q^��X�UF�\�)��+�+ж���<�jS��k:���:K��: �;}�;M*;	�5;�b=;�oB;��E;�IG;]7H;s�H;��H;�H;-�H;��H;��H;��H;��H;��H;��H;��H;u�H;P�H;��H;��H;��H;��H;��H;��H;��H;P�H;u�H;��H;��H;��H;��H;��H;��H;��H;-�H;�H;��H;s�H;]7H;�IG;��E;�oB;�b=;	�5;M*;}�; �;K��:���:�k:jS���<�+ж��+�\�)�UF��X�      ����o���W��O�ѻf���[ǐ��X��6��
���K�?<":gL�:�`�:�h;[�%;��3;�<;Y/B;��E;�[G;�GH;N�H;��H;b�H;�H;7�H;=�H;��H;�H;�H;��H;��H;��H;]�H;O�H;K�H;'�H;K�H;O�H;]�H;��H;��H;��H;�H;�H;��H;=�H;7�H;�H;b�H;��H;N�H;�GH;�[G;��E;Y/B;�<;��3;[�%;�h;�`�:gL�:?<":�K��
���6��X�[ǐ�f���O�ѻW��o���      ��n��mj���]���J�n�1�K4�k��R���U
x�gX���y�3
9���:ף�:@�;v�#;w�2;�<;�oB;7�E;��G;�dH;��H;8�H;��H;��H;��H;��H;9�H;F�H;8�H;�H;��H;��H;��H;��H;��H;��H;��H;��H;��H;�H;8�H;F�H;9�H;��H;��H;��H;��H;8�H;��H;�dH;��G;7�E;�oB;�<;w�2;v�#;@�;ף�:���:3
9��y�gX�U
x�R���k��K4�n�1���J���]��mj�      B<ͼ��ɼ�����֯�Ҷ��ㄼ��Y�-�*�I���t���X��sѺ�(�N<Q:]��:��
;v�#;��3;�b=;#C;3CF;�G;�H;��H;�H;9�H;��H;X�H;!�H;d�H;��H;b�H;5�H;O�H;	�H;��H;�H;��H;	�H;O�H;5�H;b�H;��H;d�H;!�H;X�H;��H;9�H;�H;��H;�H;�G;3CF;#C;�b=;��3;v�#;��
;]��:N<Q:�(��sѺ�X�t��I���-�*���Y�ㄼҶ���֯�������ɼ      ��'�#�$����y��  ���ۼ����+����]��X!�>ۻ�+��+�a���>:]��:@�;[�%;	�5;��>;�'D;�F;� H;8�H;[�H;��H;��H;��H;��H;k�H;��H;��H;��H;��H;h�H;K�H;m�H;K�H;h�H;��H;��H;��H;��H;k�H;��H;��H;��H;��H;[�H;8�H;� H;�F;�'D;��>;	�5;[�%;@�;]��:�>:a��+��+��>ۻ�X!���]��+�������ۼ�  �y����#�$�      �����v����w�]�c��J�Ȅ-�x��;缈沼ㄼ��;�����k��56�a��N<Q:ף�:�h;M*;��8;��@;�OE;�tG;DhH;��H;��H;�H;#�H;��H;z�H;��H;��H;��H;��H;��H;��H;��H;��H;��H;��H;��H;��H;��H;z�H;��H;#�H;�H;��H;��H;DhH;�tG;�OE;��@;��8;M*;�h;ף�:N<Q:a��56�k��������;�ㄼ�沼�;�x�Ȅ-��J�]�c���w��v��      nHͽ̪ɽ�;��"����������[�z0�p��'<ͼо��u�J���k��+��(����:�`�:}�;�/;�K<;!C;:lF;��G;�H;�H;�H;�H;A�H;T�H;��H;%�H;/�H;�H;�H;�H;��H;�H;�H;�H;/�H;%�H;��H;T�H;A�H;�H;�H;�H;�H;��G;:lF;!C;�K<;�/;}�;�`�:���:�(�+�k����u�J�о��'<ͼp��z0���[�������"���;��̪ɽ      ��-�}��|�ű�ƽUP���v���J�D����ۼ��u�J������+���sѺ3
9gL�: �;�$;#�5;�?;��D;j[G;eH;��H;��H;��H;��H;!�H;��H;T�H;n�H;Z�H;T�H;a�H;7�H;a�H;T�H;Z�H;n�H;T�H;��H;!�H;��H;��H;��H;��H;eH;j[G;��D;�?;#�5;�$; �;gL�:3
9�sѺ�+������u�J�����ۼD���J��v��UP��ƽű�|�}��-�       j�Ide�M0X�sD�\{+�z�����k㻽R���IDX������ۼо����;�>ۻ�X���y�?<":K��:��;��-;��;;�B;�yF;�H;��H;|�H;&�H;��H;��H;��H;n�H;��H;��H;��H;��H;z�H;��H;��H;��H;��H;n�H;��H;��H;��H;&�H;|�H;��H;�H;�yF;�B;��;;��-;��;K��:?<":��y��X�>ۻ��;�о����ۼ���IDX�R���k㻽���z��\{+�sD�M0X�Ide�      ��Fh��b���I���|x���O��C(�y�Īɽ����IDX�D��'<ͼㄼ�X!�t��gX��K����:�x;8�#;$H6;IQ@;�OE;��G;��H;��H;2�H;��H;��H;��H;v�H;��H;��H;��H;��H;��H;��H;��H;��H;��H;v�H;��H;��H;��H;2�H;��H;��H;��G;�OE;IQ@;$H6;8�#;�x;���:�K�gX�t���X!�ㄼ'<ͼD��IDX�����Īɽy��C(���O��|x��I��b��Fh��      /�����������;^ɰ��G����i�.�5��	�ĪɽR����J�p���沼��]�I���U
x��
���k:6��:v;��/;�,=;��C;N�F;#HH;��H;(�H;��H;$�H;��H;��H;��H;�H;�H;�H;$�H;�H;�H;�H;��H;��H;��H;$�H;��H;(�H;��H;#HH;N�F;��C;�,=;��/;v;6��:�k:�
��U
x�I�����]��沼p���J�R���Īɽ�	�.�5���i��G��^ɰ��;��徨���      �2�L�-��"�$E�����4Kɾa��w�s�.�5�y�k㻽�v��z0��;��+��-�*�R����6�jS�L�:��	;��(;6�9;�.B;�CF;YH;ժH;��H;��H;��H;w�H;��H;�H;0�H;C�H;<�H;Y�H;<�H;C�H;0�H;�H;��H;w�H;��H;��H;��H;ժH;YH;�CF;�.B;6�9;��(;��	;L�:jS��6�R���-�*��+���;�z0��v��k㻽y�.�5�w�s�a��4Kɾ����$E��"�L�-�      3s�cm�/�\�]�C�,�%����TҾa����i��C(����UP����[�x������Y�k���X���<���k:���:*� ;�5;[Q@;ptE;�G;9�H;M�H;��H;�H;J�H;l�H;$�H;c�H;s�H;X�H;��H;X�H;s�H;c�H;$�H;l�H;J�H;�H;��H;M�H;9�H;�G;ptE;[Q@;�5;*� ;���:��k:��<��X�k����Y����x���[�UP����콡C(���i�a���TҾ��,�%�]�C�/�\�cm�      �ޞ�������RF�3�W�M�-���4Kɾ�G����O�z��ƽ����Ȅ-���ۼㄼK4�[ǐ�+ж��Z:o��:�;˕1;c>;|�D;�[G;KrH;��H;j�H;f�H;'�H;u�H;)�H;i�H;��H;|�H;��H;|�H;��H;i�H;)�H;u�H;'�H;f�H;j�H;��H;KrH;�[G;|�D;c>;˕1;�;o��:�Z:+ж�[ǐ�K4�ㄼ��ۼȄ-�����ƽz����O��G��4Kɾ��M�-�3�W�RF�������      ��ſ~��Bw���ޞ�|���3�W�,�%�����^ɰ��|x�\{+�ű����J��  �Ҷ��n�1�f����+�
9s�:�;5�-;��<;��C;�G;�SH;R�H;��H;��H;��H;V�H;3�H;��H;��H;��H;��H;��H;��H;��H;3�H;V�H;��H;��H;��H;R�H;�SH;�G;��C;��<;5�-;�;s�:
9�+�f���n�1�Ҷ���  ��J���ű�\{+��|x�^ɰ�����,�%�3�W�|����ޞ�Bw��~��      ������Կp���ޞ�RF�]�C�$E��;�I��sD�|�"��]�c�y��֯���J�O�ѻ\�)���K����:Q�
;M*;��:;�C;�F;�7H;Z�H;��H;w�H;��H;?�H;:�H;��H;��H;��H;��H;��H;��H;��H;:�H;?�H;��H;w�H;��H;Z�H;�7H;�F;�C;��:;M*;Q�
;���:��K�\�)�O�ѻ��J��֯�y�]�c�"��|�sD��I���;$E�]�C�RF��ޞ�p���Կ��      ������{���ԿBw�����/�\��"����b��M0X�}���;����w����������]�W��UF�*��pȒ:1�;_�';؎9;2oB;�yF;� H;��H;8�H;�H;��H;F�H;:�H;��H;��H;��H;�H;��H;��H;��H;:�H;F�H;��H;�H;8�H;��H;� H;�yF;2oB;؎9;_�';1�;pȒ:*��UF�W�黼�]����������w��;��}��M0X�b������"�/�\����Bw���Կ{�𿖏�      $��������~�����cm�L�-�����Fh��Ide�-�̪ɽ�v��#�$���ɼ�mj�o����X�4��oĆ:�w;j�%;M�8;B;{QF;H;5�H;U�H;	�H;q�H;B�H;6�H;��H;��H;��H;$�H;��H;��H;��H;6�H;B�H;q�H;	�H;U�H;5�H;H;{QF;B;M�8;j�%;�w;oĆ:4���X�o����mj���ɼ#�$��v��̪ɽ-�Ide�Fh������L�-�cm����~���忖����      �>���8���*�O������˿�o��<�b�=\�+m־^��K�:��J�&��F�B�F���������/��������>:�r�:eo ;�I6;DA;�HF;�MH;�H;!I;�I;I;�I;mI;I;q�H;��H;+�H;��H;q�H;I;mI;�I;I;�I;!I;�H;�MH;�HF;DA;�I6;eo ;�r�:��>:�����/���������F��F�B�&���J�K�:�^��+m־=\�<�b��o���˿����O���*���8�      ��8��4��g&�0��2����<ƿ벗��>]����G�Ѿ�p���*7����"W��MR?�	}�8����s������;�G:���:!;'�6;(kA;�XF;�SH;s�H;!I;�I;�I;�I;GI;�I;e�H;��H;�H;��H;e�H;�I;GI;�I;�I;�I;!I;s�H;�SH;�XF;(kA;'�6;!;���:;�G:���s�����8��	}�MR?�"W�����*7��p��G�Ѿ����>]�벗��<ƿ2���0���g&��4�      ��*��g&��#�o�K[�jL�������M�l5��>ľ
����,��D�撐��5�;�ݼ���q
���x��wk���b:�j�:#;ۖ7;��A;�F;�cH;�I;\!I;I;pI;BI;�I;�I;!�H;x�H;��H;x�H;!�H;�I;�I;BI;pI;I;\!I;�I;�cH;�F;��A;ۖ7;#;�j�:��b:�wk���x��q
���;�ݼ�5�撐��Dὤ�,�
���>ľl5���M����jL��K[�o��#��g&�      O�0��o����˿:1��-�y���6��z �����)�l�+��ͽ!�����&���˼^�k�q���k�X��� �ѳ�:p�;)&;�9;��B;�F;�|H;�I;f!I;5I;�I;�
I;qI;FI;��H;"�H;��H;"�H;��H;FI;qI;�
I;�I;5I;f!I;�I;�|H;�F;��B;�9;)&;p�;ѳ�:�� �k�X�q���^�k���˼��&�!����ͽ+�)�l������z ���6�-�y�:1���˿���o�0��      ����2���K[忭˿�T��蟉�s�R�����E۾̗����M�~�	������j��3�"d��ɆO���׻b�/��
�����:��	;%*;l;;�iC;�&G;�H;�I;
!I;�I;�I;�	I;�I;� I;I�H;��H; �H;��H;I�H;� I;�I;�	I;�I;�I;
!I;�I;�H;�&G;�iC;l;;%*;��	;���:�
��b�/���׻ɆO�"d���3���j����~�	���M�̗���E۾���s�R�蟉��T���˿K[�2���      �˿�<ƿjL��:1��蟉��>]���)��$���ճ���{���,�j��$��Q`I��J��-��4/�S,��ʻ ��!693�:�;o.;1-=;o`D;�G;o�H;�I;@ I;aI;TI;�I;�I;��H;��H;�H;d�H;�H;��H;��H;�I;�I;TI;aI;@ I;�I;o�H;�G;o`D;1-=;o.;�;3�:�!69ʻ �S,��4/�-���J��Q`I�$��j�齞�,���{��ճ��$����)��>]�蟉�:1��jL���<ƿ      �o��벗����-�y�s�R���)�iv��>ľ�]����I�Tl�~��������&�߮Ҽ	�}�VB�!���������!:?)�:Wy;�3;li?;�[E;��G;��H;tI;�I;�I;�I;|I;�I;�H;��H;c�H;��H;c�H;��H;�H;�I;|I;�I;�I;�I;tI;��H;��G;�[E;li?;�3;Wy;?)�:��!:����!���VB�	�}�߮Ҽ��&����~���Tl���I��]���>ľiv���)�s�R�-�y����벗�      <�b��>]���M���6�����$���>ľq��q�Z�+�K9ݽW����L����/F��&�G�\�׻�;�u�Ǌ:�h;6O$;�7;y�A;IF;:BH;��H;�I;nI;xI;I;-I;�I;�H;��H;��H;�H;��H;��H;�H;�I;-I;I;xI;nI;�I;��H;:BH;IF;y�A;�7;6O$;�h;Ǌ:u칸;�\�׻&�G�/F�������L�W��K9ݽ+�q�Z�q���>ľ�$�������6���M��>]�      =\����l5��z ��E۾�ճ��]��q�Z�F?#����A����j�(��Oϼ��������Rnۺr3�9�2�:p�;z�,;��;;C�C;�G;R�H;�
I;� I;�I;GI;/
I;�I;? I;�H;�H;��H;"�H;��H;�H;�H;? I;�I;/
I;GI;�I;� I;�
I;R�H;�G;C�C;��;;z�,;p�;�2�:r3�9Rnۺ��������Oϼ(����j��A�����F?#�q�Z��]���ճ��E۾�z �l5����      +m־G�Ѿ�>ľ����̗����{���I�+����V���{�?�/�.���,��b=���һ�@�8� ���k:D�:$a;��3;Ai?;w1E;��G;p�H;7I;xI;�I;�I;&I;�I;��H;��H;��H;��H;V�H;��H;��H;��H;��H;�I;&I;�I;�I;xI;7I;p�H;��G;w1E;Ai?;��3;$a;D�:��k:8� ��@���һb=��,��.��?�/��{��V�����+���I���{�̗�������>ľG�Ѿ      ^���p��
��)�l���M���,�Tl�K9ݽ�A���{���5��J��;���T[�I?������Q��J�9�:��;:*;5�9;jjB;ۆF;�MH;��H; I;�I;�I;"I;I;@I;_�H;��H;��H;��H;j�H;��H;��H;��H;_�H;@I;I;"I;�I;�I; I;��H;�MH;ۆF;jjB;5�9;:*;��;�:J�9�Q������I?��T[�;���J����5��{��A��K9ݽTl���,���M�)�l�
���p��      K�:��*7���,�+�~�	�j��~���W����j�?�/��J���I��%�k���b.�������<Ǌ:�m�:(;nq3;2�>;8�D;t�G;S�H;I;/ I;�I;�I;�	I;�I;`�H;��H;��H;��H;��H;_�H;��H;��H;��H;��H;`�H;�I;�	I;�I;�I;/ I;I;S�H;t�G;8�D;2�>;nq3;(;�m�:<Ǌ:�����b.����%�k��I���J��?�/���j�W��~���j��~�	�+���,��*7�      �J���D��ͽ���$�������L�(��.��;��%�k����I����/��"/�,�>:���:�A;w�,;��:;>�B;�wF;�;H;��H;
I;�I;�I;BI;�I;�I;��H;s�H;5�H;o�H;��H;l�H;��H;o�H;5�H;s�H;��H;�I;�I;BI;�I;�I;
I;��H;�;H;�wF;>�B;��:;w�,;�A;���:,�>:�"/���/��I����%�k�;��.��(����L����$������ͽ�Dὼ��      &��"W��撐�!�����j�Q`I���&����Oϼ�,���T[����I��;��qk�n:j3�:� ;!&;�6;� @;D1E;�G;��H;�I;�I;OI;I;�	I;;I;u�H;��H;�H;��H;^�H;��H;D�H;��H;^�H;��H;�H;��H;u�H;;I;�	I;I;OI;�I;�I;��H;�G;D1E;� @;�6;!&;� ;j3�:n:�qk�;��I�����T[��,��Oϼ�����&�Q`I���j�!���撐�"W��      F�B�MR?��5���&��3��J��߮Ҽ/F����b=�I?�b.����/��qk����9�ճ:�;K!;m3;��=;��C;*�F;cH;��H;�I;I;�I;$I;�I;�I;D�H;��H;��H;|�H;?�H;|�H;4�H;|�H;?�H;|�H;��H;��H;D�H;�I;�I;$I;�I;I;�I;��H;cH;*�F;��C;��=;m3;K!;�;�ճ:���9�qk���/�b.��I?�b=���/F��߮Ҽ�J���3���&��5�MR?�      F��	}�;�ݼ��˼"d��-��	�}�&�G������һ�������"/�n:�ճ:#�;�a;Ģ0;�<;��B;�HF;vH;,�H;�I;zI;I;8I;Y	I;�I;�H;/�H;T�H;�H;#�H;�H;r�H;5�H;r�H;�H;#�H;�H;T�H;/�H;�H;�I;Y	I;8I;I;zI;�I;,�H;vH;�HF;��B;�<;Ģ0;�a;#�;�ճ:n:�"/���������һ���&�G�	�}�-��"d����˼;�ݼ	}�      ����8����^�k�ɆO�4/�VB�\�׻����@��Q�����,�>:j3�:�;�a;��/;>;;J�A;��E;ʾG;��H;�	I;hI;I;�I;�I;�I;� I;��H;;�H;��H;��H;��H;�H;d�H;)�H;d�H;�H;��H;��H;��H;;�H;��H;� I;�I;�I;�I;I;hI;�	I;��H;ʾG;��E;J�A;>;;��/;�a;�;j3�:,�>:����Q���@����\�׻VB�4/�ɆO�^�k���8��      ������q
�q�����׻S,��!����;�Rnۺ8� �J�9<Ǌ:���:� ;K!;Ģ0;>;;͒A;�oE;}�G;ԍH;��H;�I;9I;ZI; I;�I;oI;��H;=�H;x�H;�H;�H;��H;��H;[�H;1�H;[�H;��H;��H;�H;�H;x�H;=�H;��H;oI;�I; I;ZI;9I;�I;��H;ԍH;}�G;�oE;͒A;>;;Ģ0;K!;� ;���:<Ǌ:J�98� �Rnۺ�;�!���S,����׻q����q
���      �/��s�����x�k�X�b�/�ʻ �����u�r3�9��k:�:�m�:�A;!&;m3;�<;J�A;�oE;isG;�{H;.�H;,I;rI;CI;�I;i	I;�I;L�H;J�H;�H;��H;x�H;��H;��H;��H;l�H;\�H;l�H;��H;��H;��H;x�H;��H;�H;J�H;L�H;�I;i	I;�I;CI;rI;,I;.�H;�{H;isG;�oE;J�A;�<;m3;!&;�A;�m�:�:��k:r3�9u칉���ʻ �b�/�k�X���x�s���      ��������wk��� ��
���!69��!:Ǌ:�2�:D�:��;(;w�,;�6;��=;��B;��E;}�G;�{H;��H;zI;I;�I;XI;�
I;"I;� I;A�H;��H;4�H;��H;�H;��H;��H;��H;~�H;l�H;~�H;��H;��H;��H;�H;��H;4�H;��H;A�H;� I;"I;�
I;XI;�I;I;zI;��H;�{H;}�G;��E;��B;��=;�6;w�,;(;��;D�:�2�:Ǌ:��!:�!69�
���� ��wk����      ��>:;�G:��b:ѳ�:���:3�:?)�:�h;p�;$a;:*;nq3;��:;� @;��C;�HF;ʾG;ԍH;.�H;zI;I;CI;:I;�I;I;VI;�H;��H;��H;p�H;B�H;��H;��H;��H;	�H;��H;y�H;��H;	�H;��H;��H;��H;B�H;p�H;��H;��H;�H;VI;I;�I;:I;CI;I;zI;.�H;ԍH;ʾG;�HF;��C;� @;��:;nq3;:*;$a;p�;�h;?)�:3�:���:ѳ�:��b:;�G:      �r�:���:�j�:p�;��	;�;Wy;6O$;z�,;��3;5�9;2�>;>�B;D1E;*�F;vH;��H;��H;,I;I;CI;�I;6I;�I;�I;��H;�H;G�H;��H;��H;��H;��H;��H;��H;)�H;��H;��H;��H;)�H;��H;��H;��H;��H;��H;��H;G�H;�H;��H;�I;�I;6I;�I;CI;I;,I;��H;��H;vH;*�F;D1E;>�B;2�>;5�9;��3;z�,;6O$;Wy;�;��	;p�;�j�:���:      eo ;!;#;)&;%*;o.;�3;�7;��;;Ai?;jjB;8�D;�wF;�G;cH;,�H;�	I;�I;rI;�I;:I;6I;�I;RI;4�H;��H;��H; �H;��H;�H;��H;x�H;��H;��H;E�H;�H;��H;�H;E�H;��H;��H;x�H;��H;�H;��H; �H;��H;��H;4�H;RI;�I;6I;:I;�I;rI;�I;�	I;,�H;cH;�G;�wF;8�D;jjB;Ai?;��;;�7;�3;o.;%*;)&;#;!;      �I6;'�6;ۖ7;�9;l;;1-=;li?;y�A;C�C;w1E;ۆF;t�G;�;H;��H;��H;�I;hI;9I;CI;XI;�I;�I;RI;E�H;��H;��H;Y�H;$�H;1�H;��H;~�H;e�H;��H;�H;��H;]�H;:�H;]�H;��H;�H;��H;e�H;~�H;��H;1�H;$�H;Y�H;��H;��H;E�H;RI;�I;�I;XI;CI;9I;hI;�I;��H;��H;�;H;t�G;ۆF;w1E;C�C;y�A;li?;1-=;l;;�9;ۖ7;'�6;      DA;(kA;��A;��B;�iC;o`D;�[E;IF;�G;��G;�MH;S�H;��H;�I;�I;zI;I;ZI;�I;�
I;I;�I;4�H;��H;��H;w�H;-�H;@�H;��H;��H;`�H;u�H;��H;O�H;��H;��H;��H;��H;��H;O�H;��H;u�H;`�H;��H;��H;@�H;-�H;w�H;��H;��H;4�H;�I;I;�
I;�I;ZI;I;zI;�I;�I;��H;S�H;�MH;��G;�G;IF;�[E;o`D;�iC;��B;��A;(kA;      �HF;�XF;�F;�F;�&G;�G;��G;:BH;R�H;p�H;��H;I;
I;�I;I;I;�I; I;i	I;"I;VI;��H;��H;��H;w�H;S�H;[�H;��H;��H;j�H;X�H;��H;&�H;��H;A�H;"�H;�H;"�H;A�H;��H;&�H;��H;X�H;j�H;��H;��H;[�H;S�H;w�H;��H;��H;��H;VI;"I;i	I; I;�I;I;I;�I;
I;I;��H;p�H;R�H;:BH;��G;�G;�&G;�F;�F;�XF;      �MH;�SH;�cH;�|H;�H;o�H;��H;��H;�
I;7I; I;/ I;�I;OI;�I;8I;�I;�I;�I;� I;�H;�H;��H;Y�H;-�H;[�H;��H;��H;X�H;[�H;��H;��H;d�H;��H;��H;��H;��H;��H;��H;��H;d�H;��H;��H;[�H;X�H;��H;��H;[�H;-�H;Y�H;��H;�H;�H;� I;�I;�I;�I;8I;�I;OI;�I;/ I; I;7I;�
I;��H;��H;o�H;�H;�|H;�cH;�SH;      �H;s�H;�I;�I;�I;�I;tI;�I;� I;xI;�I;�I;�I;I;$I;Y	I;�I;oI;L�H;A�H;��H;G�H; �H;$�H;@�H;��H;��H;k�H;O�H;��H;��H;;�H;��H;|�H;9�H;
�H;�H;
�H;9�H;|�H;��H;;�H;��H;��H;O�H;k�H;��H;��H;@�H;$�H; �H;G�H;��H;A�H;L�H;oI;�I;Y	I;$I;I;�I;�I;�I;xI;� I;�I;tI;�I;�I;�I;�I;s�H;      !I;!I;\!I;f!I;
!I;@ I;�I;nI;�I;�I;�I;�I;BI;�	I;�I;�I;� I;��H;J�H;��H;��H;��H;��H;1�H;��H;��H;X�H;O�H;��H;��H;/�H;��H;M�H;��H;��H;��H;��H;��H;��H;��H;M�H;��H;/�H;��H;��H;O�H;X�H;��H;��H;1�H;��H;��H;��H;��H;J�H;��H;� I;�I;�I;�	I;BI;�I;�I;�I;�I;nI;�I;@ I;
!I;f!I;\!I;!I;      �I;�I;I;5I;�I;aI;�I;xI;GI;�I;"I;�	I;�I;;I;�I;�H;��H;=�H;�H;4�H;p�H;��H;�H;��H;��H;j�H;[�H;��H;��H;�H;��H;C�H;��H;��H;g�H;J�H;:�H;J�H;g�H;��H;��H;C�H;��H;�H;��H;��H;[�H;j�H;��H;��H;�H;��H;p�H;4�H;�H;=�H;��H;�H;�I;;I;�I;�	I;"I;�I;GI;xI;�I;aI;�I;5I;I;�I;      I;�I;pI;�I;�I;TI;�I;I;/
I;&I;I;�I;�I;u�H;D�H;/�H;;�H;x�H;��H;��H;B�H;��H;��H;~�H;`�H;X�H;��H;��H;/�H;��H;'�H;��H;v�H;<�H;	�H;��H;��H;��H;	�H;<�H;v�H;��H;'�H;��H;/�H;��H;��H;X�H;`�H;~�H;��H;��H;B�H;��H;��H;x�H;;�H;/�H;D�H;u�H;�I;�I;I;&I;/
I;I;�I;TI;�I;�I;pI;�I;      �I;�I;BI;�
I;�	I;�I;|I;-I;�I;�I;@I;`�H;��H;��H;��H;T�H;��H;�H;x�H;�H;��H;��H;x�H;e�H;u�H;��H;��H;;�H;��H;C�H;��H;R�H;"�H;��H;��H;��H;��H;��H;��H;��H;"�H;R�H;��H;C�H;��H;;�H;��H;��H;u�H;e�H;x�H;��H;��H;�H;x�H;�H;��H;T�H;��H;��H;��H;`�H;@I;�I;�I;-I;|I;�I;�	I;�
I;BI;�I;      mI;GI;�I;qI;�I;�I;�I;�I;? I;��H;_�H;��H;s�H;�H;��H;�H;��H;�H;��H;��H;��H;��H;��H;��H;��H;&�H;d�H;��H;M�H;��H;v�H;"�H;��H;��H;��H;m�H;f�H;m�H;��H;��H;��H;"�H;v�H;��H;M�H;��H;d�H;&�H;��H;��H;��H;��H;��H;��H;��H;�H;��H;�H;��H;�H;s�H;��H;_�H;��H;? I;�I;�I;�I;�I;qI;�I;GI;      I;�I;�I;FI;� I;��H;�H;�H;�H;��H;��H;��H;5�H;��H;|�H;#�H;��H;��H;��H;��H;��H;��H;��H;�H;O�H;��H;��H;|�H;��H;��H;<�H;��H;��H;n�H;V�H;J�H;9�H;J�H;V�H;n�H;��H;��H;<�H;��H;��H;|�H;��H;��H;O�H;�H;��H;��H;��H;��H;��H;��H;��H;#�H;|�H;��H;5�H;��H;��H;��H;�H;�H;�H;��H;� I;FI;�I;�I;      q�H;e�H;!�H;��H;I�H;��H;��H;��H;�H;��H;��H;��H;o�H;^�H;?�H;�H;�H;��H;��H;��H;	�H;)�H;E�H;��H;��H;A�H;��H;9�H;��H;g�H;	�H;��H;��H;V�H;1�H;&�H;(�H;&�H;1�H;V�H;��H;��H;	�H;g�H;��H;9�H;��H;A�H;��H;��H;E�H;)�H;	�H;��H;��H;��H;�H;�H;?�H;^�H;o�H;��H;��H;��H;�H;��H;��H;��H;I�H;��H;!�H;e�H;      ��H;��H;x�H;"�H;��H;�H;c�H;��H;��H;��H;��H;��H;��H;��H;|�H;r�H;d�H;[�H;l�H;~�H;��H;��H;�H;]�H;��H;"�H;��H;
�H;��H;J�H;��H;��H;m�H;J�H;&�H;
�H;�H;
�H;&�H;J�H;m�H;��H;��H;J�H;��H;
�H;��H;"�H;��H;]�H;�H;��H;��H;~�H;l�H;[�H;d�H;r�H;|�H;��H;��H;��H;��H;��H;��H;��H;c�H;�H;��H;"�H;x�H;��H;      +�H;�H;��H;��H; �H;d�H;��H;�H;"�H;V�H;j�H;_�H;l�H;D�H;4�H;5�H;)�H;1�H;\�H;l�H;y�H;��H;��H;:�H;��H;�H;��H;�H;��H;:�H;��H;��H;f�H;9�H;(�H;�H;	�H;�H;(�H;9�H;f�H;��H;��H;:�H;��H;�H;��H;�H;��H;:�H;��H;��H;y�H;l�H;\�H;1�H;)�H;5�H;4�H;D�H;l�H;_�H;j�H;V�H;"�H;�H;��H;d�H; �H;��H;��H;�H;      ��H;��H;x�H;"�H;��H;�H;c�H;��H;��H;��H;��H;��H;��H;��H;|�H;r�H;d�H;[�H;l�H;~�H;��H;��H;�H;]�H;��H;"�H;��H;
�H;��H;J�H;��H;��H;m�H;J�H;&�H;
�H;�H;
�H;&�H;J�H;m�H;��H;��H;J�H;��H;
�H;��H;"�H;��H;]�H;�H;��H;��H;~�H;l�H;[�H;d�H;r�H;|�H;��H;��H;��H;��H;��H;��H;��H;c�H;�H;��H;"�H;x�H;��H;      q�H;e�H;!�H;��H;I�H;��H;��H;��H;�H;��H;��H;��H;o�H;^�H;?�H;�H;�H;��H;��H;��H;	�H;)�H;E�H;��H;��H;A�H;��H;9�H;��H;g�H;	�H;��H;��H;V�H;1�H;&�H;(�H;&�H;1�H;V�H;��H;��H;	�H;g�H;��H;9�H;��H;A�H;��H;��H;E�H;)�H;	�H;��H;��H;��H;�H;�H;?�H;^�H;o�H;��H;��H;��H;�H;��H;��H;��H;I�H;��H;!�H;e�H;      I;�I;�I;FI;� I;��H;�H;�H;�H;��H;��H;��H;5�H;��H;|�H;#�H;��H;��H;��H;��H;��H;��H;��H;�H;O�H;��H;��H;|�H;��H;��H;<�H;��H;��H;n�H;V�H;J�H;9�H;J�H;V�H;n�H;��H;��H;<�H;��H;��H;|�H;��H;��H;O�H;�H;��H;��H;��H;��H;��H;��H;��H;#�H;|�H;��H;5�H;��H;��H;��H;�H;�H;�H;��H;� I;FI;�I;�I;      mI;GI;�I;qI;�I;�I;�I;�I;? I;��H;_�H;��H;s�H;�H;��H;�H;��H;�H;��H;��H;��H;��H;��H;��H;��H;&�H;d�H;��H;M�H;��H;v�H;"�H;��H;��H;��H;m�H;f�H;m�H;��H;��H;��H;"�H;v�H;��H;M�H;��H;d�H;&�H;��H;��H;��H;��H;��H;��H;��H;�H;��H;�H;��H;�H;s�H;��H;_�H;��H;? I;�I;�I;�I;�I;qI;�I;GI;      �I;�I;BI;�
I;�	I;�I;|I;-I;�I;�I;@I;`�H;��H;��H;��H;T�H;��H;�H;x�H;�H;��H;��H;x�H;e�H;u�H;��H;��H;;�H;��H;C�H;��H;R�H;"�H;��H;��H;��H;��H;��H;��H;��H;"�H;R�H;��H;C�H;��H;;�H;��H;��H;u�H;e�H;x�H;��H;��H;�H;x�H;�H;��H;T�H;��H;��H;��H;`�H;@I;�I;�I;-I;|I;�I;�	I;�
I;BI;�I;      I;�I;pI;�I;�I;TI;�I;I;/
I;&I;I;�I;�I;u�H;D�H;/�H;;�H;x�H;��H;��H;B�H;��H;��H;~�H;`�H;X�H;��H;��H;/�H;��H;'�H;��H;v�H;<�H;	�H;��H;��H;��H;	�H;<�H;v�H;��H;'�H;��H;/�H;��H;��H;X�H;`�H;~�H;��H;��H;B�H;��H;��H;x�H;;�H;/�H;D�H;u�H;�I;�I;I;&I;/
I;I;�I;TI;�I;�I;pI;�I;      �I;�I;I;5I;�I;aI;�I;xI;GI;�I;"I;�	I;�I;;I;�I;�H;��H;=�H;�H;4�H;p�H;��H;�H;��H;��H;j�H;[�H;��H;��H;�H;��H;C�H;��H;��H;g�H;J�H;:�H;J�H;g�H;��H;��H;C�H;��H;�H;��H;��H;[�H;j�H;��H;��H;�H;��H;p�H;4�H;�H;=�H;��H;�H;�I;;I;�I;�	I;"I;�I;GI;xI;�I;aI;�I;5I;I;�I;      !I;!I;\!I;f!I;
!I;@ I;�I;nI;�I;�I;�I;�I;BI;�	I;�I;�I;� I;��H;J�H;��H;��H;��H;��H;1�H;��H;��H;X�H;O�H;��H;��H;/�H;��H;M�H;��H;��H;��H;��H;��H;��H;��H;M�H;��H;/�H;��H;��H;O�H;X�H;��H;��H;1�H;��H;��H;��H;��H;J�H;��H;� I;�I;�I;�	I;BI;�I;�I;�I;�I;nI;�I;@ I;
!I;f!I;\!I;!I;      �H;s�H;�I;�I;�I;�I;tI;�I;� I;xI;�I;�I;�I;I;$I;Y	I;�I;oI;L�H;A�H;��H;G�H; �H;$�H;@�H;��H;��H;k�H;O�H;��H;��H;;�H;��H;|�H;9�H;
�H;�H;
�H;9�H;|�H;��H;;�H;��H;��H;O�H;k�H;��H;��H;@�H;$�H; �H;G�H;��H;A�H;L�H;oI;�I;Y	I;$I;I;�I;�I;�I;xI;� I;�I;tI;�I;�I;�I;�I;s�H;      �MH;�SH;�cH;�|H;�H;o�H;��H;��H;�
I;7I; I;/ I;�I;OI;�I;8I;�I;�I;�I;� I;�H;�H;��H;Y�H;-�H;[�H;��H;��H;X�H;[�H;��H;��H;d�H;��H;��H;��H;��H;��H;��H;��H;d�H;��H;��H;[�H;X�H;��H;��H;[�H;-�H;Y�H;��H;�H;�H;� I;�I;�I;�I;8I;�I;OI;�I;/ I; I;7I;�
I;��H;��H;o�H;�H;�|H;�cH;�SH;      �HF;�XF;�F;�F;�&G;�G;��G;:BH;R�H;p�H;��H;I;
I;�I;I;I;�I; I;i	I;"I;VI;��H;��H;��H;w�H;S�H;[�H;��H;��H;j�H;X�H;��H;&�H;��H;A�H;"�H;�H;"�H;A�H;��H;&�H;��H;X�H;j�H;��H;��H;[�H;S�H;w�H;��H;��H;��H;VI;"I;i	I; I;�I;I;I;�I;
I;I;��H;p�H;R�H;:BH;��G;�G;�&G;�F;�F;�XF;      DA;(kA;��A;��B;�iC;o`D;�[E;IF;�G;��G;�MH;S�H;��H;�I;�I;zI;I;ZI;�I;�
I;I;�I;4�H;��H;��H;w�H;-�H;@�H;��H;��H;`�H;u�H;��H;O�H;��H;��H;��H;��H;��H;O�H;��H;u�H;`�H;��H;��H;@�H;-�H;w�H;��H;��H;4�H;�I;I;�
I;�I;ZI;I;zI;�I;�I;��H;S�H;�MH;��G;�G;IF;�[E;o`D;�iC;��B;��A;(kA;      �I6;'�6;ۖ7;�9;l;;1-=;li?;y�A;C�C;w1E;ۆF;t�G;�;H;��H;��H;�I;hI;9I;CI;XI;�I;�I;RI;E�H;��H;��H;Y�H;$�H;1�H;��H;~�H;e�H;��H;�H;��H;]�H;:�H;]�H;��H;�H;��H;e�H;~�H;��H;1�H;$�H;Y�H;��H;��H;E�H;RI;�I;�I;XI;CI;9I;hI;�I;��H;��H;�;H;t�G;ۆF;w1E;C�C;y�A;li?;1-=;l;;�9;ۖ7;'�6;      eo ;!;#;)&;%*;o.;�3;�7;��;;Ai?;jjB;8�D;�wF;�G;cH;,�H;�	I;�I;rI;�I;:I;6I;�I;RI;4�H;��H;��H; �H;��H;�H;��H;x�H;��H;��H;E�H;�H;��H;�H;E�H;��H;��H;x�H;��H;�H;��H; �H;��H;��H;4�H;RI;�I;6I;:I;�I;rI;�I;�	I;,�H;cH;�G;�wF;8�D;jjB;Ai?;��;;�7;�3;o.;%*;)&;#;!;      �r�:���:�j�:p�;��	;�;Wy;6O$;z�,;��3;5�9;2�>;>�B;D1E;*�F;vH;��H;��H;,I;I;CI;�I;6I;�I;�I;��H;�H;G�H;��H;��H;��H;��H;��H;��H;)�H;��H;��H;��H;)�H;��H;��H;��H;��H;��H;��H;G�H;�H;��H;�I;�I;6I;�I;CI;I;,I;��H;��H;vH;*�F;D1E;>�B;2�>;5�9;��3;z�,;6O$;Wy;�;��	;p�;�j�:���:      ��>:;�G:��b:ѳ�:���:3�:?)�:�h;p�;$a;:*;nq3;��:;� @;��C;�HF;ʾG;ԍH;.�H;zI;I;CI;:I;�I;I;VI;�H;��H;��H;p�H;B�H;��H;��H;��H;	�H;��H;y�H;��H;	�H;��H;��H;��H;B�H;p�H;��H;��H;�H;VI;I;�I;:I;CI;I;zI;.�H;ԍH;ʾG;�HF;��C;� @;��:;nq3;:*;$a;p�;�h;?)�:3�:���:ѳ�:��b:;�G:      ��������wk��� ��
���!69��!:Ǌ:�2�:D�:��;(;w�,;�6;��=;��B;��E;}�G;�{H;��H;zI;I;�I;XI;�
I;"I;� I;A�H;��H;4�H;��H;�H;��H;��H;��H;~�H;l�H;~�H;��H;��H;��H;�H;��H;4�H;��H;A�H;� I;"I;�
I;XI;�I;I;zI;��H;�{H;}�G;��E;��B;��=;�6;w�,;(;��;D�:�2�:Ǌ:��!:�!69�
���� ��wk����      �/��s�����x�k�X�b�/�ʻ �����u�r3�9��k:�:�m�:�A;!&;m3;�<;J�A;�oE;isG;�{H;.�H;,I;rI;CI;�I;i	I;�I;L�H;J�H;�H;��H;x�H;��H;��H;��H;l�H;\�H;l�H;��H;��H;��H;x�H;��H;�H;J�H;L�H;�I;i	I;�I;CI;rI;,I;.�H;�{H;isG;�oE;J�A;�<;m3;!&;�A;�m�:�:��k:r3�9u칉���ʻ �b�/�k�X���x�s���      ������q
�q�����׻S,��!����;�Rnۺ8� �J�9<Ǌ:���:� ;K!;Ģ0;>;;͒A;�oE;}�G;ԍH;��H;�I;9I;ZI; I;�I;oI;��H;=�H;x�H;�H;�H;��H;��H;[�H;1�H;[�H;��H;��H;�H;�H;x�H;=�H;��H;oI;�I; I;ZI;9I;�I;��H;ԍH;}�G;�oE;͒A;>;;Ģ0;K!;� ;���:<Ǌ:J�98� �Rnۺ�;�!���S,����׻q����q
���      ����8����^�k�ɆO�4/�VB�\�׻����@��Q�����,�>:j3�:�;�a;��/;>;;J�A;��E;ʾG;��H;�	I;hI;I;�I;�I;�I;� I;��H;;�H;��H;��H;��H;�H;d�H;)�H;d�H;�H;��H;��H;��H;;�H;��H;� I;�I;�I;�I;I;hI;�	I;��H;ʾG;��E;J�A;>;;��/;�a;�;j3�:,�>:����Q���@����\�׻VB�4/�ɆO�^�k���8��      F��	}�;�ݼ��˼"d��-��	�}�&�G������һ�������"/�n:�ճ:#�;�a;Ģ0;�<;��B;�HF;vH;,�H;�I;zI;I;8I;Y	I;�I;�H;/�H;T�H;�H;#�H;�H;r�H;5�H;r�H;�H;#�H;�H;T�H;/�H;�H;�I;Y	I;8I;I;zI;�I;,�H;vH;�HF;��B;�<;Ģ0;�a;#�;�ճ:n:�"/���������һ���&�G�	�}�-��"d����˼;�ݼ	}�      F�B�MR?��5���&��3��J��߮Ҽ/F����b=�I?�b.����/��qk����9�ճ:�;K!;m3;��=;��C;*�F;cH;��H;�I;I;�I;$I;�I;�I;D�H;��H;��H;|�H;?�H;|�H;4�H;|�H;?�H;|�H;��H;��H;D�H;�I;�I;$I;�I;I;�I;��H;cH;*�F;��C;��=;m3;K!;�;�ճ:���9�qk���/�b.��I?�b=���/F��߮Ҽ�J���3���&��5�MR?�      &��"W��撐�!�����j�Q`I���&����Oϼ�,���T[����I��;��qk�n:j3�:� ;!&;�6;� @;D1E;�G;��H;�I;�I;OI;I;�	I;;I;u�H;��H;�H;��H;^�H;��H;D�H;��H;^�H;��H;�H;��H;u�H;;I;�	I;I;OI;�I;�I;��H;�G;D1E;� @;�6;!&;� ;j3�:n:�qk�;��I�����T[��,��Oϼ�����&�Q`I���j�!���撐�"W��      �J���D��ͽ���$�������L�(��.��;��%�k����I����/��"/�,�>:���:�A;w�,;��:;>�B;�wF;�;H;��H;
I;�I;�I;BI;�I;�I;��H;s�H;5�H;o�H;��H;l�H;��H;o�H;5�H;s�H;��H;�I;�I;BI;�I;�I;
I;��H;�;H;�wF;>�B;��:;w�,;�A;���:,�>:�"/���/��I����%�k�;��.��(����L����$������ͽ�Dὼ��      K�:��*7���,�+�~�	�j��~���W����j�?�/��J���I��%�k���b.�������<Ǌ:�m�:(;nq3;2�>;8�D;t�G;S�H;I;/ I;�I;�I;�	I;�I;`�H;��H;��H;��H;��H;_�H;��H;��H;��H;��H;`�H;�I;�	I;�I;�I;/ I;I;S�H;t�G;8�D;2�>;nq3;(;�m�:<Ǌ:�����b.����%�k��I���J��?�/���j�W��~���j��~�	�+���,��*7�      ^���p��
��)�l���M���,�Tl�K9ݽ�A���{���5��J��;���T[�I?������Q��J�9�:��;:*;5�9;jjB;ۆF;�MH;��H; I;�I;�I;"I;I;@I;_�H;��H;��H;��H;j�H;��H;��H;��H;_�H;@I;I;"I;�I;�I; I;��H;�MH;ۆF;jjB;5�9;:*;��;�:J�9�Q������I?��T[�;���J����5��{��A��K9ݽTl���,���M�)�l�
���p��      +m־G�Ѿ�>ľ����̗����{���I�+����V���{�?�/�.���,��b=���һ�@�8� ���k:D�:$a;��3;Ai?;w1E;��G;p�H;7I;xI;�I;�I;&I;�I;��H;��H;��H;��H;V�H;��H;��H;��H;��H;�I;&I;�I;�I;xI;7I;p�H;��G;w1E;Ai?;��3;$a;D�:��k:8� ��@���һb=��,��.��?�/��{��V�����+���I���{�̗�������>ľG�Ѿ      =\����l5��z ��E۾�ճ��]��q�Z�F?#����A����j�(��Oϼ��������Rnۺr3�9�2�:p�;z�,;��;;C�C;�G;R�H;�
I;� I;�I;GI;/
I;�I;? I;�H;�H;��H;"�H;��H;�H;�H;? I;�I;/
I;GI;�I;� I;�
I;R�H;�G;C�C;��;;z�,;p�;�2�:r3�9Rnۺ��������Oϼ(����j��A�����F?#�q�Z��]���ճ��E۾�z �l5����      <�b��>]���M���6�����$���>ľq��q�Z�+�K9ݽW����L����/F��&�G�\�׻�;�u�Ǌ:�h;6O$;�7;y�A;IF;:BH;��H;�I;nI;xI;I;-I;�I;�H;��H;��H;�H;��H;��H;�H;�I;-I;I;xI;nI;�I;��H;:BH;IF;y�A;�7;6O$;�h;Ǌ:u칸;�\�׻&�G�/F�������L�W��K9ݽ+�q�Z�q���>ľ�$�������6���M��>]�      �o��벗����-�y�s�R���)�iv��>ľ�]����I�Tl�~��������&�߮Ҽ	�}�VB�!���������!:?)�:Wy;�3;li?;�[E;��G;��H;tI;�I;�I;�I;|I;�I;�H;��H;c�H;��H;c�H;��H;�H;�I;|I;�I;�I;�I;tI;��H;��G;�[E;li?;�3;Wy;?)�:��!:����!���VB�	�}�߮Ҽ��&����~���Tl���I��]���>ľiv���)�s�R�-�y����벗�      �˿�<ƿjL��:1��蟉��>]���)��$���ճ���{���,�j��$��Q`I��J��-��4/�S,��ʻ ��!693�:�;o.;1-=;o`D;�G;o�H;�I;@ I;aI;TI;�I;�I;��H;��H;�H;d�H;�H;��H;��H;�I;�I;TI;aI;@ I;�I;o�H;�G;o`D;1-=;o.;�;3�:�!69ʻ �S,��4/�-���J��Q`I�$��j�齞�,���{��ճ��$����)��>]�蟉�:1��jL���<ƿ      ����2���K[忭˿�T��蟉�s�R�����E۾̗����M�~�	������j��3�"d��ɆO���׻b�/��
�����:��	;%*;l;;�iC;�&G;�H;�I;
!I;�I;�I;�	I;�I;� I;I�H;��H; �H;��H;I�H;� I;�I;�	I;�I;�I;
!I;�I;�H;�&G;�iC;l;;%*;��	;���:�
��b�/���׻ɆO�"d���3���j����~�	���M�̗���E۾���s�R�蟉��T���˿K[�2���      O�0��o����˿:1��-�y���6��z �����)�l�+��ͽ!�����&���˼^�k�q���k�X��� �ѳ�:p�;)&;�9;��B;�F;�|H;�I;f!I;5I;�I;�
I;qI;FI;��H;"�H;��H;"�H;��H;FI;qI;�
I;�I;5I;f!I;�I;�|H;�F;��B;�9;)&;p�;ѳ�:�� �k�X�q���^�k���˼��&�!����ͽ+�)�l������z ���6�-�y�:1���˿���o�0��      ��*��g&��#�o�K[�jL�������M�l5��>ľ
����,��D�撐��5�;�ݼ���q
���x��wk���b:�j�:#;ۖ7;��A;�F;�cH;�I;\!I;I;pI;BI;�I;�I;!�H;x�H;��H;x�H;!�H;�I;�I;BI;pI;I;\!I;�I;�cH;�F;��A;ۖ7;#;�j�:��b:�wk���x��q
���;�ݼ�5�撐��Dὤ�,�
���>ľl5���M����jL��K[�o��#��g&�      ��8��4��g&�0��2����<ƿ벗��>]����G�Ѿ�p���*7����"W��MR?�	}�8����s������;�G:���:!;'�6;(kA;�XF;�SH;s�H;!I;�I;�I;�I;GI;�I;e�H;��H;�H;��H;e�H;�I;GI;�I;�I;�I;!I;s�H;�SH;�XF;(kA;'�6;!;���:;�G:���s�����8��	}�MR?�"W�����*7��p��G�Ѿ����>]�벗��<ƿ2���0���g&��4�      �Aq���i���U�A:�@�����6���q���uA�a5�� ��y^Z�����A���]�����d��|",�6��8�Ѻ���9)��:e�;eX4;p�@;�UF;��H;�FI;�aI;3NI;B9I;�(I;=I;�I;�I;�I;�
I;�I;�I;�I;=I;�(I;B9I;3NI;�aI;�FI;��H;�UF;p�@;eX4;e�;)��:���98�Ѻ6��|",��d������]��A�����y^Z�� ��a5�uA�q���6�������@�A:���U���i�      ��i���b�T�O�.5�-i������������q<�����e��[
V�FE	�!���IY�s9�Z����(�S����Ⱥ��:���:(�;L�4;i�@;kgF;��H;5HI;�aI;�MI;�8I;�(I;I;~I;�I;|I;x
I;|I;�I;~I;I;�(I;�8I;�MI;�aI;5HI;��H;kgF;i�@;L�4;(�;���:��:��ȺS���(�Z���s9��IY�!��FE	�[
V��e������q<������������-i�.5�T�O���b�      ��U�T�O�B-?�(�'���F�`欿Y�{�aa/���뾙���I����e���ZN�o5��Ǩ��nH�� ��󊮺�":��:��;��5;�_A;ښF;Z�H;<LI;aI;�LI;�7I;(I;aI;I;`I;&I;&
I;&I;`I;I;aI;(I;�7I;�LI;aI;<LI;Z�H;ښF;�_A;��5;��;��:�":󊮺� ��nH�Ǩ��o5���ZN�e������I�������aa/�Y�{��欿F����(�'�B-?�T�O�      A:�.5�(�'��������dȿ���e$_���Q�Ҿؕ��
�6�����*���`=�O���)��zG��6��@����Q:�:/";�7;�%B;�F;��H;RI;�_I;�JI;D6I;�&I;ZI;7I;�I;�
I;�	I;�
I;�I;7I;ZI;�&I;D6I;�JI;�_I;RI;��H;�F;�%B;�7;/";�:��Q:@���6��zG��)��O���`=��*�����
�6�ؕ��Q�Ҿ��e$_����dȿ�������(�'�.5�      @�-i�������B�ѿf�������q<��:��a����q����Wн齅���'�ib̼�zl�/���X�v��!�:��;�&;ڪ9;LC;wLG;�H;^XI;�]I;�GI;4I;�$I;I;(I;�I;�	I;�I;�	I;�I;(I;I;�$I;4I;�GI;�]I;^XI;�H;wLG;LC;ڪ9;�&;��;!�:v���X�/���zl�ib̼��'�齅��Wн����q��a���:��q<����f���B�ѿ������-i�      �������F��dȿf���������O���u]׾w���	�I�����A��C�d�v��֮�<RH�Kkλ�$�f5����:nM;̅+;�<;"3D;�G;�I;�]I;�ZI;	DI;I1I;�"I;aI;�I;�I;�I;�I;�I;�I;�I;aI;�"I;I1I;	DI;�ZI;�]I;�I;�G;"3D;�<;̅+;nM;���:f5��$�Kkλ<RH��֮�v�C�d��A�����	�I�w���u]׾����O�����f���dȿF�ῢ��      6��������欿��������O�}x����� ���l���"��ܽ���`=�Ý��l"��R���ۺV��9�=�:�K;��0;͞>;�LE;}"H;�$I;�`I;(VI;�?I;.I;a I;\I;"I;0
I;mI;�I;mI;0
I;"I;\I;a I;.I;�?I;(VI;�`I;�$I;}"H;�LE;͞>;��0;�K;�=�:V��9�ۺ�R��l"����Ý��`=����ܽ��"��l�� �����}x���O��������欿����      q�������Y�{�e$_��q<�������}��w���6�����!��!�h��������� d��.��f_e�QL[���Z:���:�+ ;��5;�A;�UF;̃H;@I;�aI;�PI;;I;e*I;�I;+I;WI;�I;I;MI;I;�I;WI;+I;�I;e*I;;I;�PI;�aI;@I;̃H;�UF;�A;��5;�+ ;���:��Z:QL[�f_e��.��� d��������!�h�!�������6�w���}��������q<�e$_�Y�{�����      uA��q<�aa/����:�u]׾� ��w��>�BE	�����ܽ����3�r�꼰���=",�X��2��AQ�ڮ�:�L
;�e);ބ:;E?C;?G;|�H;gSI;�^I;KJI;6I;t&I;�I;�I;ZI;�I;�I;�I;�I;�I;ZI;�I;�I;t&I;6I;KJI;�^I;gSI;|�H;?G;E?C;ބ:;�e);�L
;ڮ�:AQ�2��X��=",�����r�꼠�3�ܽ������BE	�>�w��� ��u]׾�:���aa/��q<�      a5�������Q�Ҿ�a��w����l��6�BE	���Ƚk���aG����z֮�C�W����9�k����X`,:���:�;��1;n�>;_E;M�G;CI;H^I;hYI;ZCI;�0I;V"I;cI;I;#	I;-I;�I;=I;�I;-I;#	I;I;cI;V"I;�0I;ZCI;hYI;H^I;CI;M�G;_E;n�>;��1;�;���:X`,:���9�k����C�W�z֮�����aG�k����ȽBE	��6��l�w����a��Q�Ҿ������      � ���e�����ؕ����q�	�I���"���������k���ZN�c�6¼}�y��$�PR��\� ���[��:H/;K�&;w8;��A;��F;��H;?I;aI;�QI;;<I;8+I;�I;I;vI;�I;XI;9I;� I;9I;XI;�I;vI;I;�I;8+I;;<I;�QI;aI;?I;��H;��F;��A;w8;K�&;H/;�:��[�\� �PR���$�}�y�6¼c��ZN�k������������"�	�I���q�ؕ������e��      y^Z�[
V��I�
�6�������ܽ!��ܽ���aG�c��ȼ�)����(����H5����1�Z:l�:8R;/&1;��=;ПD;P�G;�H;�WI;:]I;�HI;5I;�%I;�I;�I;�	I;�I;mI;|�H;��H;|�H;mI;�I;�	I;�I;�I;�%I;5I;�HI;:]I;�WI;�H;P�G;ПD;��=;/&1;8R;l�:1�Z:���H5������(��)���ȼc��aG�ܽ��!���ܽ�����
�6��I�[
V�      ���FE	��������Wн�A����!�h���3����6¼�)��ax/�u�һB�X�%����9���:�=;\e);�_9;�%B;ۉF;�|H;�5I;v`I;�TI;�?I;�-I; I;jI;DI;�I;jI;q�H;��H;�H;��H;q�H;jI;�I;DI;jI; I;�-I;�?I;�TI;v`I;�5I;�|H;ۉF;�%B;�_9;\e);�=;���:��9%��B�X�u�һax/��)��6¼�����3�!�h��󑽢A���Wн��콹��FE	�      �A��!��e���*��齅�C�d��`=����r��z֮�}�y���(�u�һi^e������f9���:Y�;n0";B�4;�l?;E;��G;��H;�VI;�]I;(JI;�6I;'I;�I;FI;�	I;>I;7 I;��H;��H;W�H;��H;��H;7 I;>I;�	I;FI;�I;'I;�6I;(JI;�]I;�VI;��H;��G;E;�l?;B�4;n0";Y�;���:�f9����i^e�u�һ��(�}�y�z֮�r�꼠���`=�C�d�齅��*��e��!��      �]��IY��ZN��`=���'�v�Ý���������C�W��$����B�X������9�ޚ:���:��;˷0;�<;w�C;HG;�H;�>I;P`I;�SI;^?I;2.I;z I;�I;.I;�I;�I;��H;��H;&�H;��H;&�H;��H;��H;�I;�I;.I;�I;z I;2.I;^?I;�SI;P`I;�>I;�H;HG;w�C;�<;˷0;��;���:�ޚ:�9����B�X�����$�C�W���������Ý�v���'��`=��ZN��IY�      ���s9�o5��O��ib̼�֮����� d�=",����PR��H5�%���f9�ޚ:��:6�;��-;��:;KB;`UF;;JH; I;�[I;G[I;�GI;%5I;<&I;7I;�I;9	I;^I;�H;��H;��H;n�H;�H;n�H;��H;��H;�H;^I;9	I;�I;7I;<&I;%5I;�GI;G[I;�[I; I;;JH;`UF;KB;��:;��-;6�;��:�ޚ:�f9%��H5�PR�����=",�� d�����֮�ib̼O��o5��s9�      �d��Z���Ǩ���)���zl�<RH�l"��.��X��9�k�\� ������9���:���:6�;�-;�9;j`A;۹E;J�G;��H;#RI;4_I;OI;�;I;�+I;�I;MI;*I;�I;p I;��H;��H;��H;��H;|�H;��H;��H;��H;��H;p I;�I;*I;MI;�I;�+I;�;I;OI;4_I;#RI;��H;J�G;۹E;j`A;�9;�-;6�;���:���:��9���\� �9�k�X���.��l"�<RH��zl��)��Ǩ��Z���      |",��(�nH�zG�/��Kkλ�R��f_e�2�������[�1�Z:���:Y�;��;��-;�9;�A;�bE;E�G;��H;tFI;`I;�TI;bAI;�0I;#I;�I;I;�I;I;��H;b�H;��H;!�H;,�H;��H;,�H;!�H;��H;b�H;��H;I;�I;I;�I;#I;�0I;bAI;�TI;`I;tFI;��H;E�G;�bE;�A;�9;��-;��;Y�;���:1�Z:��[����2��f_e��R��Kkλ/��zG�nH��(�      6��S��� ���6���X��$��ۺQL[�AQ�X`,:�:l�:�=;n0";˷0;��:;j`A;�bE;�G;��H;�<I;N_I;�XI;FI;5I;�&I;I;�I;
I;�I;��H;�H;6�H;�H;��H;��H;S�H;��H;��H;�H;6�H;�H;��H;�I;
I;�I;I;�&I;5I;FI;�XI;N_I;�<I;��H;�G;�bE;j`A;��:;˷0;n0";�=;l�:�:X`,:AQ�QL[��ۺ�$��X��6��� ��S��      8�Ѻ��Ⱥ󊮺@��v��f5�V��9��Z:ڮ�:���:H/;8R;\e);B�4;�<;KB;۹E;E�G;��H;�9I;q^I;�ZI;?II;8I;�)I;�I;I;I;vI;$ I;��H;��H;&�H;C�H;�H;F�H;��H;F�H;�H;C�H;&�H;��H;��H;$ I;vI;I;I;�I;�)I;8I;?II;�ZI;q^I;�9I;��H;E�G;۹E;KB;�<;B�4;\e);8R;H/;���:ڮ�:��Z:V��9f5�v��@��󊮺��Ⱥ      ���9��:�":��Q:!�:���:�=�:���:�L
;�;K�&;/&1;�_9;�l?;w�C;`UF;J�G;��H;�<I;q^I;1[I;�JI;2:I;�+I;�I;I;�I;�I;`I;��H;L�H;��H;K�H;��H;��H;��H;��H;��H;��H;��H;K�H;��H;L�H;��H;`I;�I;�I;I;�I;�+I;2:I;�JI;1[I;q^I;�<I;��H;J�G;`UF;w�C;�l?;�_9;/&1;K�&;�;�L
;���:�=�:���:!�:��Q:�":��:      )��:���:��:�:��;nM;�K;�+ ;�e);��1;w8;��=;�%B;E;HG;;JH;��H;tFI;N_I;�ZI;�JI;�:I;-I;H!I;QI;+I;1I;xI;��H;��H;��H;}�H;��H;.�H;R�H;��H;z�H;��H;R�H;.�H;��H;}�H;��H;��H;��H;xI;1I;+I;QI;H!I;-I;�:I;�JI;�ZI;N_I;tFI;��H;;JH;HG;E;�%B;��=;w8;��1;�e);�+ ;�K;nM;��;�:��:���:      e�;(�;��;/";�&;̅+;��0;��5;ބ:;n�>;��A;ПD;ۉF;��G;�H; I;#RI;`I;�XI;?II;2:I;-I;�!I;I;�I;	I;BI;^�H;��H;k�H;��H;��H;�H;��H; �H;��H;p�H;��H; �H;��H;�H;��H;��H;k�H;��H;^�H;BI;	I;�I;I;�!I;-I;2:I;?II;�XI;`I;#RI; I;�H;��G;ۉF;ПD;��A;n�>;ބ:;��5;��0;̅+;�&;/";��;(�;      eX4;L�4;��5;�7;ڪ9;�<;͞>;�A;E?C;_E;��F;P�G;�|H;��H;�>I;�[I;4_I;�TI;FI;8I;�+I;H!I;I;9I;v	I;�I; �H;��H;��H;��H;��H;�H;��H;��H;��H;��H;u�H;��H;��H;��H;��H;�H;��H;��H;��H;��H; �H;�I;v	I;9I;I;H!I;�+I;8I;FI;�TI;4_I;�[I;�>I;��H;�|H;P�G;��F;_E;E?C;�A;͞>;�<;ڪ9;�7;��5;L�4;      p�@;i�@;�_A;�%B;LC;"3D;�LE;�UF;?G;M�G;��H;�H;�5I;�VI;P`I;G[I;OI;bAI;5I;�)I;�I;QI;�I;v	I;I;.�H;D�H;��H;0�H;��H;�H;��H;[�H;��H;��H;��H;r�H;��H;��H;��H;[�H;��H;�H;��H;0�H;��H;D�H;.�H;I;v	I;�I;QI;�I;�)I;5I;bAI;OI;G[I;P`I;�VI;�5I;�H;��H;M�G;?G;�UF;�LE;"3D;LC;�%B;�_A;i�@;      �UF;kgF;ښF;�F;wLG;�G;}"H;̃H;|�H;CI;?I;�WI;v`I;�]I;�SI;�GI;�;I;�0I;�&I;�I;I;+I;	I;�I;.�H;W�H;'�H;j�H;��H;�H;��H;V�H;M�H;��H;�H;��H;��H;��H;�H;��H;M�H;V�H;��H;�H;��H;j�H;'�H;W�H;.�H;�I;	I;+I;I;�I;�&I;�0I;�;I;�GI;�SI;�]I;v`I;�WI;?I;CI;|�H;̃H;}"H;�G;wLG;�F;ښF;kgF;      ��H;��H;Z�H;��H;�H;�I;�$I;@I;gSI;H^I;aI;:]I;�TI;(JI;^?I;%5I;�+I;#I;I;I;�I;1I;BI; �H;D�H;'�H;\�H;�H;7�H;|�H;7�H;�H;F�H;��H;@�H;��H;��H;��H;@�H;��H;F�H;�H;7�H;|�H;7�H;�H;\�H;'�H;D�H; �H;BI;1I;�I;I;I;#I;�+I;%5I;^?I;(JI;�TI;:]I;aI;H^I;gSI;@I;�$I;�I;�H;��H;Z�H;��H;      �FI;5HI;<LI;RI;^XI;�]I;�`I;�aI;�^I;hYI;�QI;�HI;�?I;�6I;2.I;<&I;�I;�I;�I;I;�I;xI;^�H;��H;��H;j�H;�H;�H;��H;3�H;�H;�H;p�H;��H;|�H;F�H;@�H;F�H;|�H;��H;p�H;�H;�H;3�H;��H;�H;�H;j�H;��H;��H;^�H;xI;�I;I;�I;�I;�I;<&I;2.I;�6I;�?I;�HI;�QI;hYI;�^I;�aI;�`I;�]I;^XI;RI;<LI;5HI;      �aI;�aI;aI;�_I;�]I;�ZI;(VI;�PI;KJI;ZCI;;<I;5I;�-I;'I;z I;7I;MI;I;
I;vI;`I;��H;��H;��H;0�H;��H;7�H;��H;*�H;�H;�H;B�H;��H;2�H;��H;��H;��H;��H;��H;2�H;��H;B�H;�H;�H;*�H;��H;7�H;��H;0�H;��H;��H;��H;`I;vI;
I;I;MI;7I;z I;'I;�-I;5I;;<I;ZCI;KJI;�PI;(VI;�ZI;�]I;�_I;aI;�aI;      3NI;�MI;�LI;�JI;�GI;	DI;�?I;;I;6I;�0I;8+I;�%I; I;�I;�I;�I;*I;�I;�I;$ I;��H;��H;k�H;��H;��H;�H;|�H;3�H;�H;	�H;1�H;��H;��H;��H;H�H;(�H;%�H;(�H;H�H;��H;��H;��H;1�H;	�H;�H;3�H;|�H;�H;��H;��H;k�H;��H;��H;$ I;�I;�I;*I;�I;�I;�I; I;�%I;8+I;�0I;6I;;I;�?I;	DI;�GI;�JI;�LI;�MI;      B9I;�8I;�7I;D6I;4I;I1I;.I;e*I;t&I;V"I;�I;�I;jI;FI;.I;9	I;�I;I;��H;��H;L�H;��H;��H;��H;�H;��H;7�H;�H;�H;1�H;��H;��H;d�H;�H;��H;��H;��H;��H;��H;�H;d�H;��H;��H;1�H;�H;�H;7�H;��H;�H;��H;��H;��H;L�H;��H;��H;I;�I;9	I;.I;FI;jI;�I;�I;V"I;t&I;e*I;.I;I1I;4I;D6I;�7I;�8I;      �(I;�(I;(I;�&I;�$I;�"I;a I;�I;�I;cI;I;�I;DI;�	I;�I;^I;p I;��H;�H;��H;��H;}�H;��H;�H;��H;V�H;�H;�H;B�H;��H;��H;{�H;��H;��H;z�H;U�H;>�H;U�H;z�H;��H;��H;{�H;��H;��H;B�H;�H;�H;V�H;��H;�H;��H;}�H;��H;��H;�H;��H;p I;^I;�I;�	I;DI;�I;I;cI;�I;�I;a I;�"I;�$I;�&I;(I;�(I;      =I;I;aI;ZI;I;aI;\I;+I;�I;I;vI;�	I;�I;>I;�I;�H;��H;b�H;6�H;&�H;K�H;��H;�H;��H;[�H;M�H;F�H;p�H;��H;��H;d�H;��H;��H;\�H;�H;	�H;�H;	�H;�H;\�H;��H;��H;d�H;��H;��H;p�H;F�H;M�H;[�H;��H;�H;��H;K�H;&�H;6�H;b�H;��H;�H;�I;>I;�I;�	I;vI;I;�I;+I;\I;aI;I;ZI;aI;I;      �I;~I;I;7I;(I;�I;"I;WI;ZI;#	I;�I;�I;jI;7 I;��H;��H;��H;��H;�H;C�H;��H;.�H;��H;��H;��H;��H;��H;��H;2�H;��H;�H;��H;\�H; �H;��H;��H;��H;��H;��H; �H;\�H;��H;�H;��H;2�H;��H;��H;��H;��H;��H;��H;.�H;��H;C�H;�H;��H;��H;��H;��H;7 I;jI;�I;�I;#	I;ZI;WI;"I;�I;(I;7I;I;~I;      �I;�I;`I;�I;�I;�I;0
I;�I;�I;-I;XI;mI;q�H;��H;��H;��H;��H;!�H;��H;�H;��H;R�H; �H;��H;��H;�H;@�H;|�H;��H;H�H;��H;z�H;�H;��H;��H;��H;��H;��H;��H;��H;�H;z�H;��H;H�H;��H;|�H;@�H;�H;��H;��H; �H;R�H;��H;�H;��H;!�H;��H;��H;��H;��H;q�H;mI;XI;-I;�I;�I;0
I;�I;�I;�I;`I;�I;      �I;|I;&I;�
I;�	I;�I;mI;I;�I;�I;9I;|�H;��H;��H;&�H;n�H;��H;,�H;��H;F�H;��H;��H;��H;��H;��H;��H;��H;F�H;��H;(�H;��H;U�H;	�H;��H;��H;��H;}�H;��H;��H;��H;	�H;U�H;��H;(�H;��H;F�H;��H;��H;��H;��H;��H;��H;��H;F�H;��H;,�H;��H;n�H;&�H;��H;��H;|�H;9I;�I;�I;I;mI;�I;�	I;�
I;&I;|I;      �
I;x
I;&
I;�	I;�I;�I;�I;MI;�I;=I;� I;��H;�H;W�H;��H;�H;|�H;��H;S�H;��H;��H;z�H;p�H;u�H;r�H;��H;��H;@�H;��H;%�H;��H;>�H;�H;��H;��H;}�H;��H;}�H;��H;��H;�H;>�H;��H;%�H;��H;@�H;��H;��H;r�H;u�H;p�H;z�H;��H;��H;S�H;��H;|�H;�H;��H;W�H;�H;��H;� I;=I;�I;MI;�I;�I;�I;�	I;&
I;x
I;      �I;|I;&I;�
I;�	I;�I;mI;I;�I;�I;9I;|�H;��H;��H;&�H;n�H;��H;,�H;��H;F�H;��H;��H;��H;��H;��H;��H;��H;F�H;��H;(�H;��H;U�H;	�H;��H;��H;��H;}�H;��H;��H;��H;	�H;U�H;��H;(�H;��H;F�H;��H;��H;��H;��H;��H;��H;��H;F�H;��H;,�H;��H;n�H;&�H;��H;��H;|�H;9I;�I;�I;I;mI;�I;�	I;�
I;&I;|I;      �I;�I;`I;�I;�I;�I;0
I;�I;�I;-I;XI;mI;q�H;��H;��H;��H;��H;!�H;��H;�H;��H;R�H; �H;��H;��H;�H;@�H;|�H;��H;H�H;��H;z�H;�H;��H;��H;��H;��H;��H;��H;��H;�H;z�H;��H;H�H;��H;|�H;@�H;�H;��H;��H; �H;R�H;��H;�H;��H;!�H;��H;��H;��H;��H;q�H;mI;XI;-I;�I;�I;0
I;�I;�I;�I;`I;�I;      �I;~I;I;7I;(I;�I;"I;WI;ZI;#	I;�I;�I;jI;7 I;��H;��H;��H;��H;�H;C�H;��H;.�H;��H;��H;��H;��H;��H;��H;2�H;��H;�H;��H;\�H; �H;��H;��H;��H;��H;��H; �H;\�H;��H;�H;��H;2�H;��H;��H;��H;��H;��H;��H;.�H;��H;C�H;�H;��H;��H;��H;��H;7 I;jI;�I;�I;#	I;ZI;WI;"I;�I;(I;7I;I;~I;      =I;I;aI;ZI;I;aI;\I;+I;�I;I;vI;�	I;�I;>I;�I;�H;��H;b�H;6�H;&�H;K�H;��H;�H;��H;[�H;M�H;F�H;p�H;��H;��H;d�H;��H;��H;\�H;�H;	�H;�H;	�H;�H;\�H;��H;��H;d�H;��H;��H;p�H;F�H;M�H;[�H;��H;�H;��H;K�H;&�H;6�H;b�H;��H;�H;�I;>I;�I;�	I;vI;I;�I;+I;\I;aI;I;ZI;aI;I;      �(I;�(I;(I;�&I;�$I;�"I;a I;�I;�I;cI;I;�I;DI;�	I;�I;^I;p I;��H;�H;��H;��H;}�H;��H;�H;��H;V�H;�H;�H;B�H;��H;��H;{�H;��H;��H;z�H;U�H;>�H;U�H;z�H;��H;��H;{�H;��H;��H;B�H;�H;�H;V�H;��H;�H;��H;}�H;��H;��H;�H;��H;p I;^I;�I;�	I;DI;�I;I;cI;�I;�I;a I;�"I;�$I;�&I;(I;�(I;      B9I;�8I;�7I;D6I;4I;I1I;.I;e*I;t&I;V"I;�I;�I;jI;FI;.I;9	I;�I;I;��H;��H;L�H;��H;��H;��H;�H;��H;7�H;�H;�H;1�H;��H;��H;d�H;�H;��H;��H;��H;��H;��H;�H;d�H;��H;��H;1�H;�H;�H;7�H;��H;�H;��H;��H;��H;L�H;��H;��H;I;�I;9	I;.I;FI;jI;�I;�I;V"I;t&I;e*I;.I;I1I;4I;D6I;�7I;�8I;      3NI;�MI;�LI;�JI;�GI;	DI;�?I;;I;6I;�0I;8+I;�%I; I;�I;�I;�I;*I;�I;�I;$ I;��H;��H;k�H;��H;��H;�H;|�H;3�H;�H;	�H;1�H;��H;��H;��H;H�H;(�H;%�H;(�H;H�H;��H;��H;��H;1�H;	�H;�H;3�H;|�H;�H;��H;��H;k�H;��H;��H;$ I;�I;�I;*I;�I;�I;�I; I;�%I;8+I;�0I;6I;;I;�?I;	DI;�GI;�JI;�LI;�MI;      �aI;�aI;aI;�_I;�]I;�ZI;(VI;�PI;KJI;ZCI;;<I;5I;�-I;'I;z I;7I;MI;I;
I;vI;`I;��H;��H;��H;0�H;��H;7�H;��H;*�H;�H;�H;B�H;��H;2�H;��H;��H;��H;��H;��H;2�H;��H;B�H;�H;�H;*�H;��H;7�H;��H;0�H;��H;��H;��H;`I;vI;
I;I;MI;7I;z I;'I;�-I;5I;;<I;ZCI;KJI;�PI;(VI;�ZI;�]I;�_I;aI;�aI;      �FI;5HI;<LI;RI;^XI;�]I;�`I;�aI;�^I;hYI;�QI;�HI;�?I;�6I;2.I;<&I;�I;�I;�I;I;�I;xI;^�H;��H;��H;j�H;�H;�H;��H;3�H;�H;�H;p�H;��H;|�H;F�H;@�H;F�H;|�H;��H;p�H;�H;�H;3�H;��H;�H;�H;j�H;��H;��H;^�H;xI;�I;I;�I;�I;�I;<&I;2.I;�6I;�?I;�HI;�QI;hYI;�^I;�aI;�`I;�]I;^XI;RI;<LI;5HI;      ��H;��H;Z�H;��H;�H;�I;�$I;@I;gSI;H^I;aI;:]I;�TI;(JI;^?I;%5I;�+I;#I;I;I;�I;1I;BI; �H;D�H;'�H;\�H;�H;7�H;|�H;7�H;�H;F�H;��H;@�H;��H;��H;��H;@�H;��H;F�H;�H;7�H;|�H;7�H;�H;\�H;'�H;D�H; �H;BI;1I;�I;I;I;#I;�+I;%5I;^?I;(JI;�TI;:]I;aI;H^I;gSI;@I;�$I;�I;�H;��H;Z�H;��H;      �UF;kgF;ښF;�F;wLG;�G;}"H;̃H;|�H;CI;?I;�WI;v`I;�]I;�SI;�GI;�;I;�0I;�&I;�I;I;+I;	I;�I;.�H;W�H;'�H;j�H;��H;�H;��H;V�H;M�H;��H;�H;��H;��H;��H;�H;��H;M�H;V�H;��H;�H;��H;j�H;'�H;W�H;.�H;�I;	I;+I;I;�I;�&I;�0I;�;I;�GI;�SI;�]I;v`I;�WI;?I;CI;|�H;̃H;}"H;�G;wLG;�F;ښF;kgF;      p�@;i�@;�_A;�%B;LC;"3D;�LE;�UF;?G;M�G;��H;�H;�5I;�VI;P`I;G[I;OI;bAI;5I;�)I;�I;QI;�I;v	I;I;.�H;D�H;��H;0�H;��H;�H;��H;[�H;��H;��H;��H;r�H;��H;��H;��H;[�H;��H;�H;��H;0�H;��H;D�H;.�H;I;v	I;�I;QI;�I;�)I;5I;bAI;OI;G[I;P`I;�VI;�5I;�H;��H;M�G;?G;�UF;�LE;"3D;LC;�%B;�_A;i�@;      eX4;L�4;��5;�7;ڪ9;�<;͞>;�A;E?C;_E;��F;P�G;�|H;��H;�>I;�[I;4_I;�TI;FI;8I;�+I;H!I;I;9I;v	I;�I; �H;��H;��H;��H;��H;�H;��H;��H;��H;��H;u�H;��H;��H;��H;��H;�H;��H;��H;��H;��H; �H;�I;v	I;9I;I;H!I;�+I;8I;FI;�TI;4_I;�[I;�>I;��H;�|H;P�G;��F;_E;E?C;�A;͞>;�<;ڪ9;�7;��5;L�4;      e�;(�;��;/";�&;̅+;��0;��5;ބ:;n�>;��A;ПD;ۉF;��G;�H; I;#RI;`I;�XI;?II;2:I;-I;�!I;I;�I;	I;BI;^�H;��H;k�H;��H;��H;�H;��H; �H;��H;p�H;��H; �H;��H;�H;��H;��H;k�H;��H;^�H;BI;	I;�I;I;�!I;-I;2:I;?II;�XI;`I;#RI; I;�H;��G;ۉF;ПD;��A;n�>;ބ:;��5;��0;̅+;�&;/";��;(�;      )��:���:��:�:��;nM;�K;�+ ;�e);��1;w8;��=;�%B;E;HG;;JH;��H;tFI;N_I;�ZI;�JI;�:I;-I;H!I;QI;+I;1I;xI;��H;��H;��H;}�H;��H;.�H;R�H;��H;z�H;��H;R�H;.�H;��H;}�H;��H;��H;��H;xI;1I;+I;QI;H!I;-I;�:I;�JI;�ZI;N_I;tFI;��H;;JH;HG;E;�%B;��=;w8;��1;�e);�+ ;�K;nM;��;�:��:���:      ���9��:�":��Q:!�:���:�=�:���:�L
;�;K�&;/&1;�_9;�l?;w�C;`UF;J�G;��H;�<I;q^I;1[I;�JI;2:I;�+I;�I;I;�I;�I;`I;��H;L�H;��H;K�H;��H;��H;��H;��H;��H;��H;��H;K�H;��H;L�H;��H;`I;�I;�I;I;�I;�+I;2:I;�JI;1[I;q^I;�<I;��H;J�G;`UF;w�C;�l?;�_9;/&1;K�&;�;�L
;���:�=�:���:!�:��Q:�":��:      8�Ѻ��Ⱥ󊮺@��v��f5�V��9��Z:ڮ�:���:H/;8R;\e);B�4;�<;KB;۹E;E�G;��H;�9I;q^I;�ZI;?II;8I;�)I;�I;I;I;vI;$ I;��H;��H;&�H;C�H;�H;F�H;��H;F�H;�H;C�H;&�H;��H;��H;$ I;vI;I;I;�I;�)I;8I;?II;�ZI;q^I;�9I;��H;E�G;۹E;KB;�<;B�4;\e);8R;H/;���:ڮ�:��Z:V��9f5�v��@��󊮺��Ⱥ      6��S��� ���6���X��$��ۺQL[�AQ�X`,:�:l�:�=;n0";˷0;��:;j`A;�bE;�G;��H;�<I;N_I;�XI;FI;5I;�&I;I;�I;
I;�I;��H;�H;6�H;�H;��H;��H;S�H;��H;��H;�H;6�H;�H;��H;�I;
I;�I;I;�&I;5I;FI;�XI;N_I;�<I;��H;�G;�bE;j`A;��:;˷0;n0";�=;l�:�:X`,:AQ�QL[��ۺ�$��X��6��� ��S��      |",��(�nH�zG�/��Kkλ�R��f_e�2�������[�1�Z:���:Y�;��;��-;�9;�A;�bE;E�G;��H;tFI;`I;�TI;bAI;�0I;#I;�I;I;�I;I;��H;b�H;��H;!�H;,�H;��H;,�H;!�H;��H;b�H;��H;I;�I;I;�I;#I;�0I;bAI;�TI;`I;tFI;��H;E�G;�bE;�A;�9;��-;��;Y�;���:1�Z:��[����2��f_e��R��Kkλ/��zG�nH��(�      �d��Z���Ǩ���)���zl�<RH�l"��.��X��9�k�\� ������9���:���:6�;�-;�9;j`A;۹E;J�G;��H;#RI;4_I;OI;�;I;�+I;�I;MI;*I;�I;p I;��H;��H;��H;��H;|�H;��H;��H;��H;��H;p I;�I;*I;MI;�I;�+I;�;I;OI;4_I;#RI;��H;J�G;۹E;j`A;�9;�-;6�;���:���:��9���\� �9�k�X���.��l"�<RH��zl��)��Ǩ��Z���      ���s9�o5��O��ib̼�֮����� d�=",����PR��H5�%���f9�ޚ:��:6�;��-;��:;KB;`UF;;JH; I;�[I;G[I;�GI;%5I;<&I;7I;�I;9	I;^I;�H;��H;��H;n�H;�H;n�H;��H;��H;�H;^I;9	I;�I;7I;<&I;%5I;�GI;G[I;�[I; I;;JH;`UF;KB;��:;��-;6�;��:�ޚ:�f9%��H5�PR�����=",�� d�����֮�ib̼O��o5��s9�      �]��IY��ZN��`=���'�v�Ý���������C�W��$����B�X������9�ޚ:���:��;˷0;�<;w�C;HG;�H;�>I;P`I;�SI;^?I;2.I;z I;�I;.I;�I;�I;��H;��H;&�H;��H;&�H;��H;��H;�I;�I;.I;�I;z I;2.I;^?I;�SI;P`I;�>I;�H;HG;w�C;�<;˷0;��;���:�ޚ:�9����B�X�����$�C�W���������Ý�v���'��`=��ZN��IY�      �A��!��e���*��齅�C�d��`=����r��z֮�}�y���(�u�һi^e������f9���:Y�;n0";B�4;�l?;E;��G;��H;�VI;�]I;(JI;�6I;'I;�I;FI;�	I;>I;7 I;��H;��H;W�H;��H;��H;7 I;>I;�	I;FI;�I;'I;�6I;(JI;�]I;�VI;��H;��G;E;�l?;B�4;n0";Y�;���:�f9����i^e�u�һ��(�}�y�z֮�r�꼠���`=�C�d�齅��*��e��!��      ���FE	��������Wн�A����!�h���3����6¼�)��ax/�u�һB�X�%����9���:�=;\e);�_9;�%B;ۉF;�|H;�5I;v`I;�TI;�?I;�-I; I;jI;DI;�I;jI;q�H;��H;�H;��H;q�H;jI;�I;DI;jI; I;�-I;�?I;�TI;v`I;�5I;�|H;ۉF;�%B;�_9;\e);�=;���:��9%��B�X�u�һax/��)��6¼�����3�!�h��󑽢A���Wн��콹��FE	�      y^Z�[
V��I�
�6�������ܽ!��ܽ���aG�c��ȼ�)����(����H5����1�Z:l�:8R;/&1;��=;ПD;P�G;�H;�WI;:]I;�HI;5I;�%I;�I;�I;�	I;�I;mI;|�H;��H;|�H;mI;�I;�	I;�I;�I;�%I;5I;�HI;:]I;�WI;�H;P�G;ПD;��=;/&1;8R;l�:1�Z:���H5������(��)���ȼc��aG�ܽ��!���ܽ�����
�6��I�[
V�      � ���e�����ؕ����q�	�I���"���������k���ZN�c�6¼}�y��$�PR��\� ���[��:H/;K�&;w8;��A;��F;��H;?I;aI;�QI;;<I;8+I;�I;I;vI;�I;XI;9I;� I;9I;XI;�I;vI;I;�I;8+I;;<I;�QI;aI;?I;��H;��F;��A;w8;K�&;H/;�:��[�\� �PR���$�}�y�6¼c��ZN�k������������"�	�I���q�ؕ������e��      a5�������Q�Ҿ�a��w����l��6�BE	���Ƚk���aG����z֮�C�W����9�k����X`,:���:�;��1;n�>;_E;M�G;CI;H^I;hYI;ZCI;�0I;V"I;cI;I;#	I;-I;�I;=I;�I;-I;#	I;I;cI;V"I;�0I;ZCI;hYI;H^I;CI;M�G;_E;n�>;��1;�;���:X`,:���9�k����C�W�z֮�����aG�k����ȽBE	��6��l�w����a��Q�Ҿ������      uA��q<�aa/����:�u]׾� ��w��>�BE	�����ܽ����3�r�꼰���=",�X��2��AQ�ڮ�:�L
;�e);ބ:;E?C;?G;|�H;gSI;�^I;KJI;6I;t&I;�I;�I;ZI;�I;�I;�I;�I;�I;ZI;�I;�I;t&I;6I;KJI;�^I;gSI;|�H;?G;E?C;ބ:;�e);�L
;ڮ�:AQ�2��X��=",�����r�꼠�3�ܽ������BE	�>�w��� ��u]׾�:���aa/��q<�      q�������Y�{�e$_��q<�������}��w���6�����!��!�h��������� d��.��f_e�QL[���Z:���:�+ ;��5;�A;�UF;̃H;@I;�aI;�PI;;I;e*I;�I;+I;WI;�I;I;MI;I;�I;WI;+I;�I;e*I;;I;�PI;�aI;@I;̃H;�UF;�A;��5;�+ ;���:��Z:QL[�f_e��.��� d��������!�h�!�������6�w���}��������q<�e$_�Y�{�����      6��������欿��������O�}x����� ���l���"��ܽ���`=�Ý��l"��R���ۺV��9�=�:�K;��0;͞>;�LE;}"H;�$I;�`I;(VI;�?I;.I;a I;\I;"I;0
I;mI;�I;mI;0
I;"I;\I;a I;.I;�?I;(VI;�`I;�$I;}"H;�LE;͞>;��0;�K;�=�:V��9�ۺ�R��l"����Ý��`=����ܽ��"��l�� �����}x���O��������欿����      �������F��dȿf���������O���u]׾w���	�I�����A��C�d�v��֮�<RH�Kkλ�$�f5����:nM;̅+;�<;"3D;�G;�I;�]I;�ZI;	DI;I1I;�"I;aI;�I;�I;�I;�I;�I;�I;�I;aI;�"I;I1I;	DI;�ZI;�]I;�I;�G;"3D;�<;̅+;nM;���:f5��$�Kkλ<RH��֮�v�C�d��A�����	�I�w���u]׾����O�����f���dȿF�ῢ��      @�-i�������B�ѿf�������q<��:��a����q����Wн齅���'�ib̼�zl�/���X�v��!�:��;�&;ڪ9;LC;wLG;�H;^XI;�]I;�GI;4I;�$I;I;(I;�I;�	I;�I;�	I;�I;(I;I;�$I;4I;�GI;�]I;^XI;�H;wLG;LC;ڪ9;�&;��;!�:v���X�/���zl�ib̼��'�齅��Wн����q��a���:��q<����f���B�ѿ������-i�      A:�.5�(�'��������dȿ���e$_���Q�Ҿؕ��
�6�����*���`=�O���)��zG��6��@����Q:�:/";�7;�%B;�F;��H;RI;�_I;�JI;D6I;�&I;ZI;7I;�I;�
I;�	I;�
I;�I;7I;ZI;�&I;D6I;�JI;�_I;RI;��H;�F;�%B;�7;/";�:��Q:@���6��zG��)��O���`=��*�����
�6�ؕ��Q�Ҿ��e$_����dȿ�������(�'�.5�      ��U�T�O�B-?�(�'���F�`欿Y�{�aa/���뾙���I����e���ZN�o5��Ǩ��nH�� ��󊮺�":��:��;��5;�_A;ښF;Z�H;<LI;aI;�LI;�7I;(I;aI;I;`I;&I;&
I;&I;`I;I;aI;(I;�7I;�LI;aI;<LI;Z�H;ښF;�_A;��5;��;��:�":󊮺� ��nH�Ǩ��o5���ZN�e������I�������aa/�Y�{��欿F����(�'�B-?�T�O�      ��i���b�T�O�.5�-i������������q<�����e��[
V�FE	�!���IY�s9�Z����(�S����Ⱥ��:���:(�;L�4;i�@;kgF;��H;5HI;�aI;�MI;�8I;�(I;I;~I;�I;|I;x
I;|I;�I;~I;I;�(I;�8I;�MI;�aI;5HI;��H;kgF;i�@;L�4;(�;���:��:��ȺS���(�Z���s9��IY�!��FE	�[
V��e������q<������������-i�.5�T�O���b�      ݶ��O���ά��(�_���7�w�}߿���~,b��V�*l¾Fx�c.���Ž��t�6�����*�?��N�����sx9���:��;��2;U?@;�eF;D�H;��I;��I;9{I;�ZI;�BI;#1I;�$I;�I;�I;OI;�I;�I;�$I;#1I;�BI;�ZI;9{I;��I;��I;D�H;�eF;U?@;��2;��;���:�sx9���N��*�?����6����t���Žc.�Fx�*l¾�V�~,b����}߿w���7�(�_�ά��O���      O���A���}��+Y��3�����$ڿ"����\����(���s��3�9�����p�p�p���<<����d������9}��:�;W$3;io@;yF;��H;�I;�I;�zI;sZI;yBI;�0I;t$I;EI;uI;!I;uI;EI;t$I;�0I;yBI;sZI;�zI;�I;�I;��H;yF;io@;W$3;�;}��:���9d�������<<�p��p���p�9����3��s�(�������\�"���$ڿ����3��+Y�}�A���      ά��}�8tf��lG�Ң%��p�*�ʿV����>M����S����d�ɤ�̷�9�d��
��I��@�1���������9���:N;�T4;��@;�F;A�H;�I;ܙI;�xI;�XI;bAI;�/I;�#I;�I;�I;�I;�I;�I;�#I;�/I;bAI;�XI;�xI;ܙI;�I;A�H;�F;��@;�T4;N;���:��9������@�1��I���
�9�d�̷�ɤ��d�S�������>M�V���*�ʿ�p�Ң%��lG�8tf�}�      (�_��+Y��lG�f.�w���꿭���J䂿��5���󾋰��M�N�W��V��-�Q�*�������:i!��g��*󳺑:��:�;f06;��A;uG;I;Z�I;��I;�uI;qVI;�?I;�.I;�"I;�I;'I;�I;'I;�I;�"I;�.I;�?I;qVI;�uI;��I;Z�I;I;uG;��A;f06;�;��:�:*��g��:i!�����*���-�Q�V��W��M�N���������5�J䂿�������w�f.��lG��+Y�      ��7��3�Ң%�w��<����ſ�����\�9����Ͼ����`�3����z����9�z�ἷ���z��8}�ht�K�^:�)�:Ϣ#;��8;��B;ArG;�$I;ҘI;�I;$qI;7SI;=I;�,I;1!I;oI;I;�I;I;oI;1!I;�,I;=I;7SI;$qI;�I;ҘI;�$I;ArG;��B;��8;Ϣ#;�)�:K�^:ht��8}��z����z�Ἁ�9��z����`�3�������Ͼ9����\������ſ�<��w�Ң%��3�      w�����p������ſ!��{Ps���1�-r���d���d�}I�҈Ž��}�l*�fC��W�^�RC�e�D�"N๫��:��;�);.6;;KD;f�G;lGI;ΜI;ȎI;�kI;OI;�9I;3*I;9I;�I;�I;KI;�I;�I;9I;3*I;�9I;OI;�kI;ȎI;ΜI;lGI;f�G;KD;.6;;�);��;���:"N�e�D�RC�W�^�fC��l*���}�҈Ž}I��d��d��-r����1�{Ps�!����ſ��꿀p����      }߿�$ڿ*�ʿ�������{Ps�MX:����#l¾�ǆ���7����<5��$�Q�����t��85�������:��8ȼ:��;��.;��=;�DE;�XH;�gI;G�I;ڇI;GeI;@JI;E6I;a'I;�I;I;�I;�I;�I;I;�I;a'I;E6I;@JI;GeI;ڇI;G�I;�gI;�XH;�DE;��=;��.;��;ȼ::��8������85��t�����$�Q�<5�������7��ǆ�#l¾���MX:�{Ps��������*�ʿ�$ڿ      ���"��V���J䂿��\���1�����J˾睒�C�N�y��L������c�'���Ҽ �|��z�ko��z��*�&:�N�:̧;�V4;�@;HfF;��H;.�I;B�I;UI;=^I;�DI;&2I;<$I;cI;�I;I;�I;I;�I;cI;<$I;&2I;�DI;=^I;UI;B�I;.�I;��H;HfF;�@;�V4;̧;�N�:*�&:z��ko���z� �|���Ҽc�'����L���y��C�N�睒��J˾�����1���\�J䂿V���"��      ~,b���\��>M���5�9��-r��#l¾睒�"&W��3�<Sؽ�z��fG�����I���?��̻z�-����L��:��;Ͽ&;C{9;�C;�cG;tI;]�I;r�I;ruI;�VI;O?I;�-I;� I;�I;yI;�I;�I;�I;yI;�I;� I;�-I;O?I;�VI;ruI;r�I;]�I;tI;�cG;�C;C{9;Ͽ&;��;L��:���z�-��̻�?��I�����fG��z��<Sؽ�3�"&W�睒�#l¾-r��9����5��>M���\�      �V������������Ͼ�d���ǆ�C�N��3��c�[����\�@��EC��N�o�Ъ	�s숻/�R��9K��:�g;o�/;\�=;bE;2H;�VI;ٜI;�I;�jI;�NI;G9I;)I;=I;�I;I;�I;�
I;�I;I;�I;=I;)I;G9I;�NI;�jI;�I;ٜI;�VI;2H;bE;\�=;o�/;�g;K��:R��9/�s숻Ъ	�N�o�EC��@����\�[���cཱ3�C�N��ǆ��d����Ͼ���������      *l¾(��S������������d���7�y��<Sؽ[���d�P*�kּI\����'�����S������
�:�Y;�#;Z<7;N�A;3�F;|�H;��I;	�I;րI;	`I;�FI;3I;C$I;�I;�I;vI;i	I;iI;i	I;vI;�I;�I;C$I;3I;�FI;	`I;րI;	�I;��I;|�H;3�F;N�A;Z<7;�#;�Y;�
�:�����S������'�I\��kּP*��d�[��<Sؽy����7��d���������S���(��      Fx��s��d�M�N�`�3�}I����L����z����\�P*�'�ݼe���j<<��ڻ��V��gt�u�&:���:\B;�;/;oC=;��D;��G;8I;�I;ÓI;4sI;IUI;}>I;�,I;�I;�I;yI;�	I;I;.I;I;�	I;yI;�I;�I;�,I;}>I;IUI;4sI;ÓI;�I;8I;��G;��D;oC=;�;/;\B;���:u�&:�gt���V��ڻj<<�e���'�ݼP*���\��z��L������}I�`�3�M�N��d��s�      c.��3�ɤ�W����҈Ž<5�����fG�@��kּe���9yC�?�V7}�﮼�W�x9���:&	;O�&;�:8;��A;F;ϸH;WxI;��I;�I;PeI;�JI;m6I;�&I;�I;�I;vI;/I;�I;�I;�I;/I;vI;�I;�I;�&I;m6I;�JI;PeI;�I;��I;WxI;ϸH;F;��A;�:8;O�&;&	;���:W�x9﮼�V7}�?�9yC�e���kּ@��fG����<5��҈Ž��W��ɤ��3�      ��Ž9���̷�V���z����}�$�Q�c�'����EC��I\��j<<�?��n����*U�d��:[��:-�;�&3;��>;�E;�H;};I;�I;ÔI;�uI;�WI;�@I;�.I;� I;�I;I;oI;�I;<I;�I;<I;�I;oI;I;�I;� I;�.I;�@I;�WI;�uI;ÔI;�I;};I;�H;�E;��>;�&3;-�;[��:d��:*U����n��?�j<<�I\��EC�����c�'�$�Q���}��z��V��̷�9���      ��t���p�9�d�-�Q���9�l*������Ҽ�I��N�o���'��ڻV7}���dH��߄:�k�:¿;�.;5<;�nC;^6G;��H;�I;��I;�I;<eI;^KI;7I;�&I;�I;�I;i
I;dI;�I;��H;l�H;��H;�I;dI;i
I;�I;�I;�&I;7I;^KI;<eI;�I;��I;�I;��H;^6G;�nC;5<;�.;¿;�k�:�߄:dH���V7}��ڻ��'�N�o��I����Ҽ���l*���9�-�Q�9�d���p�      6��p��
�*���z��fC���t�� �|��?�Ъ	������V�﮼�*U��߄:��:�g;7�+;�9;��A;�eF;w�H;�^I;��I;��I; rI;�UI;�?I;�-I; I;uI;(I;�I;�I;i�H;��H;�H;��H;i�H;�I;�I;(I;uI; I;�-I;�?I;�UI; rI;��I;��I;�^I;w�H;�eF;��A;�9;7�+;�g;��:�߄:*U�﮼���V����Ъ	��?� �|��t��fC��z��*����
�p�      ���p���I���������W�^�85��z��̻s숻�S��gt�W�x9d��:�k�:�g;z�*;��8;�@; �E;W'H;�7I;ߒI;3�I;o}I;�_I;�GI;�4I;z%I;�I;RI;	I;�I;��H;�H;i�H;��H;i�H;�H;��H;�I;	I;RI;�I;z%I;�4I;�GI;�_I;o}I;3�I;ߒI;�7I;W'H; �E;�@;��8;z�*;�g;�k�:d��:W�x9�gt��S�s숻�̻�z�85�W�^���������I��p��      *�?��<<�@�1�:i!��z�RC����ko��z�-�/򳺬���u�&:���:[��:¿;7�+;��8;X�@;]E;��G;eI;
�I;l�I;P�I;�hI;UOI;#;I;�*I;�I;�I;nI;EI;� I;��H;��H;d�H;��H;d�H;��H;��H;� I;EI;nI;�I;�I;�*I;#;I;UOI;�hI;P�I;l�I;
�I;eI;��G;]E;X�@;��8;7�+;¿;[��:���:u�&:����/�z�-�ko�����RC��z�:i!�@�1��<<�      �N����������g���8}�e�D����z�����R��9�
�:���:&	;-�;�.;�9;�@;]E;��G;]I;�~I;#�I;h�I;�oI;�UI;�@I;�/I;�!I;�I;I;I;�I;��H;s�H;��H;r�H;��H;r�H;��H;s�H;��H;�I;I;I;�I;�!I;�/I;�@I;�UI;�oI;h�I;#�I;�~I;]I;��G;]E;�@;�9;�.;-�;&	;���:�
�:R��9���z�����e�D��8}��g���������      ��d�����*�ht�"N�:��8*�&:L��:K��:�Y;\B;O�&;�&3;5<;��A; �E;��G;]I;w{I;��I;��I;�tI;�ZI;*EI;�3I;E%I;�I;bI;�I;I;O�H;��H;I�H;��H;��H;1�H;��H;��H;I�H;��H;O�H;I;�I;bI;�I;E%I;�3I;*EI;�ZI;�tI;��I;��I;w{I;]I;��G; �E;��A;5<;�&3;O�&;\B;�Y;K��:L��:*�&::��8"N�ht�*���d���      �sx9���9��9�:K�^:���:ȼ:�N�:��;�g;�#;�;/;�:8;��>;�nC;�eF;W'H;eI;�~I;��I;ːI;wI;�]I;RHI;�6I;(I;#I;�I;�
I;\I;b�H;]�H;h�H;L�H;��H;��H;��H;��H;��H;L�H;h�H;]�H;b�H;\I;�
I;�I;#I;(I;�6I;RHI;�]I;wI;ːI;��I;�~I;eI;W'H;�eF;�nC;��>;�:8;�;/;�#;�g;��;�N�:ȼ:���:K�^:�:��9���9      ���:}��:���:��:�)�:��;��;̧;Ͽ&;o�/;Z<7;oC=;��A;�E;^6G;w�H;�7I;
�I;#�I;��I;wI;�^I;�II;�8I;*I;I;LI;QI;�I;M I;�H;��H;*�H;N�H;��H;�H;��H;�H;��H;N�H;*�H;��H;�H;M I;�I;QI;LI;I;*I;�8I;�II;�^I;wI;��I;#�I;
�I;�7I;w�H;^6G;�E;��A;oC=;Z<7;o�/;Ͽ&;̧;��;��;�)�:��:���:}��:      ��;�;N;�;Ϣ#;�);��.;�V4;C{9;\�=;N�A;��D;F;�H;��H;�^I;ߒI;l�I;h�I;�tI;�]I;�II;>9I;6+I;VI;�I;gI;�I;4I;��H;�H;F�H;�H;{�H;p�H;��H;b�H;��H;p�H;{�H;�H;F�H;�H;��H;4I;�I;gI;�I;VI;6+I;>9I;�II;�]I;�tI;h�I;l�I;ߒI;�^I;��H;�H;F;��D;N�A;\�=;C{9;�V4;��.;�);Ϣ#;�;N;�;      ��2;W$3;�T4;f06;��8;.6;;��=;�@;�C;bE;3�F;��G;ϸH;};I;�I;��I;3�I;P�I;�oI;�ZI;RHI;�8I;6+I;�I;5I;2I;iI;�I;Y�H;t�H;q�H;:�H;L�H;��H;��H;i�H;�H;i�H;��H;��H;L�H;:�H;q�H;t�H;Y�H;�I;iI;2I;5I;�I;6+I;�8I;RHI;�ZI;�oI;P�I;3�I;��I;�I;};I;ϸH;��G;3�F;bE;�C;�@;��=;.6;;��8;f06;�T4;W$3;      U?@;io@;��@;��A;��B;KD;�DE;HfF;�cG;2H;|�H;8I;WxI;�I;��I;��I;o}I;�hI;�UI;*EI;�6I;*I;VI;5I;tI;�I;QI;��H;��H;��H;.�H;0�H;��H;}�H;��H;,�H;	�H;,�H;��H;}�H;��H;0�H;.�H;��H;��H;��H;QI;�I;tI;5I;VI;*I;�6I;*EI;�UI;�hI;o}I;��I;��I;�I;WxI;8I;|�H;2H;�cG;HfF;�DE;KD;��B;��A;��@;io@;      �eF;yF;�F;uG;ArG;f�G;�XH;��H;tI;�VI;��I;�I;��I;ÔI;�I; rI;�_I;UOI;�@I;�3I;(I;I;�I;2I;�I;jI;��H;�H;��H;b�H;?�H;r�H;#�H;9�H;|�H;�H;�H;�H;|�H;9�H;#�H;r�H;?�H;b�H;��H;�H;��H;jI;�I;2I;�I;I;(I;�3I;�@I;UOI;�_I; rI;�I;ÔI;��I;�I;��I;�VI;tI;��H;�XH;f�G;ArG;uG;�F;yF;      D�H;��H;A�H;I;�$I;lGI;�gI;.�I;]�I;ٜI;	�I;ÓI;�I;�uI;<eI;�UI;�GI;#;I;�/I;E%I;#I;LI;gI;iI;QI;��H;�H;��H;s�H;@�H;{�H; �H;��H;�H;q�H;�H;�H;�H;q�H;�H;��H; �H;{�H;@�H;s�H;��H;�H;��H;QI;iI;gI;LI;#I;E%I;�/I;#;I;�GI;�UI;<eI;�uI;�I;ÓI;	�I;ٜI;]�I;.�I;�gI;lGI;�$I;I;A�H;��H;      ��I;�I;�I;Z�I;ҘI;ΜI;G�I;B�I;r�I;�I;րI;4sI;PeI;�WI;^KI;�?I;�4I;�*I;�!I;�I;�I;QI;�I;�I;��H;�H;��H;l�H;Q�H;j�H;��H;��H;��H;�H;��H;H�H;1�H;H�H;��H;�H;��H;��H;��H;j�H;Q�H;l�H;��H;�H;��H;�I;�I;QI;�I;�I;�!I;�*I;�4I;�?I;^KI;�WI;PeI;4sI;րI;�I;r�I;B�I;G�I;ΜI;ҘI;Z�I;�I;�I;      ��I;�I;ܙI;��I;�I;ȎI;ڇI;UI;ruI;�jI;	`I;IUI;�JI;�@I;7I;�-I;z%I;�I;�I;bI;�
I;�I;4I;Y�H;��H;��H;s�H;Q�H;j�H;��H;��H;��H;��H;-�H;��H;��H;Y�H;��H;��H;-�H;��H;��H;��H;��H;j�H;Q�H;s�H;��H;��H;Y�H;4I;�I;�
I;bI;�I;�I;z%I;�-I;7I;�@I;�JI;IUI;	`I;�jI;ruI;UI;ڇI;ȎI;�I;��I;ܙI;�I;      9{I;�zI;�xI;�uI;$qI;�kI;GeI;=^I;�VI;�NI;�FI;}>I;m6I;�.I;�&I; I;�I;�I;I;�I;\I;M I;��H;t�H;��H;b�H;@�H;j�H;��H;��H;��H;��H;�H;��H;�H;��H;��H;��H;�H;��H;�H;��H;��H;��H;��H;j�H;@�H;b�H;��H;t�H;��H;M I;\I;�I;I;�I;�I; I;�&I;�.I;m6I;}>I;�FI;�NI;�VI;=^I;GeI;�kI;$qI;�uI;�xI;�zI;      �ZI;sZI;�XI;qVI;7SI;OI;@JI;�DI;O?I;G9I;3I;�,I;�&I;� I;�I;uI;RI;nI;I;I;b�H;�H;�H;q�H;.�H;?�H;{�H;��H;��H;��H;��H;��H;`�H;��H;|�H;c�H;Z�H;c�H;|�H;��H;`�H;��H;��H;��H;��H;��H;{�H;?�H;.�H;q�H;�H;�H;b�H;I;I;nI;RI;uI;�I;� I;�&I;�,I;3I;G9I;O?I;�DI;@JI;OI;7SI;qVI;�XI;sZI;      �BI;yBI;bAI;�?I;=I;�9I;E6I;&2I;�-I;)I;C$I;�I;�I;�I;�I;(I;	I;EI;�I;O�H;]�H;��H;F�H;:�H;0�H;r�H; �H;��H;��H;��H;��H;I�H;��H;U�H;�H;��H;��H;��H;�H;U�H;��H;I�H;��H;��H;��H;��H; �H;r�H;0�H;:�H;F�H;��H;]�H;O�H;�I;EI;	I;(I;�I;�I;�I;�I;C$I;)I;�-I;&2I;E6I;�9I;=I;�?I;bAI;yBI;      #1I;�0I;�/I;�.I;�,I;3*I;a'I;<$I;� I;=I;�I;�I;�I;I;i
I;�I;�I;� I;��H;��H;h�H;*�H;�H;L�H;��H;#�H;��H;��H;��H;�H;`�H;��H;9�H;��H;��H;��H;t�H;��H;��H;��H;9�H;��H;`�H;�H;��H;��H;��H;#�H;��H;L�H;�H;*�H;h�H;��H;��H;� I;�I;�I;i
I;I;�I;�I;�I;=I;� I;<$I;a'I;3*I;�,I;�.I;�/I;�0I;      �$I;t$I;�#I;�"I;1!I;9I;�I;cI;�I;�I;�I;yI;vI;oI;dI;�I;��H;��H;s�H;I�H;L�H;N�H;{�H;��H;}�H;9�H;�H;�H;-�H;��H;��H;U�H;��H;��H;b�H;@�H;)�H;@�H;b�H;��H;��H;U�H;��H;��H;-�H;�H;�H;9�H;}�H;��H;{�H;N�H;L�H;I�H;s�H;��H;��H;�I;dI;oI;vI;yI;�I;�I;�I;cI;�I;9I;1!I;�"I;�#I;t$I;      �I;EI;�I;�I;oI;�I;I;�I;yI;I;vI;�	I;/I;�I;�I;i�H;�H;��H;��H;��H;��H;��H;p�H;��H;��H;|�H;q�H;��H;��H;�H;|�H;�H;��H;b�H;�H;�H;�H;�H;�H;b�H;��H;�H;|�H;�H;��H;��H;q�H;|�H;��H;��H;p�H;��H;��H;��H;��H;��H;�H;i�H;�I;�I;/I;�	I;vI;I;yI;�I;I;�I;oI;�I;�I;EI;      �I;uI;�I;'I;I;�I;�I;I;�I;�I;i	I;I;�I;<I;��H;��H;i�H;d�H;r�H;��H;��H;�H;��H;i�H;,�H;�H;�H;H�H;��H;��H;c�H;��H;��H;@�H;�H;��H;��H;��H;�H;@�H;��H;��H;c�H;��H;��H;H�H;�H;�H;,�H;i�H;��H;�H;��H;��H;r�H;d�H;i�H;��H;��H;<I;�I;I;i	I;�I;�I;I;�I;�I;I;'I;�I;uI;      OI;!I;�I;�I;�I;KI;�I;�I;�I;�
I;iI;.I;�I;�I;l�H;�H;��H;��H;��H;1�H;��H;��H;b�H;�H;	�H;�H;�H;1�H;Y�H;��H;Z�H;��H;t�H;)�H;�H;��H;��H;��H;�H;)�H;t�H;��H;Z�H;��H;Y�H;1�H;�H;�H;	�H;�H;b�H;��H;��H;1�H;��H;��H;��H;�H;l�H;�I;�I;.I;iI;�
I;�I;�I;�I;KI;�I;�I;�I;!I;      �I;uI;�I;'I;I;�I;�I;I;�I;�I;i	I;I;�I;<I;��H;��H;i�H;d�H;r�H;��H;��H;�H;��H;i�H;,�H;�H;�H;H�H;��H;��H;c�H;��H;��H;@�H;�H;��H;��H;��H;�H;@�H;��H;��H;c�H;��H;��H;H�H;�H;�H;,�H;i�H;��H;�H;��H;��H;r�H;d�H;i�H;��H;��H;<I;�I;I;i	I;�I;�I;I;�I;�I;I;'I;�I;uI;      �I;EI;�I;�I;oI;�I;I;�I;yI;I;vI;�	I;/I;�I;�I;i�H;�H;��H;��H;��H;��H;��H;p�H;��H;��H;|�H;q�H;��H;��H;�H;|�H;�H;��H;b�H;�H;�H;�H;�H;�H;b�H;��H;�H;|�H;�H;��H;��H;q�H;|�H;��H;��H;p�H;��H;��H;��H;��H;��H;�H;i�H;�I;�I;/I;�	I;vI;I;yI;�I;I;�I;oI;�I;�I;EI;      �$I;t$I;�#I;�"I;1!I;9I;�I;cI;�I;�I;�I;yI;vI;oI;dI;�I;��H;��H;s�H;I�H;L�H;N�H;{�H;��H;}�H;9�H;�H;�H;-�H;��H;��H;U�H;��H;��H;b�H;@�H;)�H;@�H;b�H;��H;��H;U�H;��H;��H;-�H;�H;�H;9�H;}�H;��H;{�H;N�H;L�H;I�H;s�H;��H;��H;�I;dI;oI;vI;yI;�I;�I;�I;cI;�I;9I;1!I;�"I;�#I;t$I;      #1I;�0I;�/I;�.I;�,I;3*I;a'I;<$I;� I;=I;�I;�I;�I;I;i
I;�I;�I;� I;��H;��H;h�H;*�H;�H;L�H;��H;#�H;��H;��H;��H;�H;`�H;��H;9�H;��H;��H;��H;t�H;��H;��H;��H;9�H;��H;`�H;�H;��H;��H;��H;#�H;��H;L�H;�H;*�H;h�H;��H;��H;� I;�I;�I;i
I;I;�I;�I;�I;=I;� I;<$I;a'I;3*I;�,I;�.I;�/I;�0I;      �BI;yBI;bAI;�?I;=I;�9I;E6I;&2I;�-I;)I;C$I;�I;�I;�I;�I;(I;	I;EI;�I;O�H;]�H;��H;F�H;:�H;0�H;r�H; �H;��H;��H;��H;��H;I�H;��H;U�H;�H;��H;��H;��H;�H;U�H;��H;I�H;��H;��H;��H;��H; �H;r�H;0�H;:�H;F�H;��H;]�H;O�H;�I;EI;	I;(I;�I;�I;�I;�I;C$I;)I;�-I;&2I;E6I;�9I;=I;�?I;bAI;yBI;      �ZI;sZI;�XI;qVI;7SI;OI;@JI;�DI;O?I;G9I;3I;�,I;�&I;� I;�I;uI;RI;nI;I;I;b�H;�H;�H;q�H;.�H;?�H;{�H;��H;��H;��H;��H;��H;`�H;��H;|�H;c�H;Z�H;c�H;|�H;��H;`�H;��H;��H;��H;��H;��H;{�H;?�H;.�H;q�H;�H;�H;b�H;I;I;nI;RI;uI;�I;� I;�&I;�,I;3I;G9I;O?I;�DI;@JI;OI;7SI;qVI;�XI;sZI;      9{I;�zI;�xI;�uI;$qI;�kI;GeI;=^I;�VI;�NI;�FI;}>I;m6I;�.I;�&I; I;�I;�I;I;�I;\I;M I;��H;t�H;��H;b�H;@�H;j�H;��H;��H;��H;��H;�H;��H;�H;��H;��H;��H;�H;��H;�H;��H;��H;��H;��H;j�H;@�H;b�H;��H;t�H;��H;M I;\I;�I;I;�I;�I; I;�&I;�.I;m6I;}>I;�FI;�NI;�VI;=^I;GeI;�kI;$qI;�uI;�xI;�zI;      ��I;�I;ܙI;��I;�I;ȎI;ڇI;UI;ruI;�jI;	`I;IUI;�JI;�@I;7I;�-I;z%I;�I;�I;bI;�
I;�I;4I;Y�H;��H;��H;s�H;Q�H;j�H;��H;��H;��H;��H;-�H;��H;��H;Y�H;��H;��H;-�H;��H;��H;��H;��H;j�H;Q�H;s�H;��H;��H;Y�H;4I;�I;�
I;bI;�I;�I;z%I;�-I;7I;�@I;�JI;IUI;	`I;�jI;ruI;UI;ڇI;ȎI;�I;��I;ܙI;�I;      ��I;�I;�I;Z�I;ҘI;ΜI;G�I;B�I;r�I;�I;րI;4sI;PeI;�WI;^KI;�?I;�4I;�*I;�!I;�I;�I;QI;�I;�I;��H;�H;��H;l�H;Q�H;j�H;��H;��H;��H;�H;��H;H�H;1�H;H�H;��H;�H;��H;��H;��H;j�H;Q�H;l�H;��H;�H;��H;�I;�I;QI;�I;�I;�!I;�*I;�4I;�?I;^KI;�WI;PeI;4sI;րI;�I;r�I;B�I;G�I;ΜI;ҘI;Z�I;�I;�I;      D�H;��H;A�H;I;�$I;lGI;�gI;.�I;]�I;ٜI;	�I;ÓI;�I;�uI;<eI;�UI;�GI;#;I;�/I;E%I;#I;LI;gI;iI;QI;��H;�H;��H;s�H;@�H;{�H; �H;��H;�H;q�H;�H;�H;�H;q�H;�H;��H; �H;{�H;@�H;s�H;��H;�H;��H;QI;iI;gI;LI;#I;E%I;�/I;#;I;�GI;�UI;<eI;�uI;�I;ÓI;	�I;ٜI;]�I;.�I;�gI;lGI;�$I;I;A�H;��H;      �eF;yF;�F;uG;ArG;f�G;�XH;��H;tI;�VI;��I;�I;��I;ÔI;�I; rI;�_I;UOI;�@I;�3I;(I;I;�I;2I;�I;jI;��H;�H;��H;b�H;?�H;r�H;#�H;9�H;|�H;�H;�H;�H;|�H;9�H;#�H;r�H;?�H;b�H;��H;�H;��H;jI;�I;2I;�I;I;(I;�3I;�@I;UOI;�_I; rI;�I;ÔI;��I;�I;��I;�VI;tI;��H;�XH;f�G;ArG;uG;�F;yF;      U?@;io@;��@;��A;��B;KD;�DE;HfF;�cG;2H;|�H;8I;WxI;�I;��I;��I;o}I;�hI;�UI;*EI;�6I;*I;VI;5I;tI;�I;QI;��H;��H;��H;.�H;0�H;��H;}�H;��H;,�H;	�H;,�H;��H;}�H;��H;0�H;.�H;��H;��H;��H;QI;�I;tI;5I;VI;*I;�6I;*EI;�UI;�hI;o}I;��I;��I;�I;WxI;8I;|�H;2H;�cG;HfF;�DE;KD;��B;��A;��@;io@;      ��2;W$3;�T4;f06;��8;.6;;��=;�@;�C;bE;3�F;��G;ϸH;};I;�I;��I;3�I;P�I;�oI;�ZI;RHI;�8I;6+I;�I;5I;2I;iI;�I;Y�H;t�H;q�H;:�H;L�H;��H;��H;i�H;�H;i�H;��H;��H;L�H;:�H;q�H;t�H;Y�H;�I;iI;2I;5I;�I;6+I;�8I;RHI;�ZI;�oI;P�I;3�I;��I;�I;};I;ϸH;��G;3�F;bE;�C;�@;��=;.6;;��8;f06;�T4;W$3;      ��;�;N;�;Ϣ#;�);��.;�V4;C{9;\�=;N�A;��D;F;�H;��H;�^I;ߒI;l�I;h�I;�tI;�]I;�II;>9I;6+I;VI;�I;gI;�I;4I;��H;�H;F�H;�H;{�H;p�H;��H;b�H;��H;p�H;{�H;�H;F�H;�H;��H;4I;�I;gI;�I;VI;6+I;>9I;�II;�]I;�tI;h�I;l�I;ߒI;�^I;��H;�H;F;��D;N�A;\�=;C{9;�V4;��.;�);Ϣ#;�;N;�;      ���:}��:���:��:�)�:��;��;̧;Ͽ&;o�/;Z<7;oC=;��A;�E;^6G;w�H;�7I;
�I;#�I;��I;wI;�^I;�II;�8I;*I;I;LI;QI;�I;M I;�H;��H;*�H;N�H;��H;�H;��H;�H;��H;N�H;*�H;��H;�H;M I;�I;QI;LI;I;*I;�8I;�II;�^I;wI;��I;#�I;
�I;�7I;w�H;^6G;�E;��A;oC=;Z<7;o�/;Ͽ&;̧;��;��;�)�:��:���:}��:      �sx9���9��9�:K�^:���:ȼ:�N�:��;�g;�#;�;/;�:8;��>;�nC;�eF;W'H;eI;�~I;��I;ːI;wI;�]I;RHI;�6I;(I;#I;�I;�
I;\I;b�H;]�H;h�H;L�H;��H;��H;��H;��H;��H;L�H;h�H;]�H;b�H;\I;�
I;�I;#I;(I;�6I;RHI;�]I;wI;ːI;��I;�~I;eI;W'H;�eF;�nC;��>;�:8;�;/;�#;�g;��;�N�:ȼ:���:K�^:�:��9���9      ��d�����*�ht�"N�:��8*�&:L��:K��:�Y;\B;O�&;�&3;5<;��A; �E;��G;]I;w{I;��I;��I;�tI;�ZI;*EI;�3I;E%I;�I;bI;�I;I;O�H;��H;I�H;��H;��H;1�H;��H;��H;I�H;��H;O�H;I;�I;bI;�I;E%I;�3I;*EI;�ZI;�tI;��I;��I;w{I;]I;��G; �E;��A;5<;�&3;O�&;\B;�Y;K��:L��:*�&::��8"N�ht�*���d���      �N����������g���8}�e�D����z�����R��9�
�:���:&	;-�;�.;�9;�@;]E;��G;]I;�~I;#�I;h�I;�oI;�UI;�@I;�/I;�!I;�I;I;I;�I;��H;s�H;��H;r�H;��H;r�H;��H;s�H;��H;�I;I;I;�I;�!I;�/I;�@I;�UI;�oI;h�I;#�I;�~I;]I;��G;]E;�@;�9;�.;-�;&	;���:�
�:R��9���z�����e�D��8}��g���������      *�?��<<�@�1�:i!��z�RC����ko��z�-�/򳺬���u�&:���:[��:¿;7�+;��8;X�@;]E;��G;eI;
�I;l�I;P�I;�hI;UOI;#;I;�*I;�I;�I;nI;EI;� I;��H;��H;d�H;��H;d�H;��H;��H;� I;EI;nI;�I;�I;�*I;#;I;UOI;�hI;P�I;l�I;
�I;eI;��G;]E;X�@;��8;7�+;¿;[��:���:u�&:����/�z�-�ko�����RC��z�:i!�@�1��<<�      ���p���I���������W�^�85��z��̻s숻�S��gt�W�x9d��:�k�:�g;z�*;��8;�@; �E;W'H;�7I;ߒI;3�I;o}I;�_I;�GI;�4I;z%I;�I;RI;	I;�I;��H;�H;i�H;��H;i�H;�H;��H;�I;	I;RI;�I;z%I;�4I;�GI;�_I;o}I;3�I;ߒI;�7I;W'H; �E;�@;��8;z�*;�g;�k�:d��:W�x9�gt��S�s숻�̻�z�85�W�^���������I��p��      6��p��
�*���z��fC���t�� �|��?�Ъ	������V�﮼�*U��߄:��:�g;7�+;�9;��A;�eF;w�H;�^I;��I;��I; rI;�UI;�?I;�-I; I;uI;(I;�I;�I;i�H;��H;�H;��H;i�H;�I;�I;(I;uI; I;�-I;�?I;�UI; rI;��I;��I;�^I;w�H;�eF;��A;�9;7�+;�g;��:�߄:*U�﮼���V����Ъ	��?� �|��t��fC��z��*����
�p�      ��t���p�9�d�-�Q���9�l*������Ҽ�I��N�o���'��ڻV7}���dH��߄:�k�:¿;�.;5<;�nC;^6G;��H;�I;��I;�I;<eI;^KI;7I;�&I;�I;�I;i
I;dI;�I;��H;l�H;��H;�I;dI;i
I;�I;�I;�&I;7I;^KI;<eI;�I;��I;�I;��H;^6G;�nC;5<;�.;¿;�k�:�߄:dH���V7}��ڻ��'�N�o��I����Ҽ���l*���9�-�Q�9�d���p�      ��Ž9���̷�V���z����}�$�Q�c�'����EC��I\��j<<�?��n����*U�d��:[��:-�;�&3;��>;�E;�H;};I;�I;ÔI;�uI;�WI;�@I;�.I;� I;�I;I;oI;�I;<I;�I;<I;�I;oI;I;�I;� I;�.I;�@I;�WI;�uI;ÔI;�I;};I;�H;�E;��>;�&3;-�;[��:d��:*U����n��?�j<<�I\��EC�����c�'�$�Q���}��z��V��̷�9���      c.��3�ɤ�W����҈Ž<5�����fG�@��kּe���9yC�?�V7}�﮼�W�x9���:&	;O�&;�:8;��A;F;ϸH;WxI;��I;�I;PeI;�JI;m6I;�&I;�I;�I;vI;/I;�I;�I;�I;/I;vI;�I;�I;�&I;m6I;�JI;PeI;�I;��I;WxI;ϸH;F;��A;�:8;O�&;&	;���:W�x9﮼�V7}�?�9yC�e���kּ@��fG����<5��҈Ž��W��ɤ��3�      Fx��s��d�M�N�`�3�}I����L����z����\�P*�'�ݼe���j<<��ڻ��V��gt�u�&:���:\B;�;/;oC=;��D;��G;8I;�I;ÓI;4sI;IUI;}>I;�,I;�I;�I;yI;�	I;I;.I;I;�	I;yI;�I;�I;�,I;}>I;IUI;4sI;ÓI;�I;8I;��G;��D;oC=;�;/;\B;���:u�&:�gt���V��ڻj<<�e���'�ݼP*���\��z��L������}I�`�3�M�N��d��s�      *l¾(��S������������d���7�y��<Sؽ[���d�P*�kּI\����'�����S������
�:�Y;�#;Z<7;N�A;3�F;|�H;��I;	�I;րI;	`I;�FI;3I;C$I;�I;�I;vI;i	I;iI;i	I;vI;�I;�I;C$I;3I;�FI;	`I;րI;	�I;��I;|�H;3�F;N�A;Z<7;�#;�Y;�
�:�����S������'�I\��kּP*��d�[��<Sؽy����7��d���������S���(��      �V������������Ͼ�d���ǆ�C�N��3��c�[����\�@��EC��N�o�Ъ	�s숻/�R��9K��:�g;o�/;\�=;bE;2H;�VI;ٜI;�I;�jI;�NI;G9I;)I;=I;�I;I;�I;�
I;�I;I;�I;=I;)I;G9I;�NI;�jI;�I;ٜI;�VI;2H;bE;\�=;o�/;�g;K��:R��9/�s숻Ъ	�N�o�EC��@����\�[���cཱ3�C�N��ǆ��d����Ͼ���������      ~,b���\��>M���5�9��-r��#l¾睒�"&W��3�<Sؽ�z��fG�����I���?��̻z�-����L��:��;Ͽ&;C{9;�C;�cG;tI;]�I;r�I;ruI;�VI;O?I;�-I;� I;�I;yI;�I;�I;�I;yI;�I;� I;�-I;O?I;�VI;ruI;r�I;]�I;tI;�cG;�C;C{9;Ͽ&;��;L��:���z�-��̻�?��I�����fG��z��<Sؽ�3�"&W�睒�#l¾-r��9����5��>M���\�      ���"��V���J䂿��\���1�����J˾睒�C�N�y��L������c�'���Ҽ �|��z�ko��z��*�&:�N�:̧;�V4;�@;HfF;��H;.�I;B�I;UI;=^I;�DI;&2I;<$I;cI;�I;I;�I;I;�I;cI;<$I;&2I;�DI;=^I;UI;B�I;.�I;��H;HfF;�@;�V4;̧;�N�:*�&:z��ko���z� �|���Ҽc�'����L���y��C�N�睒��J˾�����1���\�J䂿V���"��      }߿�$ڿ*�ʿ�������{Ps�MX:����#l¾�ǆ���7����<5��$�Q�����t��85�������:��8ȼ:��;��.;��=;�DE;�XH;�gI;G�I;ڇI;GeI;@JI;E6I;a'I;�I;I;�I;�I;�I;I;�I;a'I;E6I;@JI;GeI;ڇI;G�I;�gI;�XH;�DE;��=;��.;��;ȼ::��8������85��t�����$�Q�<5�������7��ǆ�#l¾���MX:�{Ps��������*�ʿ�$ڿ      w�����p������ſ!��{Ps���1�-r���d���d�}I�҈Ž��}�l*�fC��W�^�RC�e�D�"N๫��:��;�);.6;;KD;f�G;lGI;ΜI;ȎI;�kI;OI;�9I;3*I;9I;�I;�I;KI;�I;�I;9I;3*I;�9I;OI;�kI;ȎI;ΜI;lGI;f�G;KD;.6;;�);��;���:"N�e�D�RC�W�^�fC��l*���}�҈Ž}I��d��d��-r����1�{Ps�!����ſ��꿀p����      ��7��3�Ң%�w��<����ſ�����\�9����Ͼ����`�3����z����9�z�ἷ���z��8}�ht�K�^:�)�:Ϣ#;��8;��B;ArG;�$I;ҘI;�I;$qI;7SI;=I;�,I;1!I;oI;I;�I;I;oI;1!I;�,I;=I;7SI;$qI;�I;ҘI;�$I;ArG;��B;��8;Ϣ#;�)�:K�^:ht��8}��z����z�Ἁ�9��z����`�3�������Ͼ9����\������ſ�<��w�Ң%��3�      (�_��+Y��lG�f.�w���꿭���J䂿��5���󾋰��M�N�W��V��-�Q�*�������:i!��g��*󳺑:��:�;f06;��A;uG;I;Z�I;��I;�uI;qVI;�?I;�.I;�"I;�I;'I;�I;'I;�I;�"I;�.I;�?I;qVI;�uI;��I;Z�I;I;uG;��A;f06;�;��:�:*��g��:i!�����*���-�Q�V��W��M�N���������5�J䂿�������w�f.��lG��+Y�      ά��}�8tf��lG�Ң%��p�*�ʿV����>M����S����d�ɤ�̷�9�d��
��I��@�1���������9���:N;�T4;��@;�F;A�H;�I;ܙI;�xI;�XI;bAI;�/I;�#I;�I;�I;�I;�I;�I;�#I;�/I;bAI;�XI;�xI;ܙI;�I;A�H;�F;��@;�T4;N;���:��9������@�1��I���
�9�d�̷�ɤ��d�S�������>M�V���*�ʿ�p�Ң%��lG�8tf�}�      O���A���}��+Y��3�����$ڿ"����\����(���s��3�9�����p�p�p���<<����d������9}��:�;W$3;io@;yF;��H;�I;�I;�zI;sZI;yBI;�0I;t$I;EI;uI;!I;uI;EI;t$I;�0I;yBI;sZI;�zI;�I;�I;��H;yF;io@;W$3;�;}��:���9d�������<<�p��p���p�9����3��s�(�������\�"���$ڿ����3��+Y�}�A���      ����,������Q���F�Q�Ù$�.���~�7�}�E(�>�׾�T���L+���սr����@L��jO�8�ͻ����l8�m�:��;U�1;��?;uF;s�H;��I;��I;��I;�uI;�VI;�@I;1I;�&I;� I;I;� I;�&I;1I;�@I;�VI;�uI;��I;��I;��I;s�H;uF;��?;U�1;��;�m�:�l8���8�ͻjO�@L����r����ս�L+��T��>�׾E(�7�}�~�.���Ù$�F�Q�Q��������,��      �,��^�� P���{��K��x �����n�����w��$���Ҿf��� (���ѽٷ��7����$�K��ɻ����8���:��;��1;@;��F;.I;�I;4�I;ŝI;�tI;OVI;�@I;�0I;�&I;� I;�I;� I;�&I;�0I;�@I;OVI;�tI;ŝI;4�I;�I;.I;��F;@;��1;��;���:��8���ɻ$�K����7�ٷ����ѽ (�f�����Ҿ�$���w�n��������x ��K��{� P��^��      ���� P�������d���;� ����㿰���#f�b��ž��z���C�ƽ40v�d5�R����o@����oj��Pu9_I�:>\;�63;@�@;�F;XI;��I;{�I;p�I;�rI;�TI;^?I;0I;&I;, I;MI;, I;&I;0I;^?I;�TI;�rI;p�I;{�I;��I;XI;�F;@�@;�63;>\;_I�:�Pu9oj�����o@�R���d5�40v�C�ƽ����z�žb��#f�������� ����;���d���� P��      Q����{���d��F�Ù$�7����ɿ,蒿��K�O���j�� Zb�H�8�����a����`���%�.� e��V�غ̨�9�W�:VW;�15;@�A;� G;[6I;��I;k�I;m�I;�oI;�RI;�=I;�.I;�$I;AI;OI;AI;�$I;�.I;�=I;�RI;�oI;m�I;k�I;��I;[6I;� G;@�A;�15;VW;�W�:̨�9V�غ e��%�.�`��������a�8���H� Zb��j��O����K�,蒿��ɿ7��Ù$��F���d��{�      F�Q��K���;�Ù$��;
��޿�����w�o,���澝���(�D������I��3�G�����N��Ǩ�1��9�����9:���:�m!;��7;۸B;}�G;
YI;L�I;��I;ّI;�kI;�OI;4;I;�,I;3#I;�I;�I;�I;3#I;�,I;4;I;�OI;�kI;ّI;��I;L�I;
YI;}�G;۸B;��7;�m!;���:��9:9���1��Ǩ��N�����3�G��I������(�D��������o,���w�����޿�;
�Ù$���;��K�      Ù$��x � ��7���޿m���ǅ����F�{�
��~����z��$���ս$���P2+���ϼWPp����J�]��*�#��:-�;�7';��:;�C;,H;�|I;?�I;��I;��I;�fI;�KI;:8I;V*I;E!I;I;GI;I;E!I;V*I;:8I;�KI;�fI;��I;��I;?�I;�|I;,H;�C;��:;�7';-�;#��:�*�J�]����WPp���ϼP2+�$�����ս�$���z��~��{�
���F�ǅ��m����޿7�� ���x �      .���������㿆�ɿ���ǅ����P�b��:�׾�`��U�H����@��a�a�!����!D�Gɻ�!������U�:�~;�H-;H{=;BBE;ȄH;)�I; �I;��I;ׂI;�`I;BGI;�4I;�'I;�I;I;pI;I;�I;�'I;�4I;BGI;�`I;ׂI;��I; �I;)�I;ȄH;BBE;H{=;�H-;�~;�U�:�����!�Gɻ!D���!��a�a��@����U�H��`��:�׾b����P�ǅ�������ɿ��㿯���      ~�n�������,蒿��w���F�b��Ȱ�����Yb�+����ѽ�%��'D4����@X��ʨ��H���轺P��9cp�:�; 93;;P@;�uF;9�H;&�I;��I;��I;�yI;�YI;3BI;�0I;�$I;eI;�I;@I;�I;eI;�$I;�0I;3BI;�YI;�yI;��I;��I;&�I;9�H;�uF;;P@; 93;�;cp�:P��9�轺�H��ʨ�@X�����'D4��%����ѽ+���Yb����Ȱ�b����F���w�,蒿����n���      7�}���w�#f���K�o,�{�
�:�׾�����k���'�lz꽥I���;V�LM�*����iO��G�mpE����c�:T� ;¾$;̳8;r�B;�G;VJI;1�I;:�I;a�I;*pI;�RI;�<I;�,I;%!I;�I;9I;�I;9I;�I;%!I;�,I;�<I;�RI;*pI;a�I;:�I;1�I;VJI;�G;r�B;̳8;¾$;T� ;c�:���mpE��G��iO�*���LM��;V��I��lz���'���k����:�׾{�
�o,���K�#f���w�      E(��$�b��O������~���`���Yb���'��U�N$��S�m�5����ϼ0�����_�����غ�0�9d��:F;�F.;3{=;bE;�[H;B�I;��I;��I;�I;%fI;&KI;7I;&(I;�I;�I;�I;DI;�I;�I;�I;&(I;7I;&KI;%fI;�I;��I;��I;B�I;�[H;bE;3{=;�F.;F;d��:�0�9��غ_������0����ϼ5��S�m�N$���U���'��Yb��`���~�����O��b���$�      >�׾��Ҿž�j��������z�U�H�+��lz�N$��0v�!2+����9���5�-ɻ34�0�����:���:Nn!;*O6;)kA;��F;��H;��I;��I;�I;k|I;�[I;~CI;%1I;�#I;�I;jI;�I;�I;�I;jI;�I;�#I;%1I;~CI;�[I;k|I;�I;��I;��I;��H;��F;)kA;*O6;Nn!;���:���:0��34�-ɻ�5�9�����!2+�0v�N$��lz�+��U�H���z������j��ž��Ҿ      �T��f�����z� Zb�(�D��$�����ѽ�I��S�m�!2+��������K��ﻙ�p�:�����9MR�:�.;��-;��<;iyD;uH;�lI;�I;��I;��I;�nI;�QI;�;I;!+I;�I;*I;OI;�I;�I;�I;OI;*I;�I;!+I;�;I;�QI;�nI;��I;��I;�I;�lI;uH;iyD;��<;��-;�.;MR�:��9:�����p��ﻍ�K������!2+�S�m��I����ѽ���$�(�D� Zb���z�f���      �L+� (���H�������ս�@���%���;V�5���������MS�������yF�)�n8o�:�;��$;^7;K�A;��F;�H;��I;��I;��I;��I;uaI;�GI;.4I;A%I;II;ZI;I;�	I; 	I;�	I;I;ZI;II;A%I;.4I;�GI;uaI;��I;��I;��I;��I;�H;��F;K�A;^7;��$;�;o�:)�n8yF⺦������MS�������5���;V��%���@����ս����H��� (�      ��ս��ѽC�ƽ8����I��$���a�a�'D4�LM���ϼ9����K�����G��\g�e�o���:�@�:�X;��1;kk>;�
E;/H;;pI;"�I;	�I;��I;!rI;�TI;>I;�,I;~I;�I;�I;�	I;/I;MI;/I;�	I;�I;�I;~I;�,I;>I;�TI;!rI;��I;	�I;"�I;;pI;/H;�
E;kk>;��1;�X;�@�:��:e�o�\g��G�������K�9����ϼLM�'D4�a�a�$����I��8���C�ƽ��ѽ      r��ٷ��40v���a�3�G�P2+�!�����*���0���5��ﻦ��\g��ହ�g:_�:�;1H-;3f;;NC;)RG;�I;�I;@�I;�I;%�I;+bI;�HI;�4I;�%I;�I;PI;�
I;�I;eI;sI;eI;�I;�
I;PI;�I;�%I;�4I;�HI;+bI;%�I;�I;@�I;�I;�I;)RG;NC;3f;;1H-;�;_�:�g:�ହ\g�������5�0��*������!��P2+�3�G���a�40v�ٷ��      ��7�d5���������ϼ��@X���iO����-ɻ��p�yF�e�o��g:^�:ZF;�*;�9;��A;�tF;<�H;�I;��I;ɺI;e�I;�oI;SSI;n=I;9,I;�I;�I;I;pI;�I;�I;� I;�I;�I;pI;I;�I;�I;9,I;n=I;SSI;�oI;e�I;ɺI;��I;�I;<�H;�tF;��A;�9;�*;ZF;^�:�g:e�o�yF⺙�p�-ɻ����iO�@X������ϼ������d5�7�      @L�����R���`����N��WPp�!D�ʨ��G�_���34�:���)�n8��:_�:ZF;�(;��7;v�@;��E;nPH;6lI;��I;�I;��I;C|I;�]I;�EI;�2I;�#I;{I;�I;		I;(I;� I;�H;h�H;�H;� I;(I;		I;�I;{I;�#I;�2I;�EI;�]I;C|I;��I;�I;��I;6lI;nPH;��E;v�@;��7;�(;ZF;_�:��:)�n8:���34�_����G�ʨ�!D�WPp��N��`���R������      jO�$�K��o@�%�.�Ǩ����Gɻ�H��mpE���غ0����9o�:�@�:�;�*;��7;�O@;�[E;H;�HI;��I;��I;)�I;|�I;ZgI;�MI;z9I;W)I;�I;�I;�
I;,I;'I;G�H;s�H;��H;s�H;G�H;'I;,I;�
I;�I;�I;W)I;z9I;�MI;ZgI;|�I;)�I;��I;��I;�HI;H;�[E;�O@;��7;�*;�;�@�:o�:��90����غmpE��H��Gɻ���Ǩ�%�.��o@�$�K�      8�ͻ�ɻ��� e��1��J�]��!��轺����0�9���:MR�:�;�X;1H-;�9;v�@;�[E;��G;Q4I;ֳI;d�I;��I;m�I;�oI;�TI;q?I;M.I;� I;�I;ZI;�I;�I;6�H;��H;,�H;��H;,�H;��H;6�H;�I;�I;ZI;�I;� I;M.I;q?I;�TI;�oI;m�I;��I;d�I;ֳI;Q4I;��G;�[E;v�@;�9;1H-;�X;�;MR�:���:�0�9����轺�!�J�]�1�� e������ɻ      �����oj�V�غ9����*�����P��9c�:d��:���:�.;��$;��1;3f;;��A;��E;H;Q4I;X�I;��I;m�I;��I;�uI;tZI;yDI;�2I;L$I;�I;�I;hI;�I;��H;t�H;7�H;��H;��H;��H;7�H;t�H;��H;�I;hI;�I;�I;L$I;�2I;yDI;tZI;�uI;��I;m�I;��I;X�I;Q4I;H;��E;��A;3f;;��1;��$;�.;���:d��:c�:P��9�����*�9���V�غoj���      �l8��8�Pu9̨�9��9:#��:�U�:cp�:T� ;F;Nn!;��-;^7;kk>;NC;�tF;nPH;�HI;ֳI;��I;кI;ԙI;�yI;�^I;aHI;e6I;}'I;vI;�I;1
I;�I;>�H;��H;��H;�H;��H;��H;��H;�H;��H;��H;>�H;�I;1
I;�I;vI;}'I;e6I;aHI;�^I;�yI;ԙI;кI;��I;ֳI;�HI;nPH;�tF;NC;kk>;^7;��-;Nn!;F;T� ;cp�:�U�:#��:��9:̨�9�Pu9��8      �m�:���:_I�:�W�:���:-�;�~;�;¾$;�F.;*O6;��<;K�A;�
E;)RG;<�H;6lI;��I;d�I;m�I;ԙI;�zI;�`I;�JI;�8I;�)I;�I;�I;�I;9I; I;�H;��H;{�H; �H;�H;��H;�H; �H;{�H;��H;�H; I;9I;�I;�I;�I;�)I;�8I;�JI;�`I;�zI;ԙI;m�I;d�I;��I;6lI;<�H;)RG;�
E;K�A;��<;*O6;�F.;¾$;�;�~;-�;���:�W�:_I�:���:      ��;��;>\;VW;�m!;�7';�H-; 93;̳8;3{=;)kA;iyD;��F;/H;�I;�I;��I;��I;��I;��I;�yI;�`I;�KI;4:I;+I;FI;8I;I;MI;� I;��H;�H;w�H;�H;�H;a�H;2�H;a�H;�H;�H;w�H;�H;��H;� I;MI;I;8I;FI;+I;4:I;�KI;�`I;�yI;��I;��I;��I;��I;�I;�I;/H;��F;iyD;)kA;3{=;̳8; 93;�H-;�7';�m!;VW;>\;��;      U�1;��1;�63;�15;��7;��:;H{=;;P@;r�B;bE;��F;uH;�H;;pI;�I;��I;�I;)�I;m�I;�uI;�^I;�JI;4:I;�+I; I;+I;�I;*I;�I;�H;��H;~�H;4�H;��H;{�H;��H;��H;��H;{�H;��H;4�H;~�H;��H;�H;�I;*I;�I;+I; I;�+I;4:I;�JI;�^I;�uI;m�I;)�I;�I;��I;�I;;pI;�H;uH;��F;bE;r�B;;P@;H{=;��:;��7;�15;�63;��1;      ��?;@;@�@;@�A;۸B;�C;BBE;�uF;�G;�[H;��H;�lI;��I;"�I;@�I;ɺI;��I;|�I;�oI;tZI;aHI;�8I;+I; I;�I;tI;�I;I;t�H;��H;��H;;�H;d�H;��H;��H;f�H;=�H;f�H;��H;��H;d�H;;�H;��H;��H;t�H;I;�I;tI;�I; I;+I;�8I;aHI;tZI;�oI;|�I;��I;ɺI;@�I;"�I;��I;�lI;��H;�[H;�G;�uF;BBE;�C;۸B;@�A;@�@;@;      uF;��F;�F;� G;}�G;,H;ȄH;9�H;VJI;B�I;��I;�I;��I;	�I;�I;e�I;C|I;ZgI;�TI;yDI;e6I;�)I;FI;+I;tI;�I;ZI;��H;��H;��H;6�H;I�H;��H;j�H;��H;$�H;��H;$�H;��H;j�H;��H;I�H;6�H;��H;��H;��H;ZI;�I;tI;+I;FI;�)I;e6I;yDI;�TI;ZgI;C|I;e�I;�I;	�I;��I;�I;��I;B�I;VJI;9�H;ȄH;,H;}�G;� G;�F;��F;      s�H;.I;XI;[6I;
YI;�|I;)�I;&�I;1�I;��I;��I;��I;��I;��I;%�I;�oI;�]I;�MI;q?I;�2I;}'I;�I;8I;�I;�I;ZI;��H;2�H;��H;@�H;1�H;s�H;&�H;#�H;��H;�H;��H;�H;��H;#�H;&�H;s�H;1�H;@�H;��H;2�H;��H;ZI;�I;�I;8I;�I;}'I;�2I;q?I;�MI;�]I;�oI;%�I;��I;��I;��I;��I;��I;1�I;&�I;)�I;�|I;
YI;[6I;XI;.I;      ��I;�I;��I;��I;L�I;?�I; �I;��I;:�I;��I;�I;��I;��I;!rI;+bI;SSI;�EI;z9I;M.I;L$I;vI;�I;I;*I;I;��H;2�H;�H;M�H;-�H;e�H;��H;��H;�H;b�H;	�H;��H;	�H;b�H;�H;��H;��H;e�H;-�H;M�H;�H;2�H;��H;I;*I;I;�I;vI;L$I;M.I;z9I;�EI;SSI;+bI;!rI;��I;��I;�I;��I;:�I;��I; �I;?�I;L�I;��I;��I;�I;      ��I;4�I;{�I;k�I;��I;��I;��I;��I;a�I;�I;k|I;�nI;uaI;�TI;�HI;n=I;�2I;W)I;� I;�I;�I;�I;MI;�I;t�H;��H;��H;M�H;8�H;a�H;��H;��H;��H;�H;��H;<�H;5�H;<�H;��H;�H;��H;��H;��H;a�H;8�H;M�H;��H;��H;t�H;�I;MI;�I;�I;�I;� I;W)I;�2I;n=I;�HI;�TI;uaI;�nI;k|I;�I;a�I;��I;��I;��I;��I;k�I;{�I;4�I;      ��I;ŝI;p�I;m�I;ّI;��I;ׂI;�yI;*pI;%fI;�[I;�QI;�GI;>I;�4I;9,I;�#I;�I;�I;�I;1
I;9I;� I;�H;��H;��H;@�H;-�H;a�H;��H;��H;��H;��H;"�H;��H;��H;c�H;��H;��H;"�H;��H;��H;��H;��H;a�H;-�H;@�H;��H;��H;�H;� I;9I;1
I;�I;�I;�I;�#I;9,I;�4I;>I;�GI;�QI;�[I;%fI;*pI;�yI;ׂI;��I;ّI;m�I;p�I;ŝI;      �uI;�tI;�rI;�oI;�kI;�fI;�`I;�YI;�RI;&KI;~CI;�;I;.4I;�,I;�%I;�I;{I;�I;ZI;hI;�I; I;��H;��H;��H;6�H;1�H;e�H;��H;��H;��H;��H;��H;c�H;�H;��H;��H;��H;�H;c�H;��H;��H;��H;��H;��H;e�H;1�H;6�H;��H;��H;��H; I;�I;hI;ZI;�I;{I;�I;�%I;�,I;.4I;�;I;~CI;&KI;�RI;�YI;�`I;�fI;�kI;�oI;�rI;�tI;      �VI;OVI;�TI;�RI;�OI;�KI;BGI;3BI;�<I;7I;%1I;!+I;A%I;~I;�I;�I;�I;�
I;�I;�I;>�H;�H;�H;~�H;;�H;I�H;s�H;��H;��H;��H;��H;��H;K�H;��H;��H;J�H;P�H;J�H;��H;��H;K�H;��H;��H;��H;��H;��H;s�H;I�H;;�H;~�H;�H;�H;>�H;�I;�I;�
I;�I;�I;�I;~I;A%I;!+I;%1I;7I;�<I;3BI;BGI;�KI;�OI;�RI;�TI;OVI;      �@I;�@I;^?I;�=I;4;I;:8I;�4I;�0I;�,I;&(I;�#I;�I;II;�I;PI;I;		I;,I;�I;��H;��H;��H;w�H;4�H;d�H;��H;&�H;��H;��H;��H;��H;K�H;��H;d�H;�H;��H;��H;��H;�H;d�H;��H;K�H;��H;��H;��H;��H;&�H;��H;d�H;4�H;w�H;��H;��H;��H;�I;,I;		I;I;PI;�I;II;�I;�#I;&(I;�,I;�0I;�4I;:8I;4;I;�=I;^?I;�@I;      1I;�0I;0I;�.I;�,I;V*I;�'I;�$I;%!I;�I;�I;*I;ZI;�I;�
I;pI;(I;'I;6�H;t�H;��H;{�H;�H;��H;��H;j�H;#�H;�H;�H;"�H;c�H;��H;d�H;��H;��H;��H;��H;��H;��H;��H;d�H;��H;c�H;"�H;�H;�H;#�H;j�H;��H;��H;�H;{�H;��H;t�H;6�H;'I;(I;pI;�
I;�I;ZI;*I;�I;�I;%!I;�$I;�'I;V*I;�,I;�.I;0I;�0I;      �&I;�&I;&I;�$I;3#I;E!I;�I;eI;�I;�I;jI;OI;I;�	I;�I;�I;� I;G�H;��H;7�H;�H; �H;�H;{�H;��H;��H;��H;b�H;��H;��H;�H;��H;�H;��H;��H;d�H;[�H;d�H;��H;��H;�H;��H;�H;��H;��H;b�H;��H;��H;��H;{�H;�H; �H;�H;7�H;��H;G�H;� I;�I;�I;�	I;I;OI;jI;�I;�I;eI;�I;E!I;3#I;�$I;&I;�&I;      � I;� I;, I;AI;�I;I;I;�I;9I;�I;�I;�I;�	I;/I;eI;�I;�H;s�H;,�H;��H;��H;�H;a�H;��H;f�H;$�H;�H;	�H;<�H;��H;��H;J�H;��H;��H;d�H;2�H;/�H;2�H;d�H;��H;��H;J�H;��H;��H;<�H;	�H;�H;$�H;f�H;��H;a�H;�H;��H;��H;,�H;s�H;�H;�I;eI;/I;�	I;�I;�I;�I;9I;�I;I;I;�I;AI;, I;� I;      I;�I;MI;OI;�I;GI;pI;@I;�I;DI;�I;�I; 	I;MI;sI;� I;h�H;��H;��H;��H;��H;��H;2�H;��H;=�H;��H;��H;��H;5�H;c�H;��H;P�H;��H;��H;[�H;/�H;�H;/�H;[�H;��H;��H;P�H;��H;c�H;5�H;��H;��H;��H;=�H;��H;2�H;��H;��H;��H;��H;��H;h�H;� I;sI;MI; 	I;�I;�I;DI;�I;@I;pI;GI;�I;OI;MI;�I;      � I;� I;, I;AI;�I;I;I;�I;9I;�I;�I;�I;�	I;/I;eI;�I;�H;s�H;,�H;��H;��H;�H;a�H;��H;f�H;$�H;�H;	�H;<�H;��H;��H;J�H;��H;��H;d�H;2�H;/�H;2�H;d�H;��H;��H;J�H;��H;��H;<�H;	�H;�H;$�H;f�H;��H;a�H;�H;��H;��H;,�H;s�H;�H;�I;eI;/I;�	I;�I;�I;�I;9I;�I;I;I;�I;AI;, I;� I;      �&I;�&I;&I;�$I;3#I;E!I;�I;eI;�I;�I;jI;OI;I;�	I;�I;�I;� I;G�H;��H;7�H;�H; �H;�H;{�H;��H;��H;��H;b�H;��H;��H;�H;��H;�H;��H;��H;d�H;[�H;d�H;��H;��H;�H;��H;�H;��H;��H;b�H;��H;��H;��H;{�H;�H; �H;�H;7�H;��H;G�H;� I;�I;�I;�	I;I;OI;jI;�I;�I;eI;�I;E!I;3#I;�$I;&I;�&I;      1I;�0I;0I;�.I;�,I;V*I;�'I;�$I;%!I;�I;�I;*I;ZI;�I;�
I;pI;(I;'I;6�H;t�H;��H;{�H;�H;��H;��H;j�H;#�H;�H;�H;"�H;c�H;��H;d�H;��H;��H;��H;��H;��H;��H;��H;d�H;��H;c�H;"�H;�H;�H;#�H;j�H;��H;��H;�H;{�H;��H;t�H;6�H;'I;(I;pI;�
I;�I;ZI;*I;�I;�I;%!I;�$I;�'I;V*I;�,I;�.I;0I;�0I;      �@I;�@I;^?I;�=I;4;I;:8I;�4I;�0I;�,I;&(I;�#I;�I;II;�I;PI;I;		I;,I;�I;��H;��H;��H;w�H;4�H;d�H;��H;&�H;��H;��H;��H;��H;K�H;��H;d�H;�H;��H;��H;��H;�H;d�H;��H;K�H;��H;��H;��H;��H;&�H;��H;d�H;4�H;w�H;��H;��H;��H;�I;,I;		I;I;PI;�I;II;�I;�#I;&(I;�,I;�0I;�4I;:8I;4;I;�=I;^?I;�@I;      �VI;OVI;�TI;�RI;�OI;�KI;BGI;3BI;�<I;7I;%1I;!+I;A%I;~I;�I;�I;�I;�
I;�I;�I;>�H;�H;�H;~�H;;�H;I�H;s�H;��H;��H;��H;��H;��H;K�H;��H;��H;J�H;P�H;J�H;��H;��H;K�H;��H;��H;��H;��H;��H;s�H;I�H;;�H;~�H;�H;�H;>�H;�I;�I;�
I;�I;�I;�I;~I;A%I;!+I;%1I;7I;�<I;3BI;BGI;�KI;�OI;�RI;�TI;OVI;      �uI;�tI;�rI;�oI;�kI;�fI;�`I;�YI;�RI;&KI;~CI;�;I;.4I;�,I;�%I;�I;{I;�I;ZI;hI;�I; I;��H;��H;��H;6�H;1�H;e�H;��H;��H;��H;��H;��H;c�H;�H;��H;��H;��H;�H;c�H;��H;��H;��H;��H;��H;e�H;1�H;6�H;��H;��H;��H; I;�I;hI;ZI;�I;{I;�I;�%I;�,I;.4I;�;I;~CI;&KI;�RI;�YI;�`I;�fI;�kI;�oI;�rI;�tI;      ��I;ŝI;p�I;m�I;ّI;��I;ׂI;�yI;*pI;%fI;�[I;�QI;�GI;>I;�4I;9,I;�#I;�I;�I;�I;1
I;9I;� I;�H;��H;��H;@�H;-�H;a�H;��H;��H;��H;��H;"�H;��H;��H;c�H;��H;��H;"�H;��H;��H;��H;��H;a�H;-�H;@�H;��H;��H;�H;� I;9I;1
I;�I;�I;�I;�#I;9,I;�4I;>I;�GI;�QI;�[I;%fI;*pI;�yI;ׂI;��I;ّI;m�I;p�I;ŝI;      ��I;4�I;{�I;k�I;��I;��I;��I;��I;a�I;�I;k|I;�nI;uaI;�TI;�HI;n=I;�2I;W)I;� I;�I;�I;�I;MI;�I;t�H;��H;��H;M�H;8�H;a�H;��H;��H;��H;�H;��H;<�H;5�H;<�H;��H;�H;��H;��H;��H;a�H;8�H;M�H;��H;��H;t�H;�I;MI;�I;�I;�I;� I;W)I;�2I;n=I;�HI;�TI;uaI;�nI;k|I;�I;a�I;��I;��I;��I;��I;k�I;{�I;4�I;      ��I;�I;��I;��I;L�I;?�I; �I;��I;:�I;��I;�I;��I;��I;!rI;+bI;SSI;�EI;z9I;M.I;L$I;vI;�I;I;*I;I;��H;2�H;�H;M�H;-�H;e�H;��H;��H;�H;b�H;	�H;��H;	�H;b�H;�H;��H;��H;e�H;-�H;M�H;�H;2�H;��H;I;*I;I;�I;vI;L$I;M.I;z9I;�EI;SSI;+bI;!rI;��I;��I;�I;��I;:�I;��I; �I;?�I;L�I;��I;��I;�I;      s�H;.I;XI;[6I;
YI;�|I;)�I;&�I;1�I;��I;��I;��I;��I;��I;%�I;�oI;�]I;�MI;q?I;�2I;}'I;�I;8I;�I;�I;ZI;��H;2�H;��H;@�H;1�H;s�H;&�H;#�H;��H;�H;��H;�H;��H;#�H;&�H;s�H;1�H;@�H;��H;2�H;��H;ZI;�I;�I;8I;�I;}'I;�2I;q?I;�MI;�]I;�oI;%�I;��I;��I;��I;��I;��I;1�I;&�I;)�I;�|I;
YI;[6I;XI;.I;      uF;��F;�F;� G;}�G;,H;ȄH;9�H;VJI;B�I;��I;�I;��I;	�I;�I;e�I;C|I;ZgI;�TI;yDI;e6I;�)I;FI;+I;tI;�I;ZI;��H;��H;��H;6�H;I�H;��H;j�H;��H;$�H;��H;$�H;��H;j�H;��H;I�H;6�H;��H;��H;��H;ZI;�I;tI;+I;FI;�)I;e6I;yDI;�TI;ZgI;C|I;e�I;�I;	�I;��I;�I;��I;B�I;VJI;9�H;ȄH;,H;}�G;� G;�F;��F;      ��?;@;@�@;@�A;۸B;�C;BBE;�uF;�G;�[H;��H;�lI;��I;"�I;@�I;ɺI;��I;|�I;�oI;tZI;aHI;�8I;+I; I;�I;tI;�I;I;t�H;��H;��H;;�H;d�H;��H;��H;f�H;=�H;f�H;��H;��H;d�H;;�H;��H;��H;t�H;I;�I;tI;�I; I;+I;�8I;aHI;tZI;�oI;|�I;��I;ɺI;@�I;"�I;��I;�lI;��H;�[H;�G;�uF;BBE;�C;۸B;@�A;@�@;@;      U�1;��1;�63;�15;��7;��:;H{=;;P@;r�B;bE;��F;uH;�H;;pI;�I;��I;�I;)�I;m�I;�uI;�^I;�JI;4:I;�+I; I;+I;�I;*I;�I;�H;��H;~�H;4�H;��H;{�H;��H;��H;��H;{�H;��H;4�H;~�H;��H;�H;�I;*I;�I;+I; I;�+I;4:I;�JI;�^I;�uI;m�I;)�I;�I;��I;�I;;pI;�H;uH;��F;bE;r�B;;P@;H{=;��:;��7;�15;�63;��1;      ��;��;>\;VW;�m!;�7';�H-; 93;̳8;3{=;)kA;iyD;��F;/H;�I;�I;��I;��I;��I;��I;�yI;�`I;�KI;4:I;+I;FI;8I;I;MI;� I;��H;�H;w�H;�H;�H;a�H;2�H;a�H;�H;�H;w�H;�H;��H;� I;MI;I;8I;FI;+I;4:I;�KI;�`I;�yI;��I;��I;��I;��I;�I;�I;/H;��F;iyD;)kA;3{=;̳8; 93;�H-;�7';�m!;VW;>\;��;      �m�:���:_I�:�W�:���:-�;�~;�;¾$;�F.;*O6;��<;K�A;�
E;)RG;<�H;6lI;��I;d�I;m�I;ԙI;�zI;�`I;�JI;�8I;�)I;�I;�I;�I;9I; I;�H;��H;{�H; �H;�H;��H;�H; �H;{�H;��H;�H; I;9I;�I;�I;�I;�)I;�8I;�JI;�`I;�zI;ԙI;m�I;d�I;��I;6lI;<�H;)RG;�
E;K�A;��<;*O6;�F.;¾$;�;�~;-�;���:�W�:_I�:���:      �l8��8�Pu9̨�9��9:#��:�U�:cp�:T� ;F;Nn!;��-;^7;kk>;NC;�tF;nPH;�HI;ֳI;��I;кI;ԙI;�yI;�^I;aHI;e6I;}'I;vI;�I;1
I;�I;>�H;��H;��H;�H;��H;��H;��H;�H;��H;��H;>�H;�I;1
I;�I;vI;}'I;e6I;aHI;�^I;�yI;ԙI;кI;��I;ֳI;�HI;nPH;�tF;NC;kk>;^7;��-;Nn!;F;T� ;cp�:�U�:#��:��9:̨�9�Pu9��8      �����oj�V�غ9����*�����P��9c�:d��:���:�.;��$;��1;3f;;��A;��E;H;Q4I;X�I;��I;m�I;��I;�uI;tZI;yDI;�2I;L$I;�I;�I;hI;�I;��H;t�H;7�H;��H;��H;��H;7�H;t�H;��H;�I;hI;�I;�I;L$I;�2I;yDI;tZI;�uI;��I;m�I;��I;X�I;Q4I;H;��E;��A;3f;;��1;��$;�.;���:d��:c�:P��9�����*�9���V�غoj���      8�ͻ�ɻ��� e��1��J�]��!��轺����0�9���:MR�:�;�X;1H-;�9;v�@;�[E;��G;Q4I;ֳI;d�I;��I;m�I;�oI;�TI;q?I;M.I;� I;�I;ZI;�I;�I;6�H;��H;,�H;��H;,�H;��H;6�H;�I;�I;ZI;�I;� I;M.I;q?I;�TI;�oI;m�I;��I;d�I;ֳI;Q4I;��G;�[E;v�@;�9;1H-;�X;�;MR�:���:�0�9����轺�!�J�]�1�� e������ɻ      jO�$�K��o@�%�.�Ǩ����Gɻ�H��mpE���غ0����9o�:�@�:�;�*;��7;�O@;�[E;H;�HI;��I;��I;)�I;|�I;ZgI;�MI;z9I;W)I;�I;�I;�
I;,I;'I;G�H;s�H;��H;s�H;G�H;'I;,I;�
I;�I;�I;W)I;z9I;�MI;ZgI;|�I;)�I;��I;��I;�HI;H;�[E;�O@;��7;�*;�;�@�:o�:��90����غmpE��H��Gɻ���Ǩ�%�.��o@�$�K�      @L�����R���`����N��WPp�!D�ʨ��G�_���34�:���)�n8��:_�:ZF;�(;��7;v�@;��E;nPH;6lI;��I;�I;��I;C|I;�]I;�EI;�2I;�#I;{I;�I;		I;(I;� I;�H;h�H;�H;� I;(I;		I;�I;{I;�#I;�2I;�EI;�]I;C|I;��I;�I;��I;6lI;nPH;��E;v�@;��7;�(;ZF;_�:��:)�n8:���34�_����G�ʨ�!D�WPp��N��`���R������      ��7�d5���������ϼ��@X���iO����-ɻ��p�yF�e�o��g:^�:ZF;�*;�9;��A;�tF;<�H;�I;��I;ɺI;e�I;�oI;SSI;n=I;9,I;�I;�I;I;pI;�I;�I;� I;�I;�I;pI;I;�I;�I;9,I;n=I;SSI;�oI;e�I;ɺI;��I;�I;<�H;�tF;��A;�9;�*;ZF;^�:�g:e�o�yF⺙�p�-ɻ����iO�@X������ϼ������d5�7�      r��ٷ��40v���a�3�G�P2+�!�����*���0���5��ﻦ��\g��ହ�g:_�:�;1H-;3f;;NC;)RG;�I;�I;@�I;�I;%�I;+bI;�HI;�4I;�%I;�I;PI;�
I;�I;eI;sI;eI;�I;�
I;PI;�I;�%I;�4I;�HI;+bI;%�I;�I;@�I;�I;�I;)RG;NC;3f;;1H-;�;_�:�g:�ହ\g�������5�0��*������!��P2+�3�G���a�40v�ٷ��      ��ս��ѽC�ƽ8����I��$���a�a�'D4�LM���ϼ9����K�����G��\g�e�o���:�@�:�X;��1;kk>;�
E;/H;;pI;"�I;	�I;��I;!rI;�TI;>I;�,I;~I;�I;�I;�	I;/I;MI;/I;�	I;�I;�I;~I;�,I;>I;�TI;!rI;��I;	�I;"�I;;pI;/H;�
E;kk>;��1;�X;�@�:��:e�o�\g��G�������K�9����ϼLM�'D4�a�a�$����I��8���C�ƽ��ѽ      �L+� (���H�������ս�@���%���;V�5���������MS�������yF�)�n8o�:�;��$;^7;K�A;��F;�H;��I;��I;��I;��I;uaI;�GI;.4I;A%I;II;ZI;I;�	I; 	I;�	I;I;ZI;II;A%I;.4I;�GI;uaI;��I;��I;��I;��I;�H;��F;K�A;^7;��$;�;o�:)�n8yF⺦������MS�������5���;V��%���@����ս����H��� (�      �T��f�����z� Zb�(�D��$�����ѽ�I��S�m�!2+��������K��ﻙ�p�:�����9MR�:�.;��-;��<;iyD;uH;�lI;�I;��I;��I;�nI;�QI;�;I;!+I;�I;*I;OI;�I;�I;�I;OI;*I;�I;!+I;�;I;�QI;�nI;��I;��I;�I;�lI;uH;iyD;��<;��-;�.;MR�:��9:�����p��ﻍ�K������!2+�S�m��I����ѽ���$�(�D� Zb���z�f���      >�׾��Ҿž�j��������z�U�H�+��lz�N$��0v�!2+����9���5�-ɻ34�0�����:���:Nn!;*O6;)kA;��F;��H;��I;��I;�I;k|I;�[I;~CI;%1I;�#I;�I;jI;�I;�I;�I;jI;�I;�#I;%1I;~CI;�[I;k|I;�I;��I;��I;��H;��F;)kA;*O6;Nn!;���:���:0��34�-ɻ�5�9�����!2+�0v�N$��lz�+��U�H���z������j��ž��Ҿ      E(��$�b��O������~���`���Yb���'��U�N$��S�m�5����ϼ0�����_�����غ�0�9d��:F;�F.;3{=;bE;�[H;B�I;��I;��I;�I;%fI;&KI;7I;&(I;�I;�I;�I;DI;�I;�I;�I;&(I;7I;&KI;%fI;�I;��I;��I;B�I;�[H;bE;3{=;�F.;F;d��:�0�9��غ_������0����ϼ5��S�m�N$���U���'��Yb��`���~�����O��b���$�      7�}���w�#f���K�o,�{�
�:�׾�����k���'�lz꽥I���;V�LM�*����iO��G�mpE����c�:T� ;¾$;̳8;r�B;�G;VJI;1�I;:�I;a�I;*pI;�RI;�<I;�,I;%!I;�I;9I;�I;9I;�I;%!I;�,I;�<I;�RI;*pI;a�I;:�I;1�I;VJI;�G;r�B;̳8;¾$;T� ;c�:���mpE��G��iO�*���LM��;V��I��lz���'���k����:�׾{�
�o,���K�#f���w�      ~�n�������,蒿��w���F�b��Ȱ�����Yb�+����ѽ�%��'D4����@X��ʨ��H���轺P��9cp�:�; 93;;P@;�uF;9�H;&�I;��I;��I;�yI;�YI;3BI;�0I;�$I;eI;�I;@I;�I;eI;�$I;�0I;3BI;�YI;�yI;��I;��I;&�I;9�H;�uF;;P@; 93;�;cp�:P��9�轺�H��ʨ�@X�����'D4��%����ѽ+���Yb����Ȱ�b����F���w�,蒿����n���      .���������㿆�ɿ���ǅ����P�b��:�׾�`��U�H����@��a�a�!����!D�Gɻ�!������U�:�~;�H-;H{=;BBE;ȄH;)�I; �I;��I;ׂI;�`I;BGI;�4I;�'I;�I;I;pI;I;�I;�'I;�4I;BGI;�`I;ׂI;��I; �I;)�I;ȄH;BBE;H{=;�H-;�~;�U�:�����!�Gɻ!D���!��a�a��@����U�H��`��:�׾b����P�ǅ�������ɿ��㿯���      Ù$��x � ��7���޿m���ǅ����F�{�
��~����z��$���ս$���P2+���ϼWPp����J�]��*�#��:-�;�7';��:;�C;,H;�|I;?�I;��I;��I;�fI;�KI;:8I;V*I;E!I;I;GI;I;E!I;V*I;:8I;�KI;�fI;��I;��I;?�I;�|I;,H;�C;��:;�7';-�;#��:�*�J�]����WPp���ϼP2+�$�����ս�$���z��~��{�
���F�ǅ��m����޿7�� ���x �      F�Q��K���;�Ù$��;
��޿�����w�o,���澝���(�D������I��3�G�����N��Ǩ�1��9�����9:���:�m!;��7;۸B;}�G;
YI;L�I;��I;ّI;�kI;�OI;4;I;�,I;3#I;�I;�I;�I;3#I;�,I;4;I;�OI;�kI;ّI;��I;L�I;
YI;}�G;۸B;��7;�m!;���:��9:9���1��Ǩ��N�����3�G��I������(�D��������o,���w�����޿�;
�Ù$���;��K�      Q����{���d��F�Ù$�7����ɿ,蒿��K�O���j�� Zb�H�8�����a����`���%�.� e��V�غ̨�9�W�:VW;�15;@�A;� G;[6I;��I;k�I;m�I;�oI;�RI;�=I;�.I;�$I;AI;OI;AI;�$I;�.I;�=I;�RI;�oI;m�I;k�I;��I;[6I;� G;@�A;�15;VW;�W�:̨�9V�غ e��%�.�`��������a�8���H� Zb��j��O����K�,蒿��ɿ7��Ù$��F���d��{�      ���� P�������d���;� ����㿰���#f�b��ž��z���C�ƽ40v�d5�R����o@����oj��Pu9_I�:>\;�63;@�@;�F;XI;��I;{�I;p�I;�rI;�TI;^?I;0I;&I;, I;MI;, I;&I;0I;^?I;�TI;�rI;p�I;{�I;��I;XI;�F;@�@;�63;>\;_I�:�Pu9oj�����o@�R���d5�40v�C�ƽ����z�žb��#f�������� ����;���d���� P��      �,��^�� P���{��K��x �����n�����w��$���Ҿf��� (���ѽٷ��7����$�K��ɻ����8���:��;��1;@;��F;.I;�I;4�I;ŝI;�tI;OVI;�@I;�0I;�&I;� I;�I;� I;�&I;�0I;�@I;OVI;�tI;ŝI;4�I;�I;.I;��F;@;��1;��;���:��8���ɻ$�K����7�ٷ����ѽ (�f�����Ҿ�$���w�n��������x ��K��{� P��^��      A(��o'���o��L�d��X1�|x�Ŀ����3�v���x����4�s��b+���'�"�ü�yY�llٻq&�<�p�Y��:_;��0;��?;�F;tI;�I;��I;H�I;��I;ucI;�JI;�8I;�-I;�&I;�$I;�&I;�-I;�8I;�JI;ucI;��I;H�I;��I;�I;tI;�F;��?;��0;_;Y��:<�p�q&�llٻ�yY�"�ü�'�b+��s����4��x��v���3����Ŀ|x��X1�d�L��o��o'��      o'���X��c^�������]]���,�N9�3g��S�����/����o��j1��hܽ���-$��l��,}U��Ի~!�{�-���:;�41;��?;m�F;N&I;��I;7�I;Z�I;ąI;�bI;]JI;�8I;E-I;�&I;�$I;�&I;E-I;�8I;]JI;�bI;ąI;Z�I;7�I;��I;N&I;m�F;��?;�41;;��:{�-�~!��Ի,}U��l���-$����hܽj1��o���྘�/�S���3g��N9���,��]]�����c^���X��      �o��c^���ē��4z�1K�e��M��$ﱿQ�v��X#���Ѿń�	�&�w�нk̀�r��������I� ǻ�5��9�
�:X�;!�2;��@;�F;:I;�I;�I;��I;��I;qaI;II;�7I;~,I;�%I;�#I;�%I;~,I;�7I;II;qaI;��I;��I;�I;�I;:I;�F;��@;!�2;X�;�
�:�9�5� ǻ��I�����r��k̀�w�н	�&�ń���Ѿ�X#�Q�v�$ﱿM��e��1K��4z��ē�c^��      L������4z���V��X1��<�pؿ����RZ��	�(���KUo����fy��?l�l�S����7������𺧽�9��:��;]�4;�sA;�1G;�WI;��I;r�I;)�I;�I;�^I;GI;A6I;+I;�$I;�"I;�$I;+I;A6I;GI;�^I;�I;)�I;r�I;��I;�WI;�1G;�sA;]�4;��;��:���9�𺘼����7�S��l�?l�fy�����KUo�(����	��RZ����pؿ�<��X1���V��4z�����      d��]]�1K��X1�Xf���kQ��R���Z58��A���נ���O���h什�Q�,���cߓ��� �W��{谺�":��:$ ;�/7; �B;`�G;{I;�I;��I;զI;]{I;Z[I;hDI;<4I;X)I;R#I;G!I;R#I;X)I;<4I;hDI;Z[I;]{I;զI;��I;�I;{I;`�G; �B;�/7;$ ;��:�":{谺W���� �cߓ�,����Q�h什����O��נ��A��Z58�R���kQ����Xf��X1�1K��]]�      �X1���,�e���<���2g��c_���U�˂�ՌȾ	ń�-�-�q��Y ��8�2�.?ټ��{�G"��n��O���u:�O ;�&;6":;[�C;!%H;1�I;D�I;��I;�I;�uI;�VI;AI;�1I;3'I;c!I;}I;c!I;3'I;�1I;AI;�VI;�uI;�I;��I;D�I;1�I;!%H;[�C;6":;�&;�O ;��u:�O��n�G"���{�.?ټ8�2�Y ��q��-�-�	ń�ՌȾ˂��U�c_��2g���<�e����,�      |x�N9�M��pؿkQ��c_��4�_��X#�p���f��<�S�{�����-l�T�-w��e�M�"�Ի��+��LT���:�d;�[,;	/=;�AE;|�H;��I;��I;��I;֕I;�nI;�QI;/=I;|.I;�$I;I;cI;I;�$I;|.I;/=I;�QI;�nI;֕I;��I;��I;��I;|�H;�AE;	/=;�[,;�d;��:�LT���+�"�Իe�M�-w��T�-l�����{�<�S��f��p���X#�4�_�c_��kQ��pؿM��N9�      Ŀ3g��$ﱿ���R����U��X#�r��d���JUo�
�#��hܽ����n<����_���҉ �;❻I�Ժ�l�9s��:�U;�2;�@;t�F;�I;�I;b�I;K�I;��I;%gI;.LI;�8I;+I;�!I;�I;�I;�I;�!I;+I;�8I;.LI;%gI;��I;K�I;b�I;�I;�I;t�F;�@;�2;�U;s��:�l�9I�Ժ;❻҉ �_�������n<�����hܽ
�#�JUo�d���r���X#��U�R������$ﱿ3g��      ���S���Q�v��RZ�Z58�˂�p��d���hoy�`1�gO��d什�`�`��6����yY���컞�T��1���u:��:\~#;.88;�B;��G;lI;-�I;"�I;L�I;��I;�^I;!FI;4I;C'I;�I;�I;)I;�I;�I;C'I;4I;!FI;�^I;��I;L�I;"�I;-�I;lI;��G;�B;.88;\~#;��:��u:�1���T���컶yY�6���`���`�d什gO��`1�hoy�d���p��˂�Z58��RZ�Q�v�S���      �3���/��X#��	��A��ՌȾ�f��JUo�`1�Ӱ���n���x��'��>ټ�@��-l�S���$��'�39�!�:;Q;!d-;�.=;�E;wH;��I;-�I;��I; �I;6uI;�VI;�?I;/I;B#I;_I;�I;TI;�I;_I;B#I;/I;�?I;�VI;6uI; �I;��I;-�I;��I;wH;�E;�.=;!d-;;Q;�!�:'�39$��S���-l��@���>ټ�'��x��n��Ӱ��`1�JUo��f��ՌȾ�A���	��X#���/�      v���ྃ�Ѿ(����נ�	ń�<�S�
�#�gO���n��R̀��2�,������>���Ի��B��#�\m:�E�:o ;��5;�EA;��F;�I;r�I;p�I;ŽI;��I;�iI;�MI;.9I;�)I;I;�I;�I;iI;�I;�I;I;�)I;.9I;�MI;�iI;��I;ŽI;p�I;r�I;�I;��F;�EA;��5;o ;�E�:\m:�#���B���Ի��>���,���2�R̀��n��gO��
�#�<�S�	ń��נ�(�����Ѿ��      �x���o��ń�KUo���O�-�-�{��hܽd什�x��2��b��yR���|U��2�����"찺�m�9��:C;��,;�g<;�qD;h$H;�I;��I;��I;&�I;&I;�]I;(EI;r2I;�$I;�I;}I;�I;QI;�I;}I;�I;�$I;r2I;(EI;�]I;&I;&�I;��I;��I;�I;h$H;�qD;�g<;��,;C;��:�m�9"찺����2���|U�yR���b���2��x�d什�hܽ{�-�-���O�KUo�ń��o��      ��4�j1�	�&������q�ཌྷ�������`��'�,��yR����]�����V��[��o�o����:{�;=~#;0�6;nsA;s�F;�I;��I;��I;��I;6�I;�oI;�RI;�<I;�+I;�I;�I;�I;`I;WI;`I;�I;�I;�I;�+I;�<I;�RI;�oI;6�I;��I;��I;��I;�I;s�F;nsA;0�6;=~#;{�;���:o�o�[���V�������]�yR��,��'��`��������q�������	�&�j1�      s�ཾhܽw�нfy��h什Y ��-l��n<�`���>ټ�𛼝|U����H᝻�2�������u:jj�:�;}61;j(>;sE;,IH;p�I;��I;��I;�I;��I;zaI;�GI;G4I;~%I;�I;�I;XI;=
I;7	I;=
I;XI;�I;�I;~%I;G4I;�GI;zaI;��I;�I;��I;��I;p�I;,IH;sE;j(>;}61;�;jj�:��u:�����2�H᝻����|U����>ټ`���n<�-l�Y ��h什fy��w�н�hܽ      b+����k̀�?l��Q�8�2�T����6����@����>��2���V���2����	 R:���:�;�[,;P;;;C;�dG;w8I;��I;U�I;��I;_�I;�pI;�SI;=I;W,I;KI;�I;�I;�	I;+I;'I;+I;�	I;�I;�I;KI;W,I;=I;�SI;�pI;_�I;��I;U�I;��I;w8I;�dG;;C;P;;�[,;�;���:	 R:���2��V���2����>��@��6������T�8�2��Q�?l�k̀���      �'��-$�r��l�,���.?ټ-w��_����yY�-l���Ի���[������	 R:���:�Q;�);��8;��A;�F;S�H;J�I;��I;��I;ɨI;$�I;�_I;GI;�3I;�$I;cI;�I;�
I;�I;*I;]I;*I;�I;�
I;�I;cI;�$I;�3I;GI;�_I;$�I;ɨI;��I;��I;J�I;S�H;�F;��A;��8;�);�Q;���:	 R:����[�������Ի-l��yY�_���-w��.?ټ,���l�r���-$�      "�ü�l������S��cߓ���{�e�M�҉ ����S�����B�"찺o�o���u:���:�Q;E�';)07;ք@;�E;�kH;N�I;��I;��I;,�I;��I;�kI;�PI;D;I;�*I;�I;�I;|I;�I;[I;CI;� I;CI;[I;�I;|I;�I;�I;�*I;D;I;�PI;�kI;��I;,�I;��I;��I;N�I;�kH;�E;ք@;)07;E�';�Q;���:��u:o�o�"찺��B�S������҉ �e�M���{�cߓ�S�������l��      �yY�,}U���I���7��� �G"�"�Ի;❻��T�$���#��m�9���:jj�:�;�);)07;D@;V\E;�#H;�jI;(�I;s�I;�I;M�I;�vI;�YI;�BI;�0I;g"I;DI;�I;EI;�I;N I;�H;�H;�H;N I;�I;EI;�I;DI;g"I;�0I;�BI;�YI;�vI;M�I;�I;s�I;(�I;�jI;�#H;V\E;D@;)07;�);�;jj�:���:�m�9�#�$���T�;❻"�ԻG"��� ���7���I�,}U�      llٻ�Ի ǻ����W���n���+�I�Ժ�1�'�39\m:��:{�;�;�[,;��8;ք@;V\E;�	H;jUI;��I;	�I;�I;}�I;#�I;�aI;}II;>6I;�&I;�I;GI;�	I;OI;O I;{�H;��H;��H;��H;{�H;O I;OI;�	I;GI;�I;�&I;>6I;}II;�aI;#�I;}�I;�I;	�I;��I;jUI;�	H;V\E;ք@;��8;�[,;�;{�;��:\m:'�39�1�I�Ժ��+��n�W������ ǻ�Ի      q&�~!��5���{谺�O��LT��l�9��u:�!�:�E�:C;=~#;}61;P;;��A;�E;�#H;jUI;,�I;��I;1�I;��I;�I;-hI;COI;7;I;+I;3I;�I;�I;�I;� I;F�H;��H;��H;�H;��H;��H;F�H;� I;�I;�I;�I;3I;+I;7;I;COI;-hI;�I;��I;1�I;��I;,�I;jUI;�#H;�E;��A;P;;}61;=~#;C;�E�:�!�:��u:�l�9�LT��O�{谺���5�~!�      <�p�{�-��9���9�":��u:��:s��:��:;Q;o ;��,;0�6;j(>;;C;�F;�kH;�jI;��I;��I;��I;4�I;��I;�lI;�SI;??I;�.I;8!I;nI;�I;�I;�I;��H;��H;��H;c�H;��H;c�H;��H;��H;��H;�I;�I;�I;nI;8!I;�.I;??I;�SI;�lI;��I;4�I;��I;��I;��I;�jI;�kH;�F;;C;j(>;0�6;��,;o ;;Q;��:s��:��:��u:�":���9�9{�-�      Y��:��:�
�:��:��:�O ;�d;�U;\~#;!d-;��5;�g<;nsA;sE;�dG;S�H;N�I;(�I;	�I;1�I;4�I;�I;"oI;aVI;BI;X1I;�#I;�I;�I;VI;�I;�H;��H;�H;f�H;?�H;��H;?�H;f�H;�H;��H;�H;�I;VI;�I;�I;�#I;X1I;BI;aVI;"oI;�I;4�I;1�I;	�I;(�I;N�I;S�H;�dG;sE;nsA;�g<;��5;!d-;\~#;�U;�d;�O ;��:��:�
�:��:      _;;X�;��;$ ;�&;�[,;�2;.88;�.=;�EA;�qD;s�F;,IH;w8I;J�I;��I;s�I;�I;��I;��I;"oI;bWI;�CI;3I;s%I;8I;�I;�	I;�I;��H;��H;��H;��H;H�H;V�H;�H;V�H;H�H;��H;��H;��H;��H;�I;�	I;�I;8I;s%I;3I;�CI;bWI;"oI;��I;��I;�I;s�I;��I;J�I;w8I;,IH;s�F;�qD;�EA;�.=;.88;�2;�[,;�&;$ ;��;X�;;      ��0;�41;!�2;]�4;�/7;6":;	/=;�@;�B;�E;��F;h$H;�I;p�I;��I;��I;��I;�I;}�I;�I;�lI;aVI;�CI;�3I;Y&I;EI;I;�
I;II;>�H;A�H;��H;��H;��H;p�H;��H;w�H;��H;p�H;��H;��H;��H;A�H;>�H;II;�
I;I;EI;Y&I;�3I;�CI;aVI;�lI;�I;}�I;�I;��I;��I;��I;p�I;�I;h$H;��F;�E;�B;�@;	/=;6":;�/7;]�4;!�2;�41;      ��?;��?;��@;�sA; �B;[�C;�AE;t�F;��G;wH;�I;�I;��I;��I;U�I;��I;,�I;M�I;#�I;-hI;�SI;BI;3I;Y&I;�I;�I;)I;�I;��H;��H;&�H;z�H;p�H;��H;��H;5�H;�H;5�H;��H;��H;p�H;z�H;&�H;��H;��H;�I;)I;�I;�I;Y&I;3I;BI;�SI;-hI;#�I;M�I;,�I;��I;U�I;��I;��I;�I;�I;wH;��G;t�F;�AE;[�C; �B;�sA;��@;��?;      �F;m�F;�F;�1G;`�G;!%H;|�H;�I;lI;��I;r�I;��I;��I;��I;��I;ɨI;��I;�vI;�aI;COI;??I;X1I;s%I;EI;�I;OI;1I; I;��H;U�H;��H;c�H;��H;4�H;e�H;��H;��H;��H;e�H;4�H;��H;c�H;��H;U�H;��H; I;1I;OI;�I;EI;s%I;X1I;??I;COI;�aI;�vI;��I;ɨI;��I;��I;��I;��I;r�I;��I;lI;�I;|�H;!%H;`�G;�1G;�F;m�F;      tI;N&I;:I;�WI;{I;1�I;��I;�I;-�I;-�I;p�I;��I;��I;�I;_�I;$�I;�kI;�YI;}II;7;I;�.I;�#I;8I;I;)I;1I; I;��H;~�H;��H;\�H;a�H;��H;��H;�H;��H;w�H;��H;�H;��H;��H;a�H;\�H;��H;~�H;��H; I;1I;)I;I;8I;�#I;�.I;7;I;}II;�YI;�kI;$�I;_�I;�I;��I;��I;p�I;-�I;-�I;�I;��I;1�I;{I;�WI;:I;N&I;      �I;��I;�I;��I;�I;D�I;��I;b�I;"�I;��I;ŽI;&�I;6�I;��I;�pI;�_I;�PI;�BI;>6I;+I;8!I;�I;�I;�
I;�I; I;��H;y�H;��H;c�H;a�H;��H;��H;��H;��H;��H;y�H;��H;��H;��H;��H;��H;a�H;c�H;��H;y�H;��H; I;�I;�
I;�I;�I;8!I;+I;>6I;�BI;�PI;�_I;�pI;��I;6�I;&�I;ŽI;��I;"�I;b�I;��I;D�I;�I;��I;�I;��I;      ��I;7�I;�I;r�I;��I;��I;��I;K�I;L�I; �I;��I;&I;�oI;zaI;�SI;GI;D;I;�0I;�&I;3I;nI;�I;�	I;II;��H;��H;~�H;��H;X�H;[�H;��H;Z�H;L�H;��H;��H;��H;��H;��H;��H;��H;L�H;Z�H;��H;[�H;X�H;��H;~�H;��H;��H;II;�	I;�I;nI;3I;�&I;�0I;D;I;GI;�SI;zaI;�oI;&I;��I; �I;L�I;K�I;��I;��I;��I;r�I;�I;7�I;      H�I;Z�I;��I;)�I;զI;�I;֕I;��I;��I;6uI;�iI;�]I;�RI;�GI;=I;�3I;�*I;g"I;�I;�I;�I;VI;�I;>�H;��H;U�H;��H;c�H;[�H;��H;6�H;�H;B�H;��H;�H;��H;��H;��H;�H;��H;B�H;�H;6�H;��H;[�H;c�H;��H;U�H;��H;>�H;�I;VI;�I;�I;�I;g"I;�*I;�3I;=I;�GI;�RI;�]I;�iI;6uI;��I;��I;֕I;�I;զI;)�I;��I;Z�I;      ��I;ąI;��I;�I;]{I;�uI;�nI;%gI;�^I;�VI;�MI;(EI;�<I;G4I;W,I;�$I;�I;DI;GI;�I;�I;�I;��H;A�H;&�H;��H;\�H;a�H;��H;6�H;�H;�H;\�H;��H;z�H;7�H;��H;7�H;z�H;��H;\�H;�H;�H;6�H;��H;a�H;\�H;��H;&�H;A�H;��H;�I;�I;�I;GI;DI;�I;�$I;W,I;G4I;�<I;(EI;�MI;�VI;�^I;%gI;�nI;�uI;]{I;�I;��I;ąI;      ucI;�bI;qaI;�^I;Z[I;�VI;�QI;.LI;!FI;�?I;.9I;r2I;�+I;~%I;KI;cI;�I;�I;�	I;�I;�I;�H;��H;��H;z�H;c�H;a�H;��H;Z�H;�H;�H;U�H;��H;,�H;��H;��H;��H;��H;��H;,�H;��H;U�H;�H;�H;Z�H;��H;a�H;c�H;z�H;��H;��H;�H;�I;�I;�	I;�I;�I;cI;KI;~%I;�+I;r2I;.9I;�?I;!FI;.LI;�QI;�VI;Z[I;�^I;qaI;�bI;      �JI;]JI;II;GI;hDI;AI;/=I;�8I;4I;/I;�)I;�$I;�I;�I;�I;�I;|I;EI;OI;� I;��H;��H;��H;��H;p�H;��H;��H;��H;L�H;B�H;\�H;��H;�H;��H;M�H;!�H;3�H;!�H;M�H;��H;�H;��H;\�H;B�H;L�H;��H;��H;��H;p�H;��H;��H;��H;��H;� I;OI;EI;|I;�I;�I;�I;�I;�$I;�)I;/I;4I;�8I;/=I;AI;hDI;GI;II;]JI;      �8I;�8I;�7I;A6I;<4I;�1I;|.I;+I;C'I;B#I;I;�I;�I;�I;�I;�
I;�I;�I;O I;F�H;��H;�H;��H;��H;��H;4�H;��H;��H;��H;��H;��H;,�H;��H;<�H;��H;��H;��H;��H;��H;<�H;��H;,�H;��H;��H;��H;��H;��H;4�H;��H;��H;��H;�H;��H;F�H;O I;�I;�I;�
I;�I;�I;�I;�I;I;B#I;C'I;+I;|.I;�1I;<4I;A6I;�7I;�8I;      �-I;E-I;~,I;+I;X)I;3'I;�$I;�!I;�I;_I;�I;}I;�I;XI;�	I;�I;[I;N I;{�H;��H;��H;f�H;H�H;p�H;��H;e�H;�H;��H;��H;�H;z�H;��H;M�H;��H;��H;��H;�H;��H;��H;��H;M�H;��H;z�H;�H;��H;��H;�H;e�H;��H;p�H;H�H;f�H;��H;��H;{�H;N I;[I;�I;�	I;XI;�I;}I;�I;_I;�I;�!I;�$I;3'I;X)I;+I;~,I;E-I;      �&I;�&I;�%I;�$I;R#I;c!I;I;�I;�I;�I;�I;�I;`I;=
I;+I;*I;CI;�H;��H;��H;c�H;?�H;V�H;��H;5�H;��H;��H;��H;��H;��H;7�H;��H;!�H;��H;��H;k�H;r�H;k�H;��H;��H;!�H;��H;7�H;��H;��H;��H;��H;��H;5�H;��H;V�H;?�H;c�H;��H;��H;�H;CI;*I;+I;=
I;`I;�I;�I;�I;�I;�I;I;c!I;R#I;�$I;�%I;�&I;      �$I;�$I;�#I;�"I;G!I;}I;cI;�I;)I;TI;iI;QI;WI;7	I;'I;]I;� I;�H;��H;�H;��H;��H;�H;w�H;�H;��H;w�H;y�H;��H;��H;��H;��H;3�H;��H;�H;r�H;w�H;r�H;�H;��H;3�H;��H;��H;��H;��H;y�H;w�H;��H;�H;w�H;�H;��H;��H;�H;��H;�H;� I;]I;'I;7	I;WI;QI;iI;TI;)I;�I;cI;}I;G!I;�"I;�#I;�$I;      �&I;�&I;�%I;�$I;R#I;c!I;I;�I;�I;�I;�I;�I;`I;=
I;+I;*I;CI;�H;��H;��H;c�H;?�H;V�H;��H;5�H;��H;��H;��H;��H;��H;7�H;��H;!�H;��H;��H;k�H;r�H;k�H;��H;��H;!�H;��H;7�H;��H;��H;��H;��H;��H;5�H;��H;V�H;?�H;c�H;��H;��H;�H;CI;*I;+I;=
I;`I;�I;�I;�I;�I;�I;I;c!I;R#I;�$I;�%I;�&I;      �-I;E-I;~,I;+I;X)I;3'I;�$I;�!I;�I;_I;�I;}I;�I;XI;�	I;�I;[I;N I;{�H;��H;��H;f�H;H�H;p�H;��H;e�H;�H;��H;��H;�H;z�H;��H;M�H;��H;��H;��H;�H;��H;��H;��H;M�H;��H;z�H;�H;��H;��H;�H;e�H;��H;p�H;H�H;f�H;��H;��H;{�H;N I;[I;�I;�	I;XI;�I;}I;�I;_I;�I;�!I;�$I;3'I;X)I;+I;~,I;E-I;      �8I;�8I;�7I;A6I;<4I;�1I;|.I;+I;C'I;B#I;I;�I;�I;�I;�I;�
I;�I;�I;O I;F�H;��H;�H;��H;��H;��H;4�H;��H;��H;��H;��H;��H;,�H;��H;<�H;��H;��H;��H;��H;��H;<�H;��H;,�H;��H;��H;��H;��H;��H;4�H;��H;��H;��H;�H;��H;F�H;O I;�I;�I;�
I;�I;�I;�I;�I;I;B#I;C'I;+I;|.I;�1I;<4I;A6I;�7I;�8I;      �JI;]JI;II;GI;hDI;AI;/=I;�8I;4I;/I;�)I;�$I;�I;�I;�I;�I;|I;EI;OI;� I;��H;��H;��H;��H;p�H;��H;��H;��H;L�H;B�H;\�H;��H;�H;��H;M�H;!�H;3�H;!�H;M�H;��H;�H;��H;\�H;B�H;L�H;��H;��H;��H;p�H;��H;��H;��H;��H;� I;OI;EI;|I;�I;�I;�I;�I;�$I;�)I;/I;4I;�8I;/=I;AI;hDI;GI;II;]JI;      ucI;�bI;qaI;�^I;Z[I;�VI;�QI;.LI;!FI;�?I;.9I;r2I;�+I;~%I;KI;cI;�I;�I;�	I;�I;�I;�H;��H;��H;z�H;c�H;a�H;��H;Z�H;�H;�H;U�H;��H;,�H;��H;��H;��H;��H;��H;,�H;��H;U�H;�H;�H;Z�H;��H;a�H;c�H;z�H;��H;��H;�H;�I;�I;�	I;�I;�I;cI;KI;~%I;�+I;r2I;.9I;�?I;!FI;.LI;�QI;�VI;Z[I;�^I;qaI;�bI;      ��I;ąI;��I;�I;]{I;�uI;�nI;%gI;�^I;�VI;�MI;(EI;�<I;G4I;W,I;�$I;�I;DI;GI;�I;�I;�I;��H;A�H;&�H;��H;\�H;a�H;��H;6�H;�H;�H;\�H;��H;z�H;7�H;��H;7�H;z�H;��H;\�H;�H;�H;6�H;��H;a�H;\�H;��H;&�H;A�H;��H;�I;�I;�I;GI;DI;�I;�$I;W,I;G4I;�<I;(EI;�MI;�VI;�^I;%gI;�nI;�uI;]{I;�I;��I;ąI;      H�I;Z�I;��I;)�I;զI;�I;֕I;��I;��I;6uI;�iI;�]I;�RI;�GI;=I;�3I;�*I;g"I;�I;�I;�I;VI;�I;>�H;��H;U�H;��H;c�H;[�H;��H;6�H;�H;B�H;��H;�H;��H;��H;��H;�H;��H;B�H;�H;6�H;��H;[�H;c�H;��H;U�H;��H;>�H;�I;VI;�I;�I;�I;g"I;�*I;�3I;=I;�GI;�RI;�]I;�iI;6uI;��I;��I;֕I;�I;զI;)�I;��I;Z�I;      ��I;7�I;�I;r�I;��I;��I;��I;K�I;L�I; �I;��I;&I;�oI;zaI;�SI;GI;D;I;�0I;�&I;3I;nI;�I;�	I;II;��H;��H;~�H;��H;X�H;[�H;��H;Z�H;L�H;��H;��H;��H;��H;��H;��H;��H;L�H;Z�H;��H;[�H;X�H;��H;~�H;��H;��H;II;�	I;�I;nI;3I;�&I;�0I;D;I;GI;�SI;zaI;�oI;&I;��I; �I;L�I;K�I;��I;��I;��I;r�I;�I;7�I;      �I;��I;�I;��I;�I;D�I;��I;b�I;"�I;��I;ŽI;&�I;6�I;��I;�pI;�_I;�PI;�BI;>6I;+I;8!I;�I;�I;�
I;�I; I;��H;y�H;��H;c�H;a�H;��H;��H;��H;��H;��H;y�H;��H;��H;��H;��H;��H;a�H;c�H;��H;y�H;��H; I;�I;�
I;�I;�I;8!I;+I;>6I;�BI;�PI;�_I;�pI;��I;6�I;&�I;ŽI;��I;"�I;b�I;��I;D�I;�I;��I;�I;��I;      tI;N&I;:I;�WI;{I;1�I;��I;�I;-�I;-�I;p�I;��I;��I;�I;_�I;$�I;�kI;�YI;}II;7;I;�.I;�#I;8I;I;)I;1I; I;��H;~�H;��H;\�H;a�H;��H;��H;�H;��H;w�H;��H;�H;��H;��H;a�H;\�H;��H;~�H;��H; I;1I;)I;I;8I;�#I;�.I;7;I;}II;�YI;�kI;$�I;_�I;�I;��I;��I;p�I;-�I;-�I;�I;��I;1�I;{I;�WI;:I;N&I;      �F;m�F;�F;�1G;`�G;!%H;|�H;�I;lI;��I;r�I;��I;��I;��I;��I;ɨI;��I;�vI;�aI;COI;??I;X1I;s%I;EI;�I;OI;1I; I;��H;U�H;��H;c�H;��H;4�H;e�H;��H;��H;��H;e�H;4�H;��H;c�H;��H;U�H;��H; I;1I;OI;�I;EI;s%I;X1I;??I;COI;�aI;�vI;��I;ɨI;��I;��I;��I;��I;r�I;��I;lI;�I;|�H;!%H;`�G;�1G;�F;m�F;      ��?;��?;��@;�sA; �B;[�C;�AE;t�F;��G;wH;�I;�I;��I;��I;U�I;��I;,�I;M�I;#�I;-hI;�SI;BI;3I;Y&I;�I;�I;)I;�I;��H;��H;&�H;z�H;p�H;��H;��H;5�H;�H;5�H;��H;��H;p�H;z�H;&�H;��H;��H;�I;)I;�I;�I;Y&I;3I;BI;�SI;-hI;#�I;M�I;,�I;��I;U�I;��I;��I;�I;�I;wH;��G;t�F;�AE;[�C; �B;�sA;��@;��?;      ��0;�41;!�2;]�4;�/7;6":;	/=;�@;�B;�E;��F;h$H;�I;p�I;��I;��I;��I;�I;}�I;�I;�lI;aVI;�CI;�3I;Y&I;EI;I;�
I;II;>�H;A�H;��H;��H;��H;p�H;��H;w�H;��H;p�H;��H;��H;��H;A�H;>�H;II;�
I;I;EI;Y&I;�3I;�CI;aVI;�lI;�I;}�I;�I;��I;��I;��I;p�I;�I;h$H;��F;�E;�B;�@;	/=;6":;�/7;]�4;!�2;�41;      _;;X�;��;$ ;�&;�[,;�2;.88;�.=;�EA;�qD;s�F;,IH;w8I;J�I;��I;s�I;�I;��I;��I;"oI;bWI;�CI;3I;s%I;8I;�I;�	I;�I;��H;��H;��H;��H;H�H;V�H;�H;V�H;H�H;��H;��H;��H;��H;�I;�	I;�I;8I;s%I;3I;�CI;bWI;"oI;��I;��I;�I;s�I;��I;J�I;w8I;,IH;s�F;�qD;�EA;�.=;.88;�2;�[,;�&;$ ;��;X�;;      Y��:��:�
�:��:��:�O ;�d;�U;\~#;!d-;��5;�g<;nsA;sE;�dG;S�H;N�I;(�I;	�I;1�I;4�I;�I;"oI;aVI;BI;X1I;�#I;�I;�I;VI;�I;�H;��H;�H;f�H;?�H;��H;?�H;f�H;�H;��H;�H;�I;VI;�I;�I;�#I;X1I;BI;aVI;"oI;�I;4�I;1�I;	�I;(�I;N�I;S�H;�dG;sE;nsA;�g<;��5;!d-;\~#;�U;�d;�O ;��:��:�
�:��:      <�p�{�-��9���9�":��u:��:s��:��:;Q;o ;��,;0�6;j(>;;C;�F;�kH;�jI;��I;��I;��I;4�I;��I;�lI;�SI;??I;�.I;8!I;nI;�I;�I;�I;��H;��H;��H;c�H;��H;c�H;��H;��H;��H;�I;�I;�I;nI;8!I;�.I;??I;�SI;�lI;��I;4�I;��I;��I;��I;�jI;�kH;�F;;C;j(>;0�6;��,;o ;;Q;��:s��:��:��u:�":���9�9{�-�      q&�~!��5���{谺�O��LT��l�9��u:�!�:�E�:C;=~#;}61;P;;��A;�E;�#H;jUI;,�I;��I;1�I;��I;�I;-hI;COI;7;I;+I;3I;�I;�I;�I;� I;F�H;��H;��H;�H;��H;��H;F�H;� I;�I;�I;�I;3I;+I;7;I;COI;-hI;�I;��I;1�I;��I;,�I;jUI;�#H;�E;��A;P;;}61;=~#;C;�E�:�!�:��u:�l�9�LT��O�{谺���5�~!�      llٻ�Ի ǻ����W���n���+�I�Ժ�1�'�39\m:��:{�;�;�[,;��8;ք@;V\E;�	H;jUI;��I;	�I;�I;}�I;#�I;�aI;}II;>6I;�&I;�I;GI;�	I;OI;O I;{�H;��H;��H;��H;{�H;O I;OI;�	I;GI;�I;�&I;>6I;}II;�aI;#�I;}�I;�I;	�I;��I;jUI;�	H;V\E;ք@;��8;�[,;�;{�;��:\m:'�39�1�I�Ժ��+��n�W������ ǻ�Ի      �yY�,}U���I���7��� �G"�"�Ի;❻��T�$���#��m�9���:jj�:�;�);)07;D@;V\E;�#H;�jI;(�I;s�I;�I;M�I;�vI;�YI;�BI;�0I;g"I;DI;�I;EI;�I;N I;�H;�H;�H;N I;�I;EI;�I;DI;g"I;�0I;�BI;�YI;�vI;M�I;�I;s�I;(�I;�jI;�#H;V\E;D@;)07;�);�;jj�:���:�m�9�#�$���T�;❻"�ԻG"��� ���7���I�,}U�      "�ü�l������S��cߓ���{�e�M�҉ ����S�����B�"찺o�o���u:���:�Q;E�';)07;ք@;�E;�kH;N�I;��I;��I;,�I;��I;�kI;�PI;D;I;�*I;�I;�I;|I;�I;[I;CI;� I;CI;[I;�I;|I;�I;�I;�*I;D;I;�PI;�kI;��I;,�I;��I;��I;N�I;�kH;�E;ք@;)07;E�';�Q;���:��u:o�o�"찺��B�S������҉ �e�M���{�cߓ�S�������l��      �'��-$�r��l�,���.?ټ-w��_����yY�-l���Ի���[������	 R:���:�Q;�);��8;��A;�F;S�H;J�I;��I;��I;ɨI;$�I;�_I;GI;�3I;�$I;cI;�I;�
I;�I;*I;]I;*I;�I;�
I;�I;cI;�$I;�3I;GI;�_I;$�I;ɨI;��I;��I;J�I;S�H;�F;��A;��8;�);�Q;���:	 R:����[�������Ի-l��yY�_���-w��.?ټ,���l�r���-$�      b+����k̀�?l��Q�8�2�T����6����@����>��2���V���2����	 R:���:�;�[,;P;;;C;�dG;w8I;��I;U�I;��I;_�I;�pI;�SI;=I;W,I;KI;�I;�I;�	I;+I;'I;+I;�	I;�I;�I;KI;W,I;=I;�SI;�pI;_�I;��I;U�I;��I;w8I;�dG;;C;P;;�[,;�;���:	 R:���2��V���2����>��@��6������T�8�2��Q�?l�k̀���      s�ཾhܽw�нfy��h什Y ��-l��n<�`���>ټ�𛼝|U����H᝻�2�������u:jj�:�;}61;j(>;sE;,IH;p�I;��I;��I;�I;��I;zaI;�GI;G4I;~%I;�I;�I;XI;=
I;7	I;=
I;XI;�I;�I;~%I;G4I;�GI;zaI;��I;�I;��I;��I;p�I;,IH;sE;j(>;}61;�;jj�:��u:�����2�H᝻����|U����>ټ`���n<�-l�Y ��h什fy��w�н�hܽ      ��4�j1�	�&������q�ཌྷ�������`��'�,��yR����]�����V��[��o�o����:{�;=~#;0�6;nsA;s�F;�I;��I;��I;��I;6�I;�oI;�RI;�<I;�+I;�I;�I;�I;`I;WI;`I;�I;�I;�I;�+I;�<I;�RI;�oI;6�I;��I;��I;��I;�I;s�F;nsA;0�6;=~#;{�;���:o�o�[���V�������]�yR��,��'��`��������q�������	�&�j1�      �x���o��ń�KUo���O�-�-�{��hܽd什�x��2��b��yR���|U��2�����"찺�m�9��:C;��,;�g<;�qD;h$H;�I;��I;��I;&�I;&I;�]I;(EI;r2I;�$I;�I;}I;�I;QI;�I;}I;�I;�$I;r2I;(EI;�]I;&I;&�I;��I;��I;�I;h$H;�qD;�g<;��,;C;��:�m�9"찺����2���|U�yR���b���2��x�d什�hܽ{�-�-���O�KUo�ń��o��      v���ྃ�Ѿ(����נ�	ń�<�S�
�#�gO���n��R̀��2�,������>���Ի��B��#�\m:�E�:o ;��5;�EA;��F;�I;r�I;p�I;ŽI;��I;�iI;�MI;.9I;�)I;I;�I;�I;iI;�I;�I;I;�)I;.9I;�MI;�iI;��I;ŽI;p�I;r�I;�I;��F;�EA;��5;o ;�E�:\m:�#���B���Ի��>���,���2�R̀��n��gO��
�#�<�S�	ń��נ�(�����Ѿ��      �3���/��X#��	��A��ՌȾ�f��JUo�`1�Ӱ���n���x��'��>ټ�@��-l�S���$��'�39�!�:;Q;!d-;�.=;�E;wH;��I;-�I;��I; �I;6uI;�VI;�?I;/I;B#I;_I;�I;TI;�I;_I;B#I;/I;�?I;�VI;6uI; �I;��I;-�I;��I;wH;�E;�.=;!d-;;Q;�!�:'�39$��S���-l��@���>ټ�'��x��n��Ӱ��`1�JUo��f��ՌȾ�A���	��X#���/�      ���S���Q�v��RZ�Z58�˂�p��d���hoy�`1�gO��d什�`�`��6����yY���컞�T��1���u:��:\~#;.88;�B;��G;lI;-�I;"�I;L�I;��I;�^I;!FI;4I;C'I;�I;�I;)I;�I;�I;C'I;4I;!FI;�^I;��I;L�I;"�I;-�I;lI;��G;�B;.88;\~#;��:��u:�1���T���컶yY�6���`���`�d什gO��`1�hoy�d���p��˂�Z58��RZ�Q�v�S���      Ŀ3g��$ﱿ���R����U��X#�r��d���JUo�
�#��hܽ����n<����_���҉ �;❻I�Ժ�l�9s��:�U;�2;�@;t�F;�I;�I;b�I;K�I;��I;%gI;.LI;�8I;+I;�!I;�I;�I;�I;�!I;+I;�8I;.LI;%gI;��I;K�I;b�I;�I;�I;t�F;�@;�2;�U;s��:�l�9I�Ժ;❻҉ �_�������n<�����hܽ
�#�JUo�d���r���X#��U�R������$ﱿ3g��      |x�N9�M��pؿkQ��c_��4�_��X#�p���f��<�S�{�����-l�T�-w��e�M�"�Ի��+��LT���:�d;�[,;	/=;�AE;|�H;��I;��I;��I;֕I;�nI;�QI;/=I;|.I;�$I;I;cI;I;�$I;|.I;/=I;�QI;�nI;֕I;��I;��I;��I;|�H;�AE;	/=;�[,;�d;��:�LT���+�"�Իe�M�-w��T�-l�����{�<�S��f��p���X#�4�_�c_��kQ��pؿM��N9�      �X1���,�e���<���2g��c_���U�˂�ՌȾ	ń�-�-�q��Y ��8�2�.?ټ��{�G"��n��O���u:�O ;�&;6":;[�C;!%H;1�I;D�I;��I;�I;�uI;�VI;AI;�1I;3'I;c!I;}I;c!I;3'I;�1I;AI;�VI;�uI;�I;��I;D�I;1�I;!%H;[�C;6":;�&;�O ;��u:�O��n�G"���{�.?ټ8�2�Y ��q��-�-�	ń�ՌȾ˂��U�c_��2g���<�e����,�      d��]]�1K��X1�Xf���kQ��R���Z58��A���נ���O���h什�Q�,���cߓ��� �W��{谺�":��:$ ;�/7; �B;`�G;{I;�I;��I;զI;]{I;Z[I;hDI;<4I;X)I;R#I;G!I;R#I;X)I;<4I;hDI;Z[I;]{I;զI;��I;�I;{I;`�G; �B;�/7;$ ;��:�":{谺W���� �cߓ�,����Q�h什����O��נ��A��Z58�R���kQ����Xf��X1�1K��]]�      L������4z���V��X1��<�pؿ����RZ��	�(���KUo����fy��?l�l�S����7������𺧽�9��:��;]�4;�sA;�1G;�WI;��I;r�I;)�I;�I;�^I;GI;A6I;+I;�$I;�"I;�$I;+I;A6I;GI;�^I;�I;)�I;r�I;��I;�WI;�1G;�sA;]�4;��;��:���9�𺘼����7�S��l�?l�fy�����KUo�(����	��RZ����pؿ�<��X1���V��4z�����      �o��c^���ē��4z�1K�e��M��$ﱿQ�v��X#���Ѿń�	�&�w�нk̀�r��������I� ǻ�5��9�
�:X�;!�2;��@;�F;:I;�I;�I;��I;��I;qaI;II;�7I;~,I;�%I;�#I;�%I;~,I;�7I;II;qaI;��I;��I;�I;�I;:I;�F;��@;!�2;X�;�
�:�9�5� ǻ��I�����r��k̀�w�н	�&�ń���Ѿ�X#�Q�v�$ﱿM��e��1K��4z��ē�c^��      o'���X��c^�������]]���,�N9�3g��S�����/����o��j1��hܽ���-$��l��,}U��Ի~!�{�-���:;�41;��?;m�F;N&I;��I;7�I;Z�I;ąI;�bI;]JI;�8I;E-I;�&I;�$I;�&I;E-I;�8I;]JI;�bI;ąI;Z�I;7�I;��I;N&I;m�F;��?;�41;;��:{�-�~!��Ի,}U��l���-$����hܽj1��o���྘�/�S���3g��N9���,��]]�����c^���X��      j����������΢��+�j��5���	���ȿ%8����7�D�꾂S���7�3但L��-�)��ƼE�\���ݻ�+�!wɸ��:?w;��0;��?;~�F;+I;��I;�I;�I;H�I;�gI;NI;�;I;�/I;�(I;�&I;�(I;�/I;�;I;NI;�gI;H�I;�I;�I;��I;+I;~�F;��?;��0;?w;��:!wɸ�+���ݻE�\��Ƽ-�)��L��3��7��S��D�꾧�7�%8����ȿ��	��5�+�j�΢����������      ��������B��Z�����c�321�#X��ÿhڇ�q�3��s��7��74�i�Gى���&�-Nüq�X�>�ػ��%���J�Ё�:�a;{�0;��?;9�F;�1I;�I;c�I;
�I;m�I;xgI;�MI;R;I;�/I;~(I;�&I;~(I;�/I;R;I;�MI;xgI;m�I;
�I;c�I;�I;�1I;9�F;��?;{�0;�a;Ё�:��J���%�>�ػq�X�-Nü��&�Gى�i�74��7���s�q�3�hڇ��ÿ#X�321���c�Z����B�����      �����B����C��s�P���#�I�������x|��'�YD־�X��s�)�&Խ�Ă�\<�]_���-M�j ˻^���8ё�:�;J2;/u@;��F;�EI;��I;,�I;F�I;%�I;�eI;ZLI;c:I;�.I;�'I;�%I;�'I;�.I;c:I;ZLI;�eI;%�I;F�I;,�I;��I;�EI;��F;/u@;J2;�;ё�:�8^��j ˻�-M�]_��\<��Ă�&Խs�)��X��YD־�'��x|����I�����#�s�P�C�����B��      ΢��Z���C���/]��5�L���,ݿ)8��nm_��K��t��Y�s�'>�����J�o��3��۩��:��T�������9�d�:�;;�^4;&gA;:7G;�cI;%�I;P�I;w�I;��I;KcI;7JI;�8I;m-I;�&I;�$I;�&I;m-I;�8I;7JI;KcI;��I;w�I;P�I;%�I;�cI;:7G;&gA;�^4;�;;�d�:��9����T���:��۩��3�J�o�����'>�Y�s��t���K�nm_�)8���,ݿL���5��/]�C��Z���      +�j���c�s�P��5���o��E���gڇ�Dv<�&���q���_S��������+T��� �P$��+H#�V���o3����:ȯ�:R�;77;��B;��G;׆I;7�I;��I;�I;��I;�_I;fGI;�6I;�+I;+%I;#I;+%I;�+I;�6I;fGI;�_I;��I;�I;��I;7�I;׆I;��G;��B;77;R�;ȯ�:��:o3��V���+H#�P$���� �+T���������_S�q��&���Dv<�gڇ�E���o�����5�s�P���c�      �5�321���#�L��o���ÿ�ҕ�Z������̾�X����0�3�8W����5��zܼ������k�s��Y\�_�n:���:��%;��9;��C;.H;2�I;1�I;%�I;��I;�zI;.[I;�CI;�3I;L)I;8#I;8!I;8#I;L)I;�3I;�CI;.[I;�zI;��I;%�I;1�I;2�I;.H;��C;��9;��%;���:_�n:�Y\�k�s��������zܼ��5�8W��3佃�0��X����̾���Z��ҕ��ÿo��L����#�321�      ��	�#X�I����,ݿE����ҕ� �d��'�?��#���{�W����t���C�o��G��*���Q�'�ػ�0�+�~���:��;N,;q=;WAE;��H;��I;��I;h�I;�I;�sI;�UI;�?I;�0I;�&I;� I;�I;� I;�&I;�0I;�?I;�UI;�sI;�I;h�I;��I;��I;��H;WAE;q=;N,;��;��:+�~��0�'�ػ�Q��*���G�C�o�t������{�W�#���?�꾊'� �d��ҕ�E����,ݿI���#X�      ��ȿ�ÿ���)8��gڇ�Z��'�����l8��Y�s�0�&�`�9{??�W�A琼�G#��7���Vܺ��9U�:��;9K2;c@;��F;I;��I;��I;p�I;d�I;�kI;�OI;u;I;-I;�#I;DI;eI;DI;�#I;-I;u;I;�OI;�kI;d�I;p�I;��I;��I;I;��F;c@;9K2;��;U�:��9�Vܺ�7���G#�A琼W�{??�9`�0�&�Y�s�l8�������'�Z�gڇ�)8������ÿ      %8��hڇ��x|�nm_�Dv<����?��l8��'6~�r74��l������Inc�G��_��2�\�@:�TZ�� >���n:\��:#;�8;ݿB;��G;�wI;��I;��I;��I;��I;ZcI;�II;�6I;5)I;W I;mI;�I;mI;W I;5)I;�6I;�II;ZcI;��I;��I;��I;��I;�wI;��G;ݿB;�8;#;\��:��n:� >�TZ�@:�2�\�_��G��Inc������l��r74�'6~�l8��?�꾎��Dv<�nm_��x|�hڇ�      ��7�q�3��'��K�&�����̾#���Y�s�r74����*N���|��)�^zܼZ��� � ��O���D9뇹:.�;-;%=;�E;!�H;o�I;N�I;��I;ȤI;<zI;�ZI;�BI;q1I;2%I;�I;II;�I;II;�I;2%I;q1I;�BI;�ZI;<zI;ȤI;��I;N�I;o�I;!�H;�E;%=;-;.�;뇹:D9O��� ��� �Z��^zܼ�)��|�*N�����r74�Y�s�#�����̾&����K��'�q�3�      D���s�YD־�t��q���X��{�W�0�&��l��*N���Ă�|�5�׃���Q��#�A���ػ��G�&/�;f:`�:ĕ;y�5;�8A;]�F;�)I;��I;��I;+�I;~�I;RnI;�QI;�;I;4,I;� I;bI;I;�I;I;bI;� I;4,I;�;I;�QI;RnI;~�I;+�I;��I;��I;�)I;]�F;�8A;y�5;ĕ;`�:;f:&/���G���ػ#�A��Q��׃��|�5��Ă�*N���l��0�&�{�W��X��q���t��YD־�s�      �S���7���X��Y�s��_S���0����`ང����|�|�5����۩��X�fc �����5����9#��:��;�,;�K<;vnD;'-H;�I;��I;��I;u�I;q�I;ZbI;|HI;�4I;�&I;fI;�I;�I;�I;�I;�I;fI;�&I;�4I;|HI;ZbI;q�I;u�I;��I;��I;�I;'-H;vnD;�K<;�,;��;#��:��9�5�����fc ��X�۩����|�5��|�����`ས����0��_S�Y�s��X���7��      �7�74�s�)�'>����3�t���9Inc��)�׃��۩��a�1R�ܒ��$O�c�ȸ&��:��;�#;��6;gA;��F;�I;Y�I;��I;0�I;��I;�tI;�VI;�?I;%.I;|!I;3I;I;�I;xI;�I;I;3I;|!I;%.I;�?I;�VI;�tI;��I;0�I;��I;Y�I;�I;��F;gA;��6;�#;��;&��:c�ȸ$O�ܒ��1R��a�۩�׃���)�Inc�9t���3����'>�s�)�74�      3�i�&Խ��������8W��C�o�{??�G��^zܼ�Q���X�1R�/7�������Ϲ��n:�k�:"=;��0;�>;KE;rRH;d�I;��I;�I;[�I;y�I;�eI;DKI;�6I;'I;%I;I;{I;8I;Y
I;8I;{I;I;%I;'I;�6I;DKI;�eI;y�I;[�I;�I;��I;d�I;rRH;KE;�>;��0;"=;�k�:��n:��Ϲ���/7��1R��X��Q��^zܼG��{??�C�o�8W����������&Խi�      �L��Gى��Ă�J�o�+T���5��G�W�_��Z��#�A�fc �ܒ��������:�J:uj�:�d;3,;��:;#4C;+kG;DI;�I;��I;��I;��I;�uI;�WI;b@I;�.I;,!I;�I;�I;�
I;I;eI;I;�
I;�I;�I;,!I;�.I;b@I;�WI;�uI;��I;��I;��I;�I;DI;+kG;#4C;��:;3,;�d;uj�::�J:������ܒ��fc �#�A�Z��_��W��G���5�+T�J�o��Ă�Gى�      -�)���&�\<��3��� ��zܼ�*��A琼2�\�� ���ػ���$O���Ϲ:�J:{h�:v�;��(;�d8;��A;+�F;��H;>�I;��I;!�I;�I;}�I;zdI;�JI;46I;�&I;I;'I;�I;{I;�I;@I;�I;{I;�I;'I;I;�&I;46I;�JI;zdI;}�I;�I;!�I;��I;>�I;��H;+�F;��A;�d8;��(;v�;{h�::�J:��Ϲ$O������ػ� �2�\�A琼�*���zܼ�� ��3�\<���&�      �Ƽ-Nü]_���۩�P$������Q��G#�@:� ����G��5��c�ȸ��n:uj�:v�;+�';�7;�u@;<�E;.uH;�I;��I;��I;]�I;��I;�pI;�TI;I>I;�,I;�I;,I;�I;�I;ZI;I;7I;I;ZI;�I;�I;,I;�I;�,I;I>I;�TI;�pI;��I;]�I;��I;��I;�I;.uH;<�E;�u@;�7;+�';v�;uj�:��n:c�ȸ�5����G� ��@:�G#��Q����P$���۩�]_��-Nü      E�\�q�X��-M��:�+H#����'�ػ�7��TZ�O���&/���9&��:�k�:�d;��(;�7;�@;;\E;�,H;OvI;��I;��I;��I;ܡI;�{I;�]I;�EI;3I;b$I;�I;�I;\	I;UI;7I;@�H;��H;@�H;7I;UI;\	I;�I;�I;b$I;3I;�EI;�]I;�{I;ܡI;��I;��I;��I;OvI;�,H;;\E;�@;�7;��(;�d;�k�:&��:��9&/�O���TZ��7��'�ػ���+H#��:��-M�q�X�      ��ݻ>�ػj ˻�T��V���k�s��0��Vܺ� >�D9;f:#��:��;"=;3,;�d8;�u@;;\E;IH;aI;*�I;��I;X�I;��I;y�I;fI;MI;�8I;)I;~I;�I;I;II;I;Z�H;��H;��H;��H;Z�H;I;II;I;�I;~I;)I;�8I;MI;fI;y�I;��I;X�I;��I;*�I;aI;IH;;\E;�u@;�d8;3,;"=;��;#��:;f:D9� >��Vܺ�0�k�s�V����T��j ˻>�ػ      �+���%�^�����o3���Y\�+�~���9��n:뇹:`�:��;�#;��0;��:;��A;<�E;�,H;aI;��I;��I;��I;"�I;͌I;�lI;SI; >I;I-I;�I;kI;I;tI;�I;�H;��H;�H;��H;�H;��H;�H;�I;tI;I;kI;�I;I-I; >I;SI;�lI;͌I;"�I;��I;��I;��I;aI;�,H;<�E;��A;��:;��0;�#;��;`�:뇹:��n:��9+�~��Y\�o3�����^����%�      !wɸ��J��8��9��:_�n:��:U�:\��:.�;ĕ;�,;��6;�>;#4C;+�F;.uH;OvI;*�I;��I;P�I;޷I;o�I;�qI;�WI;JBI;1I;<#I;�I;�I;�I;XI;Q�H;@�H;��H;��H;��H;��H;��H;@�H;Q�H;XI;�I;�I;�I;<#I;1I;JBI;�WI;�qI;o�I;޷I;P�I;��I;*�I;OvI;.uH;+�F;#4C;�>;��6;�,;ĕ;.�;\��:U�:��:_�n:��:��9�8��J�      ��:Ё�:ё�:�d�:ȯ�:���:��;��;#;-;y�5;�K<;gA;KE;+kG;��H;�I;��I;��I;��I;޷I;	�I;	tI;�ZI;hEI;�3I;�%I;FI;�I;c	I;~I;��H;�H;��H;��H;��H;x�H;��H;��H;��H;�H;��H;~I;c	I;�I;FI;�%I;�3I;hEI;�ZI;	tI;	�I;޷I;��I;��I;��I;�I;��H;+kG;KE;gA;�K<;y�5;-;#;��;��;���:ȯ�:�d�:ё�:Ё�:      ?w;�a;�;�;;R�;��%;N,;9K2;�8;%=;�8A;vnD;��F;rRH;DI;>�I;��I;��I;X�I;"�I;o�I;	tI;v[I;�FI;�5I;�'I;�I;TI;�
I;]I;V�H;��H;]�H;�H;��H;��H;��H;��H;��H;�H;]�H;��H;V�H;]I;�
I;TI;�I;�'I;�5I;�FI;v[I;	tI;o�I;"�I;X�I;��I;��I;>�I;DI;rRH;��F;vnD;�8A;%=;�8;9K2;N,;��%;R�;�;;�;�a;      ��0;{�0;J2;�^4;77;��9;q=;c@;ݿB;�E;]�F;'-H;�I;d�I;�I;��I;��I;��I;��I;͌I;�qI;�ZI;�FI;36I;�(I;I;iI;�I;@I;��H;��H;��H;
�H; �H;��H;�H;��H;�H;��H; �H;
�H;��H;��H;��H;@I;�I;iI;I;�(I;36I;�FI;�ZI;�qI;͌I;��I;��I;��I;��I;�I;d�I;�I;'-H;]�F;�E;ݿB;c@;q=;��9;77;�^4;J2;{�0;      ��?;��?;/u@;&gA;��B;��C;WAE;��F;��G;!�H;�)I;�I;Y�I;��I;��I;!�I;]�I;ܡI;y�I;�lI;�WI;hEI;�5I;�(I;qI;�I;HI;�I;� I;D�H;��H;��H;��H;7�H;�H;v�H;=�H;v�H;�H;7�H;��H;��H;��H;D�H;� I;�I;HI;�I;qI;�(I;�5I;hEI;�WI;�lI;y�I;ܡI;]�I;!�I;��I;��I;Y�I;�I;�)I;!�H;��G;��F;WAE;��C;��B;&gA;/u@;��?;      ~�F;9�F;��F;:7G;��G;.H;��H;I;�wI;o�I;��I;��I;��I;�I;��I;�I;��I;�{I;fI;SI;JBI;�3I;�'I;I;�I;�I;CI;� I;{�H;��H;�H;��H;��H;��H;��H; �H;��H; �H;��H;��H;��H;��H;�H;��H;{�H;� I;CI;�I;�I;I;�'I;�3I;JBI;SI;fI;�{I;��I;�I;��I;�I;��I;��I;��I;o�I;�wI;I;��H;.H;��G;:7G;��F;9�F;      +I;�1I;�EI;�cI;׆I;2�I;��I;��I;��I;N�I;��I;��I;0�I;[�I;��I;}�I;�pI;�]I;MI; >I;1I;�%I;�I;iI;HI;CI;� I;��H;�H;	�H;��H;��H;E�H;)�H;3�H;��H;��H;��H;3�H;)�H;E�H;��H;��H;	�H;�H;��H;� I;CI;HI;iI;�I;�%I;1I; >I;MI;�]I;�pI;}�I;��I;[�I;0�I;��I;��I;N�I;��I;��I;��I;2�I;׆I;�cI;�EI;�1I;      ��I;�I;��I;%�I;7�I;1�I;��I;��I;��I;��I;+�I;u�I;��I;y�I;�uI;zdI;�TI;�EI;�8I;I-I;<#I;FI;TI;�I;�I;� I;��H;?�H;'�H;��H;��H;�H;��H;��H;(�H;��H;��H;��H;(�H;��H;��H;�H;��H;��H;'�H;?�H;��H;� I;�I;�I;TI;FI;<#I;I-I;�8I;�EI;�TI;zdI;�uI;y�I;��I;u�I;+�I;��I;��I;��I;��I;1�I;7�I;%�I;��I;�I;      �I;c�I;,�I;P�I;��I;%�I;h�I;p�I;��I;ȤI;~�I;q�I;�tI;�eI;�WI;�JI;I>I;3I;)I;�I;�I;�I;�
I;@I;� I;{�H;�H;'�H;��H;��H;��H;��H;[�H;��H;A�H;��H;��H;��H;A�H;��H;[�H;��H;��H;��H;��H;'�H;�H;{�H;� I;@I;�
I;�I;�I;�I;)I;3I;I>I;�JI;�WI;�eI;�tI;q�I;~�I;ȤI;��I;p�I;h�I;%�I;��I;P�I;,�I;c�I;      �I;
�I;F�I;w�I;�I;��I;�I;d�I;��I;<zI;RnI;ZbI;�VI;DKI;b@I;46I;�,I;b$I;~I;kI;�I;c	I;]I;��H;D�H;��H;	�H;��H;��H;��H;��H;O�H;f�H;��H;'�H;��H;��H;��H;'�H;��H;f�H;O�H;��H;��H;��H;��H;	�H;��H;D�H;��H;]I;c	I;�I;kI;~I;b$I;�,I;46I;b@I;DKI;�VI;ZbI;RnI;<zI;��I;d�I;�I;��I;�I;w�I;F�I;
�I;      H�I;m�I;%�I;��I;��I;�zI;�sI;�kI;ZcI;�ZI;�QI;|HI;�?I;�6I;�.I;�&I;�I;�I;�I;I;�I;~I;V�H;��H;��H;�H;��H;��H;��H;��H;C�H;>�H;��H;��H;p�H;N�H;5�H;N�H;p�H;��H;��H;>�H;C�H;��H;��H;��H;��H;�H;��H;��H;V�H;~I;�I;I;�I;�I;�I;�&I;�.I;�6I;�?I;|HI;�QI;�ZI;ZcI;�kI;�sI;�zI;��I;��I;%�I;m�I;      �gI;xgI;�eI;KcI;�_I;.[I;�UI;�OI;�II;�BI;�;I;�4I;%.I;'I;,!I;I;,I;�I;I;tI;XI;��H;��H;��H;��H;��H;��H;�H;��H;O�H;>�H;��H;��H;8�H;��H;��H;��H;��H;��H;8�H;��H;��H;>�H;O�H;��H;�H;��H;��H;��H;��H;��H;��H;XI;tI;I;�I;,I;I;,!I;'I;%.I;�4I;�;I;�BI;�II;�OI;�UI;.[I;�_I;KcI;�eI;xgI;      NI;�MI;ZLI;7JI;fGI;�CI;�?I;u;I;�6I;q1I;4,I;�&I;|!I;%I;�I;'I;�I;\	I;II;�I;Q�H;�H;]�H;
�H;��H;��H;E�H;��H;[�H;f�H;��H;��H;�H;��H;{�H;;�H;2�H;;�H;{�H;��H;�H;��H;��H;f�H;[�H;��H;E�H;��H;��H;
�H;]�H;�H;Q�H;�I;II;\	I;�I;'I;�I;%I;|!I;�&I;4,I;q1I;�6I;u;I;�?I;�CI;fGI;7JI;ZLI;�MI;      �;I;R;I;c:I;�8I;�6I;�3I;�0I;-I;5)I;2%I;� I;fI;3I;I;�I;�I;�I;UI;I;�H;@�H;��H;�H; �H;7�H;��H;)�H;��H;��H;��H;��H;8�H;��H;W�H;�H;��H;��H;��H;�H;W�H;��H;8�H;��H;��H;��H;��H;)�H;��H;7�H; �H;�H;��H;@�H;�H;I;UI;�I;�I;�I;I;3I;fI;� I;2%I;5)I;-I;�0I;�3I;�6I;�8I;c:I;R;I;      �/I;�/I;�.I;m-I;�+I;L)I;�&I;�#I;W I;�I;bI;�I;I;{I;�
I;{I;ZI;7I;Z�H;��H;��H;��H;��H;��H;�H;��H;3�H;(�H;A�H;'�H;p�H;��H;{�H;�H;��H;��H;��H;��H;��H;�H;{�H;��H;p�H;'�H;A�H;(�H;3�H;��H;�H;��H;��H;��H;��H;��H;Z�H;7I;ZI;{I;�
I;{I;I;�I;bI;�I;W I;�#I;�&I;L)I;�+I;m-I;�.I;�/I;      �(I;~(I;�'I;�&I;+%I;8#I;� I;DI;mI;II;I;�I;�I;8I;I;�I;I;@�H;��H;�H;��H;��H;��H;�H;v�H; �H;��H;��H;��H;��H;N�H;��H;;�H;��H;��H;o�H;i�H;o�H;��H;��H;;�H;��H;N�H;��H;��H;��H;��H; �H;v�H;�H;��H;��H;��H;�H;��H;@�H;I;�I;I;8I;�I;�I;I;II;mI;DI;� I;8#I;+%I;�&I;�'I;~(I;      �&I;�&I;�%I;�$I;#I;8!I;�I;eI;�I;�I;�I;�I;xI;Y
I;eI;@I;7I;��H;��H;��H;��H;x�H;��H;��H;=�H;��H;��H;��H;��H;��H;5�H;��H;2�H;��H;��H;i�H;L�H;i�H;��H;��H;2�H;��H;5�H;��H;��H;��H;��H;��H;=�H;��H;��H;x�H;��H;��H;��H;��H;7I;@I;eI;Y
I;xI;�I;�I;�I;�I;eI;�I;8!I;#I;�$I;�%I;�&I;      �(I;~(I;�'I;�&I;+%I;8#I;� I;DI;mI;II;I;�I;�I;8I;I;�I;I;@�H;��H;�H;��H;��H;��H;�H;v�H; �H;��H;��H;��H;��H;N�H;��H;;�H;��H;��H;o�H;i�H;o�H;��H;��H;;�H;��H;N�H;��H;��H;��H;��H; �H;v�H;�H;��H;��H;��H;�H;��H;@�H;I;�I;I;8I;�I;�I;I;II;mI;DI;� I;8#I;+%I;�&I;�'I;~(I;      �/I;�/I;�.I;m-I;�+I;L)I;�&I;�#I;W I;�I;bI;�I;I;{I;�
I;{I;ZI;7I;Z�H;��H;��H;��H;��H;��H;�H;��H;3�H;(�H;A�H;'�H;p�H;��H;{�H;�H;��H;��H;��H;��H;��H;�H;{�H;��H;p�H;'�H;A�H;(�H;3�H;��H;�H;��H;��H;��H;��H;��H;Z�H;7I;ZI;{I;�
I;{I;I;�I;bI;�I;W I;�#I;�&I;L)I;�+I;m-I;�.I;�/I;      �;I;R;I;c:I;�8I;�6I;�3I;�0I;-I;5)I;2%I;� I;fI;3I;I;�I;�I;�I;UI;I;�H;@�H;��H;�H; �H;7�H;��H;)�H;��H;��H;��H;��H;8�H;��H;W�H;�H;��H;��H;��H;�H;W�H;��H;8�H;��H;��H;��H;��H;)�H;��H;7�H; �H;�H;��H;@�H;�H;I;UI;�I;�I;�I;I;3I;fI;� I;2%I;5)I;-I;�0I;�3I;�6I;�8I;c:I;R;I;      NI;�MI;ZLI;7JI;fGI;�CI;�?I;u;I;�6I;q1I;4,I;�&I;|!I;%I;�I;'I;�I;\	I;II;�I;Q�H;�H;]�H;
�H;��H;��H;E�H;��H;[�H;f�H;��H;��H;�H;��H;{�H;;�H;2�H;;�H;{�H;��H;�H;��H;��H;f�H;[�H;��H;E�H;��H;��H;
�H;]�H;�H;Q�H;�I;II;\	I;�I;'I;�I;%I;|!I;�&I;4,I;q1I;�6I;u;I;�?I;�CI;fGI;7JI;ZLI;�MI;      �gI;xgI;�eI;KcI;�_I;.[I;�UI;�OI;�II;�BI;�;I;�4I;%.I;'I;,!I;I;,I;�I;I;tI;XI;��H;��H;��H;��H;��H;��H;�H;��H;O�H;>�H;��H;��H;8�H;��H;��H;��H;��H;��H;8�H;��H;��H;>�H;O�H;��H;�H;��H;��H;��H;��H;��H;��H;XI;tI;I;�I;,I;I;,!I;'I;%.I;�4I;�;I;�BI;�II;�OI;�UI;.[I;�_I;KcI;�eI;xgI;      H�I;m�I;%�I;��I;��I;�zI;�sI;�kI;ZcI;�ZI;�QI;|HI;�?I;�6I;�.I;�&I;�I;�I;�I;I;�I;~I;V�H;��H;��H;�H;��H;��H;��H;��H;C�H;>�H;��H;��H;p�H;N�H;5�H;N�H;p�H;��H;��H;>�H;C�H;��H;��H;��H;��H;�H;��H;��H;V�H;~I;�I;I;�I;�I;�I;�&I;�.I;�6I;�?I;|HI;�QI;�ZI;ZcI;�kI;�sI;�zI;��I;��I;%�I;m�I;      �I;
�I;F�I;w�I;�I;��I;�I;d�I;��I;<zI;RnI;ZbI;�VI;DKI;b@I;46I;�,I;b$I;~I;kI;�I;c	I;]I;��H;D�H;��H;	�H;��H;��H;��H;��H;O�H;f�H;��H;'�H;��H;��H;��H;'�H;��H;f�H;O�H;��H;��H;��H;��H;	�H;��H;D�H;��H;]I;c	I;�I;kI;~I;b$I;�,I;46I;b@I;DKI;�VI;ZbI;RnI;<zI;��I;d�I;�I;��I;�I;w�I;F�I;
�I;      �I;c�I;,�I;P�I;��I;%�I;h�I;p�I;��I;ȤI;~�I;q�I;�tI;�eI;�WI;�JI;I>I;3I;)I;�I;�I;�I;�
I;@I;� I;{�H;�H;'�H;��H;��H;��H;��H;[�H;��H;A�H;��H;��H;��H;A�H;��H;[�H;��H;��H;��H;��H;'�H;�H;{�H;� I;@I;�
I;�I;�I;�I;)I;3I;I>I;�JI;�WI;�eI;�tI;q�I;~�I;ȤI;��I;p�I;h�I;%�I;��I;P�I;,�I;c�I;      ��I;�I;��I;%�I;7�I;1�I;��I;��I;��I;��I;+�I;u�I;��I;y�I;�uI;zdI;�TI;�EI;�8I;I-I;<#I;FI;TI;�I;�I;� I;��H;?�H;'�H;��H;��H;�H;��H;��H;(�H;��H;��H;��H;(�H;��H;��H;�H;��H;��H;'�H;?�H;��H;� I;�I;�I;TI;FI;<#I;I-I;�8I;�EI;�TI;zdI;�uI;y�I;��I;u�I;+�I;��I;��I;��I;��I;1�I;7�I;%�I;��I;�I;      +I;�1I;�EI;�cI;׆I;2�I;��I;��I;��I;N�I;��I;��I;0�I;[�I;��I;}�I;�pI;�]I;MI; >I;1I;�%I;�I;iI;HI;CI;� I;��H;�H;	�H;��H;��H;E�H;)�H;3�H;��H;��H;��H;3�H;)�H;E�H;��H;��H;	�H;�H;��H;� I;CI;HI;iI;�I;�%I;1I; >I;MI;�]I;�pI;}�I;��I;[�I;0�I;��I;��I;N�I;��I;��I;��I;2�I;׆I;�cI;�EI;�1I;      ~�F;9�F;��F;:7G;��G;.H;��H;I;�wI;o�I;��I;��I;��I;�I;��I;�I;��I;�{I;fI;SI;JBI;�3I;�'I;I;�I;�I;CI;� I;{�H;��H;�H;��H;��H;��H;��H; �H;��H; �H;��H;��H;��H;��H;�H;��H;{�H;� I;CI;�I;�I;I;�'I;�3I;JBI;SI;fI;�{I;��I;�I;��I;�I;��I;��I;��I;o�I;�wI;I;��H;.H;��G;:7G;��F;9�F;      ��?;��?;/u@;&gA;��B;��C;WAE;��F;��G;!�H;�)I;�I;Y�I;��I;��I;!�I;]�I;ܡI;y�I;�lI;�WI;hEI;�5I;�(I;qI;�I;HI;�I;� I;D�H;��H;��H;��H;7�H;�H;v�H;=�H;v�H;�H;7�H;��H;��H;��H;D�H;� I;�I;HI;�I;qI;�(I;�5I;hEI;�WI;�lI;y�I;ܡI;]�I;!�I;��I;��I;Y�I;�I;�)I;!�H;��G;��F;WAE;��C;��B;&gA;/u@;��?;      ��0;{�0;J2;�^4;77;��9;q=;c@;ݿB;�E;]�F;'-H;�I;d�I;�I;��I;��I;��I;��I;͌I;�qI;�ZI;�FI;36I;�(I;I;iI;�I;@I;��H;��H;��H;
�H; �H;��H;�H;��H;�H;��H; �H;
�H;��H;��H;��H;@I;�I;iI;I;�(I;36I;�FI;�ZI;�qI;͌I;��I;��I;��I;��I;�I;d�I;�I;'-H;]�F;�E;ݿB;c@;q=;��9;77;�^4;J2;{�0;      ?w;�a;�;�;;R�;��%;N,;9K2;�8;%=;�8A;vnD;��F;rRH;DI;>�I;��I;��I;X�I;"�I;o�I;	tI;v[I;�FI;�5I;�'I;�I;TI;�
I;]I;V�H;��H;]�H;�H;��H;��H;��H;��H;��H;�H;]�H;��H;V�H;]I;�
I;TI;�I;�'I;�5I;�FI;v[I;	tI;o�I;"�I;X�I;��I;��I;>�I;DI;rRH;��F;vnD;�8A;%=;�8;9K2;N,;��%;R�;�;;�;�a;      ��:Ё�:ё�:�d�:ȯ�:���:��;��;#;-;y�5;�K<;gA;KE;+kG;��H;�I;��I;��I;��I;޷I;	�I;	tI;�ZI;hEI;�3I;�%I;FI;�I;c	I;~I;��H;�H;��H;��H;��H;x�H;��H;��H;��H;�H;��H;~I;c	I;�I;FI;�%I;�3I;hEI;�ZI;	tI;	�I;޷I;��I;��I;��I;�I;��H;+kG;KE;gA;�K<;y�5;-;#;��;��;���:ȯ�:�d�:ё�:Ё�:      !wɸ��J��8��9��:_�n:��:U�:\��:.�;ĕ;�,;��6;�>;#4C;+�F;.uH;OvI;*�I;��I;P�I;޷I;o�I;�qI;�WI;JBI;1I;<#I;�I;�I;�I;XI;Q�H;@�H;��H;��H;��H;��H;��H;@�H;Q�H;XI;�I;�I;�I;<#I;1I;JBI;�WI;�qI;o�I;޷I;P�I;��I;*�I;OvI;.uH;+�F;#4C;�>;��6;�,;ĕ;.�;\��:U�:��:_�n:��:��9�8��J�      �+���%�^�����o3���Y\�+�~���9��n:뇹:`�:��;�#;��0;��:;��A;<�E;�,H;aI;��I;��I;��I;"�I;͌I;�lI;SI; >I;I-I;�I;kI;I;tI;�I;�H;��H;�H;��H;�H;��H;�H;�I;tI;I;kI;�I;I-I; >I;SI;�lI;͌I;"�I;��I;��I;��I;aI;�,H;<�E;��A;��:;��0;�#;��;`�:뇹:��n:��9+�~��Y\�o3�����^����%�      ��ݻ>�ػj ˻�T��V���k�s��0��Vܺ� >�D9;f:#��:��;"=;3,;�d8;�u@;;\E;IH;aI;*�I;��I;X�I;��I;y�I;fI;MI;�8I;)I;~I;�I;I;II;I;Z�H;��H;��H;��H;Z�H;I;II;I;�I;~I;)I;�8I;MI;fI;y�I;��I;X�I;��I;*�I;aI;IH;;\E;�u@;�d8;3,;"=;��;#��:;f:D9� >��Vܺ�0�k�s�V����T��j ˻>�ػ      E�\�q�X��-M��:�+H#����'�ػ�7��TZ�O���&/���9&��:�k�:�d;��(;�7;�@;;\E;�,H;OvI;��I;��I;��I;ܡI;�{I;�]I;�EI;3I;b$I;�I;�I;\	I;UI;7I;@�H;��H;@�H;7I;UI;\	I;�I;�I;b$I;3I;�EI;�]I;�{I;ܡI;��I;��I;��I;OvI;�,H;;\E;�@;�7;��(;�d;�k�:&��:��9&/�O���TZ��7��'�ػ���+H#��:��-M�q�X�      �Ƽ-Nü]_���۩�P$������Q��G#�@:� ����G��5��c�ȸ��n:uj�:v�;+�';�7;�u@;<�E;.uH;�I;��I;��I;]�I;��I;�pI;�TI;I>I;�,I;�I;,I;�I;�I;ZI;I;7I;I;ZI;�I;�I;,I;�I;�,I;I>I;�TI;�pI;��I;]�I;��I;��I;�I;.uH;<�E;�u@;�7;+�';v�;uj�:��n:c�ȸ�5����G� ��@:�G#��Q����P$���۩�]_��-Nü      -�)���&�\<��3��� ��zܼ�*��A琼2�\�� ���ػ���$O���Ϲ:�J:{h�:v�;��(;�d8;��A;+�F;��H;>�I;��I;!�I;�I;}�I;zdI;�JI;46I;�&I;I;'I;�I;{I;�I;@I;�I;{I;�I;'I;I;�&I;46I;�JI;zdI;}�I;�I;!�I;��I;>�I;��H;+�F;��A;�d8;��(;v�;{h�::�J:��Ϲ$O������ػ� �2�\�A琼�*���zܼ�� ��3�\<���&�      �L��Gى��Ă�J�o�+T���5��G�W�_��Z��#�A�fc �ܒ��������:�J:uj�:�d;3,;��:;#4C;+kG;DI;�I;��I;��I;��I;�uI;�WI;b@I;�.I;,!I;�I;�I;�
I;I;eI;I;�
I;�I;�I;,!I;�.I;b@I;�WI;�uI;��I;��I;��I;�I;DI;+kG;#4C;��:;3,;�d;uj�::�J:������ܒ��fc �#�A�Z��_��W��G���5�+T�J�o��Ă�Gى�      3�i�&Խ��������8W��C�o�{??�G��^zܼ�Q���X�1R�/7�������Ϲ��n:�k�:"=;��0;�>;KE;rRH;d�I;��I;�I;[�I;y�I;�eI;DKI;�6I;'I;%I;I;{I;8I;Y
I;8I;{I;I;%I;'I;�6I;DKI;�eI;y�I;[�I;�I;��I;d�I;rRH;KE;�>;��0;"=;�k�:��n:��Ϲ���/7��1R��X��Q��^zܼG��{??�C�o�8W����������&Խi�      �7�74�s�)�'>����3�t���9Inc��)�׃��۩��a�1R�ܒ��$O�c�ȸ&��:��;�#;��6;gA;��F;�I;Y�I;��I;0�I;��I;�tI;�VI;�?I;%.I;|!I;3I;I;�I;xI;�I;I;3I;|!I;%.I;�?I;�VI;�tI;��I;0�I;��I;Y�I;�I;��F;gA;��6;�#;��;&��:c�ȸ$O�ܒ��1R��a�۩�׃���)�Inc�9t���3����'>�s�)�74�      �S���7���X��Y�s��_S���0����`ང����|�|�5����۩��X�fc �����5����9#��:��;�,;�K<;vnD;'-H;�I;��I;��I;u�I;q�I;ZbI;|HI;�4I;�&I;fI;�I;�I;�I;�I;�I;fI;�&I;�4I;|HI;ZbI;q�I;u�I;��I;��I;�I;'-H;vnD;�K<;�,;��;#��:��9�5�����fc ��X�۩����|�5��|�����`ས����0��_S�Y�s��X���7��      D���s�YD־�t��q���X��{�W�0�&��l��*N���Ă�|�5�׃���Q��#�A���ػ��G�&/�;f:`�:ĕ;y�5;�8A;]�F;�)I;��I;��I;+�I;~�I;RnI;�QI;�;I;4,I;� I;bI;I;�I;I;bI;� I;4,I;�;I;�QI;RnI;~�I;+�I;��I;��I;�)I;]�F;�8A;y�5;ĕ;`�:;f:&/���G���ػ#�A��Q��׃��|�5��Ă�*N���l��0�&�{�W��X��q���t��YD־�s�      ��7�q�3��'��K�&�����̾#���Y�s�r74����*N���|��)�^zܼZ��� � ��O���D9뇹:.�;-;%=;�E;!�H;o�I;N�I;��I;ȤI;<zI;�ZI;�BI;q1I;2%I;�I;II;�I;II;�I;2%I;q1I;�BI;�ZI;<zI;ȤI;��I;N�I;o�I;!�H;�E;%=;-;.�;뇹:D9O��� ��� �Z��^zܼ�)��|�*N�����r74�Y�s�#�����̾&����K��'�q�3�      %8��hڇ��x|�nm_�Dv<����?��l8��'6~�r74��l������Inc�G��_��2�\�@:�TZ�� >���n:\��:#;�8;ݿB;��G;�wI;��I;��I;��I;��I;ZcI;�II;�6I;5)I;W I;mI;�I;mI;W I;5)I;�6I;�II;ZcI;��I;��I;��I;��I;�wI;��G;ݿB;�8;#;\��:��n:� >�TZ�@:�2�\�_��G��Inc������l��r74�'6~�l8��?�꾎��Dv<�nm_��x|�hڇ�      ��ȿ�ÿ���)8��gڇ�Z��'�����l8��Y�s�0�&�`�9{??�W�A琼�G#��7���Vܺ��9U�:��;9K2;c@;��F;I;��I;��I;p�I;d�I;�kI;�OI;u;I;-I;�#I;DI;eI;DI;�#I;-I;u;I;�OI;�kI;d�I;p�I;��I;��I;I;��F;c@;9K2;��;U�:��9�Vܺ�7���G#�A琼W�{??�9`�0�&�Y�s�l8�������'�Z�gڇ�)8������ÿ      ��	�#X�I����,ݿE����ҕ� �d��'�?��#���{�W����t���C�o��G��*���Q�'�ػ�0�+�~���:��;N,;q=;WAE;��H;��I;��I;h�I;�I;�sI;�UI;�?I;�0I;�&I;� I;�I;� I;�&I;�0I;�?I;�UI;�sI;�I;h�I;��I;��I;��H;WAE;q=;N,;��;��:+�~��0�'�ػ�Q��*���G�C�o�t������{�W�#���?�꾊'� �d��ҕ�E����,ݿI���#X�      �5�321���#�L��o���ÿ�ҕ�Z������̾�X����0�3�8W����5��zܼ������k�s��Y\�_�n:���:��%;��9;��C;.H;2�I;1�I;%�I;��I;�zI;.[I;�CI;�3I;L)I;8#I;8!I;8#I;L)I;�3I;�CI;.[I;�zI;��I;%�I;1�I;2�I;.H;��C;��9;��%;���:_�n:�Y\�k�s��������zܼ��5�8W��3佃�0��X����̾���Z��ҕ��ÿo��L����#�321�      +�j���c�s�P��5���o��E���gڇ�Dv<�&���q���_S��������+T��� �P$��+H#�V���o3����:ȯ�:R�;77;��B;��G;׆I;7�I;��I;�I;��I;�_I;fGI;�6I;�+I;+%I;#I;+%I;�+I;�6I;fGI;�_I;��I;�I;��I;7�I;׆I;��G;��B;77;R�;ȯ�:��:o3��V���+H#�P$���� �+T���������_S�q��&���Dv<�gڇ�E���o�����5�s�P���c�      ΢��Z���C���/]��5�L���,ݿ)8��nm_��K��t��Y�s�'>�����J�o��3��۩��:��T�������9�d�:�;;�^4;&gA;:7G;�cI;%�I;P�I;w�I;��I;KcI;7JI;�8I;m-I;�&I;�$I;�&I;m-I;�8I;7JI;KcI;��I;w�I;P�I;%�I;�cI;:7G;&gA;�^4;�;;�d�:��9����T���:��۩��3�J�o�����'>�Y�s��t���K�nm_�)8���,ݿL���5��/]�C��Z���      �����B����C��s�P���#�I�������x|��'�YD־�X��s�)�&Խ�Ă�\<�]_���-M�j ˻^���8ё�:�;J2;/u@;��F;�EI;��I;,�I;F�I;%�I;�eI;ZLI;c:I;�.I;�'I;�%I;�'I;�.I;c:I;ZLI;�eI;%�I;F�I;,�I;��I;�EI;��F;/u@;J2;�;ё�:�8^��j ˻�-M�]_��\<��Ă�&Խs�)��X��YD־�'��x|����I�����#�s�P�C�����B��      ��������B��Z�����c�321�#X��ÿhڇ�q�3��s��7��74�i�Gى���&�-Nüq�X�>�ػ��%���J�Ё�:�a;{�0;��?;9�F;�1I;�I;c�I;
�I;m�I;xgI;�MI;R;I;�/I;~(I;�&I;~(I;�/I;R;I;�MI;xgI;m�I;
�I;c�I;�I;�1I;9�F;��?;{�0;�a;Ё�:��J���%�>�ػq�X�-Nü��&�Gى�i�74��7���s�q�3�hڇ��ÿ#X�321���c�Z����B�����      A(��o'���o��L�d��X1�|x�Ŀ����3�v���x����4�s��b+���'�"�ü�yY�llٻq&�>�p�Y��:_;��0;��?;�F;tI;�I;��I;H�I;��I;ucI;�JI;�8I;�-I;�&I;�$I;�&I;�-I;�8I;�JI;ucI;��I;H�I;��I;�I;tI;�F;��?;��0;_;Y��:>�p�q&�llٻ�yY�"�ü�'�b+��s����4��x��v���3����Ŀ|x��X1�d�L��o��o'��      o'���X��c^�������]]���,�N9�3g��S�����/����o��j1��hܽ���-$��l��,}U��Ի~!���-���:;�41;��?;m�F;N&I;��I;7�I;Z�I;ąI;�bI;]JI;�8I;E-I;�&I;�$I;�&I;E-I;�8I;]JI;�bI;ąI;Z�I;7�I;��I;N&I;m�F;��?;�41;;��:��-�~!��Ի,}U��l���-$����hܽj1��o���྘�/�S���3g��N9���,��]]�����c^���X��      �o��c^���ē��4z�1K�e��M��$ﱿQ�v��X#���Ѿń�	�&�w�нk̀�r��������I� ǻ�5��9�
�:X�;!�2;��@;�F;:I;�I;�I;��I;��I;qaI;II;�7I;~,I;�%I;�#I;�%I;~,I;�7I;II;qaI;��I;��I;�I;�I;:I;�F;��@;!�2;X�;�
�:�9�5� ǻ��I�����r��k̀�w�н	�&�ń���Ѿ�X#�Q�v�$ﱿM��e��1K��4z��ē�c^��      L������4z���V��X1��<�pؿ����RZ��	�(���KUo����fy��?l�l�S����7������𺧽�9��:��;]�4;�sA;�1G;�WI;��I;r�I;)�I;�I;�^I;GI;A6I;+I;�$I;�"I;�$I;+I;A6I;GI;�^I;�I;)�I;r�I;��I;�WI;�1G;�sA;]�4;��;��:���9�𺘼����7�S��l�?l�fy�����KUo�(����	��RZ����pؿ�<��X1���V��4z�����      d��]]�1K��X1�Xf���kQ��R���Z58��A���נ���O���h什�Q�,���cߓ��� �W��|谺�":��:$ ;�/7; �B;`�G;{I;�I;��I;զI;]{I;Z[I;hDI;<4I;X)I;R#I;G!I;R#I;X)I;<4I;hDI;Z[I;]{I;զI;��I;�I;{I;`�G; �B;�/7;$ ;��:�":|谺W���� �cߓ�,����Q�h什����O��נ��A��Z58�R���kQ����Xf��X1�1K��]]�      �X1���,�e���<���2g��c_���U�˂�ՌȾ	ń�-�-�q��Y ��8�2�.?ټ��{�G"��n��O���u:�O ;�&;6":;[�C;!%H;1�I;D�I;��I;�I;�uI;�VI;AI;�1I;3'I;c!I;}I;c!I;3'I;�1I;AI;�VI;�uI;�I;��I;D�I;1�I;!%H;[�C;6":;�&;�O ;��u:�O��n�G"���{�.?ټ8�2�Y ��q��-�-�	ń�ՌȾ˂��U�c_��2g���<�e����,�      |x�N9�M��pؿkQ��c_��4�_��X#�p���f��<�S�{�����-l�T�-w��e�M�"�Ի��+��LT���:�d;�[,;	/=;�AE;|�H;��I;��I;��I;֕I;�nI;�QI;/=I;|.I;�$I;I;cI;I;�$I;|.I;/=I;�QI;�nI;֕I;��I;��I;��I;|�H;�AE;	/=;�[,;�d;��:�LT���+�"�Իe�M�-w��T�-l�����{�<�S��f��p���X#�4�_�c_��kQ��pؿM��N9�      Ŀ3g��$ﱿ���R����U��X#�r��d���JUo�
�#��hܽ����n<����_���҉ �;❻I�Ժ�l�9s��:�U;�2;�@;t�F;�I;�I;b�I;K�I;��I;%gI;.LI;�8I;+I;�!I;�I;�I;�I;�!I;+I;�8I;.LI;%gI;��I;K�I;b�I;�I;�I;t�F;�@;�2;�U;s��:�l�9I�Ժ;❻҉ �_�������n<�����hܽ
�#�JUo�d���r���X#��U�R������$ﱿ3g��      ���S���Q�v��RZ�Z58�˂�p��d���hoy�`1�gO��d什�`�`��6����yY���컞�T��1���u:��:\~#;.88;�B;��G;lI;-�I;"�I;L�I;��I;�^I;!FI;4I;C'I;�I;�I;)I;�I;�I;C'I;4I;!FI;�^I;��I;L�I;"�I;-�I;lI;��G;�B;.88;\~#;��:��u:�1���T���컶yY�6���`���`�d什gO��`1�hoy�d���p��˂�Z58��RZ�Q�v�S���      �3���/��X#��	��A��ՌȾ�f��JUo�`1�Ӱ���n���x��'��>ټ�@��-l�S���$��&�39�!�:;Q;!d-;�.=;�E;wH;��I;-�I;��I; �I;6uI;�VI;�?I;/I;B#I;_I;�I;TI;�I;_I;B#I;/I;�?I;�VI;6uI; �I;��I;-�I;��I;wH;�E;�.=;!d-;;Q;�!�:&�39$��S���-l��@���>ټ�'��x��n��Ӱ��`1�JUo��f��ՌȾ�A���	��X#���/�      v���ྃ�Ѿ(����נ�	ń�<�S�
�#�gO���n��R̀��2�,������>���Ի��B��#�[m:�E�:o ;��5;�EA;��F;�I;r�I;p�I;ŽI;��I;�iI;�MI;.9I;�)I;I;�I;�I;iI;�I;�I;I;�)I;.9I;�MI;�iI;��I;ŽI;p�I;r�I;�I;��F;�EA;��5;o ;�E�:[m:�#���B���Ի��>���,���2�R̀��n��gO��
�#�<�S�	ń��נ�(�����Ѿ��      �x���o��ń�KUo���O�-�-�{��hܽd什�x��2��b��yR���|U��2�����"찺�m�9��:C;��,;�g<;�qD;h$H;�I;��I;��I;&�I;&I;�]I;(EI;r2I;�$I;�I;}I;�I;QI;�I;}I;�I;�$I;r2I;(EI;�]I;&I;&�I;��I;��I;�I;h$H;�qD;�g<;��,;C;��:�m�9"찺����2���|U�yR���b���2��x�d什�hܽ{�-�-���O�KUo�ń��o��      ��4�j1�	�&������q�ཌྷ�������`��'�,��yR����]�����V��[��q�o����:{�;=~#;0�6;nsA;s�F;�I;��I;��I;��I;6�I;�oI;�RI;�<I;�+I;�I;�I;�I;`I;WI;`I;�I;�I;�I;�+I;�<I;�RI;�oI;6�I;��I;��I;��I;�I;s�F;nsA;0�6;=~#;{�;���:q�o�[���V�������]�yR��,��'��`��������q�������	�&�j1�      s�ཾhܽw�нfy��h什Y ��-l��n<�`���>ټ�𛼝|U����H᝻�2�������u:jj�:�;}61;j(>;sE;,IH;p�I;��I;��I;�I;��I;zaI;�GI;G4I;~%I;�I;�I;XI;<
I;7	I;<
I;XI;�I;�I;~%I;G4I;�GI;zaI;��I;�I;��I;��I;p�I;,IH;sE;j(>;}61;�;jj�:��u:�����2�H᝻����|U����>ټ`���n<�-l�Y ��h什fy��w�н�hܽ      b+����k̀�?l��Q�8�2�T����6����@����>��2���V���2���� R:���:�;�[,;P;;;C;�dG;w8I;��I;U�I;��I;_�I;�pI;�SI;=I;W,I;KI;�I;�I;�	I;+I;'I;+I;�	I;�I;�I;KI;W,I;=I;�SI;�pI;_�I;��I;U�I;��I;w8I;�dG;;C;P;;�[,;�;���: R:���2��V���2����>��@��6������T�8�2��Q�?l�k̀���      �'��-$�r��l�,���.?ټ-w��_����yY�-l���Ի���[������ R:���:�Q;�);��8;��A;�F;S�H;J�I;��I;��I;ȨI;$�I;�_I;GI;�3I;�$I;cI;�I;�
I;�I;*I;]I;*I;�I;�
I;�I;cI;�$I;�3I;GI;�_I;$�I;ȨI;��I;��I;J�I;S�H;�F;��A;��8;�);�Q;���: R:����[�������Ի-l��yY�_���-w��.?ټ,���l�r���-$�      "�ü�l������S��cߓ���{�e�M�҉ ����S�����B�"찺q�o���u:���:�Q;D�';)07;ք@;�E;�kH;N�I;��I;��I;,�I;��I;�kI;�PI;D;I;�*I;�I;�I;|I;�I;[I;CI;� I;CI;[I;�I;|I;�I;�I;�*I;D;I;�PI;�kI;��I;,�I;��I;��I;N�I;�kH;�E;ք@;)07;D�';�Q;���:��u:q�o�"찺��B�S������҉ �e�M���{�cߓ�S�������l��      �yY�,}U���I���7��� �G"�"�Ի;❻��T�$���#��m�9���:jj�:�;�);)07;D@;V\E;�#H;�jI;(�I;s�I;�I;L�I;�vI;�YI;�BI;�0I;g"I;DI;�I;EI;�I;N I;�H;�H;�H;N I;�I;EI;�I;DI;g"I;�0I;�BI;�YI;�vI;L�I;�I;s�I;(�I;�jI;�#H;V\E;D@;)07;�);�;jj�:���:�m�9�#�$���T�;❻"�ԻG"��� ���7���I�,}U�      llٻ�Ի ǻ����W���n���+�I�Ժ�1�&�39[m:��:{�;�;�[,;��8;ք@;V\E;�	H;jUI;��I;	�I;�I;}�I;#�I;�aI;}II;>6I;�&I;�I;GI;�	I;OI;O I;{�H;��H;��H;��H;{�H;O I;OI;�	I;GI;�I;�&I;>6I;}II;�aI;#�I;}�I;�I;	�I;��I;jUI;�	H;V\E;ք@;��8;�[,;�;{�;��:[m:&�39�1�I�Ժ��+��n�W������ ǻ�Ի      q&�~!��5���|谺�O��LT��l�9��u:�!�:�E�:C;=~#;}61;P;;��A;�E;�#H;jUI;,�I;��I;1�I;��I;�I;-hI;COI;7;I;+I;3I;�I;�I;�I;� I;F�H;��H;��H;�H;��H;��H;F�H;� I;�I;�I;�I;3I;+I;7;I;COI;-hI;�I;��I;1�I;��I;,�I;jUI;�#H;�E;��A;P;;}61;=~#;C;�E�:�!�:��u:�l�9�LT��O�|谺���5�~!�      >�p���-��9���9�":��u:��:s��:��:;Q;o ;��,;0�6;j(>;;C;�F;�kH;�jI;��I;��I;��I;4�I;��I;�lI;�SI;??I;�.I;8!I;nI;�I;�I;�I;��H;��H;��H;c�H;��H;c�H;��H;��H;��H;�I;�I;�I;nI;8!I;�.I;??I;�SI;�lI;��I;4�I;��I;��I;��I;�jI;�kH;�F;;C;j(>;0�6;��,;o ;;Q;��:s��:��:��u:�":���9�9��-�      Y��:��:�
�:��:��:�O ;�d;�U;\~#;!d-;��5;�g<;nsA;sE;�dG;S�H;N�I;(�I;	�I;1�I;4�I;�I;"oI;aVI;BI;X1I;�#I;�I;�I;VI;�I;�H;��H;�H;f�H;?�H;��H;?�H;f�H;�H;��H;�H;�I;VI;�I;�I;�#I;X1I;BI;aVI;"oI;�I;4�I;1�I;	�I;(�I;N�I;S�H;�dG;sE;nsA;�g<;��5;!d-;\~#;�U;�d;�O ;��:��:�
�:��:      _;;X�;��;$ ;�&;�[,;�2;.88;�.=;�EA;�qD;s�F;,IH;w8I;J�I;��I;s�I;�I;��I;��I;"oI;bWI;�CI;3I;s%I;8I;�I;�	I;�I;��H;��H;��H;��H;H�H;V�H;�H;V�H;H�H;��H;��H;��H;��H;�I;�	I;�I;8I;s%I;3I;�CI;bWI;"oI;��I;��I;�I;s�I;��I;J�I;w8I;,IH;s�F;�qD;�EA;�.=;.88;�2;�[,;�&;$ ;��;X�;;      ��0;�41;!�2;]�4;�/7;6":;	/=;�@;�B;�E;��F;h$H;�I;p�I;��I;��I;��I;�I;}�I;�I;�lI;aVI;�CI;�3I;Y&I;EI;I;�
I;II;>�H;A�H;��H;��H;��H;p�H;��H;w�H;��H;p�H;��H;��H;��H;A�H;>�H;II;�
I;I;EI;Y&I;�3I;�CI;aVI;�lI;�I;}�I;�I;��I;��I;��I;p�I;�I;h$H;��F;�E;�B;�@;	/=;6":;�/7;]�4;!�2;�41;      ��?;��?;��@;�sA; �B;[�C;�AE;t�F;��G;wH;�I;�I;��I;��I;U�I;��I;,�I;L�I;#�I;-hI;�SI;BI;3I;Y&I;�I;�I;)I;�I;��H;��H;&�H;z�H;p�H;��H;��H;5�H;�H;5�H;��H;��H;p�H;z�H;&�H;��H;��H;�I;)I;�I;�I;Y&I;3I;BI;�SI;-hI;#�I;L�I;,�I;��I;U�I;��I;��I;�I;�I;wH;��G;t�F;�AE;[�C; �B;�sA;��@;��?;      �F;m�F;�F;�1G;`�G;!%H;|�H;�I;lI;��I;r�I;��I;��I;��I;��I;ȨI;��I;�vI;�aI;COI;??I;X1I;s%I;EI;�I;OI;1I; I;��H;U�H;��H;c�H;��H;4�H;e�H;��H;��H;��H;e�H;4�H;��H;c�H;��H;U�H;��H; I;1I;OI;�I;EI;s%I;X1I;??I;COI;�aI;�vI;��I;ȨI;��I;��I;��I;��I;r�I;��I;lI;�I;|�H;!%H;`�G;�1G;�F;m�F;      tI;N&I;:I;�WI;{I;1�I;��I;�I;-�I;-�I;p�I;��I;��I;�I;_�I;$�I;�kI;�YI;}II;7;I;�.I;�#I;8I;I;)I;1I; I;��H;~�H;��H;\�H;a�H;��H;��H;�H;��H;w�H;��H;�H;��H;��H;a�H;\�H;��H;~�H;��H; I;1I;)I;I;8I;�#I;�.I;7;I;}II;�YI;�kI;$�I;_�I;�I;��I;��I;p�I;-�I;-�I;�I;��I;1�I;{I;�WI;:I;N&I;      �I;��I;�I;��I;�I;D�I;��I;b�I;"�I;��I;ŽI;&�I;6�I;��I;�pI;�_I;�PI;�BI;>6I;+I;8!I;�I;�I;�
I;�I; I;��H;y�H;��H;c�H;a�H;��H;��H;��H;��H;��H;y�H;��H;��H;��H;��H;��H;a�H;c�H;��H;y�H;��H; I;�I;�
I;�I;�I;8!I;+I;>6I;�BI;�PI;�_I;�pI;��I;6�I;&�I;ŽI;��I;"�I;b�I;��I;D�I;�I;��I;�I;��I;      ��I;7�I;�I;r�I;��I;��I;��I;K�I;L�I; �I;��I;&I;�oI;zaI;�SI;GI;D;I;�0I;�&I;3I;nI;�I;�	I;II;��H;��H;~�H;��H;X�H;[�H;��H;Z�H;L�H;��H;��H;��H;��H;��H;��H;��H;L�H;Z�H;��H;[�H;X�H;��H;~�H;��H;��H;II;�	I;�I;nI;3I;�&I;�0I;D;I;GI;�SI;zaI;�oI;&I;��I; �I;L�I;K�I;��I;��I;��I;r�I;�I;7�I;      H�I;Z�I;��I;)�I;զI;�I;֕I;��I;��I;6uI;�iI;�]I;�RI;�GI;=I;�3I;�*I;g"I;�I;�I;�I;VI;�I;>�H;��H;U�H;��H;c�H;[�H;��H;6�H;�H;B�H;��H;�H;��H;��H;��H;�H;��H;B�H;�H;6�H;��H;[�H;c�H;��H;U�H;��H;>�H;�I;VI;�I;�I;�I;g"I;�*I;�3I;=I;�GI;�RI;�]I;�iI;6uI;��I;��I;֕I;�I;զI;)�I;��I;Z�I;      ��I;ąI;��I;�I;]{I;�uI;�nI;%gI;�^I;�VI;�MI;(EI;�<I;G4I;W,I;�$I;�I;DI;GI;�I;�I;�I;��H;A�H;&�H;��H;\�H;a�H;��H;6�H;�H;�H;\�H;��H;z�H;7�H;��H;7�H;z�H;��H;\�H;�H;�H;6�H;��H;a�H;\�H;��H;&�H;A�H;��H;�I;�I;�I;GI;DI;�I;�$I;W,I;G4I;�<I;(EI;�MI;�VI;�^I;%gI;�nI;�uI;]{I;�I;��I;ąI;      ucI;�bI;qaI;�^I;Z[I;�VI;�QI;.LI;!FI;�?I;.9I;r2I;�+I;~%I;KI;cI;�I;�I;�	I;�I;�I;�H;��H;��H;z�H;c�H;a�H;��H;Z�H;�H;�H;U�H;��H;,�H;��H;��H;��H;��H;��H;,�H;��H;U�H;�H;�H;Z�H;��H;a�H;c�H;z�H;��H;��H;�H;�I;�I;�	I;�I;�I;cI;KI;~%I;�+I;r2I;.9I;�?I;!FI;.LI;�QI;�VI;Z[I;�^I;qaI;�bI;      �JI;]JI;II;GI;hDI;AI;/=I;�8I;4I;/I;�)I;�$I;�I;�I;�I;�I;|I;EI;OI;� I;��H;��H;��H;��H;p�H;��H;��H;��H;L�H;B�H;\�H;��H;�H;��H;M�H;!�H;3�H;!�H;M�H;��H;�H;��H;\�H;B�H;L�H;��H;��H;��H;p�H;��H;��H;��H;��H;� I;OI;EI;|I;�I;�I;�I;�I;�$I;�)I;/I;4I;�8I;/=I;AI;hDI;GI;II;]JI;      �8I;�8I;�7I;A6I;<4I;�1I;|.I;+I;C'I;B#I;I;�I;�I;�I;�I;�
I;�I;�I;O I;F�H;��H;�H;��H;��H;��H;4�H;��H;��H;��H;��H;��H;,�H;��H;<�H;��H;��H;��H;��H;��H;<�H;��H;,�H;��H;��H;��H;��H;��H;4�H;��H;��H;��H;�H;��H;F�H;O I;�I;�I;�
I;�I;�I;�I;�I;I;B#I;C'I;+I;|.I;�1I;<4I;A6I;�7I;�8I;      �-I;E-I;~,I;+I;X)I;3'I;�$I;�!I;�I;_I;�I;}I;�I;XI;�	I;�I;[I;N I;{�H;��H;��H;f�H;H�H;p�H;��H;e�H;�H;��H;��H;�H;z�H;��H;M�H;��H;��H;��H;�H;��H;��H;��H;M�H;��H;z�H;�H;��H;��H;�H;e�H;��H;p�H;H�H;f�H;��H;��H;{�H;N I;[I;�I;�	I;XI;�I;}I;�I;_I;�I;�!I;�$I;3'I;X)I;+I;~,I;E-I;      �&I;�&I;�%I;�$I;R#I;c!I;I;�I;�I;�I;�I;�I;`I;<
I;+I;*I;CI;�H;��H;��H;c�H;?�H;V�H;��H;5�H;��H;��H;��H;��H;��H;7�H;��H;!�H;��H;��H;k�H;r�H;k�H;��H;��H;!�H;��H;7�H;��H;��H;��H;��H;��H;5�H;��H;V�H;?�H;c�H;��H;��H;�H;CI;*I;+I;<
I;`I;�I;�I;�I;�I;�I;I;c!I;R#I;�$I;�%I;�&I;      �$I;�$I;�#I;�"I;G!I;}I;cI;�I;)I;TI;iI;QI;WI;7	I;'I;]I;� I;�H;��H;�H;��H;��H;�H;w�H;�H;��H;w�H;y�H;��H;��H;��H;��H;3�H;��H;�H;r�H;w�H;r�H;�H;��H;3�H;��H;��H;��H;��H;y�H;w�H;��H;�H;w�H;�H;��H;��H;�H;��H;�H;� I;]I;'I;7	I;WI;QI;iI;TI;)I;�I;cI;}I;G!I;�"I;�#I;�$I;      �&I;�&I;�%I;�$I;R#I;c!I;I;�I;�I;�I;�I;�I;`I;<
I;+I;*I;CI;�H;��H;��H;c�H;?�H;V�H;��H;5�H;��H;��H;��H;��H;��H;7�H;��H;!�H;��H;��H;k�H;r�H;k�H;��H;��H;!�H;��H;7�H;��H;��H;��H;��H;��H;5�H;��H;V�H;?�H;c�H;��H;��H;�H;CI;*I;+I;<
I;`I;�I;�I;�I;�I;�I;I;c!I;R#I;�$I;�%I;�&I;      �-I;E-I;~,I;+I;X)I;3'I;�$I;�!I;�I;_I;�I;}I;�I;XI;�	I;�I;[I;N I;{�H;��H;��H;f�H;H�H;p�H;��H;e�H;�H;��H;��H;�H;z�H;��H;M�H;��H;��H;��H;�H;��H;��H;��H;M�H;��H;z�H;�H;��H;��H;�H;e�H;��H;p�H;H�H;f�H;��H;��H;{�H;N I;[I;�I;�	I;XI;�I;}I;�I;_I;�I;�!I;�$I;3'I;X)I;+I;~,I;E-I;      �8I;�8I;�7I;A6I;<4I;�1I;|.I;+I;C'I;B#I;I;�I;�I;�I;�I;�
I;�I;�I;O I;F�H;��H;�H;��H;��H;��H;4�H;��H;��H;��H;��H;��H;,�H;��H;<�H;��H;��H;��H;��H;��H;<�H;��H;,�H;��H;��H;��H;��H;��H;4�H;��H;��H;��H;�H;��H;F�H;O I;�I;�I;�
I;�I;�I;�I;�I;I;B#I;C'I;+I;|.I;�1I;<4I;A6I;�7I;�8I;      �JI;]JI;II;GI;hDI;AI;/=I;�8I;4I;/I;�)I;�$I;�I;�I;�I;�I;|I;EI;OI;� I;��H;��H;��H;��H;p�H;��H;��H;��H;L�H;B�H;\�H;��H;�H;��H;M�H;!�H;3�H;!�H;M�H;��H;�H;��H;\�H;B�H;L�H;��H;��H;��H;p�H;��H;��H;��H;��H;� I;OI;EI;|I;�I;�I;�I;�I;�$I;�)I;/I;4I;�8I;/=I;AI;hDI;GI;II;]JI;      ucI;�bI;qaI;�^I;Z[I;�VI;�QI;.LI;!FI;�?I;.9I;r2I;�+I;~%I;KI;cI;�I;�I;�	I;�I;�I;�H;��H;��H;z�H;c�H;a�H;��H;Z�H;�H;�H;U�H;��H;,�H;��H;��H;��H;��H;��H;,�H;��H;U�H;�H;�H;Z�H;��H;a�H;c�H;z�H;��H;��H;�H;�I;�I;�	I;�I;�I;cI;KI;~%I;�+I;r2I;.9I;�?I;!FI;.LI;�QI;�VI;Z[I;�^I;qaI;�bI;      ��I;ąI;��I;�I;]{I;�uI;�nI;%gI;�^I;�VI;�MI;(EI;�<I;G4I;W,I;�$I;�I;DI;GI;�I;�I;�I;��H;A�H;&�H;��H;\�H;a�H;��H;6�H;�H;�H;\�H;��H;z�H;7�H;��H;7�H;z�H;��H;\�H;�H;�H;6�H;��H;a�H;\�H;��H;&�H;A�H;��H;�I;�I;�I;GI;DI;�I;�$I;W,I;G4I;�<I;(EI;�MI;�VI;�^I;%gI;�nI;�uI;]{I;�I;��I;ąI;      H�I;Z�I;��I;)�I;զI;�I;֕I;��I;��I;6uI;�iI;�]I;�RI;�GI;=I;�3I;�*I;g"I;�I;�I;�I;VI;�I;>�H;��H;U�H;��H;c�H;[�H;��H;6�H;�H;B�H;��H;�H;��H;��H;��H;�H;��H;B�H;�H;6�H;��H;[�H;c�H;��H;U�H;��H;>�H;�I;VI;�I;�I;�I;g"I;�*I;�3I;=I;�GI;�RI;�]I;�iI;6uI;��I;��I;֕I;�I;զI;)�I;��I;Z�I;      ��I;7�I;�I;r�I;��I;��I;��I;K�I;L�I; �I;��I;&I;�oI;zaI;�SI;GI;D;I;�0I;�&I;3I;nI;�I;�	I;II;��H;��H;~�H;��H;X�H;[�H;��H;Z�H;L�H;��H;��H;��H;��H;��H;��H;��H;L�H;Z�H;��H;[�H;X�H;��H;~�H;��H;��H;II;�	I;�I;nI;3I;�&I;�0I;D;I;GI;�SI;zaI;�oI;&I;��I; �I;L�I;K�I;��I;��I;��I;r�I;�I;7�I;      �I;��I;�I;��I;�I;D�I;��I;b�I;"�I;��I;ŽI;&�I;6�I;��I;�pI;�_I;�PI;�BI;>6I;+I;8!I;�I;�I;�
I;�I; I;��H;y�H;��H;c�H;a�H;��H;��H;��H;��H;��H;y�H;��H;��H;��H;��H;��H;a�H;c�H;��H;y�H;��H; I;�I;�
I;�I;�I;8!I;+I;>6I;�BI;�PI;�_I;�pI;��I;6�I;&�I;ŽI;��I;"�I;b�I;��I;D�I;�I;��I;�I;��I;      tI;N&I;:I;�WI;{I;1�I;��I;�I;-�I;-�I;p�I;��I;��I;�I;_�I;$�I;�kI;�YI;}II;7;I;�.I;�#I;8I;I;)I;1I; I;��H;~�H;��H;\�H;a�H;��H;��H;�H;��H;w�H;��H;�H;��H;��H;a�H;\�H;��H;~�H;��H; I;1I;)I;I;8I;�#I;�.I;7;I;}II;�YI;�kI;$�I;_�I;�I;��I;��I;p�I;-�I;-�I;�I;��I;1�I;{I;�WI;:I;N&I;      �F;m�F;�F;�1G;`�G;!%H;|�H;�I;lI;��I;r�I;��I;��I;��I;��I;ȨI;��I;�vI;�aI;COI;??I;X1I;s%I;EI;�I;OI;1I; I;��H;U�H;��H;c�H;��H;4�H;e�H;��H;��H;��H;e�H;4�H;��H;c�H;��H;U�H;��H; I;1I;OI;�I;EI;s%I;X1I;??I;COI;�aI;�vI;��I;ȨI;��I;��I;��I;��I;r�I;��I;lI;�I;|�H;!%H;`�G;�1G;�F;m�F;      ��?;��?;��@;�sA; �B;[�C;�AE;t�F;��G;wH;�I;�I;��I;��I;U�I;��I;,�I;L�I;#�I;-hI;�SI;BI;3I;Y&I;�I;�I;)I;�I;��H;��H;&�H;z�H;p�H;��H;��H;5�H;�H;5�H;��H;��H;p�H;z�H;&�H;��H;��H;�I;)I;�I;�I;Y&I;3I;BI;�SI;-hI;#�I;L�I;,�I;��I;U�I;��I;��I;�I;�I;wH;��G;t�F;�AE;[�C; �B;�sA;��@;��?;      ��0;�41;!�2;]�4;�/7;6":;	/=;�@;�B;�E;��F;h$H;�I;p�I;��I;��I;��I;�I;}�I;�I;�lI;aVI;�CI;�3I;Y&I;EI;I;�
I;II;>�H;A�H;��H;��H;��H;p�H;��H;w�H;��H;p�H;��H;��H;��H;A�H;>�H;II;�
I;I;EI;Y&I;�3I;�CI;aVI;�lI;�I;}�I;�I;��I;��I;��I;p�I;�I;h$H;��F;�E;�B;�@;	/=;6":;�/7;]�4;!�2;�41;      _;;X�;��;$ ;�&;�[,;�2;.88;�.=;�EA;�qD;s�F;,IH;w8I;J�I;��I;s�I;�I;��I;��I;"oI;bWI;�CI;3I;s%I;8I;�I;�	I;�I;��H;��H;��H;��H;H�H;V�H;�H;V�H;H�H;��H;��H;��H;��H;�I;�	I;�I;8I;s%I;3I;�CI;bWI;"oI;��I;��I;�I;s�I;��I;J�I;w8I;,IH;s�F;�qD;�EA;�.=;.88;�2;�[,;�&;$ ;��;X�;;      Y��:��:�
�:��:��:�O ;�d;�U;\~#;!d-;��5;�g<;nsA;sE;�dG;S�H;N�I;(�I;	�I;1�I;4�I;�I;"oI;aVI;BI;X1I;�#I;�I;�I;VI;�I;�H;��H;�H;f�H;?�H;��H;?�H;f�H;�H;��H;�H;�I;VI;�I;�I;�#I;X1I;BI;aVI;"oI;�I;4�I;1�I;	�I;(�I;N�I;S�H;�dG;sE;nsA;�g<;��5;!d-;\~#;�U;�d;�O ;��:��:�
�:��:      >�p���-��9���9�":��u:��:s��:��:;Q;o ;��,;0�6;j(>;;C;�F;�kH;�jI;��I;��I;��I;4�I;��I;�lI;�SI;??I;�.I;8!I;nI;�I;�I;�I;��H;��H;��H;c�H;��H;c�H;��H;��H;��H;�I;�I;�I;nI;8!I;�.I;??I;�SI;�lI;��I;4�I;��I;��I;��I;�jI;�kH;�F;;C;j(>;0�6;��,;o ;;Q;��:s��:��:��u:�":���9�9��-�      q&�~!��5���|谺�O��LT��l�9��u:�!�:�E�:C;=~#;}61;P;;��A;�E;�#H;jUI;,�I;��I;1�I;��I;�I;-hI;COI;7;I;+I;3I;�I;�I;�I;� I;F�H;��H;��H;�H;��H;��H;F�H;� I;�I;�I;�I;3I;+I;7;I;COI;-hI;�I;��I;1�I;��I;,�I;jUI;�#H;�E;��A;P;;}61;=~#;C;�E�:�!�:��u:�l�9�LT��O�|谺���5�~!�      llٻ�Ի ǻ����W���n���+�I�Ժ�1�&�39[m:��:{�;�;�[,;��8;ք@;V\E;�	H;jUI;��I;	�I;�I;}�I;#�I;�aI;}II;>6I;�&I;�I;GI;�	I;OI;O I;{�H;��H;��H;��H;{�H;O I;OI;�	I;GI;�I;�&I;>6I;}II;�aI;#�I;}�I;�I;	�I;��I;jUI;�	H;V\E;ք@;��8;�[,;�;{�;��:[m:&�39�1�I�Ժ��+��n�W������ ǻ�Ի      �yY�,}U���I���7��� �G"�"�Ի;❻��T�$���#��m�9���:jj�:�;�);)07;D@;V\E;�#H;�jI;(�I;s�I;�I;L�I;�vI;�YI;�BI;�0I;g"I;DI;�I;EI;�I;N I;�H;�H;�H;N I;�I;EI;�I;DI;g"I;�0I;�BI;�YI;�vI;L�I;�I;s�I;(�I;�jI;�#H;V\E;D@;)07;�);�;jj�:���:�m�9�#�$���T�;❻"�ԻG"��� ���7���I�,}U�      "�ü�l������S��cߓ���{�e�M�҉ ����S�����B�"찺q�o���u:���:�Q;D�';)07;ք@;�E;�kH;N�I;��I;��I;,�I;��I;�kI;�PI;D;I;�*I;�I;�I;|I;�I;[I;CI;� I;CI;[I;�I;|I;�I;�I;�*I;D;I;�PI;�kI;��I;,�I;��I;��I;N�I;�kH;�E;ք@;)07;D�';�Q;���:��u:q�o�"찺��B�S������҉ �e�M���{�cߓ�S�������l��      �'��-$�r��l�,���.?ټ-w��_����yY�-l���Ի���[������ R:���:�Q;�);��8;��A;�F;S�H;J�I;��I;��I;ȨI;$�I;�_I;GI;�3I;�$I;cI;�I;�
I;�I;*I;]I;*I;�I;�
I;�I;cI;�$I;�3I;GI;�_I;$�I;ȨI;��I;��I;J�I;S�H;�F;��A;��8;�);�Q;���: R:����[�������Ի-l��yY�_���-w��.?ټ,���l�r���-$�      b+����k̀�?l��Q�8�2�T����6����@����>��2���V���2���� R:���:�;�[,;P;;;C;�dG;w8I;��I;U�I;��I;_�I;�pI;�SI;=I;W,I;KI;�I;�I;�	I;+I;'I;+I;�	I;�I;�I;KI;W,I;=I;�SI;�pI;_�I;��I;U�I;��I;w8I;�dG;;C;P;;�[,;�;���: R:���2��V���2����>��@��6������T�8�2��Q�?l�k̀���      s�ཾhܽw�нfy��h什Y ��-l��n<�`���>ټ�𛼝|U����H᝻�2�������u:jj�:�;}61;j(>;sE;,IH;p�I;��I;��I;�I;��I;zaI;�GI;G4I;~%I;�I;�I;XI;<
I;7	I;<
I;XI;�I;�I;~%I;G4I;�GI;zaI;��I;�I;��I;��I;p�I;,IH;sE;j(>;}61;�;jj�:��u:�����2�H᝻����|U����>ټ`���n<�-l�Y ��h什fy��w�н�hܽ      ��4�j1�	�&������q�ཌྷ�������`��'�,��yR����]�����V��[��q�o����:{�;=~#;0�6;nsA;s�F;�I;��I;��I;��I;6�I;�oI;�RI;�<I;�+I;�I;�I;�I;`I;WI;`I;�I;�I;�I;�+I;�<I;�RI;�oI;6�I;��I;��I;��I;�I;s�F;nsA;0�6;=~#;{�;���:q�o�[���V�������]�yR��,��'��`��������q�������	�&�j1�      �x���o��ń�KUo���O�-�-�{��hܽd什�x��2��b��yR���|U��2�����"찺�m�9��:C;��,;�g<;�qD;h$H;�I;��I;��I;&�I;&I;�]I;(EI;r2I;�$I;�I;}I;�I;QI;�I;}I;�I;�$I;r2I;(EI;�]I;&I;&�I;��I;��I;�I;h$H;�qD;�g<;��,;C;��:�m�9"찺����2���|U�yR���b���2��x�d什�hܽ{�-�-���O�KUo�ń��o��      v���ྃ�Ѿ(����נ�	ń�<�S�
�#�gO���n��R̀��2�,������>���Ի��B��#�[m:�E�:o ;��5;�EA;��F;�I;r�I;p�I;ŽI;��I;�iI;�MI;.9I;�)I;I;�I;�I;iI;�I;�I;I;�)I;.9I;�MI;�iI;��I;ŽI;p�I;r�I;�I;��F;�EA;��5;o ;�E�:[m:�#���B���Ի��>���,���2�R̀��n��gO��
�#�<�S�	ń��נ�(�����Ѿ��      �3���/��X#��	��A��ՌȾ�f��JUo�`1�Ӱ���n���x��'��>ټ�@��-l�S���$��&�39�!�:;Q;!d-;�.=;�E;wH;��I;-�I;��I; �I;6uI;�VI;�?I;/I;B#I;_I;�I;TI;�I;_I;B#I;/I;�?I;�VI;6uI; �I;��I;-�I;��I;wH;�E;�.=;!d-;;Q;�!�:&�39$��S���-l��@���>ټ�'��x��n��Ӱ��`1�JUo��f��ՌȾ�A���	��X#���/�      ���S���Q�v��RZ�Z58�˂�p��d���hoy�`1�gO��d什�`�`��6����yY���컞�T��1���u:��:\~#;.88;�B;��G;lI;-�I;"�I;L�I;��I;�^I;!FI;4I;C'I;�I;�I;)I;�I;�I;C'I;4I;!FI;�^I;��I;L�I;"�I;-�I;lI;��G;�B;.88;\~#;��:��u:�1���T���컶yY�6���`���`�d什gO��`1�hoy�d���p��˂�Z58��RZ�Q�v�S���      Ŀ3g��$ﱿ���R����U��X#�r��d���JUo�
�#��hܽ����n<����_���҉ �;❻I�Ժ�l�9s��:�U;�2;�@;t�F;�I;�I;b�I;K�I;��I;%gI;.LI;�8I;+I;�!I;�I;�I;�I;�!I;+I;�8I;.LI;%gI;��I;K�I;b�I;�I;�I;t�F;�@;�2;�U;s��:�l�9I�Ժ;❻҉ �_�������n<�����hܽ
�#�JUo�d���r���X#��U�R������$ﱿ3g��      |x�N9�M��pؿkQ��c_��4�_��X#�p���f��<�S�{�����-l�T�-w��e�M�"�Ի��+��LT���:�d;�[,;	/=;�AE;|�H;��I;��I;��I;֕I;�nI;�QI;/=I;|.I;�$I;I;cI;I;�$I;|.I;/=I;�QI;�nI;֕I;��I;��I;��I;|�H;�AE;	/=;�[,;�d;��:�LT���+�"�Իe�M�-w��T�-l�����{�<�S��f��p���X#�4�_�c_��kQ��pؿM��N9�      �X1���,�e���<���2g��c_���U�˂�ՌȾ	ń�-�-�q��Y ��8�2�.?ټ��{�G"��n��O���u:�O ;�&;6":;[�C;!%H;1�I;D�I;��I;�I;�uI;�VI;AI;�1I;3'I;c!I;}I;c!I;3'I;�1I;AI;�VI;�uI;�I;��I;D�I;1�I;!%H;[�C;6":;�&;�O ;��u:�O��n�G"���{�.?ټ8�2�Y ��q��-�-�	ń�ՌȾ˂��U�c_��2g���<�e����,�      d��]]�1K��X1�Xf���kQ��R���Z58��A���נ���O���h什�Q�,���cߓ��� �W��|谺�":��:$ ;�/7; �B;`�G;{I;�I;��I;զI;]{I;Z[I;hDI;<4I;X)I;R#I;G!I;R#I;X)I;<4I;hDI;Z[I;]{I;զI;��I;�I;{I;`�G; �B;�/7;$ ;��:�":|谺W���� �cߓ�,����Q�h什����O��נ��A��Z58�R���kQ����Xf��X1�1K��]]�      L������4z���V��X1��<�pؿ����RZ��	�(���KUo����fy��?l�l�S����7������𺧽�9��:��;]�4;�sA;�1G;�WI;��I;r�I;)�I;�I;�^I;GI;A6I;+I;�$I;�"I;�$I;+I;A6I;GI;�^I;�I;)�I;r�I;��I;�WI;�1G;�sA;]�4;��;��:���9�𺘼����7�S��l�?l�fy�����KUo�(����	��RZ����pؿ�<��X1���V��4z�����      �o��c^���ē��4z�1K�e��M��$ﱿQ�v��X#���Ѿń�	�&�w�нk̀�r��������I� ǻ�5��9�
�:X�;!�2;��@;�F;:I;�I;�I;��I;��I;qaI;II;�7I;~,I;�%I;�#I;�%I;~,I;�7I;II;qaI;��I;��I;�I;�I;:I;�F;��@;!�2;X�;�
�:�9�5� ǻ��I�����r��k̀�w�н	�&�ń���Ѿ�X#�Q�v�$ﱿM��e��1K��4z��ē�c^��      o'���X��c^�������]]���,�N9�3g��S�����/����o��j1��hܽ���-$��l��,}U��Ի~!���-���:;�41;��?;m�F;N&I;��I;7�I;Z�I;ąI;�bI;]JI;�8I;E-I;�&I;�$I;�&I;E-I;�8I;]JI;�bI;ąI;Z�I;7�I;��I;N&I;m�F;��?;�41;;��:��-�~!��Ի,}U��l���-$����hܽj1��o���྘�/�S���3g��N9���,��]]�����c^���X��      ����,������Q���F�Q�Ù$�.���~�7�}�E(�>�׾�T���L+���սr����@L��jO�8�ͻ����l8�m�:��;U�1;��?;uF;s�H;��I;��I;��I;�uI;�VI;�@I;1I;�&I;� I;I;� I;�&I;1I;�@I;�VI;�uI;��I;��I;��I;s�H;uF;��?;U�1;��;�m�:�l8���8�ͻjO�@L����r����ս�L+��T��>�׾E(�7�}�~�.���Ù$�F�Q�Q��������,��      �,��^�� P���{��K��x �����n�����w��$���Ҿf��� (���ѽٷ��7����$�K��ɻ�� ��8���:��;��1;@;��F;.I;�I;4�I;ŝI;�tI;OVI;�@I;�0I;�&I;� I;�I;� I;�&I;�0I;�@I;OVI;�tI;ŝI;4�I;�I;.I;��F;@;��1;��;���: ��8���ɻ$�K����7�ٷ����ѽ (�f�����Ҿ�$���w�n��������x ��K��{� P��^��      ���� P�������d���;� ����㿰���#f�b��ž��z���C�ƽ40v�d5�R����o@����oj��Pu9_I�:>\;�63;@�@;�F;XI;��I;{�I;p�I;�rI;�TI;^?I;0I;&I;, I;MI;, I;&I;0I;^?I;�TI;�rI;p�I;{�I;��I;XI;�F;@�@;�63;>\;_I�:�Pu9oj�����o@�R���d5�40v�C�ƽ����z�žb��#f�������� ����;���d���� P��      Q����{���d��F�Ù$�7����ɿ,蒿��K�O���j�� Zb�H�8�����a����`���%�.� e��V�غ˨�9�W�:VW;�15;@�A;� G;[6I;��I;k�I;m�I;�oI;�RI;�=I;�.I;�$I;AI;OI;AI;�$I;�.I;�=I;�RI;�oI;m�I;k�I;��I;[6I;� G;@�A;�15;VW;�W�:˨�9V�غ e��%�.�`��������a�8���H� Zb��j��O����K�,蒿��ɿ7��Ù$��F���d��{�      F�Q��K���;�Ù$��;
��޿�����w�o,���澝���(�D������I��3�G�����N��Ǩ�1��9�����9:���:�m!;��7;۸B;}�G;
YI;L�I;��I;ّI;�kI;�OI;4;I;�,I;3#I;�I;�I;�I;3#I;�,I;4;I;�OI;�kI;ّI;��I;L�I;
YI;}�G;۸B;��7;�m!;���:��9:9���1��Ǩ��N�����3�G��I������(�D��������o,���w�����޿�;
�Ù$���;��K�      Ù$��x � ��7���޿m���ǅ����F�{�
��~����z��$���ս$���P2+���ϼWPp����J�]��*�#��:-�;�7';��:;�C;,H;�|I;?�I;��I;��I;�fI;�KI;:8I;V*I;E!I;I;GI;I;E!I;V*I;:8I;�KI;�fI;��I;��I;?�I;�|I;,H;�C;��:;�7';-�;#��:�*�J�]����WPp���ϼP2+�$�����ս�$���z��~��{�
���F�ǅ��m����޿7�� ���x �      .���������㿆�ɿ���ǅ����P�b��:�׾�`��U�H����@��a�a�!����!D�Gɻ�!������U�:�~;�H-;H{=;BBE;ȄH;)�I; �I;��I;ւI;�`I;BGI;�4I;�'I;�I; I;pI; I;�I;�'I;�4I;BGI;�`I;ւI;��I; �I;)�I;ȄH;BBE;H{=;�H-;�~;�U�:�����!�Gɻ!D���!��a�a��@����U�H��`��:�׾b����P�ǅ�������ɿ��㿯���      ~�n�������,蒿��w���F�b��Ȱ�����Yb�+����ѽ�%��'D4����@X��ʨ��H���轺P��9cp�:�; 93;;P@;�uF;9�H;&�I;��I;��I;�yI;�YI;3BI;�0I;�$I;eI;�I;@I;�I;eI;�$I;�0I;3BI;�YI;�yI;��I;��I;&�I;9�H;�uF;;P@; 93;�;cp�:P��9�轺�H��ʨ�@X�����'D4��%����ѽ+���Yb����Ȱ�b����F���w�,蒿����n���      7�}���w�#f���K�o,�{�
�:�׾�����k���'�lz꽥I���;V�LM�*����iO��G�mpE����c�:T� ;��$;̳8;r�B;�G;VJI;1�I;:�I;a�I;*pI;�RI;�<I;�,I;%!I;�I;9I;�I;9I;�I;%!I;�,I;�<I;�RI;*pI;a�I;:�I;1�I;VJI;�G;r�B;̳8;��$;T� ;c�:���mpE��G��iO�*���LM��;V��I��lz���'���k����:�׾{�
�o,���K�#f���w�      E(��$�b��O������~���`���Yb���'��U�N$��S�m�5����ϼ0�����_�����غ�0�9d��:F;�F.;3{=;bE;�[H;B�I;��I;��I;�I;%fI;&KI;7I;&(I;�I;�I;�I;DI;�I;�I;�I;&(I;7I;&KI;%fI;�I;��I;��I;B�I;�[H;bE;3{=;�F.;F;d��:�0�9��غ_������0����ϼ5��S�m�N$���U���'��Yb��`���~�����O��b���$�      >�׾��Ҿž�j��������z�U�H�+��lz�N$��0v�!2+����9���5�-ɻ34�0�����:���:Nn!;*O6;)kA;��F;��H;��I;��I;�I;k|I;�[I;~CI;%1I;�#I;�I;jI;�I;�I;�I;jI;�I;�#I;%1I;~CI;�[I;k|I;�I;��I;��I;��H;��F;)kA;*O6;Nn!;���:���:0��34�-ɻ�5�9�����!2+�0v�N$��lz�+��U�H���z������j��ž��Ҿ      �T��f�����z� Zb�(�D��$�����ѽ�I��S�m�!2+��������K��ﻙ�p�:�����9MR�:�.;��-;��<;iyD;uH;�lI;�I;��I;��I;�nI;�QI;�;I;!+I;�I;*I;OI;�I;�I;�I;OI;*I;�I;!+I;�;I;�QI;�nI;��I;��I;�I;�lI;uH;iyD;��<;��-;�.;MR�:��9:�����p��ﻍ�K������!2+�S�m��I����ѽ���$�(�D� Zb���z�f���      �L+� (���H�������ս�@���%���;V�5���������MS�������yF�%�n8o�:�;��$;^7;K�A;��F;�H;��I;��I;��I;��I;uaI;�GI;.4I;A%I;II;ZI;I;�	I; 	I;�	I;I;ZI;II;A%I;.4I;�GI;uaI;��I;��I;��I;��I;�H;��F;K�A;^7;��$;�;o�:%�n8yF⺦������MS�������5���;V��%���@����ս����H��� (�      ��ս��ѽC�ƽ8����I��$���a�a�'D4�LM���ϼ9����K�����G��]g�f�o���:�@�:�X;��1;kk>;�
E;/H;;pI;"�I;	�I;��I;!rI;�TI;>I;�,I;~I;�I;�I;�	I;/I;MI;/I;�	I;�I;�I;~I;�,I;>I;�TI;!rI;��I;	�I;"�I;;pI;/H;�
E;kk>;��1;�X;�@�:��:f�o�]g��G�������K�9����ϼLM�'D4�a�a�$����I��8���C�ƽ��ѽ      r��ٷ��40v���a�3�G�P2+�!�����*���0���5��ﻦ��]g��ହ�g:_�:�;1H-;3f;;NC;)RG;�I;�I;@�I;�I;%�I;+bI;�HI;�4I;�%I;�I;PI;�
I;�I;eI;sI;eI;�I;�
I;PI;�I;�%I;�4I;�HI;+bI;%�I;�I;@�I;�I;�I;)RG;NC;3f;;1H-;�;_�:�g:�ହ]g�������5�0��*������!��P2+�3�G���a�40v�ٷ��      ��7�d5���������ϼ��@X���iO����-ɻ��p�yF�f�o��g:^�:ZF;�*;�9;��A;�tF;<�H;�I;��I;ɺI;e�I;�oI;SSI;n=I;9,I;�I;�I;I;pI;�I;�I;� I;�I;�I;pI;I;�I;�I;9,I;n=I;SSI;�oI;e�I;ɺI;��I;�I;<�H;�tF;��A;�9;�*;ZF;^�:�g:f�o�yF⺙�p�-ɻ����iO�@X������ϼ������d5�7�      @L�����R���`����N��WPp�!D�ʨ��G�_���34�:���%�n8��:_�:ZF;�(;��7;v�@;��E;nPH;6lI;��I;�I;��I;C|I;�]I;�EI;�2I;�#I;{I;�I;		I;(I;� I;�H;h�H;�H;� I;(I;		I;�I;{I;�#I;�2I;�EI;�]I;C|I;��I;�I;��I;6lI;nPH;��E;v�@;��7;�(;ZF;_�:��:%�n8:���34�_����G�ʨ�!D�WPp��N��`���R������      jO�$�K��o@�%�.�Ǩ����Gɻ�H��mpE���غ0����9o�:�@�:�;�*;��7;�O@;�[E;H;�HI;��I;��I;)�I;|�I;ZgI;�MI;z9I;W)I;�I;�I;�
I;,I;'I;G�H;s�H;��H;s�H;G�H;'I;,I;�
I;�I;�I;W)I;z9I;�MI;ZgI;|�I;)�I;��I;��I;�HI;H;�[E;�O@;��7;�*;�;�@�:o�:��90����غmpE��H��Gɻ���Ǩ�%�.��o@�$�K�      8�ͻ�ɻ��� e��1��J�]��!��轺����0�9���:MR�:�;�X;1H-;�9;v�@;�[E;��G;Q4I;ֳI;d�I;��I;m�I;�oI;�TI;q?I;M.I;� I;�I;ZI;�I;�I;6�H;��H;,�H;��H;,�H;��H;6�H;�I;�I;ZI;�I;� I;M.I;q?I;�TI;�oI;m�I;��I;d�I;ֳI;Q4I;��G;�[E;v�@;�9;1H-;�X;�;MR�:���:�0�9����轺�!�J�]�1�� e������ɻ      �����oj�V�غ9����*�����P��9c�:d��:���:�.;��$;��1;3f;;��A;��E;H;Q4I;X�I;��I;m�I;��I;�uI;tZI;yDI;�2I;L$I;�I;�I;hI;�I;��H;t�H;7�H;��H;��H;��H;7�H;t�H;��H;�I;hI;�I;�I;L$I;�2I;yDI;tZI;�uI;��I;m�I;��I;X�I;Q4I;H;��E;��A;3f;;��1;��$;�.;���:d��:c�:P��9�����*�9���V�غoj���      �l8 ��8�Pu9˨�9��9:#��:�U�:cp�:T� ;F;Nn!;��-;^7;kk>;NC;�tF;nPH;�HI;ֳI;��I;кI;ԙI;�yI;�^I;aHI;e6I;}'I;vI;�I;1
I;�I;>�H;��H;��H;�H;��H;��H;��H;�H;��H;��H;>�H;�I;1
I;�I;vI;}'I;e6I;aHI;�^I;�yI;ԙI;кI;��I;ֳI;�HI;nPH;�tF;NC;kk>;^7;��-;Nn!;F;T� ;cp�:�U�:#��:��9:˨�9�Pu9 ��8      �m�:���:_I�:�W�:���:-�;�~;�;��$;�F.;*O6;��<;K�A;�
E;)RG;<�H;6lI;��I;d�I;m�I;ԙI;�zI;�`I;�JI;�8I;�)I;�I;�I;�I;9I; I;�H;��H;{�H; �H;�H;��H;�H; �H;{�H;��H;�H; I;9I;�I;�I;�I;�)I;�8I;�JI;�`I;�zI;ԙI;m�I;d�I;��I;6lI;<�H;)RG;�
E;K�A;��<;*O6;�F.;��$;�;�~;-�;���:�W�:_I�:���:      ��;��;>\;VW;�m!;�7';�H-; 93;̳8;3{=;)kA;iyD;��F;/H;�I;�I;��I;��I;��I;��I;�yI;�`I;�KI;4:I;+I;FI;8I;I;MI;� I;��H;�H;w�H;�H;�H;a�H;2�H;a�H;�H;�H;w�H;�H;��H;� I;MI;I;8I;FI;+I;4:I;�KI;�`I;�yI;��I;��I;��I;��I;�I;�I;/H;��F;iyD;)kA;3{=;̳8; 93;�H-;�7';�m!;VW;>\;��;      U�1;��1;�63;�15;��7;��:;H{=;;P@;r�B;bE;��F;uH;�H;;pI;�I;��I;�I;)�I;m�I;�uI;�^I;�JI;4:I;�+I; I;+I;�I;*I;�I;�H;��H;~�H;4�H;��H;{�H;��H;��H;��H;{�H;��H;4�H;~�H;��H;�H;�I;*I;�I;+I; I;�+I;4:I;�JI;�^I;�uI;m�I;)�I;�I;��I;�I;;pI;�H;uH;��F;bE;r�B;;P@;H{=;��:;��7;�15;�63;��1;      ��?;@;@�@;@�A;۸B;�C;BBE;�uF;�G;�[H;��H;�lI;��I;"�I;@�I;ɺI;��I;|�I;�oI;tZI;aHI;�8I;+I; I;�I;tI;�I;I;t�H;��H;��H;;�H;d�H;��H;��H;f�H;=�H;f�H;��H;��H;d�H;;�H;��H;��H;t�H;I;�I;tI;�I; I;+I;�8I;aHI;tZI;�oI;|�I;��I;ɺI;@�I;"�I;��I;�lI;��H;�[H;�G;�uF;BBE;�C;۸B;@�A;@�@;@;      uF;��F;�F;� G;}�G;,H;ȄH;9�H;VJI;B�I;��I;�I;��I;	�I;�I;e�I;C|I;ZgI;�TI;yDI;e6I;�)I;FI;+I;tI;�I;ZI;��H;��H;��H;6�H;I�H;��H;j�H;��H;$�H;��H;$�H;��H;j�H;��H;I�H;6�H;��H;��H;��H;ZI;�I;tI;+I;FI;�)I;e6I;yDI;�TI;ZgI;C|I;e�I;�I;	�I;��I;�I;��I;B�I;VJI;9�H;ȄH;,H;}�G;� G;�F;��F;      s�H;.I;XI;[6I;
YI;�|I;)�I;&�I;1�I;��I;��I;��I;��I;��I;%�I;�oI;�]I;�MI;q?I;�2I;}'I;�I;8I;�I;�I;ZI;��H;2�H;��H;@�H;1�H;s�H;&�H;#�H;��H;�H;��H;�H;��H;#�H;&�H;s�H;1�H;@�H;��H;2�H;��H;ZI;�I;�I;8I;�I;}'I;�2I;q?I;�MI;�]I;�oI;%�I;��I;��I;��I;��I;��I;1�I;&�I;)�I;�|I;
YI;[6I;XI;.I;      ��I;�I;��I;��I;L�I;?�I; �I;��I;:�I;��I;�I;��I;��I;!rI;+bI;SSI;�EI;z9I;M.I;L$I;vI;�I;I;*I;I;��H;2�H;�H;M�H;-�H;e�H;��H;��H;�H;b�H;	�H;��H;	�H;b�H;�H;��H;��H;e�H;-�H;M�H;�H;2�H;��H;I;*I;I;�I;vI;L$I;M.I;z9I;�EI;SSI;+bI;!rI;��I;��I;�I;��I;:�I;��I; �I;?�I;L�I;��I;��I;�I;      ��I;4�I;{�I;k�I;��I;��I;��I;��I;a�I;�I;k|I;�nI;uaI;�TI;�HI;n=I;�2I;W)I;� I;�I;�I;�I;MI;�I;t�H;��H;��H;M�H;8�H;a�H;��H;��H;��H;�H;��H;<�H;5�H;<�H;��H;�H;��H;��H;��H;a�H;8�H;M�H;��H;��H;t�H;�I;MI;�I;�I;�I;� I;W)I;�2I;n=I;�HI;�TI;uaI;�nI;k|I;�I;a�I;��I;��I;��I;��I;k�I;{�I;4�I;      ��I;ŝI;p�I;m�I;ّI;��I;ւI;�yI;*pI;%fI;�[I;�QI;�GI;>I;�4I;9,I;�#I;�I;�I;�I;1
I;9I;� I;�H;��H;��H;@�H;-�H;a�H;��H;��H;��H;��H;"�H;��H;��H;c�H;��H;��H;"�H;��H;��H;��H;��H;a�H;-�H;@�H;��H;��H;�H;� I;9I;1
I;�I;�I;�I;�#I;9,I;�4I;>I;�GI;�QI;�[I;%fI;*pI;�yI;ւI;��I;ّI;m�I;p�I;ŝI;      �uI;�tI;�rI;�oI;�kI;�fI;�`I;�YI;�RI;&KI;~CI;�;I;.4I;�,I;�%I;�I;{I;�I;ZI;hI;�I; I;��H;��H;��H;6�H;1�H;e�H;��H;��H;��H;��H;��H;c�H;�H;��H;��H;��H;�H;c�H;��H;��H;��H;��H;��H;e�H;1�H;6�H;��H;��H;��H; I;�I;hI;ZI;�I;{I;�I;�%I;�,I;.4I;�;I;~CI;&KI;�RI;�YI;�`I;�fI;�kI;�oI;�rI;�tI;      �VI;OVI;�TI;�RI;�OI;�KI;BGI;3BI;�<I;7I;%1I;!+I;A%I;~I;�I;�I;�I;�
I;�I;�I;>�H;�H;�H;~�H;;�H;I�H;s�H;��H;��H;��H;��H;��H;K�H;��H;��H;J�H;P�H;J�H;��H;��H;K�H;��H;��H;��H;��H;��H;s�H;I�H;;�H;~�H;�H;�H;>�H;�I;�I;�
I;�I;�I;�I;~I;A%I;!+I;%1I;7I;�<I;3BI;BGI;�KI;�OI;�RI;�TI;OVI;      �@I;�@I;^?I;�=I;4;I;:8I;�4I;�0I;�,I;&(I;�#I;�I;II;�I;PI;I;		I;,I;�I;��H;��H;��H;w�H;4�H;d�H;��H;&�H;��H;��H;��H;��H;K�H;��H;d�H;�H;��H;��H;��H;�H;d�H;��H;K�H;��H;��H;��H;��H;&�H;��H;d�H;4�H;w�H;��H;��H;��H;�I;,I;		I;I;PI;�I;II;�I;�#I;&(I;�,I;�0I;�4I;:8I;4;I;�=I;^?I;�@I;      1I;�0I;0I;�.I;�,I;V*I;�'I;�$I;%!I;�I;�I;*I;ZI;�I;�
I;pI;(I;'I;6�H;t�H;��H;{�H;�H;��H;��H;j�H;#�H;�H;�H;"�H;c�H;��H;d�H;��H;��H;��H;��H;��H;��H;��H;d�H;��H;c�H;"�H;�H;�H;#�H;j�H;��H;��H;�H;{�H;��H;t�H;6�H;'I;(I;pI;�
I;�I;ZI;*I;�I;�I;%!I;�$I;�'I;V*I;�,I;�.I;0I;�0I;      �&I;�&I;&I;�$I;3#I;E!I;�I;eI;�I;�I;jI;OI;I;�	I;�I;�I;� I;G�H;��H;7�H;�H; �H;�H;{�H;��H;��H;��H;b�H;��H;��H;�H;��H;�H;��H;��H;d�H;[�H;d�H;��H;��H;�H;��H;�H;��H;��H;b�H;��H;��H;��H;{�H;�H; �H;�H;7�H;��H;G�H;� I;�I;�I;�	I;I;OI;jI;�I;�I;eI;�I;E!I;3#I;�$I;&I;�&I;      � I;� I;, I;AI;�I;I; I;�I;9I;�I;�I;�I;�	I;/I;eI;�I;�H;s�H;,�H;��H;��H;�H;a�H;��H;f�H;$�H;�H;	�H;<�H;��H;��H;J�H;��H;��H;d�H;2�H;/�H;2�H;d�H;��H;��H;J�H;��H;��H;<�H;	�H;�H;$�H;f�H;��H;a�H;�H;��H;��H;,�H;s�H;�H;�I;eI;/I;�	I;�I;�I;�I;9I;�I; I;I;�I;AI;, I;� I;      I;�I;MI;OI;�I;GI;pI;@I;�I;DI;�I;�I; 	I;MI;sI;� I;h�H;��H;��H;��H;��H;��H;2�H;��H;=�H;��H;��H;��H;5�H;c�H;��H;P�H;��H;��H;[�H;/�H;�H;/�H;[�H;��H;��H;P�H;��H;c�H;5�H;��H;��H;��H;=�H;��H;2�H;��H;��H;��H;��H;��H;h�H;� I;sI;MI; 	I;�I;�I;DI;�I;@I;pI;GI;�I;OI;MI;�I;      � I;� I;, I;AI;�I;I; I;�I;9I;�I;�I;�I;�	I;/I;eI;�I;�H;s�H;,�H;��H;��H;�H;a�H;��H;f�H;$�H;�H;	�H;<�H;��H;��H;J�H;��H;��H;d�H;2�H;/�H;2�H;d�H;��H;��H;J�H;��H;��H;<�H;	�H;�H;$�H;f�H;��H;a�H;�H;��H;��H;,�H;s�H;�H;�I;eI;/I;�	I;�I;�I;�I;9I;�I; I;I;�I;AI;, I;� I;      �&I;�&I;&I;�$I;3#I;E!I;�I;eI;�I;�I;jI;OI;I;�	I;�I;�I;� I;G�H;��H;7�H;�H; �H;�H;{�H;��H;��H;��H;b�H;��H;��H;�H;��H;�H;��H;��H;d�H;[�H;d�H;��H;��H;�H;��H;�H;��H;��H;b�H;��H;��H;��H;{�H;�H; �H;�H;7�H;��H;G�H;� I;�I;�I;�	I;I;OI;jI;�I;�I;eI;�I;E!I;3#I;�$I;&I;�&I;      1I;�0I;0I;�.I;�,I;V*I;�'I;�$I;%!I;�I;�I;*I;ZI;�I;�
I;pI;(I;'I;6�H;t�H;��H;{�H;�H;��H;��H;j�H;#�H;�H;�H;"�H;c�H;��H;d�H;��H;��H;��H;��H;��H;��H;��H;d�H;��H;c�H;"�H;�H;�H;#�H;j�H;��H;��H;�H;{�H;��H;t�H;6�H;'I;(I;pI;�
I;�I;ZI;*I;�I;�I;%!I;�$I;�'I;V*I;�,I;�.I;0I;�0I;      �@I;�@I;^?I;�=I;4;I;:8I;�4I;�0I;�,I;&(I;�#I;�I;II;�I;PI;I;		I;,I;�I;��H;��H;��H;w�H;4�H;d�H;��H;&�H;��H;��H;��H;��H;K�H;��H;d�H;�H;��H;��H;��H;�H;d�H;��H;K�H;��H;��H;��H;��H;&�H;��H;d�H;4�H;w�H;��H;��H;��H;�I;,I;		I;I;PI;�I;II;�I;�#I;&(I;�,I;�0I;�4I;:8I;4;I;�=I;^?I;�@I;      �VI;OVI;�TI;�RI;�OI;�KI;BGI;3BI;�<I;7I;%1I;!+I;A%I;~I;�I;�I;�I;�
I;�I;�I;>�H;�H;�H;~�H;;�H;I�H;s�H;��H;��H;��H;��H;��H;K�H;��H;��H;J�H;P�H;J�H;��H;��H;K�H;��H;��H;��H;��H;��H;s�H;I�H;;�H;~�H;�H;�H;>�H;�I;�I;�
I;�I;�I;�I;~I;A%I;!+I;%1I;7I;�<I;3BI;BGI;�KI;�OI;�RI;�TI;OVI;      �uI;�tI;�rI;�oI;�kI;�fI;�`I;�YI;�RI;&KI;~CI;�;I;.4I;�,I;�%I;�I;{I;�I;ZI;hI;�I; I;��H;��H;��H;6�H;1�H;e�H;��H;��H;��H;��H;��H;c�H;�H;��H;��H;��H;�H;c�H;��H;��H;��H;��H;��H;e�H;1�H;6�H;��H;��H;��H; I;�I;hI;ZI;�I;{I;�I;�%I;�,I;.4I;�;I;~CI;&KI;�RI;�YI;�`I;�fI;�kI;�oI;�rI;�tI;      ��I;ŝI;p�I;m�I;ّI;��I;ւI;�yI;*pI;%fI;�[I;�QI;�GI;>I;�4I;9,I;�#I;�I;�I;�I;1
I;9I;� I;�H;��H;��H;@�H;-�H;a�H;��H;��H;��H;��H;"�H;��H;��H;c�H;��H;��H;"�H;��H;��H;��H;��H;a�H;-�H;@�H;��H;��H;�H;� I;9I;1
I;�I;�I;�I;�#I;9,I;�4I;>I;�GI;�QI;�[I;%fI;*pI;�yI;ւI;��I;ّI;m�I;p�I;ŝI;      ��I;4�I;{�I;k�I;��I;��I;��I;��I;a�I;�I;k|I;�nI;uaI;�TI;�HI;n=I;�2I;W)I;� I;�I;�I;�I;MI;�I;t�H;��H;��H;M�H;8�H;a�H;��H;��H;��H;�H;��H;<�H;5�H;<�H;��H;�H;��H;��H;��H;a�H;8�H;M�H;��H;��H;t�H;�I;MI;�I;�I;�I;� I;W)I;�2I;n=I;�HI;�TI;uaI;�nI;k|I;�I;a�I;��I;��I;��I;��I;k�I;{�I;4�I;      ��I;�I;��I;��I;L�I;?�I; �I;��I;:�I;��I;�I;��I;��I;!rI;+bI;SSI;�EI;z9I;M.I;L$I;vI;�I;I;*I;I;��H;2�H;�H;M�H;-�H;e�H;��H;��H;�H;b�H;	�H;��H;	�H;b�H;�H;��H;��H;e�H;-�H;M�H;�H;2�H;��H;I;*I;I;�I;vI;L$I;M.I;z9I;�EI;SSI;+bI;!rI;��I;��I;�I;��I;:�I;��I; �I;?�I;L�I;��I;��I;�I;      s�H;.I;XI;[6I;
YI;�|I;)�I;&�I;1�I;��I;��I;��I;��I;��I;%�I;�oI;�]I;�MI;q?I;�2I;}'I;�I;8I;�I;�I;ZI;��H;2�H;��H;@�H;1�H;s�H;&�H;#�H;��H;�H;��H;�H;��H;#�H;&�H;s�H;1�H;@�H;��H;2�H;��H;ZI;�I;�I;8I;�I;}'I;�2I;q?I;�MI;�]I;�oI;%�I;��I;��I;��I;��I;��I;1�I;&�I;)�I;�|I;
YI;[6I;XI;.I;      uF;��F;�F;� G;}�G;,H;ȄH;9�H;VJI;B�I;��I;�I;��I;	�I;�I;e�I;C|I;ZgI;�TI;yDI;e6I;�)I;FI;+I;tI;�I;ZI;��H;��H;��H;6�H;I�H;��H;j�H;��H;$�H;��H;$�H;��H;j�H;��H;I�H;6�H;��H;��H;��H;ZI;�I;tI;+I;FI;�)I;e6I;yDI;�TI;ZgI;C|I;e�I;�I;	�I;��I;�I;��I;B�I;VJI;9�H;ȄH;,H;}�G;� G;�F;��F;      ��?;@;@�@;@�A;۸B;�C;BBE;�uF;�G;�[H;��H;�lI;��I;"�I;@�I;ɺI;��I;|�I;�oI;tZI;aHI;�8I;+I; I;�I;tI;�I;I;t�H;��H;��H;;�H;d�H;��H;��H;f�H;=�H;f�H;��H;��H;d�H;;�H;��H;��H;t�H;I;�I;tI;�I; I;+I;�8I;aHI;tZI;�oI;|�I;��I;ɺI;@�I;"�I;��I;�lI;��H;�[H;�G;�uF;BBE;�C;۸B;@�A;@�@;@;      U�1;��1;�63;�15;��7;��:;H{=;;P@;r�B;bE;��F;uH;�H;;pI;�I;��I;�I;)�I;m�I;�uI;�^I;�JI;4:I;�+I; I;+I;�I;*I;�I;�H;��H;~�H;4�H;��H;{�H;��H;��H;��H;{�H;��H;4�H;~�H;��H;�H;�I;*I;�I;+I; I;�+I;4:I;�JI;�^I;�uI;m�I;)�I;�I;��I;�I;;pI;�H;uH;��F;bE;r�B;;P@;H{=;��:;��7;�15;�63;��1;      ��;��;>\;VW;�m!;�7';�H-; 93;̳8;3{=;)kA;iyD;��F;/H;�I;�I;��I;��I;��I;��I;�yI;�`I;�KI;4:I;+I;FI;8I;I;MI;� I;��H;�H;w�H;�H;�H;a�H;2�H;a�H;�H;�H;w�H;�H;��H;� I;MI;I;8I;FI;+I;4:I;�KI;�`I;�yI;��I;��I;��I;��I;�I;�I;/H;��F;iyD;)kA;3{=;̳8; 93;�H-;�7';�m!;VW;>\;��;      �m�:���:_I�:�W�:���:-�;�~;�;��$;�F.;*O6;��<;K�A;�
E;)RG;<�H;6lI;��I;d�I;m�I;ԙI;�zI;�`I;�JI;�8I;�)I;�I;�I;�I;9I; I;�H;��H;{�H; �H;�H;��H;�H; �H;{�H;��H;�H; I;9I;�I;�I;�I;�)I;�8I;�JI;�`I;�zI;ԙI;m�I;d�I;��I;6lI;<�H;)RG;�
E;K�A;��<;*O6;�F.;��$;�;�~;-�;���:�W�:_I�:���:      �l8 ��8�Pu9˨�9��9:#��:�U�:cp�:T� ;F;Nn!;��-;^7;kk>;NC;�tF;nPH;�HI;ֳI;��I;кI;ԙI;�yI;�^I;aHI;e6I;}'I;vI;�I;1
I;�I;>�H;��H;��H;�H;��H;��H;��H;�H;��H;��H;>�H;�I;1
I;�I;vI;}'I;e6I;aHI;�^I;�yI;ԙI;кI;��I;ֳI;�HI;nPH;�tF;NC;kk>;^7;��-;Nn!;F;T� ;cp�:�U�:#��:��9:˨�9�Pu9 ��8      �����oj�V�غ9����*�����P��9c�:d��:���:�.;��$;��1;3f;;��A;��E;H;Q4I;X�I;��I;m�I;��I;�uI;tZI;yDI;�2I;L$I;�I;�I;hI;�I;��H;t�H;7�H;��H;��H;��H;7�H;t�H;��H;�I;hI;�I;�I;L$I;�2I;yDI;tZI;�uI;��I;m�I;��I;X�I;Q4I;H;��E;��A;3f;;��1;��$;�.;���:d��:c�:P��9�����*�9���V�غoj���      8�ͻ�ɻ��� e��1��J�]��!��轺����0�9���:MR�:�;�X;1H-;�9;v�@;�[E;��G;Q4I;ֳI;d�I;��I;m�I;�oI;�TI;q?I;M.I;� I;�I;ZI;�I;�I;6�H;��H;,�H;��H;,�H;��H;6�H;�I;�I;ZI;�I;� I;M.I;q?I;�TI;�oI;m�I;��I;d�I;ֳI;Q4I;��G;�[E;v�@;�9;1H-;�X;�;MR�:���:�0�9����轺�!�J�]�1�� e������ɻ      jO�$�K��o@�%�.�Ǩ����Gɻ�H��mpE���غ0����9o�:�@�:�;�*;��7;�O@;�[E;H;�HI;��I;��I;)�I;|�I;ZgI;�MI;z9I;W)I;�I;�I;�
I;,I;'I;G�H;s�H;��H;s�H;G�H;'I;,I;�
I;�I;�I;W)I;z9I;�MI;ZgI;|�I;)�I;��I;��I;�HI;H;�[E;�O@;��7;�*;�;�@�:o�:��90����غmpE��H��Gɻ���Ǩ�%�.��o@�$�K�      @L�����R���`����N��WPp�!D�ʨ��G�_���34�:���%�n8��:_�:ZF;�(;��7;v�@;��E;nPH;6lI;��I;�I;��I;C|I;�]I;�EI;�2I;�#I;{I;�I;		I;(I;� I;�H;h�H;�H;� I;(I;		I;�I;{I;�#I;�2I;�EI;�]I;C|I;��I;�I;��I;6lI;nPH;��E;v�@;��7;�(;ZF;_�:��:%�n8:���34�_����G�ʨ�!D�WPp��N��`���R������      ��7�d5���������ϼ��@X���iO����-ɻ��p�yF�f�o��g:^�:ZF;�*;�9;��A;�tF;<�H;�I;��I;ɺI;e�I;�oI;SSI;n=I;9,I;�I;�I;I;pI;�I;�I;� I;�I;�I;pI;I;�I;�I;9,I;n=I;SSI;�oI;e�I;ɺI;��I;�I;<�H;�tF;��A;�9;�*;ZF;^�:�g:f�o�yF⺙�p�-ɻ����iO�@X������ϼ������d5�7�      r��ٷ��40v���a�3�G�P2+�!�����*���0���5��ﻦ��]g��ହ�g:_�:�;1H-;3f;;NC;)RG;�I;�I;@�I;�I;%�I;+bI;�HI;�4I;�%I;�I;PI;�
I;�I;eI;sI;eI;�I;�
I;PI;�I;�%I;�4I;�HI;+bI;%�I;�I;@�I;�I;�I;)RG;NC;3f;;1H-;�;_�:�g:�ହ]g�������5�0��*������!��P2+�3�G���a�40v�ٷ��      ��ս��ѽC�ƽ8����I��$���a�a�'D4�LM���ϼ9����K�����G��]g�f�o���:�@�:�X;��1;kk>;�
E;/H;;pI;"�I;	�I;��I;!rI;�TI;>I;�,I;~I;�I;�I;�	I;/I;MI;/I;�	I;�I;�I;~I;�,I;>I;�TI;!rI;��I;	�I;"�I;;pI;/H;�
E;kk>;��1;�X;�@�:��:f�o�]g��G�������K�9����ϼLM�'D4�a�a�$����I��8���C�ƽ��ѽ      �L+� (���H�������ս�@���%���;V�5���������MS�������yF�%�n8o�:�;��$;^7;K�A;��F;�H;��I;��I;��I;��I;uaI;�GI;.4I;A%I;II;ZI;I;�	I; 	I;�	I;I;ZI;II;A%I;.4I;�GI;uaI;��I;��I;��I;��I;�H;��F;K�A;^7;��$;�;o�:%�n8yF⺦������MS�������5���;V��%���@����ս����H��� (�      �T��f�����z� Zb�(�D��$�����ѽ�I��S�m�!2+��������K��ﻙ�p�:�����9MR�:�.;��-;��<;iyD;uH;�lI;�I;��I;��I;�nI;�QI;�;I;!+I;�I;*I;OI;�I;�I;�I;OI;*I;�I;!+I;�;I;�QI;�nI;��I;��I;�I;�lI;uH;iyD;��<;��-;�.;MR�:��9:�����p��ﻍ�K������!2+�S�m��I����ѽ���$�(�D� Zb���z�f���      >�׾��Ҿž�j��������z�U�H�+��lz�N$��0v�!2+����9���5�-ɻ34�0�����:���:Nn!;*O6;)kA;��F;��H;��I;��I;�I;k|I;�[I;~CI;%1I;�#I;�I;jI;�I;�I;�I;jI;�I;�#I;%1I;~CI;�[I;k|I;�I;��I;��I;��H;��F;)kA;*O6;Nn!;���:���:0��34�-ɻ�5�9�����!2+�0v�N$��lz�+��U�H���z������j��ž��Ҿ      E(��$�b��O������~���`���Yb���'��U�N$��S�m�5����ϼ0�����_�����غ�0�9d��:F;�F.;3{=;bE;�[H;B�I;��I;��I;�I;%fI;&KI;7I;&(I;�I;�I;�I;DI;�I;�I;�I;&(I;7I;&KI;%fI;�I;��I;��I;B�I;�[H;bE;3{=;�F.;F;d��:�0�9��غ_������0����ϼ5��S�m�N$���U���'��Yb��`���~�����O��b���$�      7�}���w�#f���K�o,�{�
�:�׾�����k���'�lz꽥I���;V�LM�*����iO��G�mpE����c�:T� ;��$;̳8;r�B;�G;VJI;1�I;:�I;a�I;*pI;�RI;�<I;�,I;%!I;�I;9I;�I;9I;�I;%!I;�,I;�<I;�RI;*pI;a�I;:�I;1�I;VJI;�G;r�B;̳8;��$;T� ;c�:���mpE��G��iO�*���LM��;V��I��lz���'���k����:�׾{�
�o,���K�#f���w�      ~�n�������,蒿��w���F�b��Ȱ�����Yb�+����ѽ�%��'D4����@X��ʨ��H���轺P��9cp�:�; 93;;P@;�uF;9�H;&�I;��I;��I;�yI;�YI;3BI;�0I;�$I;eI;�I;@I;�I;eI;�$I;�0I;3BI;�YI;�yI;��I;��I;&�I;9�H;�uF;;P@; 93;�;cp�:P��9�轺�H��ʨ�@X�����'D4��%����ѽ+���Yb����Ȱ�b����F���w�,蒿����n���      .���������㿆�ɿ���ǅ����P�b��:�׾�`��U�H����@��a�a�!����!D�Gɻ�!������U�:�~;�H-;H{=;BBE;ȄH;)�I; �I;��I;ւI;�`I;BGI;�4I;�'I;�I; I;pI; I;�I;�'I;�4I;BGI;�`I;ւI;��I; �I;)�I;ȄH;BBE;H{=;�H-;�~;�U�:�����!�Gɻ!D���!��a�a��@����U�H��`��:�׾b����P�ǅ�������ɿ��㿯���      Ù$��x � ��7���޿m���ǅ����F�{�
��~����z��$���ս$���P2+���ϼWPp����J�]��*�#��:-�;�7';��:;�C;,H;�|I;?�I;��I;��I;�fI;�KI;:8I;V*I;E!I;I;GI;I;E!I;V*I;:8I;�KI;�fI;��I;��I;?�I;�|I;,H;�C;��:;�7';-�;#��:�*�J�]����WPp���ϼP2+�$�����ս�$���z��~��{�
���F�ǅ��m����޿7�� ���x �      F�Q��K���;�Ù$��;
��޿�����w�o,���澝���(�D������I��3�G�����N��Ǩ�1��9�����9:���:�m!;��7;۸B;}�G;
YI;L�I;��I;ّI;�kI;�OI;4;I;�,I;3#I;�I;�I;�I;3#I;�,I;4;I;�OI;�kI;ّI;��I;L�I;
YI;}�G;۸B;��7;�m!;���:��9:9���1��Ǩ��N�����3�G��I������(�D��������o,���w�����޿�;
�Ù$���;��K�      Q����{���d��F�Ù$�7����ɿ,蒿��K�O���j�� Zb�H�8�����a����`���%�.� e��V�غ˨�9�W�:VW;�15;@�A;� G;[6I;��I;k�I;m�I;�oI;�RI;�=I;�.I;�$I;AI;OI;AI;�$I;�.I;�=I;�RI;�oI;m�I;k�I;��I;[6I;� G;@�A;�15;VW;�W�:˨�9V�غ e��%�.�`��������a�8���H� Zb��j��O����K�,蒿��ɿ7��Ù$��F���d��{�      ���� P�������d���;� ����㿰���#f�b��ž��z���C�ƽ40v�d5�R����o@����oj��Pu9_I�:>\;�63;@�@;�F;XI;��I;{�I;p�I;�rI;�TI;^?I;0I;&I;, I;MI;, I;&I;0I;^?I;�TI;�rI;p�I;{�I;��I;XI;�F;@�@;�63;>\;_I�:�Pu9oj�����o@�R���d5�40v�C�ƽ����z�žb��#f�������� ����;���d���� P��      �,��^�� P���{��K��x �����n�����w��$���Ҿf��� (���ѽٷ��7����$�K��ɻ�� ��8���:��;��1;@;��F;.I;�I;4�I;ŝI;�tI;OVI;�@I;�0I;�&I;� I;�I;� I;�&I;�0I;�@I;OVI;�tI;ŝI;4�I;�I;.I;��F;@;��1;��;���: ��8���ɻ$�K����7�ٷ����ѽ (�f�����Ҿ�$���w�n��������x ��K��{� P��^��      ݶ��O���ά��(�_���7�w�}߿���~,b��V�*l¾Fx�c.���Ž��t�6�����*�?��N�����sx9���:��;��2;U?@;�eF;D�H;��I;��I;9{I;�ZI;�BI;#1I;�$I;�I;�I;NI;�I;�I;�$I;#1I;�BI;�ZI;9{I;��I;��I;D�H;�eF;U?@;��2;��;���:�sx9���N��*�?����6����t���Žc.�Fx�*l¾�V�~,b����}߿w���7�(�_�ά��O���      O���A���}��+Y��3�����$ڿ"����\����(���s��3�9�����p�p�p���<<����d������9}��:�;V$3;io@;yF;��H;�I;�I;�zI;sZI;yBI;�0I;t$I;EI;uI; I;uI;EI;t$I;�0I;yBI;sZI;�zI;�I;�I;��H;yF;io@;V$3;�;}��:���9d�������<<�p��p���p�9����3��s�(�������\�"���$ڿ����3��+Y�}�A���      ά��}�8tf��lG�Ң%��p�*�ʿV����>M����S����d�ɤ�̷�9�d��
��I��@�1���������9���:N;�T4;��@;�F;A�H;�I;ܙI;�xI;�XI;bAI;�/I;�#I;�I;�I;�I;�I;�I;�#I;�/I;bAI;�XI;�xI;ܙI;�I;A�H;�F;��@;�T4;N;���:��9������@�1��I���
�9�d�̷�ɤ��d�S�������>M�V���*�ʿ�p�Ң%��lG�8tf�}�      (�_��+Y��lG�f.�w���꿭���J䂿��5���󾋰��M�N�W��V��-�Q�*�������:i!��g��+󳺑:��:�;f06;��A;uG;I;Z�I;��I;�uI;qVI;�?I;�.I;�"I;�I;'I;�I;'I;�I;�"I;�.I;�?I;qVI;�uI;��I;Z�I;I;uG;��A;f06;�;��:�:+��g��:i!�����*���-�Q�V��W��M�N���������5�J䂿�������w�f.��lG��+Y�      ��7��3�Ң%�w��<����ſ�����\�9����Ͼ����`�3����z����9�z�ἷ���z��8}�ht�J�^:�)�:Ϣ#;��8;��B;ArG;�$I;јI;�I;$qI;7SI;=I;�,I;1!I;oI;I;�I;I;oI;1!I;�,I;=I;7SI;$qI;�I;јI;�$I;ArG;��B;��8;Ϣ#;�)�:J�^:ht��8}��z����z�Ἁ�9��z����`�3�������Ͼ9����\������ſ�<��w�Ң%��3�      w�����p������ſ!��{Ps���1�-r���d���d�}I�҈Ž��}�l*�fC��W�^�RC�e�D�#N๫��:��;�);.6;;KD;e�G;kGI;ΜI;ȎI;�kI;OI;�9I;3*I;9I;�I;�I;KI;�I;�I;9I;3*I;�9I;OI;�kI;ȎI;ΜI;kGI;e�G;KD;.6;;�);��;���:#N�e�D�RC�W�^�fC��l*���}�҈Ž}I��d��d��-r����1�{Ps�!����ſ��꿀p����      }߿�$ڿ*�ʿ�������{Ps�MX:����#l¾�ǆ���7����<5��$�Q�����t��85�������7��8ȼ:��;��.;��=;�DE;�XH;�gI;G�I;ڇI;GeI;@JI;E6I;a'I;�I;I;�I;�I;�I;I;�I;a'I;E6I;@JI;GeI;ڇI;G�I;�gI;�XH;�DE;��=;��.;��;ȼ:7��8������85��t�����$�Q�<5�������7��ǆ�#l¾���MX:�{Ps��������*�ʿ�$ڿ      ���"��V���J䂿��\���1�����J˾睒�C�N�y��L������c�'���Ҽ �|��z�ko��z��*�&:�N�:̧;�V4;�@;HfF;��H;.�I;B�I;UI;=^I;�DI;&2I;<$I;cI;�I;I;�I;I;�I;cI;<$I;&2I;�DI;=^I;UI;B�I;.�I;��H;HfF;�@;�V4;̧;�N�:*�&:z��ko���z� �|���Ҽc�'����L���y��C�N�睒��J˾�����1���\�J䂿V���"��      ~,b���\��>M���5�9��-r��#l¾睒�"&W��3�<Sؽ�z��fG�����I���?��̻z�-����L��:��;Ͽ&;C{9;�C;�cG;tI;]�I;r�I;ruI;�VI;O?I;�-I;� I;�I;yI;�I;�I;�I;yI;�I;� I;�-I;O?I;�VI;ruI;r�I;]�I;tI;�cG;�C;C{9;Ͽ&;��;L��:���z�-��̻�?��I�����fG��z��<Sؽ�3�"&W�睒�#l¾-r��9����5��>M���\�      �V������������Ͼ�d���ǆ�C�N��3��c�[����\�@��EC��N�o�Ъ	�s숻/�Q��9K��:�g;o�/;\�=;bE;2H;�VI;ٜI;�I;�jI;�NI;G9I;)I;=I;�I;I;�I;�
I;�I;I;�I;=I;)I;G9I;�NI;�jI;�I;ٜI;�VI;2H;bE;\�=;o�/;�g;K��:Q��9/�s숻Ъ	�N�o�EC��@����\�[���cཱ3�C�N��ǆ��d����Ͼ���������      *l¾(��S������������d���7�y��<Sؽ[���d�P*�kּI\����'�����S������
�:�Y;�#;Z<7;N�A;2�F;|�H;��I;	�I;րI;	`I;�FI;3I;C$I;�I;�I;vI;i	I;iI;i	I;vI;�I;�I;C$I;3I;�FI;	`I;րI;	�I;��I;|�H;2�F;N�A;Z<7;�#;�Y;�
�:�����S������'�I\��kּP*��d�[��<Sؽy����7��d���������S���(��      Fx��s��d�M�N�`�3�}I����L����z����\�P*�'�ݼe���j<<��ڻ��V��gt�u�&:���:\B;�;/;oC=;��D;��G;8I;�I;ÓI;4sI;IUI;}>I;�,I;�I;�I;yI;�	I;I;.I;I;�	I;yI;�I;�I;�,I;}>I;IUI;4sI;ÓI;�I;8I;��G;��D;oC=;�;/;\B;���:u�&:�gt���V��ڻj<<�e���'�ݼP*���\��z��L������}I�`�3�M�N��d��s�      c.��3�ɤ�W����҈Ž<5�����fG�@��kּe���9yC�?�W7}�﮼�U�x9���:&	;O�&;�:8;��A;F;ϸH;WxI;��I;�I;PeI;�JI;m6I;�&I;�I;�I;uI;/I;�I;�I;�I;/I;uI;�I;�I;�&I;m6I;�JI;PeI;�I;��I;WxI;ϸH;F;��A;�:8;O�&;&	;���:U�x9﮼�W7}�?�9yC�e���kּ@��fG����<5��҈Ž��W��ɤ��3�      ��Ž9���̷�V���z����}�$�Q�c�'����EC��I\��j<<�?��n����0U�d��:[��:-�;�&3;��>;�E;�H;};I;�I;ÔI;�uI;�WI;�@I;�.I;� I;�I;I;oI;�I;<I;�I;<I;�I;oI;I;�I;� I;�.I;�@I;�WI;�uI;ÔI;�I;};I;�H;�E;��>;�&3;-�;[��:d��:0U����n��?�j<<�I\��EC�����c�'�$�Q���}��z��V��̷�9���      ��t���p�9�d�-�Q���9�l*������Ҽ�I��N�o���'��ڻW7}���eH��߄:�k�:¿;�.;5<;�nC;^6G;��H;�I;��I;�I;<eI;^KI;7I;�&I;�I;�I;i
I;dI;�I;��H;l�H;��H;�I;dI;i
I;�I;�I;�&I;7I;^KI;<eI;�I;��I;�I;��H;^6G;�nC;5<;�.;¿;�k�:�߄:eH���W7}��ڻ��'�N�o��I����Ҽ���l*���9�-�Q�9�d���p�      6��p��
�*���z��fC���t�� �|��?�Ъ	������V�﮼�0U��߄:��:�g;6�+;�9;��A;�eF;w�H;�^I;��I;��I; rI;�UI;�?I;�-I; I;uI;(I;�I;�I;i�H;��H;�H;��H;i�H;�I;�I;(I;uI; I;�-I;�?I;�UI; rI;��I;��I;�^I;w�H;�eF;��A;�9;6�+;�g;��:�߄:0U�﮼���V����Ъ	��?� �|��t��fC��z��*����
�p�      ���p���I���������W�^�85��z��̻s숻�S��gt�U�x9d��:�k�:�g;z�*;�8;�@; �E;W'H;�7I;ߒI;3�I;o}I;�_I;�GI;�4I;y%I;�I;RI;	I;�I;��H;�H;i�H;��H;i�H;�H;��H;�I;	I;RI;�I;y%I;�4I;�GI;�_I;o}I;3�I;ߒI;�7I;W'H; �E;�@;�8;z�*;�g;�k�:d��:U�x9�gt��S�s숻�̻�z�85�W�^���������I��p��      *�?��<<�@�1�:i!��z�RC����ko��z�-�/򳺬���u�&:���:[��:¿;6�+;�8;W�@;]E;��G;eI;
�I;l�I;P�I;�hI;UOI;#;I;�*I;�I;�I;nI;EI;� I;��H;��H;d�H;��H;d�H;��H;��H;� I;EI;nI;�I;�I;�*I;#;I;UOI;�hI;P�I;l�I;
�I;eI;��G;]E;W�@;�8;6�+;¿;[��:���:u�&:����/�z�-�ko�����RC��z�:i!�@�1��<<�      �N����������g���8}�e�D����z�����Q��9�
�:���:&	;-�;�.;�9;�@;]E;��G;]I;�~I;#�I;g�I;�oI;�UI;�@I;�/I;�!I;�I;I;I;�I;��H;s�H;��H;r�H;��H;r�H;��H;s�H;��H;�I;I;I;�I;�!I;�/I;�@I;�UI;�oI;g�I;#�I;�~I;]I;��G;]E;�@;�9;�.;-�;&	;���:�
�:Q��9���z�����e�D��8}��g���������      ��d�����+�ht�#N�7��8*�&:L��:K��:�Y;\B;O�&;�&3;5<;��A; �E;��G;]I;w{I;��I;��I;�tI;�ZI;*EI;�3I;E%I;�I;bI;�I;I;O�H;��H;I�H;��H;��H;1�H;��H;��H;I�H;��H;O�H;I;�I;bI;�I;E%I;�3I;*EI;�ZI;�tI;��I;��I;w{I;]I;��G; �E;��A;5<;�&3;O�&;\B;�Y;K��:L��:*�&:7��8#N�ht�+���d���      �sx9���9��9�:J�^:���:ȼ:�N�:��;�g;�#;�;/;�:8;��>;�nC;�eF;W'H;eI;�~I;��I;ːI;wI;�]I;RHI;�6I;(I;#I;�I;�
I;\I;b�H;]�H;h�H;L�H;��H;��H;��H;��H;��H;L�H;h�H;]�H;b�H;\I;�
I;�I;#I;(I;�6I;RHI;�]I;wI;ːI;��I;�~I;eI;W'H;�eF;�nC;��>;�:8;�;/;�#;�g;��;�N�:ȼ:���:J�^:�:��9���9      ���:}��:���:��:�)�:��;��;̧;Ͽ&;o�/;Z<7;oC=;��A;�E;^6G;w�H;�7I;
�I;#�I;��I;wI;�^I;�II;�8I;*I;I;LI;QI;�I;M I;�H;��H;*�H;M�H;��H;�H;��H;�H;��H;M�H;*�H;��H;�H;M I;�I;QI;LI;I;*I;�8I;�II;�^I;wI;��I;#�I;
�I;�7I;w�H;^6G;�E;��A;oC=;Z<7;o�/;Ͽ&;̧;��;��;�)�:��:���:}��:      ��;�;N;�;Ϣ#;�);��.;�V4;C{9;\�=;N�A;��D;F;�H;��H;�^I;ߒI;l�I;g�I;�tI;�]I;�II;>9I;6+I;VI;�I;gI;�I;4I;��H;�H;F�H;�H;{�H;p�H;��H;b�H;��H;p�H;{�H;�H;F�H;�H;��H;4I;�I;gI;�I;VI;6+I;>9I;�II;�]I;�tI;g�I;l�I;ߒI;�^I;��H;�H;F;��D;N�A;\�=;C{9;�V4;��.;�);Ϣ#;�;N;�;      ��2;V$3;�T4;f06;��8;.6;;��=;�@;�C;bE;2�F;��G;ϸH;};I;�I;��I;3�I;P�I;�oI;�ZI;RHI;�8I;6+I;�I;5I;2I;iI;�I;Y�H;t�H;q�H;:�H;L�H;��H;��H;i�H;�H;i�H;��H;��H;L�H;:�H;q�H;t�H;Y�H;�I;iI;2I;5I;�I;6+I;�8I;RHI;�ZI;�oI;P�I;3�I;��I;�I;};I;ϸH;��G;2�F;bE;�C;�@;��=;.6;;��8;f06;�T4;V$3;      U?@;io@;��@;��A;��B;KD;�DE;HfF;�cG;2H;|�H;8I;WxI;�I;��I;��I;o}I;�hI;�UI;*EI;�6I;*I;VI;5I;tI;�I;QI;��H;��H;��H;.�H;0�H;��H;}�H;��H;,�H;	�H;,�H;��H;}�H;��H;0�H;.�H;��H;��H;��H;QI;�I;tI;5I;VI;*I;�6I;*EI;�UI;�hI;o}I;��I;��I;�I;WxI;8I;|�H;2H;�cG;HfF;�DE;KD;��B;��A;��@;io@;      �eF;yF;�F;uG;ArG;e�G;�XH;��H;tI;�VI;��I;�I;��I;ÔI;�I; rI;�_I;UOI;�@I;�3I;(I;I;�I;2I;�I;jI;��H;�H;��H;b�H;?�H;q�H;#�H;9�H;|�H;�H;�H;�H;|�H;9�H;#�H;q�H;?�H;b�H;��H;�H;��H;jI;�I;2I;�I;I;(I;�3I;�@I;UOI;�_I; rI;�I;ÔI;��I;�I;��I;�VI;tI;��H;�XH;e�G;ArG;uG;�F;yF;      D�H;��H;A�H;I;�$I;kGI;�gI;.�I;]�I;ٜI;	�I;ÓI;�I;�uI;<eI;�UI;�GI;#;I;�/I;E%I;#I;LI;gI;iI;QI;��H;�H;��H;s�H;@�H;{�H; �H;��H;�H;q�H;�H;�H;�H;q�H;�H;��H; �H;{�H;@�H;s�H;��H;�H;��H;QI;iI;gI;LI;#I;E%I;�/I;#;I;�GI;�UI;<eI;�uI;�I;ÓI;	�I;ٜI;]�I;.�I;�gI;kGI;�$I;I;A�H;��H;      ��I;�I;�I;Z�I;јI;ΜI;G�I;B�I;r�I;�I;րI;4sI;PeI;�WI;^KI;�?I;�4I;�*I;�!I;�I;�I;QI;�I;�I;��H;�H;��H;l�H;Q�H;j�H;��H;��H;��H;�H;��H;H�H;1�H;H�H;��H;�H;��H;��H;��H;j�H;Q�H;l�H;��H;�H;��H;�I;�I;QI;�I;�I;�!I;�*I;�4I;�?I;^KI;�WI;PeI;4sI;րI;�I;r�I;B�I;G�I;ΜI;јI;Z�I;�I;�I;      ��I;�I;ܙI;��I;�I;ȎI;ڇI;UI;ruI;�jI;	`I;IUI;�JI;�@I;7I;�-I;y%I;�I;�I;bI;�
I;�I;4I;Y�H;��H;��H;s�H;Q�H;j�H;��H;��H;��H;��H;-�H;��H;��H;Y�H;��H;��H;-�H;��H;��H;��H;��H;j�H;Q�H;s�H;��H;��H;Y�H;4I;�I;�
I;bI;�I;�I;y%I;�-I;7I;�@I;�JI;IUI;	`I;�jI;ruI;UI;ڇI;ȎI;�I;��I;ܙI;�I;      9{I;�zI;�xI;�uI;$qI;�kI;GeI;=^I;�VI;�NI;�FI;}>I;m6I;�.I;�&I; I;�I;�I;I;�I;\I;M I;��H;t�H;��H;b�H;@�H;j�H;��H;��H;��H;��H;�H;��H;�H;��H;��H;��H;�H;��H;�H;��H;��H;��H;��H;j�H;@�H;b�H;��H;t�H;��H;M I;\I;�I;I;�I;�I; I;�&I;�.I;m6I;}>I;�FI;�NI;�VI;=^I;GeI;�kI;$qI;�uI;�xI;�zI;      �ZI;sZI;�XI;qVI;7SI;OI;@JI;�DI;O?I;G9I;3I;�,I;�&I;� I;�I;uI;RI;nI;I;I;b�H;�H;�H;q�H;.�H;?�H;{�H;��H;��H;��H;��H;��H;`�H;��H;|�H;c�H;Z�H;c�H;|�H;��H;`�H;��H;��H;��H;��H;��H;{�H;?�H;.�H;q�H;�H;�H;b�H;I;I;nI;RI;uI;�I;� I;�&I;�,I;3I;G9I;O?I;�DI;@JI;OI;7SI;qVI;�XI;sZI;      �BI;yBI;bAI;�?I;=I;�9I;E6I;&2I;�-I;)I;C$I;�I;�I;�I;�I;(I;	I;EI;�I;O�H;]�H;��H;F�H;:�H;0�H;q�H; �H;��H;��H;��H;��H;I�H;��H;U�H;�H;��H;��H;��H;�H;U�H;��H;I�H;��H;��H;��H;��H; �H;q�H;0�H;:�H;F�H;��H;]�H;O�H;�I;EI;	I;(I;�I;�I;�I;�I;C$I;)I;�-I;&2I;E6I;�9I;=I;�?I;bAI;yBI;      #1I;�0I;�/I;�.I;�,I;3*I;a'I;<$I;� I;=I;�I;�I;�I;I;i
I;�I;�I;� I;��H;��H;h�H;*�H;�H;L�H;��H;#�H;��H;��H;��H;�H;`�H;��H;9�H;��H;��H;��H;t�H;��H;��H;��H;9�H;��H;`�H;�H;��H;��H;��H;#�H;��H;L�H;�H;*�H;h�H;��H;��H;� I;�I;�I;i
I;I;�I;�I;�I;=I;� I;<$I;a'I;3*I;�,I;�.I;�/I;�0I;      �$I;t$I;�#I;�"I;1!I;9I;�I;cI;�I;�I;�I;yI;uI;oI;dI;�I;��H;��H;s�H;I�H;L�H;M�H;{�H;��H;}�H;9�H;�H;�H;-�H;��H;��H;U�H;��H;��H;b�H;@�H;)�H;@�H;b�H;��H;��H;U�H;��H;��H;-�H;�H;�H;9�H;}�H;��H;{�H;M�H;L�H;I�H;s�H;��H;��H;�I;dI;oI;uI;yI;�I;�I;�I;cI;�I;9I;1!I;�"I;�#I;t$I;      �I;EI;�I;�I;oI;�I;I;�I;yI;I;vI;�	I;/I;�I;�I;i�H;�H;��H;��H;��H;��H;��H;p�H;��H;��H;|�H;q�H;��H;��H;�H;|�H;�H;��H;b�H;�H;�H;�H;�H;�H;b�H;��H;�H;|�H;�H;��H;��H;q�H;|�H;��H;��H;p�H;��H;��H;��H;��H;��H;�H;i�H;�I;�I;/I;�	I;vI;I;yI;�I;I;�I;oI;�I;�I;EI;      �I;uI;�I;'I;I;�I;�I;I;�I;�I;i	I;I;�I;<I;��H;��H;i�H;d�H;r�H;��H;��H;�H;��H;i�H;,�H;�H;�H;H�H;��H;��H;c�H;��H;��H;@�H;�H;��H;��H;��H;�H;@�H;��H;��H;c�H;��H;��H;H�H;�H;�H;,�H;i�H;��H;�H;��H;��H;r�H;d�H;i�H;��H;��H;<I;�I;I;i	I;�I;�I;I;�I;�I;I;'I;�I;uI;      NI; I;�I;�I;�I;KI;�I;�I;�I;�
I;iI;.I;�I;�I;l�H;�H;��H;��H;��H;1�H;��H;��H;b�H;�H;	�H;�H;�H;1�H;Y�H;��H;Z�H;��H;t�H;)�H;�H;��H;��H;��H;�H;)�H;t�H;��H;Z�H;��H;Y�H;1�H;�H;�H;	�H;�H;b�H;��H;��H;1�H;��H;��H;��H;�H;l�H;�I;�I;.I;iI;�
I;�I;�I;�I;KI;�I;�I;�I; I;      �I;uI;�I;'I;I;�I;�I;I;�I;�I;i	I;I;�I;<I;��H;��H;i�H;d�H;r�H;��H;��H;�H;��H;i�H;,�H;�H;�H;H�H;��H;��H;c�H;��H;��H;@�H;�H;��H;��H;��H;�H;@�H;��H;��H;c�H;��H;��H;H�H;�H;�H;,�H;i�H;��H;�H;��H;��H;r�H;d�H;i�H;��H;��H;<I;�I;I;i	I;�I;�I;I;�I;�I;I;'I;�I;uI;      �I;EI;�I;�I;oI;�I;I;�I;yI;I;vI;�	I;/I;�I;�I;i�H;�H;��H;��H;��H;��H;��H;p�H;��H;��H;|�H;q�H;��H;��H;�H;|�H;�H;��H;b�H;�H;�H;�H;�H;�H;b�H;��H;�H;|�H;�H;��H;��H;q�H;|�H;��H;��H;p�H;��H;��H;��H;��H;��H;�H;i�H;�I;�I;/I;�	I;vI;I;yI;�I;I;�I;oI;�I;�I;EI;      �$I;t$I;�#I;�"I;1!I;9I;�I;cI;�I;�I;�I;yI;uI;oI;dI;�I;��H;��H;s�H;I�H;L�H;M�H;{�H;��H;}�H;9�H;�H;�H;-�H;��H;��H;U�H;��H;��H;b�H;@�H;)�H;@�H;b�H;��H;��H;U�H;��H;��H;-�H;�H;�H;9�H;}�H;��H;{�H;M�H;L�H;I�H;s�H;��H;��H;�I;dI;oI;uI;yI;�I;�I;�I;cI;�I;9I;1!I;�"I;�#I;t$I;      #1I;�0I;�/I;�.I;�,I;3*I;a'I;<$I;� I;=I;�I;�I;�I;I;i
I;�I;�I;� I;��H;��H;h�H;*�H;�H;L�H;��H;#�H;��H;��H;��H;�H;`�H;��H;9�H;��H;��H;��H;t�H;��H;��H;��H;9�H;��H;`�H;�H;��H;��H;��H;#�H;��H;L�H;�H;*�H;h�H;��H;��H;� I;�I;�I;i
I;I;�I;�I;�I;=I;� I;<$I;a'I;3*I;�,I;�.I;�/I;�0I;      �BI;yBI;bAI;�?I;=I;�9I;E6I;&2I;�-I;)I;C$I;�I;�I;�I;�I;(I;	I;EI;�I;O�H;]�H;��H;F�H;:�H;0�H;q�H; �H;��H;��H;��H;��H;I�H;��H;U�H;�H;��H;��H;��H;�H;U�H;��H;I�H;��H;��H;��H;��H; �H;q�H;0�H;:�H;F�H;��H;]�H;O�H;�I;EI;	I;(I;�I;�I;�I;�I;C$I;)I;�-I;&2I;E6I;�9I;=I;�?I;bAI;yBI;      �ZI;sZI;�XI;qVI;7SI;OI;@JI;�DI;O?I;G9I;3I;�,I;�&I;� I;�I;uI;RI;nI;I;I;b�H;�H;�H;q�H;.�H;?�H;{�H;��H;��H;��H;��H;��H;`�H;��H;|�H;c�H;Z�H;c�H;|�H;��H;`�H;��H;��H;��H;��H;��H;{�H;?�H;.�H;q�H;�H;�H;b�H;I;I;nI;RI;uI;�I;� I;�&I;�,I;3I;G9I;O?I;�DI;@JI;OI;7SI;qVI;�XI;sZI;      9{I;�zI;�xI;�uI;$qI;�kI;GeI;=^I;�VI;�NI;�FI;}>I;m6I;�.I;�&I; I;�I;�I;I;�I;\I;M I;��H;t�H;��H;b�H;@�H;j�H;��H;��H;��H;��H;�H;��H;�H;��H;��H;��H;�H;��H;�H;��H;��H;��H;��H;j�H;@�H;b�H;��H;t�H;��H;M I;\I;�I;I;�I;�I; I;�&I;�.I;m6I;}>I;�FI;�NI;�VI;=^I;GeI;�kI;$qI;�uI;�xI;�zI;      ��I;�I;ܙI;��I;�I;ȎI;ڇI;UI;ruI;�jI;	`I;IUI;�JI;�@I;7I;�-I;y%I;�I;�I;bI;�
I;�I;4I;Y�H;��H;��H;s�H;Q�H;j�H;��H;��H;��H;��H;-�H;��H;��H;Y�H;��H;��H;-�H;��H;��H;��H;��H;j�H;Q�H;s�H;��H;��H;Y�H;4I;�I;�
I;bI;�I;�I;y%I;�-I;7I;�@I;�JI;IUI;	`I;�jI;ruI;UI;ڇI;ȎI;�I;��I;ܙI;�I;      ��I;�I;�I;Z�I;јI;ΜI;G�I;B�I;r�I;�I;րI;4sI;PeI;�WI;^KI;�?I;�4I;�*I;�!I;�I;�I;QI;�I;�I;��H;�H;��H;l�H;Q�H;j�H;��H;��H;��H;�H;��H;H�H;1�H;H�H;��H;�H;��H;��H;��H;j�H;Q�H;l�H;��H;�H;��H;�I;�I;QI;�I;�I;�!I;�*I;�4I;�?I;^KI;�WI;PeI;4sI;րI;�I;r�I;B�I;G�I;ΜI;јI;Z�I;�I;�I;      D�H;��H;A�H;I;�$I;kGI;�gI;.�I;]�I;ٜI;	�I;ÓI;�I;�uI;<eI;�UI;�GI;#;I;�/I;E%I;#I;LI;gI;iI;QI;��H;�H;��H;s�H;@�H;{�H; �H;��H;�H;q�H;�H;�H;�H;q�H;�H;��H; �H;{�H;@�H;s�H;��H;�H;��H;QI;iI;gI;LI;#I;E%I;�/I;#;I;�GI;�UI;<eI;�uI;�I;ÓI;	�I;ٜI;]�I;.�I;�gI;kGI;�$I;I;A�H;��H;      �eF;yF;�F;uG;ArG;e�G;�XH;��H;tI;�VI;��I;�I;��I;ÔI;�I; rI;�_I;UOI;�@I;�3I;(I;I;�I;2I;�I;jI;��H;�H;��H;b�H;?�H;q�H;#�H;9�H;|�H;�H;�H;�H;|�H;9�H;#�H;q�H;?�H;b�H;��H;�H;��H;jI;�I;2I;�I;I;(I;�3I;�@I;UOI;�_I; rI;�I;ÔI;��I;�I;��I;�VI;tI;��H;�XH;e�G;ArG;uG;�F;yF;      U?@;io@;��@;��A;��B;KD;�DE;HfF;�cG;2H;|�H;8I;WxI;�I;��I;��I;o}I;�hI;�UI;*EI;�6I;*I;VI;5I;tI;�I;QI;��H;��H;��H;.�H;0�H;��H;}�H;��H;,�H;	�H;,�H;��H;}�H;��H;0�H;.�H;��H;��H;��H;QI;�I;tI;5I;VI;*I;�6I;*EI;�UI;�hI;o}I;��I;��I;�I;WxI;8I;|�H;2H;�cG;HfF;�DE;KD;��B;��A;��@;io@;      ��2;V$3;�T4;f06;��8;.6;;��=;�@;�C;bE;2�F;��G;ϸH;};I;�I;��I;3�I;P�I;�oI;�ZI;RHI;�8I;6+I;�I;5I;2I;iI;�I;Y�H;t�H;q�H;:�H;L�H;��H;��H;i�H;�H;i�H;��H;��H;L�H;:�H;q�H;t�H;Y�H;�I;iI;2I;5I;�I;6+I;�8I;RHI;�ZI;�oI;P�I;3�I;��I;�I;};I;ϸH;��G;2�F;bE;�C;�@;��=;.6;;��8;f06;�T4;V$3;      ��;�;N;�;Ϣ#;�);��.;�V4;C{9;\�=;N�A;��D;F;�H;��H;�^I;ߒI;l�I;g�I;�tI;�]I;�II;>9I;6+I;VI;�I;gI;�I;4I;��H;�H;F�H;�H;{�H;p�H;��H;b�H;��H;p�H;{�H;�H;F�H;�H;��H;4I;�I;gI;�I;VI;6+I;>9I;�II;�]I;�tI;g�I;l�I;ߒI;�^I;��H;�H;F;��D;N�A;\�=;C{9;�V4;��.;�);Ϣ#;�;N;�;      ���:}��:���:��:�)�:��;��;̧;Ͽ&;o�/;Z<7;oC=;��A;�E;^6G;w�H;�7I;
�I;#�I;��I;wI;�^I;�II;�8I;*I;I;LI;QI;�I;M I;�H;��H;*�H;M�H;��H;�H;��H;�H;��H;M�H;*�H;��H;�H;M I;�I;QI;LI;I;*I;�8I;�II;�^I;wI;��I;#�I;
�I;�7I;w�H;^6G;�E;��A;oC=;Z<7;o�/;Ͽ&;̧;��;��;�)�:��:���:}��:      �sx9���9��9�:J�^:���:ȼ:�N�:��;�g;�#;�;/;�:8;��>;�nC;�eF;W'H;eI;�~I;��I;ːI;wI;�]I;RHI;�6I;(I;#I;�I;�
I;\I;b�H;]�H;h�H;L�H;��H;��H;��H;��H;��H;L�H;h�H;]�H;b�H;\I;�
I;�I;#I;(I;�6I;RHI;�]I;wI;ːI;��I;�~I;eI;W'H;�eF;�nC;��>;�:8;�;/;�#;�g;��;�N�:ȼ:���:J�^:�:��9���9      ��d�����+�ht�#N�7��8*�&:L��:K��:�Y;\B;O�&;�&3;5<;��A; �E;��G;]I;w{I;��I;��I;�tI;�ZI;*EI;�3I;E%I;�I;bI;�I;I;O�H;��H;I�H;��H;��H;1�H;��H;��H;I�H;��H;O�H;I;�I;bI;�I;E%I;�3I;*EI;�ZI;�tI;��I;��I;w{I;]I;��G; �E;��A;5<;�&3;O�&;\B;�Y;K��:L��:*�&:7��8#N�ht�+���d���      �N����������g���8}�e�D����z�����Q��9�
�:���:&	;-�;�.;�9;�@;]E;��G;]I;�~I;#�I;g�I;�oI;�UI;�@I;�/I;�!I;�I;I;I;�I;��H;s�H;��H;r�H;��H;r�H;��H;s�H;��H;�I;I;I;�I;�!I;�/I;�@I;�UI;�oI;g�I;#�I;�~I;]I;��G;]E;�@;�9;�.;-�;&	;���:�
�:Q��9���z�����e�D��8}��g���������      *�?��<<�@�1�:i!��z�RC����ko��z�-�/򳺬���u�&:���:[��:¿;6�+;�8;W�@;]E;��G;eI;
�I;l�I;P�I;�hI;UOI;#;I;�*I;�I;�I;nI;EI;� I;��H;��H;d�H;��H;d�H;��H;��H;� I;EI;nI;�I;�I;�*I;#;I;UOI;�hI;P�I;l�I;
�I;eI;��G;]E;W�@;�8;6�+;¿;[��:���:u�&:����/�z�-�ko�����RC��z�:i!�@�1��<<�      ���p���I���������W�^�85��z��̻s숻�S��gt�U�x9d��:�k�:�g;z�*;�8;�@; �E;W'H;�7I;ߒI;3�I;o}I;�_I;�GI;�4I;y%I;�I;RI;	I;�I;��H;�H;i�H;��H;i�H;�H;��H;�I;	I;RI;�I;y%I;�4I;�GI;�_I;o}I;3�I;ߒI;�7I;W'H; �E;�@;�8;z�*;�g;�k�:d��:U�x9�gt��S�s숻�̻�z�85�W�^���������I��p��      6��p��
�*���z��fC���t�� �|��?�Ъ	������V�﮼�0U��߄:��:�g;6�+;�9;��A;�eF;w�H;�^I;��I;��I; rI;�UI;�?I;�-I; I;uI;(I;�I;�I;i�H;��H;�H;��H;i�H;�I;�I;(I;uI; I;�-I;�?I;�UI; rI;��I;��I;�^I;w�H;�eF;��A;�9;6�+;�g;��:�߄:0U�﮼���V����Ъ	��?� �|��t��fC��z��*����
�p�      ��t���p�9�d�-�Q���9�l*������Ҽ�I��N�o���'��ڻW7}���eH��߄:�k�:¿;�.;5<;�nC;^6G;��H;�I;��I;�I;<eI;^KI;7I;�&I;�I;�I;i
I;dI;�I;��H;l�H;��H;�I;dI;i
I;�I;�I;�&I;7I;^KI;<eI;�I;��I;�I;��H;^6G;�nC;5<;�.;¿;�k�:�߄:eH���W7}��ڻ��'�N�o��I����Ҽ���l*���9�-�Q�9�d���p�      ��Ž9���̷�V���z����}�$�Q�c�'����EC��I\��j<<�?��n����0U�d��:[��:-�;�&3;��>;�E;�H;};I;�I;ÔI;�uI;�WI;�@I;�.I;� I;�I;I;oI;�I;<I;�I;<I;�I;oI;I;�I;� I;�.I;�@I;�WI;�uI;ÔI;�I;};I;�H;�E;��>;�&3;-�;[��:d��:0U����n��?�j<<�I\��EC�����c�'�$�Q���}��z��V��̷�9���      c.��3�ɤ�W����҈Ž<5�����fG�@��kּe���9yC�?�W7}�﮼�U�x9���:&	;O�&;�:8;��A;F;ϸH;WxI;��I;�I;PeI;�JI;m6I;�&I;�I;�I;uI;/I;�I;�I;�I;/I;uI;�I;�I;�&I;m6I;�JI;PeI;�I;��I;WxI;ϸH;F;��A;�:8;O�&;&	;���:U�x9﮼�W7}�?�9yC�e���kּ@��fG����<5��҈Ž��W��ɤ��3�      Fx��s��d�M�N�`�3�}I����L����z����\�P*�'�ݼe���j<<��ڻ��V��gt�u�&:���:\B;�;/;oC=;��D;��G;8I;�I;ÓI;4sI;IUI;}>I;�,I;�I;�I;yI;�	I;I;.I;I;�	I;yI;�I;�I;�,I;}>I;IUI;4sI;ÓI;�I;8I;��G;��D;oC=;�;/;\B;���:u�&:�gt���V��ڻj<<�e���'�ݼP*���\��z��L������}I�`�3�M�N��d��s�      *l¾(��S������������d���7�y��<Sؽ[���d�P*�kּI\����'�����S������
�:�Y;�#;Z<7;N�A;2�F;|�H;��I;	�I;րI;	`I;�FI;3I;C$I;�I;�I;vI;i	I;iI;i	I;vI;�I;�I;C$I;3I;�FI;	`I;րI;	�I;��I;|�H;2�F;N�A;Z<7;�#;�Y;�
�:�����S������'�I\��kּP*��d�[��<Sؽy����7��d���������S���(��      �V������������Ͼ�d���ǆ�C�N��3��c�[����\�@��EC��N�o�Ъ	�s숻/�Q��9K��:�g;o�/;\�=;bE;2H;�VI;ٜI;�I;�jI;�NI;G9I;)I;=I;�I;I;�I;�
I;�I;I;�I;=I;)I;G9I;�NI;�jI;�I;ٜI;�VI;2H;bE;\�=;o�/;�g;K��:Q��9/�s숻Ъ	�N�o�EC��@����\�[���cཱ3�C�N��ǆ��d����Ͼ���������      ~,b���\��>M���5�9��-r��#l¾睒�"&W��3�<Sؽ�z��fG�����I���?��̻z�-����L��:��;Ͽ&;C{9;�C;�cG;tI;]�I;r�I;ruI;�VI;O?I;�-I;� I;�I;yI;�I;�I;�I;yI;�I;� I;�-I;O?I;�VI;ruI;r�I;]�I;tI;�cG;�C;C{9;Ͽ&;��;L��:���z�-��̻�?��I�����fG��z��<Sؽ�3�"&W�睒�#l¾-r��9����5��>M���\�      ���"��V���J䂿��\���1�����J˾睒�C�N�y��L������c�'���Ҽ �|��z�ko��z��*�&:�N�:̧;�V4;�@;HfF;��H;.�I;B�I;UI;=^I;�DI;&2I;<$I;cI;�I;I;�I;I;�I;cI;<$I;&2I;�DI;=^I;UI;B�I;.�I;��H;HfF;�@;�V4;̧;�N�:*�&:z��ko���z� �|���Ҽc�'����L���y��C�N�睒��J˾�����1���\�J䂿V���"��      }߿�$ڿ*�ʿ�������{Ps�MX:����#l¾�ǆ���7����<5��$�Q�����t��85�������7��8ȼ:��;��.;��=;�DE;�XH;�gI;G�I;ڇI;GeI;@JI;E6I;a'I;�I;I;�I;�I;�I;I;�I;a'I;E6I;@JI;GeI;ڇI;G�I;�gI;�XH;�DE;��=;��.;��;ȼ:7��8������85��t�����$�Q�<5�������7��ǆ�#l¾���MX:�{Ps��������*�ʿ�$ڿ      w�����p������ſ!��{Ps���1�-r���d���d�}I�҈Ž��}�l*�fC��W�^�RC�e�D�#N๫��:��;�);.6;;KD;e�G;kGI;ΜI;ȎI;�kI;OI;�9I;3*I;9I;�I;�I;KI;�I;�I;9I;3*I;�9I;OI;�kI;ȎI;ΜI;kGI;e�G;KD;.6;;�);��;���:#N�e�D�RC�W�^�fC��l*���}�҈Ž}I��d��d��-r����1�{Ps�!����ſ��꿀p����      ��7��3�Ң%�w��<����ſ�����\�9����Ͼ����`�3����z����9�z�ἷ���z��8}�ht�J�^:�)�:Ϣ#;��8;��B;ArG;�$I;јI;�I;$qI;7SI;=I;�,I;1!I;oI;I;�I;I;oI;1!I;�,I;=I;7SI;$qI;�I;јI;�$I;ArG;��B;��8;Ϣ#;�)�:J�^:ht��8}��z����z�Ἁ�9��z����`�3�������Ͼ9����\������ſ�<��w�Ң%��3�      (�_��+Y��lG�f.�w���꿭���J䂿��5���󾋰��M�N�W��V��-�Q�*�������:i!��g��+󳺑:��:�;f06;��A;uG;I;Z�I;��I;�uI;qVI;�?I;�.I;�"I;�I;'I;�I;'I;�I;�"I;�.I;�?I;qVI;�uI;��I;Z�I;I;uG;��A;f06;�;��:�:+��g��:i!�����*���-�Q�V��W��M�N���������5�J䂿�������w�f.��lG��+Y�      ά��}�8tf��lG�Ң%��p�*�ʿV����>M����S����d�ɤ�̷�9�d��
��I��@�1���������9���:N;�T4;��@;�F;A�H;�I;ܙI;�xI;�XI;bAI;�/I;�#I;�I;�I;�I;�I;�I;�#I;�/I;bAI;�XI;�xI;ܙI;�I;A�H;�F;��@;�T4;N;���:��9������@�1��I���
�9�d�̷�ɤ��d�S�������>M�V���*�ʿ�p�Ң%��lG�8tf�}�      O���A���}��+Y��3�����$ڿ"����\����(���s��3�9�����p�p�p���<<����d������9}��:�;V$3;io@;yF;��H;�I;�I;�zI;sZI;yBI;�0I;t$I;EI;uI; I;uI;EI;t$I;�0I;yBI;sZI;�zI;�I;�I;��H;yF;io@;V$3;�;}��:���9d�������<<�p��p���p�9����3��s�(�������\�"���$ڿ����3��+Y�}�A���      �Aq���i���U�A:�@�����6���q���uA�a5�� ��y^Z�����A���]�����d��|",�6��8�Ѻ���9)��:e�;eX4;p�@;�UF;��H;�FI;�aI;2NI;B9I;�(I;=I;�I;�I;�I;�
I;�I;�I;�I;=I;�(I;B9I;2NI;�aI;�FI;��H;�UF;p�@;eX4;e�;)��:���98�Ѻ6��|",��d������]��A�����y^Z�� ��a5�uA�q���6�������@�A:���U���i�      ��i���b�T�O�.5�-i������������q<�����e��[
V�FE	�!���IY�s9�Z����(� S����Ⱥ��:���:(�;L�4;h�@;kgF;��H;4HI;�aI;�MI;�8I;�(I;I;~I;�I;{I;x
I;{I;�I;~I;I;�(I;�8I;�MI;�aI;4HI;��H;kgF;h�@;L�4;(�;���:��:��Ⱥ S���(�Z���s9��IY�!��FE	�[
V��e������q<������������-i�.5�T�O���b�      ��U�T�O�B-?�(�'���F�`欿Y�{�aa/���뾙���I����e���ZN�o5��Ǩ��nH�� ��󊮺ߧ":��:��;��5;�_A;ښF;Z�H;<LI;aI;�LI;�7I;(I;aI;I;`I;&I;&
I;&I;`I;I;aI;(I;�7I;�LI;aI;<LI;Z�H;ښF;�_A;��5;��;��:ߧ":󊮺� ��nH�Ǩ��o5���ZN�e������I�������aa/�Y�{��欿F����(�'�B-?�T�O�      A:�.5�(�'��������dȿ���e$_���Q�Ҿؕ��
�6�����*���`=�P���)��zG��6��@����Q:�:/";�7;�%B;�F;��H;RI;�_I;�JI;D6I;�&I;ZI;7I;�I;�
I;�	I;�
I;�I;7I;ZI;�&I;D6I;�JI;�_I;RI;��H;�F;�%B;�7;/";�:��Q:@���6��zG��)��P���`=��*�����
�6�ؕ��Q�Ҿ��e$_����dȿ�������(�'�.5�      @�-i�������B�ѿf�������q<��:��a����q����Wн齅���'�ib̼�zl�/���X�w��!�:��;�&;ڪ9;LC;wLG;�H;^XI;�]I;�GI;4I;�$I;I;(I;�I;�	I;�I;�	I;�I;(I;I;�$I;4I;�GI;�]I;^XI;�H;wLG;LC;ڪ9;�&;��;!�:w���X�/���zl�ib̼��'�齅��Wн����q��a���:��q<����f���B�ѿ������-i�      �������F��dȿf���������O���u]׾w���	�I�����A��C�d�v��֮�<RH�Kkλ�$�h5����:nM;˅+;�<;"3D;�G;�I;�]I;�ZI;	DI;I1I;�"I;aI;�I;�I;�I;�I;�I;�I;�I;aI;�"I;I1I;	DI;�ZI;�]I;�I;�G;"3D;�<;˅+;nM;���:h5��$�Kkλ<RH��֮�v�C�d��A�����	�I�w���u]׾����O�����f���dȿF�ῢ��      6��������欿��������O�}x����� ���l���"��ܽ���`=�Ý��l"��R���ۺU��9�=�:�K;��0;͞>;�LE;}"H;�$I;�`I;(VI;�?I;.I;` I;\I;"I;0
I;mI;�I;mI;0
I;"I;\I;` I;.I;�?I;(VI;�`I;�$I;}"H;�LE;͞>;��0;�K;�=�:U��9�ۺ�R��l"����Ý��`=����ܽ��"��l�� �����}x���O��������欿����      q�������Y�{�e$_��q<�������}��w���6�����!��!�h��������� d��.��f_e�QL[���Z:���:�+ ;��5;�A;�UF;̃H;@I;�aI;�PI;;I;e*I;�I;+I;WI;�I;I;MI;I;�I;WI;+I;�I;e*I;;I;�PI;�aI;@I;̃H;�UF;�A;��5;�+ ;���:��Z:QL[�f_e��.��� d��������!�h�!�������6�w���}��������q<�e$_�Y�{�����      uA��q<�aa/����:�u]׾� ��w��>�BE	�����ܽ����3�r�꼰���=",�X��3��"AQ�ڮ�:�L
;�e);ބ:;D?C;?G;|�H;gSI;�^I;KJI;6I;t&I;�I;�I;ZI;�I;�I;�I;�I;�I;ZI;�I;�I;t&I;6I;KJI;�^I;gSI;|�H;?G;D?C;ބ:;�e);�L
;ڮ�:"AQ�3��X��=",�����r�꼠�3�ܽ������BE	�>�w��� ��u]׾�:���aa/��q<�      a5�������Q�Ҿ�a��w����l��6�BE	���Ƚk���aG����z֮�C�W����9�k����W`,:���:�;��1;n�>;^E;M�G;CI;H^I;hYI;ZCI;�0I;V"I;cI;I;#	I;-I;�I;=I;�I;-I;#	I;I;cI;V"I;�0I;ZCI;hYI;H^I;CI;M�G;^E;n�>;��1;�;���:W`,:���9�k����C�W�z֮�����aG�k����ȽBE	��6��l�w����a��Q�Ҿ������      � ���e�����ؕ����q�	�I���"���������k���ZN�c�6¼}�y��$�PR��\� ��[��:G/;K�&;w8;��A;��F;��H;?I;aI;�QI;;<I;7+I;�I;I;vI;�I;XI;9I;� I;9I;XI;�I;vI;I;�I;7+I;;<I;�QI;aI;?I;��H;��F;��A;w8;K�&;G/;�:�[�\� �PR���$�}�y�6¼c��ZN�k������������"�	�I���q�ؕ������e��      y^Z�[
V��I�
�6�������ܽ!��ܽ���aG�c��ȼ�)����(����H5����1�Z:l�:8R;/&1;��=;ПD;P�G;�H;�WI;:]I;�HI;5I;�%I;�I;�I;�	I;�I;mI;|�H;��H;|�H;mI;�I;�	I;�I;�I;�%I;5I;�HI;:]I;�WI;�H;P�G;ПD;��=;/&1;8R;l�:1�Z:���H5������(��)���ȼc��aG�ܽ��!���ܽ�����
�6��I�[
V�      ���FE	��������Wн�A����!�h���3����6¼�)��ax/�u�һC�X�%����9���:�=;\e);�_9;�%B;ډF;�|H;�5I;v`I;�TI;�?I;�-I; I;jI;DI;�I;jI;q�H;��H;�H;��H;q�H;jI;�I;DI;jI; I;�-I;�?I;�TI;v`I;�5I;�|H;ډF;�%B;�_9;\e);�=;���:��9%��C�X�u�һax/��)��6¼�����3�!�h��󑽢A���Wн��콹��FE	�      �A��!��e���*��齅�C�d��`=����r��z֮�}�y���(�u�һj^e������f9���:Y�;n0";B�4;�l?;E;��G;��H;�VI;�]I;(JI;�6I;'I;�I;FI;�	I;>I;7 I;��H;��H;W�H;��H;��H;7 I;>I;�	I;FI;�I;'I;�6I;(JI;�]I;�VI;��H;��G;E;�l?;B�4;n0";Y�;���:�f9����j^e�u�һ��(�}�y�z֮�r�꼠���`=�C�d�齅��*��e��!��      �]��IY��ZN��`=���'�v�Ý���������C�W��$����C�X������9�ޚ:���:��;˷0;�<;v�C;HG;�H;�>I;P`I;�SI;^?I;2.I;z I;�I;.I;�I;�I;��H;��H;&�H;��H;&�H;��H;��H;�I;�I;.I;�I;z I;2.I;^?I;�SI;P`I;�>I;�H;HG;v�C;�<;˷0;��;���:�ޚ:�9����C�X�����$�C�W���������Ý�v���'��`=��ZN��IY�      ���s9�o5��P��ib̼�֮����� d�=",����PR��H5�%���f9�ޚ:��:6�;��-;��:;KB;`UF;;JH; I;�[I;G[I;�GI;%5I;<&I;7I;�I;9	I;^I;�H;��H;��H;n�H;�H;n�H;��H;��H;�H;^I;9	I;�I;7I;<&I;%5I;�GI;G[I;�[I; I;;JH;`UF;KB;��:;��-;6�;��:�ޚ:�f9%��H5�PR�����=",�� d�����֮�ib̼P��o5��s9�      �d��Z���Ǩ���)���zl�<RH�l"��.��X��9�k�\� ������9���:���:6�;�-;�9;j`A;۹E;J�G;��H;#RI;4_I;OI;�;I;�+I;�I;MI;*I;�I;p I;��H;��H;��H;��H;|�H;��H;��H;��H;��H;p I;�I;*I;MI;�I;�+I;�;I;OI;4_I;#RI;��H;J�G;۹E;j`A;�9;�-;6�;���:���:��9���\� �9�k�X���.��l"�<RH��zl��)��Ǩ��Z���      |",��(�nH�zG�/��Kkλ�R��f_e�3������[�1�Z:���:Y�;��;��-;�9;�A;�bE;E�G;��H;tFI;`I;�TI;bAI;�0I;#I;�I;I;�I;I;��H;b�H;��H;!�H;,�H;��H;,�H;!�H;��H;b�H;��H;I;�I;I;�I;#I;�0I;bAI;�TI;`I;tFI;��H;E�G;�bE;�A;�9;��-;��;Y�;���:1�Z:�[����3��f_e��R��Kkλ/��zG�nH��(�      6�� S��� ���6���X��$��ۺQL[�"AQ�W`,:�:l�:�=;n0";˷0;��:;j`A;�bE;�G;��H;�<I;N_I;�XI;FI;5I;�&I;I;�I;
I;�I;��H;�H;6�H;�H;��H;��H;S�H;��H;��H;�H;6�H;�H;��H;�I;
I;�I;I;�&I;5I;FI;�XI;N_I;�<I;��H;�G;�bE;j`A;��:;˷0;n0";�=;l�:�:W`,:"AQ�QL[��ۺ�$��X��6��� �� S��      8�Ѻ��Ⱥ󊮺@��w��h5�U��9��Z:ڮ�:���:G/;8R;\e);B�4;�<;KB;۹E;E�G;��H;�9I;q^I;�ZI;?II;8I;�)I;�I;I;I;vI;$ I;��H;��H;&�H;C�H;�H;F�H;��H;F�H;�H;C�H;&�H;��H;��H;$ I;vI;I;I;�I;�)I;8I;?II;�ZI;q^I;�9I;��H;E�G;۹E;KB;�<;B�4;\e);8R;G/;���:ڮ�:��Z:U��9h5�w��@��󊮺��Ⱥ      ���9��:ߧ":��Q:!�:���:�=�:���:�L
;�;K�&;/&1;�_9;�l?;v�C;`UF;J�G;��H;�<I;q^I;1[I;�JI;2:I;�+I;�I;I;�I;�I;`I;��H;L�H;��H;K�H;��H;��H;��H;��H;��H;��H;��H;K�H;��H;L�H;��H;`I;�I;�I;I;�I;�+I;2:I;�JI;1[I;q^I;�<I;��H;J�G;`UF;v�C;�l?;�_9;/&1;K�&;�;�L
;���:�=�:���:!�:��Q:ߧ":��:      )��:���:��:�:��;nM;�K;�+ ;�e);��1;w8;��=;�%B;E;HG;;JH;��H;tFI;N_I;�ZI;�JI;�:I;-I;H!I;QI;+I;0I;xI;��H;��H;��H;}�H;��H;.�H;R�H;��H;y�H;��H;R�H;.�H;��H;}�H;��H;��H;��H;xI;0I;+I;QI;H!I;-I;�:I;�JI;�ZI;N_I;tFI;��H;;JH;HG;E;�%B;��=;w8;��1;�e);�+ ;�K;nM;��;�:��:���:      e�;(�;��;/";�&;˅+;��0;��5;ބ:;n�>;��A;ПD;ډF;��G;�H; I;#RI;`I;�XI;?II;2:I;-I;�!I;I;�I;	I;BI;^�H;��H;j�H;��H;��H;�H;��H; �H;��H;p�H;��H; �H;��H;�H;��H;��H;j�H;��H;^�H;BI;	I;�I;I;�!I;-I;2:I;?II;�XI;`I;#RI; I;�H;��G;ډF;ПD;��A;n�>;ބ:;��5;��0;˅+;�&;/";��;(�;      eX4;L�4;��5;�7;ڪ9;�<;͞>;�A;D?C;^E;��F;P�G;�|H;��H;�>I;�[I;4_I;�TI;FI;8I;�+I;H!I;I;9I;v	I;�I; �H;��H;��H;��H;��H;�H;��H;��H;��H;��H;u�H;��H;��H;��H;��H;�H;��H;��H;��H;��H; �H;�I;v	I;9I;I;H!I;�+I;8I;FI;�TI;4_I;�[I;�>I;��H;�|H;P�G;��F;^E;D?C;�A;͞>;�<;ڪ9;�7;��5;L�4;      p�@;h�@;�_A;�%B;LC;"3D;�LE;�UF;?G;M�G;��H;�H;�5I;�VI;P`I;G[I;OI;bAI;5I;�)I;�I;QI;�I;v	I;I;.�H;D�H;��H;0�H;��H;�H;��H;[�H;��H;��H;��H;r�H;��H;��H;��H;[�H;��H;�H;��H;0�H;��H;D�H;.�H;I;v	I;�I;QI;�I;�)I;5I;bAI;OI;G[I;P`I;�VI;�5I;�H;��H;M�G;?G;�UF;�LE;"3D;LC;�%B;�_A;h�@;      �UF;kgF;ښF;�F;wLG;�G;}"H;̃H;|�H;CI;?I;�WI;v`I;�]I;�SI;�GI;�;I;�0I;�&I;�I;I;+I;	I;�I;.�H;W�H;'�H;j�H;��H;�H;��H;V�H;L�H;��H;�H;��H;��H;��H;�H;��H;L�H;V�H;��H;�H;��H;j�H;'�H;W�H;.�H;�I;	I;+I;I;�I;�&I;�0I;�;I;�GI;�SI;�]I;v`I;�WI;?I;CI;|�H;̃H;}"H;�G;wLG;�F;ښF;kgF;      ��H;��H;Z�H;��H;�H;�I;�$I;@I;gSI;H^I;aI;:]I;�TI;(JI;^?I;%5I;�+I;#I;I;I;�I;0I;BI; �H;D�H;'�H;\�H;�H;7�H;|�H;7�H;�H;F�H;��H;@�H;��H;��H;��H;@�H;��H;F�H;�H;7�H;|�H;7�H;�H;\�H;'�H;D�H; �H;BI;0I;�I;I;I;#I;�+I;%5I;^?I;(JI;�TI;:]I;aI;H^I;gSI;@I;�$I;�I;�H;��H;Z�H;��H;      �FI;4HI;<LI;RI;^XI;�]I;�`I;�aI;�^I;hYI;�QI;�HI;�?I;�6I;2.I;<&I;�I;�I;�I;I;�I;xI;^�H;��H;��H;j�H;�H;�H;��H;3�H;�H;�H;p�H;��H;|�H;F�H;@�H;F�H;|�H;��H;p�H;�H;�H;3�H;��H;�H;�H;j�H;��H;��H;^�H;xI;�I;I;�I;�I;�I;<&I;2.I;�6I;�?I;�HI;�QI;hYI;�^I;�aI;�`I;�]I;^XI;RI;<LI;4HI;      �aI;�aI;aI;�_I;�]I;�ZI;(VI;�PI;KJI;ZCI;;<I;5I;�-I;'I;z I;7I;MI;I;
I;vI;`I;��H;��H;��H;0�H;��H;7�H;��H;*�H;�H;�H;B�H;��H;2�H;��H;��H;��H;��H;��H;2�H;��H;B�H;�H;�H;*�H;��H;7�H;��H;0�H;��H;��H;��H;`I;vI;
I;I;MI;7I;z I;'I;�-I;5I;;<I;ZCI;KJI;�PI;(VI;�ZI;�]I;�_I;aI;�aI;      2NI;�MI;�LI;�JI;�GI;	DI;�?I;;I;6I;�0I;7+I;�%I; I;�I;�I;�I;*I;�I;�I;$ I;��H;��H;j�H;��H;��H;�H;|�H;3�H;�H;�H;1�H;��H;��H;��H;H�H;(�H;%�H;(�H;H�H;��H;��H;��H;1�H;�H;�H;3�H;|�H;�H;��H;��H;j�H;��H;��H;$ I;�I;�I;*I;�I;�I;�I; I;�%I;7+I;�0I;6I;;I;�?I;	DI;�GI;�JI;�LI;�MI;      B9I;�8I;�7I;D6I;4I;I1I;.I;e*I;t&I;V"I;�I;�I;jI;FI;.I;9	I;�I;I;��H;��H;L�H;��H;��H;��H;�H;��H;7�H;�H;�H;1�H;��H;��H;d�H;�H;��H;��H;��H;��H;��H;�H;d�H;��H;��H;1�H;�H;�H;7�H;��H;�H;��H;��H;��H;L�H;��H;��H;I;�I;9	I;.I;FI;jI;�I;�I;V"I;t&I;e*I;.I;I1I;4I;D6I;�7I;�8I;      �(I;�(I;(I;�&I;�$I;�"I;` I;�I;�I;cI;I;�I;DI;�	I;�I;^I;p I;��H;�H;��H;��H;}�H;��H;�H;��H;V�H;�H;�H;B�H;��H;��H;{�H;��H;��H;z�H;T�H;>�H;T�H;z�H;��H;��H;{�H;��H;��H;B�H;�H;�H;V�H;��H;�H;��H;}�H;��H;��H;�H;��H;p I;^I;�I;�	I;DI;�I;I;cI;�I;�I;` I;�"I;�$I;�&I;(I;�(I;      =I;I;aI;ZI;I;aI;\I;+I;�I;I;vI;�	I;�I;>I;�I;�H;��H;b�H;6�H;&�H;K�H;��H;�H;��H;[�H;L�H;F�H;p�H;��H;��H;d�H;��H;��H;\�H;�H;	�H;�H;	�H;�H;\�H;��H;��H;d�H;��H;��H;p�H;F�H;L�H;[�H;��H;�H;��H;K�H;&�H;6�H;b�H;��H;�H;�I;>I;�I;�	I;vI;I;�I;+I;\I;aI;I;ZI;aI;I;      �I;~I;I;7I;(I;�I;"I;WI;ZI;#	I;�I;�I;jI;7 I;��H;��H;��H;��H;�H;C�H;��H;.�H;��H;��H;��H;��H;��H;��H;2�H;��H;�H;��H;\�H; �H;��H;��H;��H;��H;��H; �H;\�H;��H;�H;��H;2�H;��H;��H;��H;��H;��H;��H;.�H;��H;C�H;�H;��H;��H;��H;��H;7 I;jI;�I;�I;#	I;ZI;WI;"I;�I;(I;7I;I;~I;      �I;�I;`I;�I;�I;�I;0
I;�I;�I;-I;XI;mI;q�H;��H;��H;��H;��H;!�H;��H;�H;��H;R�H; �H;��H;��H;�H;@�H;|�H;��H;H�H;��H;z�H;�H;��H;��H;��H;��H;��H;��H;��H;�H;z�H;��H;H�H;��H;|�H;@�H;�H;��H;��H; �H;R�H;��H;�H;��H;!�H;��H;��H;��H;��H;q�H;mI;XI;-I;�I;�I;0
I;�I;�I;�I;`I;�I;      �I;{I;&I;�
I;�	I;�I;mI;I;�I;�I;9I;|�H;��H;��H;&�H;n�H;��H;,�H;��H;F�H;��H;��H;��H;��H;��H;��H;��H;F�H;��H;(�H;��H;T�H;	�H;��H;��H;��H;}�H;��H;��H;��H;	�H;T�H;��H;(�H;��H;F�H;��H;��H;��H;��H;��H;��H;��H;F�H;��H;,�H;��H;n�H;&�H;��H;��H;|�H;9I;�I;�I;I;mI;�I;�	I;�
I;&I;{I;      �
I;x
I;&
I;�	I;�I;�I;�I;MI;�I;=I;� I;��H;�H;W�H;��H;�H;|�H;��H;S�H;��H;��H;y�H;p�H;u�H;r�H;��H;��H;@�H;��H;%�H;��H;>�H;�H;��H;��H;}�H;��H;}�H;��H;��H;�H;>�H;��H;%�H;��H;@�H;��H;��H;r�H;u�H;p�H;y�H;��H;��H;S�H;��H;|�H;�H;��H;W�H;�H;��H;� I;=I;�I;MI;�I;�I;�I;�	I;&
I;x
I;      �I;{I;&I;�
I;�	I;�I;mI;I;�I;�I;9I;|�H;��H;��H;&�H;n�H;��H;,�H;��H;F�H;��H;��H;��H;��H;��H;��H;��H;F�H;��H;(�H;��H;T�H;	�H;��H;��H;��H;}�H;��H;��H;��H;	�H;T�H;��H;(�H;��H;F�H;��H;��H;��H;��H;��H;��H;��H;F�H;��H;,�H;��H;n�H;&�H;��H;��H;|�H;9I;�I;�I;I;mI;�I;�	I;�
I;&I;{I;      �I;�I;`I;�I;�I;�I;0
I;�I;�I;-I;XI;mI;q�H;��H;��H;��H;��H;!�H;��H;�H;��H;R�H; �H;��H;��H;�H;@�H;|�H;��H;H�H;��H;z�H;�H;��H;��H;��H;��H;��H;��H;��H;�H;z�H;��H;H�H;��H;|�H;@�H;�H;��H;��H; �H;R�H;��H;�H;��H;!�H;��H;��H;��H;��H;q�H;mI;XI;-I;�I;�I;0
I;�I;�I;�I;`I;�I;      �I;~I;I;7I;(I;�I;"I;WI;ZI;#	I;�I;�I;jI;7 I;��H;��H;��H;��H;�H;C�H;��H;.�H;��H;��H;��H;��H;��H;��H;2�H;��H;�H;��H;\�H; �H;��H;��H;��H;��H;��H; �H;\�H;��H;�H;��H;2�H;��H;��H;��H;��H;��H;��H;.�H;��H;C�H;�H;��H;��H;��H;��H;7 I;jI;�I;�I;#	I;ZI;WI;"I;�I;(I;7I;I;~I;      =I;I;aI;ZI;I;aI;\I;+I;�I;I;vI;�	I;�I;>I;�I;�H;��H;b�H;6�H;&�H;K�H;��H;�H;��H;[�H;L�H;F�H;p�H;��H;��H;d�H;��H;��H;\�H;�H;	�H;�H;	�H;�H;\�H;��H;��H;d�H;��H;��H;p�H;F�H;L�H;[�H;��H;�H;��H;K�H;&�H;6�H;b�H;��H;�H;�I;>I;�I;�	I;vI;I;�I;+I;\I;aI;I;ZI;aI;I;      �(I;�(I;(I;�&I;�$I;�"I;` I;�I;�I;cI;I;�I;DI;�	I;�I;^I;p I;��H;�H;��H;��H;}�H;��H;�H;��H;V�H;�H;�H;B�H;��H;��H;{�H;��H;��H;z�H;T�H;>�H;T�H;z�H;��H;��H;{�H;��H;��H;B�H;�H;�H;V�H;��H;�H;��H;}�H;��H;��H;�H;��H;p I;^I;�I;�	I;DI;�I;I;cI;�I;�I;` I;�"I;�$I;�&I;(I;�(I;      B9I;�8I;�7I;D6I;4I;I1I;.I;e*I;t&I;V"I;�I;�I;jI;FI;.I;9	I;�I;I;��H;��H;L�H;��H;��H;��H;�H;��H;7�H;�H;�H;1�H;��H;��H;d�H;�H;��H;��H;��H;��H;��H;�H;d�H;��H;��H;1�H;�H;�H;7�H;��H;�H;��H;��H;��H;L�H;��H;��H;I;�I;9	I;.I;FI;jI;�I;�I;V"I;t&I;e*I;.I;I1I;4I;D6I;�7I;�8I;      2NI;�MI;�LI;�JI;�GI;	DI;�?I;;I;6I;�0I;7+I;�%I; I;�I;�I;�I;*I;�I;�I;$ I;��H;��H;j�H;��H;��H;�H;|�H;3�H;�H;�H;1�H;��H;��H;��H;H�H;(�H;%�H;(�H;H�H;��H;��H;��H;1�H;�H;�H;3�H;|�H;�H;��H;��H;j�H;��H;��H;$ I;�I;�I;*I;�I;�I;�I; I;�%I;7+I;�0I;6I;;I;�?I;	DI;�GI;�JI;�LI;�MI;      �aI;�aI;aI;�_I;�]I;�ZI;(VI;�PI;KJI;ZCI;;<I;5I;�-I;'I;z I;7I;MI;I;
I;vI;`I;��H;��H;��H;0�H;��H;7�H;��H;*�H;�H;�H;B�H;��H;2�H;��H;��H;��H;��H;��H;2�H;��H;B�H;�H;�H;*�H;��H;7�H;��H;0�H;��H;��H;��H;`I;vI;
I;I;MI;7I;z I;'I;�-I;5I;;<I;ZCI;KJI;�PI;(VI;�ZI;�]I;�_I;aI;�aI;      �FI;4HI;<LI;RI;^XI;�]I;�`I;�aI;�^I;hYI;�QI;�HI;�?I;�6I;2.I;<&I;�I;�I;�I;I;�I;xI;^�H;��H;��H;j�H;�H;�H;��H;3�H;�H;�H;p�H;��H;|�H;F�H;@�H;F�H;|�H;��H;p�H;�H;�H;3�H;��H;�H;�H;j�H;��H;��H;^�H;xI;�I;I;�I;�I;�I;<&I;2.I;�6I;�?I;�HI;�QI;hYI;�^I;�aI;�`I;�]I;^XI;RI;<LI;4HI;      ��H;��H;Z�H;��H;�H;�I;�$I;@I;gSI;H^I;aI;:]I;�TI;(JI;^?I;%5I;�+I;#I;I;I;�I;0I;BI; �H;D�H;'�H;\�H;�H;7�H;|�H;7�H;�H;F�H;��H;@�H;��H;��H;��H;@�H;��H;F�H;�H;7�H;|�H;7�H;�H;\�H;'�H;D�H; �H;BI;0I;�I;I;I;#I;�+I;%5I;^?I;(JI;�TI;:]I;aI;H^I;gSI;@I;�$I;�I;�H;��H;Z�H;��H;      �UF;kgF;ښF;�F;wLG;�G;}"H;̃H;|�H;CI;?I;�WI;v`I;�]I;�SI;�GI;�;I;�0I;�&I;�I;I;+I;	I;�I;.�H;W�H;'�H;j�H;��H;�H;��H;V�H;L�H;��H;�H;��H;��H;��H;�H;��H;L�H;V�H;��H;�H;��H;j�H;'�H;W�H;.�H;�I;	I;+I;I;�I;�&I;�0I;�;I;�GI;�SI;�]I;v`I;�WI;?I;CI;|�H;̃H;}"H;�G;wLG;�F;ښF;kgF;      p�@;h�@;�_A;�%B;LC;"3D;�LE;�UF;?G;M�G;��H;�H;�5I;�VI;P`I;G[I;OI;bAI;5I;�)I;�I;QI;�I;v	I;I;.�H;D�H;��H;0�H;��H;�H;��H;[�H;��H;��H;��H;r�H;��H;��H;��H;[�H;��H;�H;��H;0�H;��H;D�H;.�H;I;v	I;�I;QI;�I;�)I;5I;bAI;OI;G[I;P`I;�VI;�5I;�H;��H;M�G;?G;�UF;�LE;"3D;LC;�%B;�_A;h�@;      eX4;L�4;��5;�7;ڪ9;�<;͞>;�A;D?C;^E;��F;P�G;�|H;��H;�>I;�[I;4_I;�TI;FI;8I;�+I;H!I;I;9I;v	I;�I; �H;��H;��H;��H;��H;�H;��H;��H;��H;��H;u�H;��H;��H;��H;��H;�H;��H;��H;��H;��H; �H;�I;v	I;9I;I;H!I;�+I;8I;FI;�TI;4_I;�[I;�>I;��H;�|H;P�G;��F;^E;D?C;�A;͞>;�<;ڪ9;�7;��5;L�4;      e�;(�;��;/";�&;˅+;��0;��5;ބ:;n�>;��A;ПD;ډF;��G;�H; I;#RI;`I;�XI;?II;2:I;-I;�!I;I;�I;	I;BI;^�H;��H;j�H;��H;��H;�H;��H; �H;��H;p�H;��H; �H;��H;�H;��H;��H;j�H;��H;^�H;BI;	I;�I;I;�!I;-I;2:I;?II;�XI;`I;#RI; I;�H;��G;ډF;ПD;��A;n�>;ބ:;��5;��0;˅+;�&;/";��;(�;      )��:���:��:�:��;nM;�K;�+ ;�e);��1;w8;��=;�%B;E;HG;;JH;��H;tFI;N_I;�ZI;�JI;�:I;-I;H!I;QI;+I;0I;xI;��H;��H;��H;}�H;��H;.�H;R�H;��H;y�H;��H;R�H;.�H;��H;}�H;��H;��H;��H;xI;0I;+I;QI;H!I;-I;�:I;�JI;�ZI;N_I;tFI;��H;;JH;HG;E;�%B;��=;w8;��1;�e);�+ ;�K;nM;��;�:��:���:      ���9��:ߧ":��Q:!�:���:�=�:���:�L
;�;K�&;/&1;�_9;�l?;v�C;`UF;J�G;��H;�<I;q^I;1[I;�JI;2:I;�+I;�I;I;�I;�I;`I;��H;L�H;��H;K�H;��H;��H;��H;��H;��H;��H;��H;K�H;��H;L�H;��H;`I;�I;�I;I;�I;�+I;2:I;�JI;1[I;q^I;�<I;��H;J�G;`UF;v�C;�l?;�_9;/&1;K�&;�;�L
;���:�=�:���:!�:��Q:ߧ":��:      8�Ѻ��Ⱥ󊮺@��w��h5�U��9��Z:ڮ�:���:G/;8R;\e);B�4;�<;KB;۹E;E�G;��H;�9I;q^I;�ZI;?II;8I;�)I;�I;I;I;vI;$ I;��H;��H;&�H;C�H;�H;F�H;��H;F�H;�H;C�H;&�H;��H;��H;$ I;vI;I;I;�I;�)I;8I;?II;�ZI;q^I;�9I;��H;E�G;۹E;KB;�<;B�4;\e);8R;G/;���:ڮ�:��Z:U��9h5�w��@��󊮺��Ⱥ      6�� S��� ���6���X��$��ۺQL[�"AQ�W`,:�:l�:�=;n0";˷0;��:;j`A;�bE;�G;��H;�<I;N_I;�XI;FI;5I;�&I;I;�I;
I;�I;��H;�H;6�H;�H;��H;��H;S�H;��H;��H;�H;6�H;�H;��H;�I;
I;�I;I;�&I;5I;FI;�XI;N_I;�<I;��H;�G;�bE;j`A;��:;˷0;n0";�=;l�:�:W`,:"AQ�QL[��ۺ�$��X��6��� �� S��      |",��(�nH�zG�/��Kkλ�R��f_e�3������[�1�Z:���:Y�;��;��-;�9;�A;�bE;E�G;��H;tFI;`I;�TI;bAI;�0I;#I;�I;I;�I;I;��H;b�H;��H;!�H;,�H;��H;,�H;!�H;��H;b�H;��H;I;�I;I;�I;#I;�0I;bAI;�TI;`I;tFI;��H;E�G;�bE;�A;�9;��-;��;Y�;���:1�Z:�[����3��f_e��R��Kkλ/��zG�nH��(�      �d��Z���Ǩ���)���zl�<RH�l"��.��X��9�k�\� ������9���:���:6�;�-;�9;j`A;۹E;J�G;��H;#RI;4_I;OI;�;I;�+I;�I;MI;*I;�I;p I;��H;��H;��H;��H;|�H;��H;��H;��H;��H;p I;�I;*I;MI;�I;�+I;�;I;OI;4_I;#RI;��H;J�G;۹E;j`A;�9;�-;6�;���:���:��9���\� �9�k�X���.��l"�<RH��zl��)��Ǩ��Z���      ���s9�o5��P��ib̼�֮����� d�=",����PR��H5�%���f9�ޚ:��:6�;��-;��:;KB;`UF;;JH; I;�[I;G[I;�GI;%5I;<&I;7I;�I;9	I;^I;�H;��H;��H;n�H;�H;n�H;��H;��H;�H;^I;9	I;�I;7I;<&I;%5I;�GI;G[I;�[I; I;;JH;`UF;KB;��:;��-;6�;��:�ޚ:�f9%��H5�PR�����=",�� d�����֮�ib̼P��o5��s9�      �]��IY��ZN��`=���'�v�Ý���������C�W��$����C�X������9�ޚ:���:��;˷0;�<;v�C;HG;�H;�>I;P`I;�SI;^?I;2.I;z I;�I;.I;�I;�I;��H;��H;&�H;��H;&�H;��H;��H;�I;�I;.I;�I;z I;2.I;^?I;�SI;P`I;�>I;�H;HG;v�C;�<;˷0;��;���:�ޚ:�9����C�X�����$�C�W���������Ý�v���'��`=��ZN��IY�      �A��!��e���*��齅�C�d��`=����r��z֮�}�y���(�u�һj^e������f9���:Y�;n0";B�4;�l?;E;��G;��H;�VI;�]I;(JI;�6I;'I;�I;FI;�	I;>I;7 I;��H;��H;W�H;��H;��H;7 I;>I;�	I;FI;�I;'I;�6I;(JI;�]I;�VI;��H;��G;E;�l?;B�4;n0";Y�;���:�f9����j^e�u�һ��(�}�y�z֮�r�꼠���`=�C�d�齅��*��e��!��      ���FE	��������Wн�A����!�h���3����6¼�)��ax/�u�һC�X�%����9���:�=;\e);�_9;�%B;ډF;�|H;�5I;v`I;�TI;�?I;�-I; I;jI;DI;�I;jI;q�H;��H;�H;��H;q�H;jI;�I;DI;jI; I;�-I;�?I;�TI;v`I;�5I;�|H;ډF;�%B;�_9;\e);�=;���:��9%��C�X�u�һax/��)��6¼�����3�!�h��󑽢A���Wн��콹��FE	�      y^Z�[
V��I�
�6�������ܽ!��ܽ���aG�c��ȼ�)����(����H5����1�Z:l�:8R;/&1;��=;ПD;P�G;�H;�WI;:]I;�HI;5I;�%I;�I;�I;�	I;�I;mI;|�H;��H;|�H;mI;�I;�	I;�I;�I;�%I;5I;�HI;:]I;�WI;�H;P�G;ПD;��=;/&1;8R;l�:1�Z:���H5������(��)���ȼc��aG�ܽ��!���ܽ�����
�6��I�[
V�      � ���e�����ؕ����q�	�I���"���������k���ZN�c�6¼}�y��$�PR��\� ��[��:G/;K�&;w8;��A;��F;��H;?I;aI;�QI;;<I;7+I;�I;I;vI;�I;XI;9I;� I;9I;XI;�I;vI;I;�I;7+I;;<I;�QI;aI;?I;��H;��F;��A;w8;K�&;G/;�:�[�\� �PR���$�}�y�6¼c��ZN�k������������"�	�I���q�ؕ������e��      a5�������Q�Ҿ�a��w����l��6�BE	���Ƚk���aG����z֮�C�W����9�k����W`,:���:�;��1;n�>;^E;M�G;CI;H^I;hYI;ZCI;�0I;V"I;cI;I;#	I;-I;�I;=I;�I;-I;#	I;I;cI;V"I;�0I;ZCI;hYI;H^I;CI;M�G;^E;n�>;��1;�;���:W`,:���9�k����C�W�z֮�����aG�k����ȽBE	��6��l�w����a��Q�Ҿ������      uA��q<�aa/����:�u]׾� ��w��>�BE	�����ܽ����3�r�꼰���=",�X��3��"AQ�ڮ�:�L
;�e);ބ:;D?C;?G;|�H;gSI;�^I;KJI;6I;t&I;�I;�I;ZI;�I;�I;�I;�I;�I;ZI;�I;�I;t&I;6I;KJI;�^I;gSI;|�H;?G;D?C;ބ:;�e);�L
;ڮ�:"AQ�3��X��=",�����r�꼠�3�ܽ������BE	�>�w��� ��u]׾�:���aa/��q<�      q�������Y�{�e$_��q<�������}��w���6�����!��!�h��������� d��.��f_e�QL[���Z:���:�+ ;��5;�A;�UF;̃H;@I;�aI;�PI;;I;e*I;�I;+I;WI;�I;I;MI;I;�I;WI;+I;�I;e*I;;I;�PI;�aI;@I;̃H;�UF;�A;��5;�+ ;���:��Z:QL[�f_e��.��� d��������!�h�!�������6�w���}��������q<�e$_�Y�{�����      6��������欿��������O�}x����� ���l���"��ܽ���`=�Ý��l"��R���ۺU��9�=�:�K;��0;͞>;�LE;}"H;�$I;�`I;(VI;�?I;.I;` I;\I;"I;0
I;mI;�I;mI;0
I;"I;\I;` I;.I;�?I;(VI;�`I;�$I;}"H;�LE;͞>;��0;�K;�=�:U��9�ۺ�R��l"����Ý��`=����ܽ��"��l�� �����}x���O��������欿����      �������F��dȿf���������O���u]׾w���	�I�����A��C�d�v��֮�<RH�Kkλ�$�h5����:nM;˅+;�<;"3D;�G;�I;�]I;�ZI;	DI;I1I;�"I;aI;�I;�I;�I;�I;�I;�I;�I;aI;�"I;I1I;	DI;�ZI;�]I;�I;�G;"3D;�<;˅+;nM;���:h5��$�Kkλ<RH��֮�v�C�d��A�����	�I�w���u]׾����O�����f���dȿF�ῢ��      @�-i�������B�ѿf�������q<��:��a����q����Wн齅���'�ib̼�zl�/���X�w��!�:��;�&;ڪ9;LC;wLG;�H;^XI;�]I;�GI;4I;�$I;I;(I;�I;�	I;�I;�	I;�I;(I;I;�$I;4I;�GI;�]I;^XI;�H;wLG;LC;ڪ9;�&;��;!�:w���X�/���zl�ib̼��'�齅��Wн����q��a���:��q<����f���B�ѿ������-i�      A:�.5�(�'��������dȿ���e$_���Q�Ҿؕ��
�6�����*���`=�P���)��zG��6��@����Q:�:/";�7;�%B;�F;��H;RI;�_I;�JI;D6I;�&I;ZI;7I;�I;�
I;�	I;�
I;�I;7I;ZI;�&I;D6I;�JI;�_I;RI;��H;�F;�%B;�7;/";�:��Q:@���6��zG��)��P���`=��*�����
�6�ؕ��Q�Ҿ��e$_����dȿ�������(�'�.5�      ��U�T�O�B-?�(�'���F�`欿Y�{�aa/���뾙���I����e���ZN�o5��Ǩ��nH�� ��󊮺ߧ":��:��;��5;�_A;ښF;Z�H;<LI;aI;�LI;�7I;(I;aI;I;`I;&I;&
I;&I;`I;I;aI;(I;�7I;�LI;aI;<LI;Z�H;ښF;�_A;��5;��;��:ߧ":󊮺� ��nH�Ǩ��o5���ZN�e������I�������aa/�Y�{��欿F����(�'�B-?�T�O�      ��i���b�T�O�.5�-i������������q<�����e��[
V�FE	�!���IY�s9�Z����(� S����Ⱥ��:���:(�;L�4;h�@;kgF;��H;4HI;�aI;�MI;�8I;�(I;I;~I;�I;{I;x
I;{I;�I;~I;I;�(I;�8I;�MI;�aI;4HI;��H;kgF;h�@;L�4;(�;���:��:��Ⱥ S���(�Z���s9��IY�!��FE	�[
V��e������q<������������-i�.5�T�O���b�      �>���8���*�O������˿�o��<�b�=\�+m־^��K�:��J�&��F�B�F���������/��������>:�r�:eo ;�I6;DA;�HF;�MH;�H;!I;�I;I;�I;mI;I;q�H;��H;+�H;��H;q�H;I;mI;�I;I;�I;!I;�H;�MH;�HF;DA;�I6;eo ;�r�:��>:�����/���������F��F�B�&���J�K�:�^��+m־=\�<�b��o���˿����O���*���8�      ��8��4��g&�0��2����<ƿ벗��>]����G�Ѿ�p���*7����"W��MR?�	}�8����s������:�G:���:!;'�6;(kA;�XF;�SH;s�H;!I;�I;�I;�I;FI;�I;e�H;��H;�H;��H;e�H;�I;FI;�I;�I;�I;!I;s�H;�SH;�XF;(kA;'�6;!;���::�G:���s�����8��	}�MR?�"W�����*7��p��G�Ѿ����>]�벗��<ƿ2���0���g&��4�      ��*��g&��#�o�K[�jL�������M�l5��>ľ
����,��D�撐��5�;�ݼ���q
���x��wk���b:�j�:#;ۖ7;��A;�F;�cH;�I;\!I;I;pI;BI;�I;�I;!�H;x�H;��H;x�H;!�H;�I;�I;BI;pI;I;\!I;�I;�cH;�F;��A;ۖ7;#;�j�:��b:�wk���x��q
���;�ݼ�5�撐��Dὤ�,�
���>ľl5���M����jL��K[�o��#��g&�      O�0��o����˿:1��-�y���6��z �����)�l�+��ͽ!�����&���˼_�k�q���k�X��� �ѳ�:p�;)&;�9;��B;�F;�|H;�I;f!I;5I;�I;�
I;qI;FI;��H;"�H;��H;"�H;��H;FI;qI;�
I;�I;5I;f!I;�I;�|H;�F;��B;�9;)&;p�;ѳ�:�� �k�X�q���_�k���˼��&�!����ͽ+�)�l������z ���6�-�y�:1���˿���o�0��      ����2���K[忭˿�T��蟉�s�R�����E۾̗����M�~�	������j��3�"d��ɆO���׻b�/��
�����:��	;%*;l;;�iC;�&G;�H;�I;
!I;�I;�I;�	I;�I;� I;I�H;��H; �H;��H;I�H;� I;�I;�	I;�I;�I;
!I;�I;�H;�&G;�iC;l;;%*;��	;���:�
��b�/���׻ɆO�"d���3���j����~�	���M�̗���E۾���s�R�蟉��T���˿K[�2���      �˿�<ƿjL��:1��蟉��>]���)��$���ճ���{���,�j��$��Q`I��J��-��4/�S,��ʻ ��!69
3�:�;o.;0-=;o`D;�G;o�H;�I;@ I;aI;TI;�I;�I;��H;��H;�H;d�H;�H;��H;��H;�I;�I;TI;aI;@ I;�I;o�H;�G;o`D;0-=;o.;�;
3�:�!69ʻ �S,��4/�-���J��Q`I�$��j�齞�,���{��ճ��$����)��>]�蟉�:1��jL���<ƿ      �o��벗����-�y�s�R���)�iv��>ľ�]����I�Tl�~��������&�߮Ҽ	�}�VB�!���������!:?)�:Vy;�3;li?;�[E;��G;��H;tI;�I;�I;�I;|I;�I;�H;��H;c�H;��H;c�H;��H;�H;�I;|I;�I;�I;�I;tI;��H;��G;�[E;li?;�3;Vy;?)�:��!:����!���VB�	�}�߮Ҽ��&����~���Tl���I��]���>ľiv���)�s�R�-�y����벗�      <�b��>]���M���6�����$���>ľq��q�Z�+�K9ݽW����L����/F��&�G�\�׻�;�u�Ǌ:�h;6O$;�7;y�A;IF;:BH;��H;�I;nI;xI;I;-I;�I;�H;��H;��H;�H;��H;��H;�H;�I;-I;I;xI;nI;�I;��H;:BH;IF;y�A;�7;6O$;�h;Ǌ:u칸;�\�׻&�G�/F�������L�W��K9ݽ+�q�Z�q���>ľ�$�������6���M��>]�      =\����l5��z ��E۾�ճ��]��q�Z�F?#����A����j�(��Oϼ��������Rnۺq3�9�2�:p�;y�,;��;;C�C;�G;R�H;�
I;� I;�I;GI;.
I;�I;? I;�H;�H;��H;"�H;��H;�H;�H;? I;�I;.
I;GI;�I;� I;�
I;R�H;�G;C�C;��;;y�,;p�;�2�:q3�9Rnۺ��������Oϼ(����j��A�����F?#�q�Z��]���ճ��E۾�z �l5����      +m־G�Ѿ�>ľ����̗����{���I�+����V���{�?�/�.���,��b=���һ�@�9� ���k:C�:$a;��3;Ai?;w1E;��G;p�H;7I;wI;�I;�I;&I;�I;��H;��H;��H;��H;V�H;��H;��H;��H;��H;�I;&I;�I;�I;wI;7I;p�H;��G;w1E;Ai?;��3;$a;C�:��k:9� ��@���һb=��,��.��?�/��{��V�����+���I���{�̗�������>ľG�Ѿ      ^���p��
��)�l���M���,�Tl�K9ݽ�A���{���5��J��;���T[�I?������Q��J�9�:��;:*;5�9;jjB;ۆF;�MH;��H; I;�I;�I;"I;I;@I;_�H;��H;��H;��H;j�H;��H;��H;��H;_�H;@I;I;"I;�I;�I; I;��H;�MH;ۆF;jjB;5�9;:*;��;�:J�9�Q������I?��T[�;���J����5��{��A��K9ݽTl���,���M�)�l�
���p��      K�:��*7���,�+�~�	�j��~���W����j�?�/��J���I��%�k���b.�������<Ǌ:�m�:(;nq3;2�>;8�D;t�G;S�H;I;/ I;�I;�I;�	I;�I;`�H;��H;��H;��H;��H;_�H;��H;��H;��H;��H;`�H;�I;�	I;�I;�I;/ I;I;S�H;t�G;8�D;2�>;nq3;(;�m�:<Ǌ:�����b.����%�k��I���J��?�/���j�W��~���j��~�	�+���,��*7�      �J���D��ͽ���$�������L�(��.��;��%�k����I����/��"/�+�>:���:�A;w�,;��:;>�B;�wF;�;H;��H;
I;�I;�I;AI;�I;�I;��H;s�H;5�H;o�H;��H;l�H;��H;o�H;5�H;s�H;��H;�I;�I;AI;�I;�I;
I;��H;�;H;�wF;>�B;��:;w�,;�A;���:+�>:�"/���/��I����%�k�;��.��(����L����$������ͽ�Dὼ��      &��"W��撐�!�����j�Q`I���&����Oϼ�,���T[����I��;��qk�n:i3�:� ;!&;�6;� @;D1E;�G;��H;�I;�I;OI;I;�	I;;I;u�H;��H;�H;��H;^�H;��H;D�H;��H;^�H;��H;�H;��H;u�H;;I;�	I;I;OI;�I;�I;��H;�G;D1E;� @;�6;!&;� ;i3�:n:�qk�;��I�����T[��,��Oϼ�����&�Q`I���j�!���撐�"W��      F�B�MR?��5���&��3��J��߮Ҽ/F����b=�I?�b.����/��qk����9�ճ:�;K!;m3;��=;��C;*�F;cH;��H;�I;I;�I;$I;�I;�I;D�H;��H;��H;|�H;?�H;|�H;3�H;|�H;?�H;|�H;��H;��H;D�H;�I;�I;$I;�I;I;�I;��H;cH;*�F;��C;��=;m3;K!;�;�ճ:���9�qk���/�b.��I?�b=���/F��߮Ҽ�J���3���&��5�MR?�      F��	}�;�ݼ��˼"d��-��	�}�&�G������һ�������"/�n:�ճ:#�;�a;Ģ0;�<;��B;�HF;vH;,�H;�I;zI;I;8I;Y	I;�I;�H;/�H;T�H;�H;#�H;�H;r�H;5�H;r�H;�H;#�H;�H;T�H;/�H;�H;�I;Y	I;8I;I;zI;�I;,�H;vH;�HF;��B;�<;Ģ0;�a;#�;�ճ:n:�"/���������һ���&�G�	�}�-��"d����˼;�ݼ	}�      ����8����_�k�ɆO�4/�VB�\�׻����@��Q�����+�>:i3�:�;�a;��/;=;;J�A;��E;ʾG;��H;�	I;hI;I;�I;�I;�I;� I;��H;;�H;��H;��H;��H;�H;d�H;)�H;d�H;�H;��H;��H;��H;;�H;��H;� I;�I;�I;�I;I;hI;�	I;��H;ʾG;��E;J�A;=;;��/;�a;�;i3�:+�>:����Q���@����\�׻VB�4/�ɆO�_�k���8��      ������q
�q�����׻S,��!����;�Rnۺ9� �J�9<Ǌ:���:� ;K!;Ģ0;=;;͒A;�oE;}�G;ԍH;��H;�I;9I;ZI; I;�I;oI;��H;=�H;x�H;�H;�H;��H;��H;[�H;1�H;[�H;��H;��H;�H;�H;x�H;=�H;��H;oI;�I; I;ZI;9I;�I;��H;ԍH;}�G;�oE;͒A;=;;Ģ0;K!;� ;���:<Ǌ:J�99� �Rnۺ�;�!���S,����׻q����q
���      �/��s�����x�k�X�b�/�ʻ �����u�q3�9��k:�:�m�:�A;!&;m3;�<;J�A;�oE;isG;�{H;.�H;,I;rI;CI;�I;i	I;�I;L�H;I�H;�H;��H;x�H;��H;��H;��H;l�H;\�H;l�H;��H;��H;��H;x�H;��H;�H;I�H;L�H;�I;i	I;�I;CI;rI;,I;.�H;�{H;isG;�oE;J�A;�<;m3;!&;�A;�m�:�:��k:q3�9u칉���ʻ �b�/�k�X���x�s���      ��������wk��� ��
���!69��!:Ǌ:�2�:C�:��;(;w�,;�6;��=;��B;��E;}�G;�{H;��H;zI;I;�I;WI;�
I;"I;� I;A�H;��H;4�H;��H;�H;��H;��H;��H;~�H;l�H;~�H;��H;��H;��H;�H;��H;4�H;��H;A�H;� I;"I;�
I;WI;�I;I;zI;��H;�{H;}�G;��E;��B;��=;�6;w�,;(;��;C�:�2�:Ǌ:��!:�!69�
���� ��wk����      ��>::�G:��b:ѳ�:���:
3�:?)�:�h;p�;$a;:*;nq3;��:;� @;��C;�HF;ʾG;ԍH;.�H;zI;I;CI;9I;�I;I;VI;�H;��H;��H;p�H;B�H;��H;��H;��H;	�H;��H;y�H;��H;	�H;��H;��H;��H;B�H;p�H;��H;��H;�H;VI;I;�I;9I;CI;I;zI;.�H;ԍH;ʾG;�HF;��C;� @;��:;nq3;:*;$a;p�;�h;?)�:
3�:���:ѳ�:��b::�G:      �r�:���:�j�:p�;��	;�;Vy;6O$;y�,;��3;5�9;2�>;>�B;D1E;*�F;vH;��H;��H;,I;I;CI;�I;6I;�I;�I;��H;�H;G�H;��H;��H;��H;��H;��H;��H;)�H;��H;��H;��H;)�H;��H;��H;��H;��H;��H;��H;G�H;�H;��H;�I;�I;6I;�I;CI;I;,I;��H;��H;vH;*�F;D1E;>�B;2�>;5�9;��3;y�,;6O$;Vy;�;��	;p�;�j�:���:      eo ;!;#;)&;%*;o.;�3;�7;��;;Ai?;jjB;8�D;�wF;�G;cH;,�H;�	I;�I;rI;�I;9I;6I;�I;RI;4�H;��H;��H; �H;��H;�H;��H;x�H;��H;��H;E�H;�H;��H;�H;E�H;��H;��H;x�H;��H;�H;��H; �H;��H;��H;4�H;RI;�I;6I;9I;�I;rI;�I;�	I;,�H;cH;�G;�wF;8�D;jjB;Ai?;��;;�7;�3;o.;%*;)&;#;!;      �I6;'�6;ۖ7;�9;l;;0-=;li?;y�A;C�C;w1E;ۆF;t�G;�;H;��H;��H;�I;hI;9I;CI;WI;�I;�I;RI;E�H;��H;��H;Y�H;$�H;1�H;��H;~�H;e�H;��H;�H;��H;]�H;:�H;]�H;��H;�H;��H;e�H;~�H;��H;1�H;$�H;Y�H;��H;��H;E�H;RI;�I;�I;WI;CI;9I;hI;�I;��H;��H;�;H;t�G;ۆF;w1E;C�C;y�A;li?;0-=;l;;�9;ۖ7;'�6;      DA;(kA;��A;��B;�iC;o`D;�[E;IF;�G;��G;�MH;S�H;��H;�I;�I;zI;I;ZI;�I;�
I;I;�I;4�H;��H;��H;w�H;-�H;@�H;��H;��H;`�H;u�H;��H;O�H;��H;��H;��H;��H;��H;O�H;��H;u�H;`�H;��H;��H;@�H;-�H;w�H;��H;��H;4�H;�I;I;�
I;�I;ZI;I;zI;�I;�I;��H;S�H;�MH;��G;�G;IF;�[E;o`D;�iC;��B;��A;(kA;      �HF;�XF;�F;�F;�&G;�G;��G;:BH;R�H;p�H;��H;I;
I;�I;I;I;�I; I;i	I;"I;VI;��H;��H;��H;w�H;S�H;[�H;��H;��H;i�H;X�H;��H;&�H;��H;@�H;"�H;�H;"�H;@�H;��H;&�H;��H;X�H;i�H;��H;��H;[�H;S�H;w�H;��H;��H;��H;VI;"I;i	I; I;�I;I;I;�I;
I;I;��H;p�H;R�H;:BH;��G;�G;�&G;�F;�F;�XF;      �MH;�SH;�cH;�|H;�H;o�H;��H;��H;�
I;7I; I;/ I;�I;OI;�I;8I;�I;�I;�I;� I;�H;�H;��H;Y�H;-�H;[�H;��H;��H;X�H;[�H;��H;��H;d�H;��H;��H;��H;��H;��H;��H;��H;d�H;��H;��H;[�H;X�H;��H;��H;[�H;-�H;Y�H;��H;�H;�H;� I;�I;�I;�I;8I;�I;OI;�I;/ I; I;7I;�
I;��H;��H;o�H;�H;�|H;�cH;�SH;      �H;s�H;�I;�I;�I;�I;tI;�I;� I;wI;�I;�I;�I;I;$I;Y	I;�I;oI;L�H;A�H;��H;G�H; �H;$�H;@�H;��H;��H;k�H;O�H;��H;��H;;�H;��H;|�H;9�H;
�H;�H;
�H;9�H;|�H;��H;;�H;��H;��H;O�H;k�H;��H;��H;@�H;$�H; �H;G�H;��H;A�H;L�H;oI;�I;Y	I;$I;I;�I;�I;�I;wI;� I;�I;tI;�I;�I;�I;�I;s�H;      !I;!I;\!I;f!I;
!I;@ I;�I;nI;�I;�I;�I;�I;AI;�	I;�I;�I;� I;��H;I�H;��H;��H;��H;��H;1�H;��H;��H;X�H;O�H;��H;��H;/�H;��H;M�H;��H;��H;��H;��H;��H;��H;��H;M�H;��H;/�H;��H;��H;O�H;X�H;��H;��H;1�H;��H;��H;��H;��H;I�H;��H;� I;�I;�I;�	I;AI;�I;�I;�I;�I;nI;�I;@ I;
!I;f!I;\!I;!I;      �I;�I;I;5I;�I;aI;�I;xI;GI;�I;"I;�	I;�I;;I;�I;�H;��H;=�H;�H;4�H;p�H;��H;�H;��H;��H;i�H;[�H;��H;��H;�H;��H;C�H;��H;��H;g�H;J�H;:�H;J�H;g�H;��H;��H;C�H;��H;�H;��H;��H;[�H;i�H;��H;��H;�H;��H;p�H;4�H;�H;=�H;��H;�H;�I;;I;�I;�	I;"I;�I;GI;xI;�I;aI;�I;5I;I;�I;      I;�I;pI;�I;�I;TI;�I;I;.
I;&I;I;�I;�I;u�H;D�H;/�H;;�H;x�H;��H;��H;B�H;��H;��H;~�H;`�H;X�H;��H;��H;/�H;��H;'�H;��H;v�H;<�H;	�H;��H;��H;��H;	�H;<�H;v�H;��H;'�H;��H;/�H;��H;��H;X�H;`�H;~�H;��H;��H;B�H;��H;��H;x�H;;�H;/�H;D�H;u�H;�I;�I;I;&I;.
I;I;�I;TI;�I;�I;pI;�I;      �I;�I;BI;�
I;�	I;�I;|I;-I;�I;�I;@I;`�H;��H;��H;��H;T�H;��H;�H;x�H;�H;��H;��H;x�H;e�H;u�H;��H;��H;;�H;��H;C�H;��H;R�H;!�H;��H;��H;��H;��H;��H;��H;��H;!�H;R�H;��H;C�H;��H;;�H;��H;��H;u�H;e�H;x�H;��H;��H;�H;x�H;�H;��H;T�H;��H;��H;��H;`�H;@I;�I;�I;-I;|I;�I;�	I;�
I;BI;�I;      mI;FI;�I;qI;�I;�I;�I;�I;? I;��H;_�H;��H;s�H;�H;��H;�H;��H;�H;��H;��H;��H;��H;��H;��H;��H;&�H;d�H;��H;M�H;��H;v�H;!�H;��H;��H;��H;m�H;f�H;m�H;��H;��H;��H;!�H;v�H;��H;M�H;��H;d�H;&�H;��H;��H;��H;��H;��H;��H;��H;�H;��H;�H;��H;�H;s�H;��H;_�H;��H;? I;�I;�I;�I;�I;qI;�I;FI;      I;�I;�I;FI;� I;��H;�H;�H;�H;��H;��H;��H;5�H;��H;|�H;#�H;��H;��H;��H;��H;��H;��H;��H;�H;O�H;��H;��H;|�H;��H;��H;<�H;��H;��H;n�H;V�H;J�H;9�H;J�H;V�H;n�H;��H;��H;<�H;��H;��H;|�H;��H;��H;O�H;�H;��H;��H;��H;��H;��H;��H;��H;#�H;|�H;��H;5�H;��H;��H;��H;�H;�H;�H;��H;� I;FI;�I;�I;      q�H;e�H;!�H;��H;I�H;��H;��H;��H;�H;��H;��H;��H;o�H;^�H;?�H;�H;�H;��H;��H;��H;	�H;)�H;E�H;��H;��H;@�H;��H;9�H;��H;g�H;	�H;��H;��H;V�H;1�H;&�H;(�H;&�H;1�H;V�H;��H;��H;	�H;g�H;��H;9�H;��H;@�H;��H;��H;E�H;)�H;	�H;��H;��H;��H;�H;�H;?�H;^�H;o�H;��H;��H;��H;�H;��H;��H;��H;I�H;��H;!�H;e�H;      ��H;��H;x�H;"�H;��H;�H;c�H;��H;��H;��H;��H;��H;��H;��H;|�H;r�H;d�H;[�H;l�H;~�H;��H;��H;�H;]�H;��H;"�H;��H;
�H;��H;J�H;��H;��H;m�H;J�H;&�H;
�H;�H;
�H;&�H;J�H;m�H;��H;��H;J�H;��H;
�H;��H;"�H;��H;]�H;�H;��H;��H;~�H;l�H;[�H;d�H;r�H;|�H;��H;��H;��H;��H;��H;��H;��H;c�H;�H;��H;"�H;x�H;��H;      +�H;�H;��H;��H; �H;d�H;��H;�H;"�H;V�H;j�H;_�H;l�H;D�H;3�H;5�H;)�H;1�H;\�H;l�H;y�H;��H;��H;:�H;��H;�H;��H;�H;��H;:�H;��H;��H;f�H;9�H;(�H;�H;	�H;�H;(�H;9�H;f�H;��H;��H;:�H;��H;�H;��H;�H;��H;:�H;��H;��H;y�H;l�H;\�H;1�H;)�H;5�H;3�H;D�H;l�H;_�H;j�H;V�H;"�H;�H;��H;d�H; �H;��H;��H;�H;      ��H;��H;x�H;"�H;��H;�H;c�H;��H;��H;��H;��H;��H;��H;��H;|�H;r�H;d�H;[�H;l�H;~�H;��H;��H;�H;]�H;��H;"�H;��H;
�H;��H;J�H;��H;��H;m�H;J�H;&�H;
�H;�H;
�H;&�H;J�H;m�H;��H;��H;J�H;��H;
�H;��H;"�H;��H;]�H;�H;��H;��H;~�H;l�H;[�H;d�H;r�H;|�H;��H;��H;��H;��H;��H;��H;��H;c�H;�H;��H;"�H;x�H;��H;      q�H;e�H;!�H;��H;I�H;��H;��H;��H;�H;��H;��H;��H;o�H;^�H;?�H;�H;�H;��H;��H;��H;	�H;)�H;E�H;��H;��H;@�H;��H;9�H;��H;g�H;	�H;��H;��H;V�H;1�H;&�H;(�H;&�H;1�H;V�H;��H;��H;	�H;g�H;��H;9�H;��H;@�H;��H;��H;E�H;)�H;	�H;��H;��H;��H;�H;�H;?�H;^�H;o�H;��H;��H;��H;�H;��H;��H;��H;I�H;��H;!�H;e�H;      I;�I;�I;FI;� I;��H;�H;�H;�H;��H;��H;��H;5�H;��H;|�H;#�H;��H;��H;��H;��H;��H;��H;��H;�H;O�H;��H;��H;|�H;��H;��H;<�H;��H;��H;n�H;V�H;J�H;9�H;J�H;V�H;n�H;��H;��H;<�H;��H;��H;|�H;��H;��H;O�H;�H;��H;��H;��H;��H;��H;��H;��H;#�H;|�H;��H;5�H;��H;��H;��H;�H;�H;�H;��H;� I;FI;�I;�I;      mI;FI;�I;qI;�I;�I;�I;�I;? I;��H;_�H;��H;s�H;�H;��H;�H;��H;�H;��H;��H;��H;��H;��H;��H;��H;&�H;d�H;��H;M�H;��H;v�H;!�H;��H;��H;��H;m�H;f�H;m�H;��H;��H;��H;!�H;v�H;��H;M�H;��H;d�H;&�H;��H;��H;��H;��H;��H;��H;��H;�H;��H;�H;��H;�H;s�H;��H;_�H;��H;? I;�I;�I;�I;�I;qI;�I;FI;      �I;�I;BI;�
I;�	I;�I;|I;-I;�I;�I;@I;`�H;��H;��H;��H;T�H;��H;�H;x�H;�H;��H;��H;x�H;e�H;u�H;��H;��H;;�H;��H;C�H;��H;R�H;!�H;��H;��H;��H;��H;��H;��H;��H;!�H;R�H;��H;C�H;��H;;�H;��H;��H;u�H;e�H;x�H;��H;��H;�H;x�H;�H;��H;T�H;��H;��H;��H;`�H;@I;�I;�I;-I;|I;�I;�	I;�
I;BI;�I;      I;�I;pI;�I;�I;TI;�I;I;.
I;&I;I;�I;�I;u�H;D�H;/�H;;�H;x�H;��H;��H;B�H;��H;��H;~�H;`�H;X�H;��H;��H;/�H;��H;'�H;��H;v�H;<�H;	�H;��H;��H;��H;	�H;<�H;v�H;��H;'�H;��H;/�H;��H;��H;X�H;`�H;~�H;��H;��H;B�H;��H;��H;x�H;;�H;/�H;D�H;u�H;�I;�I;I;&I;.
I;I;�I;TI;�I;�I;pI;�I;      �I;�I;I;5I;�I;aI;�I;xI;GI;�I;"I;�	I;�I;;I;�I;�H;��H;=�H;�H;4�H;p�H;��H;�H;��H;��H;i�H;[�H;��H;��H;�H;��H;C�H;��H;��H;g�H;J�H;:�H;J�H;g�H;��H;��H;C�H;��H;�H;��H;��H;[�H;i�H;��H;��H;�H;��H;p�H;4�H;�H;=�H;��H;�H;�I;;I;�I;�	I;"I;�I;GI;xI;�I;aI;�I;5I;I;�I;      !I;!I;\!I;f!I;
!I;@ I;�I;nI;�I;�I;�I;�I;AI;�	I;�I;�I;� I;��H;I�H;��H;��H;��H;��H;1�H;��H;��H;X�H;O�H;��H;��H;/�H;��H;M�H;��H;��H;��H;��H;��H;��H;��H;M�H;��H;/�H;��H;��H;O�H;X�H;��H;��H;1�H;��H;��H;��H;��H;I�H;��H;� I;�I;�I;�	I;AI;�I;�I;�I;�I;nI;�I;@ I;
!I;f!I;\!I;!I;      �H;s�H;�I;�I;�I;�I;tI;�I;� I;wI;�I;�I;�I;I;$I;Y	I;�I;oI;L�H;A�H;��H;G�H; �H;$�H;@�H;��H;��H;k�H;O�H;��H;��H;;�H;��H;|�H;9�H;
�H;�H;
�H;9�H;|�H;��H;;�H;��H;��H;O�H;k�H;��H;��H;@�H;$�H; �H;G�H;��H;A�H;L�H;oI;�I;Y	I;$I;I;�I;�I;�I;wI;� I;�I;tI;�I;�I;�I;�I;s�H;      �MH;�SH;�cH;�|H;�H;o�H;��H;��H;�
I;7I; I;/ I;�I;OI;�I;8I;�I;�I;�I;� I;�H;�H;��H;Y�H;-�H;[�H;��H;��H;X�H;[�H;��H;��H;d�H;��H;��H;��H;��H;��H;��H;��H;d�H;��H;��H;[�H;X�H;��H;��H;[�H;-�H;Y�H;��H;�H;�H;� I;�I;�I;�I;8I;�I;OI;�I;/ I; I;7I;�
I;��H;��H;o�H;�H;�|H;�cH;�SH;      �HF;�XF;�F;�F;�&G;�G;��G;:BH;R�H;p�H;��H;I;
I;�I;I;I;�I; I;i	I;"I;VI;��H;��H;��H;w�H;S�H;[�H;��H;��H;i�H;X�H;��H;&�H;��H;@�H;"�H;�H;"�H;@�H;��H;&�H;��H;X�H;i�H;��H;��H;[�H;S�H;w�H;��H;��H;��H;VI;"I;i	I; I;�I;I;I;�I;
I;I;��H;p�H;R�H;:BH;��G;�G;�&G;�F;�F;�XF;      DA;(kA;��A;��B;�iC;o`D;�[E;IF;�G;��G;�MH;S�H;��H;�I;�I;zI;I;ZI;�I;�
I;I;�I;4�H;��H;��H;w�H;-�H;@�H;��H;��H;`�H;u�H;��H;O�H;��H;��H;��H;��H;��H;O�H;��H;u�H;`�H;��H;��H;@�H;-�H;w�H;��H;��H;4�H;�I;I;�
I;�I;ZI;I;zI;�I;�I;��H;S�H;�MH;��G;�G;IF;�[E;o`D;�iC;��B;��A;(kA;      �I6;'�6;ۖ7;�9;l;;0-=;li?;y�A;C�C;w1E;ۆF;t�G;�;H;��H;��H;�I;hI;9I;CI;WI;�I;�I;RI;E�H;��H;��H;Y�H;$�H;1�H;��H;~�H;e�H;��H;�H;��H;]�H;:�H;]�H;��H;�H;��H;e�H;~�H;��H;1�H;$�H;Y�H;��H;��H;E�H;RI;�I;�I;WI;CI;9I;hI;�I;��H;��H;�;H;t�G;ۆF;w1E;C�C;y�A;li?;0-=;l;;�9;ۖ7;'�6;      eo ;!;#;)&;%*;o.;�3;�7;��;;Ai?;jjB;8�D;�wF;�G;cH;,�H;�	I;�I;rI;�I;9I;6I;�I;RI;4�H;��H;��H; �H;��H;�H;��H;x�H;��H;��H;E�H;�H;��H;�H;E�H;��H;��H;x�H;��H;�H;��H; �H;��H;��H;4�H;RI;�I;6I;9I;�I;rI;�I;�	I;,�H;cH;�G;�wF;8�D;jjB;Ai?;��;;�7;�3;o.;%*;)&;#;!;      �r�:���:�j�:p�;��	;�;Vy;6O$;y�,;��3;5�9;2�>;>�B;D1E;*�F;vH;��H;��H;,I;I;CI;�I;6I;�I;�I;��H;�H;G�H;��H;��H;��H;��H;��H;��H;)�H;��H;��H;��H;)�H;��H;��H;��H;��H;��H;��H;G�H;�H;��H;�I;�I;6I;�I;CI;I;,I;��H;��H;vH;*�F;D1E;>�B;2�>;5�9;��3;y�,;6O$;Vy;�;��	;p�;�j�:���:      ��>::�G:��b:ѳ�:���:
3�:?)�:�h;p�;$a;:*;nq3;��:;� @;��C;�HF;ʾG;ԍH;.�H;zI;I;CI;9I;�I;I;VI;�H;��H;��H;p�H;B�H;��H;��H;��H;	�H;��H;y�H;��H;	�H;��H;��H;��H;B�H;p�H;��H;��H;�H;VI;I;�I;9I;CI;I;zI;.�H;ԍH;ʾG;�HF;��C;� @;��:;nq3;:*;$a;p�;�h;?)�:
3�:���:ѳ�:��b::�G:      ��������wk��� ��
���!69��!:Ǌ:�2�:C�:��;(;w�,;�6;��=;��B;��E;}�G;�{H;��H;zI;I;�I;WI;�
I;"I;� I;A�H;��H;4�H;��H;�H;��H;��H;��H;~�H;l�H;~�H;��H;��H;��H;�H;��H;4�H;��H;A�H;� I;"I;�
I;WI;�I;I;zI;��H;�{H;}�G;��E;��B;��=;�6;w�,;(;��;C�:�2�:Ǌ:��!:�!69�
���� ��wk����      �/��s�����x�k�X�b�/�ʻ �����u�q3�9��k:�:�m�:�A;!&;m3;�<;J�A;�oE;isG;�{H;.�H;,I;rI;CI;�I;i	I;�I;L�H;I�H;�H;��H;x�H;��H;��H;��H;l�H;\�H;l�H;��H;��H;��H;x�H;��H;�H;I�H;L�H;�I;i	I;�I;CI;rI;,I;.�H;�{H;isG;�oE;J�A;�<;m3;!&;�A;�m�:�:��k:q3�9u칉���ʻ �b�/�k�X���x�s���      ������q
�q�����׻S,��!����;�Rnۺ9� �J�9<Ǌ:���:� ;K!;Ģ0;=;;͒A;�oE;}�G;ԍH;��H;�I;9I;ZI; I;�I;oI;��H;=�H;x�H;�H;�H;��H;��H;[�H;1�H;[�H;��H;��H;�H;�H;x�H;=�H;��H;oI;�I; I;ZI;9I;�I;��H;ԍH;}�G;�oE;͒A;=;;Ģ0;K!;� ;���:<Ǌ:J�99� �Rnۺ�;�!���S,����׻q����q
���      ����8����_�k�ɆO�4/�VB�\�׻����@��Q�����+�>:i3�:�;�a;��/;=;;J�A;��E;ʾG;��H;�	I;hI;I;�I;�I;�I;� I;��H;;�H;��H;��H;��H;�H;d�H;)�H;d�H;�H;��H;��H;��H;;�H;��H;� I;�I;�I;�I;I;hI;�	I;��H;ʾG;��E;J�A;=;;��/;�a;�;i3�:+�>:����Q���@����\�׻VB�4/�ɆO�_�k���8��      F��	}�;�ݼ��˼"d��-��	�}�&�G������һ�������"/�n:�ճ:#�;�a;Ģ0;�<;��B;�HF;vH;,�H;�I;zI;I;8I;Y	I;�I;�H;/�H;T�H;�H;#�H;�H;r�H;5�H;r�H;�H;#�H;�H;T�H;/�H;�H;�I;Y	I;8I;I;zI;�I;,�H;vH;�HF;��B;�<;Ģ0;�a;#�;�ճ:n:�"/���������һ���&�G�	�}�-��"d����˼;�ݼ	}�      F�B�MR?��5���&��3��J��߮Ҽ/F����b=�I?�b.����/��qk����9�ճ:�;K!;m3;��=;��C;*�F;cH;��H;�I;I;�I;$I;�I;�I;D�H;��H;��H;|�H;?�H;|�H;3�H;|�H;?�H;|�H;��H;��H;D�H;�I;�I;$I;�I;I;�I;��H;cH;*�F;��C;��=;m3;K!;�;�ճ:���9�qk���/�b.��I?�b=���/F��߮Ҽ�J���3���&��5�MR?�      &��"W��撐�!�����j�Q`I���&����Oϼ�,���T[����I��;��qk�n:i3�:� ;!&;�6;� @;D1E;�G;��H;�I;�I;OI;I;�	I;;I;u�H;��H;�H;��H;^�H;��H;D�H;��H;^�H;��H;�H;��H;u�H;;I;�	I;I;OI;�I;�I;��H;�G;D1E;� @;�6;!&;� ;i3�:n:�qk�;��I�����T[��,��Oϼ�����&�Q`I���j�!���撐�"W��      �J���D��ͽ���$�������L�(��.��;��%�k����I����/��"/�+�>:���:�A;w�,;��:;>�B;�wF;�;H;��H;
I;�I;�I;AI;�I;�I;��H;s�H;5�H;o�H;��H;l�H;��H;o�H;5�H;s�H;��H;�I;�I;AI;�I;�I;
I;��H;�;H;�wF;>�B;��:;w�,;�A;���:+�>:�"/���/��I����%�k�;��.��(����L����$������ͽ�Dὼ��      K�:��*7���,�+�~�	�j��~���W����j�?�/��J���I��%�k���b.�������<Ǌ:�m�:(;nq3;2�>;8�D;t�G;S�H;I;/ I;�I;�I;�	I;�I;`�H;��H;��H;��H;��H;_�H;��H;��H;��H;��H;`�H;�I;�	I;�I;�I;/ I;I;S�H;t�G;8�D;2�>;nq3;(;�m�:<Ǌ:�����b.����%�k��I���J��?�/���j�W��~���j��~�	�+���,��*7�      ^���p��
��)�l���M���,�Tl�K9ݽ�A���{���5��J��;���T[�I?������Q��J�9�:��;:*;5�9;jjB;ۆF;�MH;��H; I;�I;�I;"I;I;@I;_�H;��H;��H;��H;j�H;��H;��H;��H;_�H;@I;I;"I;�I;�I; I;��H;�MH;ۆF;jjB;5�9;:*;��;�:J�9�Q������I?��T[�;���J����5��{��A��K9ݽTl���,���M�)�l�
���p��      +m־G�Ѿ�>ľ����̗����{���I�+����V���{�?�/�.���,��b=���һ�@�9� ���k:C�:$a;��3;Ai?;w1E;��G;p�H;7I;wI;�I;�I;&I;�I;��H;��H;��H;��H;V�H;��H;��H;��H;��H;�I;&I;�I;�I;wI;7I;p�H;��G;w1E;Ai?;��3;$a;C�:��k:9� ��@���һb=��,��.��?�/��{��V�����+���I���{�̗�������>ľG�Ѿ      =\����l5��z ��E۾�ճ��]��q�Z�F?#����A����j�(��Oϼ��������Rnۺq3�9�2�:p�;y�,;��;;C�C;�G;R�H;�
I;� I;�I;GI;.
I;�I;? I;�H;�H;��H;"�H;��H;�H;�H;? I;�I;.
I;GI;�I;� I;�
I;R�H;�G;C�C;��;;y�,;p�;�2�:q3�9Rnۺ��������Oϼ(����j��A�����F?#�q�Z��]���ճ��E۾�z �l5����      <�b��>]���M���6�����$���>ľq��q�Z�+�K9ݽW����L����/F��&�G�\�׻�;�u�Ǌ:�h;6O$;�7;y�A;IF;:BH;��H;�I;nI;xI;I;-I;�I;�H;��H;��H;�H;��H;��H;�H;�I;-I;I;xI;nI;�I;��H;:BH;IF;y�A;�7;6O$;�h;Ǌ:u칸;�\�׻&�G�/F�������L�W��K9ݽ+�q�Z�q���>ľ�$�������6���M��>]�      �o��벗����-�y�s�R���)�iv��>ľ�]����I�Tl�~��������&�߮Ҽ	�}�VB�!���������!:?)�:Vy;�3;li?;�[E;��G;��H;tI;�I;�I;�I;|I;�I;�H;��H;c�H;��H;c�H;��H;�H;�I;|I;�I;�I;�I;tI;��H;��G;�[E;li?;�3;Vy;?)�:��!:����!���VB�	�}�߮Ҽ��&����~���Tl���I��]���>ľiv���)�s�R�-�y����벗�      �˿�<ƿjL��:1��蟉��>]���)��$���ճ���{���,�j��$��Q`I��J��-��4/�S,��ʻ ��!69
3�:�;o.;0-=;o`D;�G;o�H;�I;@ I;aI;TI;�I;�I;��H;��H;�H;d�H;�H;��H;��H;�I;�I;TI;aI;@ I;�I;o�H;�G;o`D;0-=;o.;�;
3�:�!69ʻ �S,��4/�-���J��Q`I�$��j�齞�,���{��ճ��$����)��>]�蟉�:1��jL���<ƿ      ����2���K[忭˿�T��蟉�s�R�����E۾̗����M�~�	������j��3�"d��ɆO���׻b�/��
�����:��	;%*;l;;�iC;�&G;�H;�I;
!I;�I;�I;�	I;�I;� I;I�H;��H; �H;��H;I�H;� I;�I;�	I;�I;�I;
!I;�I;�H;�&G;�iC;l;;%*;��	;���:�
��b�/���׻ɆO�"d���3���j����~�	���M�̗���E۾���s�R�蟉��T���˿K[�2���      O�0��o����˿:1��-�y���6��z �����)�l�+��ͽ!�����&���˼_�k�q���k�X��� �ѳ�:p�;)&;�9;��B;�F;�|H;�I;f!I;5I;�I;�
I;qI;FI;��H;"�H;��H;"�H;��H;FI;qI;�
I;�I;5I;f!I;�I;�|H;�F;��B;�9;)&;p�;ѳ�:�� �k�X�q���_�k���˼��&�!����ͽ+�)�l������z ���6�-�y�:1���˿���o�0��      ��*��g&��#�o�K[�jL�������M�l5��>ľ
����,��D�撐��5�;�ݼ���q
���x��wk���b:�j�:#;ۖ7;��A;�F;�cH;�I;\!I;I;pI;BI;�I;�I;!�H;x�H;��H;x�H;!�H;�I;�I;BI;pI;I;\!I;�I;�cH;�F;��A;ۖ7;#;�j�:��b:�wk���x��q
���;�ݼ�5�撐��Dὤ�,�
���>ľl5���M����jL��K[�o��#��g&�      ��8��4��g&�0��2����<ƿ벗��>]����G�Ѿ�p���*7����"W��MR?�	}�8����s������:�G:���:!;'�6;(kA;�XF;�SH;s�H;!I;�I;�I;�I;FI;�I;e�H;��H;�H;��H;e�H;�I;FI;�I;�I;�I;!I;s�H;�SH;�XF;(kA;'�6;!;���::�G:���s�����8��	}�MR?�"W�����*7��p��G�Ѿ����>]�벗��<ƿ2���0���g&��4�      ���$������꿥�ſ�ޞ�3s��2�/����� j���nHͽ������'�B<ͼ��n������Q^�0.��:�V;�R%;~n8;��A;nCF;�H;��H;��H;��H;L�H;>�H;C�H;��H;��H;��H;+�H;��H;��H;��H;C�H;>�H;L�H;��H;��H;��H;�H;nCF;��A;~n8;�R%;�V;�:0.��Q^�������n�B<ͼ��'�����nHͽ�� j���/����2�3s��ޞ���ſ������$�      $��������~�����cm�L�-�����Fh��Ide�-�̪ɽ�v��#�$���ɼ�mj�o����X�5��nĆ:�w;i�%;M�8;B;{QF;H;5�H;U�H;	�H;p�H;B�H;6�H;��H;��H;��H;$�H;��H;��H;��H;6�H;B�H;p�H;	�H;U�H;5�H;H;{QF;B;M�8;i�%;�w;nĆ:5���X�o����mj���ɼ#�$��v��̪ɽ-�Ide�Fh������L�-�cm����~���忖����      ������{���ԿBw�����/�\��"����b��M0X�}���;����w����������]�W��UF�+��pȒ:1�;_�';؎9;2oB;�yF;� H;��H;7�H;�H;��H;F�H;:�H;��H;��H;��H;�H;��H;��H;��H;:�H;F�H;��H;�H;7�H;��H;� H;�yF;2oB;؎9;_�';1�;pȒ:+��UF�W�黼�]����������w��;��}��M0X�b������"�/�\����Bw���Կ{�𿖏�      ������Կp���ޞ�RF�]�C�$E��;�I��sD�|�"��]�c�y��֯���J�O�ѻ\�)���K����:Q�
;M*;��:;�C;�F;�7H;Z�H;��H;w�H;��H;>�H;:�H;��H;��H;��H;��H;��H;��H;��H;:�H;>�H;��H;w�H;��H;Z�H;�7H;�F;�C;��:;M*;Q�
;���:��K�\�)�O�ѻ��J��֯�y�]�c�"��|�sD��I���;$E�]�C�RF��ޞ�p���Կ��      ��ſ~��Bw���ޞ�|���3�W�,�%�����^ɰ��|x�\{+�ű����J��  �Ҷ��n�1�f����+�
9r�:�;5�-;��<;��C;�G;�SH;Q�H;��H;��H;��H;V�H;3�H;��H;��H;��H;��H;��H;��H;��H;3�H;V�H;��H;��H;��H;Q�H;�SH;�G;��C;��<;5�-;�;r�:
9�+�f���n�1�Ҷ���  ��J���ű�\{+��|x�^ɰ�����,�%�3�W�|����ޞ�Bw��~��      �ޞ�������RF�3�W�M�-���4Kɾ�G����O�z��ƽ����Ȅ-���ۼㄼL4�[ǐ�+ж��Z:o��:�;ʕ1;
c>;|�D;�[G;KrH;��H;i�H;e�H;'�H;u�H;)�H;h�H;��H;|�H;��H;|�H;��H;h�H;)�H;u�H;'�H;e�H;i�H;��H;KrH;�[G;|�D;
c>;ʕ1;�;o��:�Z:+ж�[ǐ�L4�ㄼ��ۼȄ-�����ƽz����O��G��4Kɾ��M�-�3�W�RF�������      3s�cm�/�\�]�C�,�%����TҾa����i��C(����UP����[�x������Y�k���X���<���k:���:)� ;�5;ZQ@;otE;�G;9�H;L�H;��H;�H;I�H;l�H;$�H;c�H;s�H;X�H;��H;X�H;s�H;c�H;$�H;l�H;I�H;�H;��H;L�H;9�H;�G;otE;ZQ@;�5;)� ;���:��k:��<��X�k����Y����x���[�UP����콡C(���i�a���TҾ��,�%�]�C�/�\�cm�      �2�L�-��"�$E�����4Kɾa��w�s�.�5�y�k㻽�v��z0��;��+��-�*�R����6�jS�L�:��	;��(;6�9;�.B;�CF;YH;ժH;��H;��H;��H;w�H;��H;�H;0�H;C�H;<�H;Y�H;<�H;C�H;0�H;�H;��H;w�H;��H;��H;��H;ժH;YH;�CF;�.B;6�9;��(;��	;L�:jS��6�R���-�*��+���;�z0��v��k㻽y�.�5�w�s�a��4Kɾ����$E��"�L�-�      /�����������;^ɰ��G����i�.�5��	�ĪɽR����J�p���沼��]�I���U
x��
���k:6��:v;��/;�,=;��C;N�F;#HH;��H;(�H;��H;#�H;��H;��H;��H;�H;�H;�H;$�H;�H;�H;�H;��H;��H;��H;#�H;��H;(�H;��H;#HH;N�F;��C;�,=;��/;v;6��:�k:�
��U
x�I�����]��沼p���J�R���Īɽ�	�.�5���i��G��^ɰ��;��徨���      ��Fh��b���I���|x���O��C(�y�Īɽ����IDX�D��'<ͼㄼ�X!�t��hX��K����:�x;7�#;$H6;IQ@;�OE;��G;��H;��H;2�H;��H;��H;��H;v�H;��H;��H;��H;��H;��H;��H;��H;��H;��H;v�H;��H;��H;��H;2�H;��H;��H;��G;�OE;IQ@;$H6;7�#;�x;���:�K�hX�t���X!�ㄼ'<ͼD��IDX�����Īɽy��C(���O��|x��I��b��Fh��       j�Ide�M0X�sD�\{+�z�����k㻽R���IDX������ۼо����;�>ۻ�X���y�><":J��:��;��-;��;;�B;�yF;�H;��H;|�H;&�H;��H;��H;��H;n�H;��H;��H;��H;��H;z�H;��H;��H;��H;��H;n�H;��H;��H;��H;&�H;|�H;��H;�H;�yF;�B;��;;��-;��;J��:><":��y��X�>ۻ��;�о����ۼ���IDX�R���k㻽���z��\{+�sD�M0X�Ide�      ��-�}��|�ű�ƽUP���v���J�D����ۼ��u�J������+���sѺ0
9gL�:�;�$;#�5;�?;��D;j[G;eH;��H;��H;��H;��H;!�H;��H;T�H;n�H;Y�H;T�H;a�H;7�H;a�H;T�H;Y�H;n�H;T�H;��H;!�H;��H;��H;��H;��H;eH;j[G;��D;�?;#�5;�$;�;gL�:0
9�sѺ�+������u�J�����ۼD���J��v��UP��ƽű�|�}��-�      nHͽ̪ɽ�;��"����������[�z0�p��'<ͼо��u�J���k��+��(����:�`�:}�;�/;�K<;!C;9lF;��G;�H;�H;�H;�H;A�H;T�H;��H;%�H;/�H;�H;�H;�H;��H;�H;�H;�H;/�H;%�H;��H;T�H;A�H;�H;�H;�H;�H;��G;9lF;!C;�K<;�/;}�;�`�:���:�(�+�k����u�J�о��'<ͼp��z0���[�������"���;��̪ɽ      �����v����w�]�c��J�Ȅ-�x��;缈沼ㄼ��;�����k��56�c��N<Q:ף�:�h;M*;��8;��@;�OE;�tG;DhH;��H;��H;�H;#�H;��H;y�H;��H;��H;��H;��H;��H;��H;��H;��H;��H;��H;��H;��H;��H;y�H;��H;#�H;�H;��H;��H;DhH;�tG;�OE;��@;��8;M*;�h;ף�:N<Q:c��56�k��������;�ㄼ�沼�;�x�Ȅ-��J�]�c���w��v��      ��'�#�$����y��  ���ۼ����+����]��X!�>ۻ�+��+�c���>:]��:@�;Z�%;	�5;��>;�'D;�F;� H;8�H;[�H;��H;��H;��H;��H;k�H;��H;��H;��H;��H;h�H;K�H;m�H;K�H;h�H;��H;��H;��H;��H;k�H;��H;��H;��H;��H;[�H;8�H;� H;�F;�'D;��>;	�5;Z�%;@�;]��:�>:c��+��+��>ۻ�X!���]��+�������ۼ�  �y����#�$�      B<ͼ��ɼ�����֯�Ҷ��ㄼ��Y�-�*�I���t���X��sѺ�(�N<Q:]��:��
;v�#;��3;�b=;#C;3CF;�G;�H;��H;�H;9�H;��H;X�H;!�H;d�H;��H;b�H;5�H;O�H;	�H;��H;�H;��H;	�H;O�H;5�H;b�H;��H;d�H;!�H;X�H;��H;9�H;�H;��H;�H;�G;3CF;#C;�b=;��3;v�#;��
;]��:N<Q:�(��sѺ�X�t��I���-�*���Y�ㄼҶ���֯�������ɼ      ��n��mj���]���J�n�1�L4�k��R���U
x�hX���y�0
9���:ף�:@�;v�#;w�2;�<;�oB;7�E;��G;�dH;��H;8�H;��H;��H;��H;��H;9�H;F�H;8�H;�H;��H;��H;��H;��H;��H;��H;��H;��H;��H;�H;8�H;F�H;9�H;��H;��H;��H;��H;8�H;��H;�dH;��G;7�E;�oB;�<;w�2;v�#;@�;ף�:���:0
9��y�hX�U
x�R���k��L4�n�1���J���]��mj�      ����o���W��O�ѻf���[ǐ��X��6��
���K�><":gL�:�`�:�h;Z�%;��3;�<;Y/B;��E;�[G;�GH;N�H;��H;a�H;�H;7�H;=�H;��H;�H;�H;��H;��H;��H;]�H;O�H;K�H;'�H;K�H;O�H;]�H;��H;��H;��H;�H;�H;��H;=�H;7�H;�H;a�H;��H;N�H;�GH;�[G;��E;Y/B;�<;��3;Z�%;�h;�`�:gL�:><":�K��
���6��X�[ǐ�f���O�ѻW��o���      �Q^��X�UF�\�)��+�+ж���<�jS��k:���:J��:�;}�;M*;	�5;�b=;�oB;��E;�IG;]7H;s�H;��H;�H;-�H;��H;��H;��H;��H;��H;��H;��H;u�H;P�H;��H;��H;��H;��H;��H;��H;��H;P�H;u�H;��H;��H;��H;��H;��H;��H;��H;-�H;�H;��H;s�H;]7H;�IG;��E;�oB;�b=;	�5;M*;}�;�;J��:���:�k:jS���<�+ж��+�\�)�UF��X�      0.�5��+�깙�K�
9�Z:��k:L�:6��:�x;��;�$;�/;��8;��>;#C;7�E;�[G;]7H;ͤH;�H;&�H;��H;5�H;��H;P�H;��H;��H;��H;z�H;5�H;�H;��H;��H;��H;��H;u�H;��H;��H;��H;��H;�H;5�H;z�H;��H;��H;��H;P�H;��H;5�H;��H;&�H;�H;ͤH;]7H;�[G;7�E;#C;��>;��8;�/;�$;��;�x;6��:L�:��k:�Z:
9��K�+��5��      �:nĆ:pȒ:���:r�:o��:���:��	;v;7�#;��-;#�5;�K<;��@;�'D;3CF;��G;�GH;s�H;�H;��H;P�H;��H;\�H;#�H;��H;��H;��H;[�H;�H;��H;��H;m�H;[�H;*�H;�H;�H;�H;*�H;[�H;m�H;��H;��H;�H;[�H;��H;��H;��H;#�H;\�H;��H;P�H;��H;�H;s�H;�GH;��G;3CF;�'D;��@;�K<;#�5;��-;7�#;v;��	;���:o��:r�:���:pȒ:nĆ:      �V;�w;1�;Q�
;�;�;)� ;��(;��/;$H6;��;;�?;!C;�OE;�F;�G;�dH;N�H;��H;&�H;P�H;��H;1�H;��H;f�H;�H;��H;b�H;��H;��H;��H;B�H;�H;�H;��H;��H;��H;��H;��H;�H;�H;B�H;��H;��H;��H;b�H;��H;�H;f�H;��H;1�H;��H;P�H;&�H;��H;N�H;�dH;�G;�F;�OE;!C;�?;��;;$H6;��/;��(;)� ;�;�;Q�
;1�;�w;      �R%;i�%;_�';M*;5�-;ʕ1;�5;6�9;�,=;IQ@;�B;��D;9lF;�tG;� H;�H;��H;��H;�H;��H;��H;1�H;�H;b�H;��H;r�H;5�H;��H;��H;��H;�H;��H;��H;��H;}�H;e�H;L�H;e�H;}�H;��H;��H;��H;�H;��H;��H;��H;5�H;r�H;��H;b�H;�H;1�H;��H;��H;�H;��H;��H;�H;� H;�tG;9lF;��D;�B;IQ@;�,=;6�9;�5;ʕ1;5�-;M*;_�';i�%;      ~n8;M�8;؎9;��:;��<;
c>;ZQ@;�.B;��C;�OE;�yF;j[G;��G;DhH;8�H;��H;8�H;a�H;-�H;5�H;\�H;��H;b�H;k�H;j�H;D�H;��H;��H;e�H;	�H;��H;��H;Y�H;(�H;"�H;�H;��H;�H;"�H;(�H;Y�H;��H;��H;	�H;e�H;��H;��H;D�H;j�H;k�H;b�H;��H;\�H;5�H;-�H;a�H;8�H;��H;8�H;DhH;��G;j[G;�yF;�OE;��C;�.B;ZQ@;
c>;��<;��:;؎9;M�8;      ��A;B;2oB;�C;��C;|�D;otE;�CF;N�F;��G;�H;eH;�H;��H;[�H;�H;��H;�H;��H;��H;#�H;f�H;��H;j�H;-�H;��H;��H;i�H; �H;��H;r�H;@�H;�H;��H;��H;��H;��H;��H;��H;��H;�H;@�H;r�H;��H; �H;i�H;��H;��H;-�H;j�H;��H;f�H;#�H;��H;��H;�H;��H;�H;[�H;��H;�H;eH;�H;��G;N�F;�CF;otE;|�D;��C;�C;2oB;B;      nCF;{QF;�yF;�F;�G;�[G;�G;YH;#HH;��H;��H;��H;�H;��H;��H;9�H;��H;7�H;��H;P�H;��H;�H;r�H;D�H;��H;��H;_�H;��H;��H;a�H;�H;��H;��H;��H;o�H;\�H;n�H;\�H;o�H;��H;��H;��H;�H;a�H;��H;��H;_�H;��H;��H;D�H;r�H;�H;��H;P�H;��H;7�H;��H;9�H;��H;��H;�H;��H;��H;��H;#HH;YH;�G;�[G;�G;�F;�yF;{QF;      �H;H;� H;�7H;�SH;KrH;9�H;ժH;��H;��H;|�H;��H;�H;�H;��H;��H;��H;=�H;��H;��H;��H;��H;5�H;��H;��H;_�H;��H;��H;H�H;�H;��H;��H;b�H;D�H;(�H;�H;�H;�H;(�H;D�H;b�H;��H;��H;�H;H�H;��H;��H;_�H;��H;��H;5�H;��H;��H;��H;��H;=�H;��H;��H;��H;�H;�H;��H;|�H;��H;��H;ժH;9�H;KrH;�SH;�7H;� H;H;      ��H;5�H;��H;Z�H;Q�H;��H;L�H;��H;(�H;2�H;&�H;��H;�H;#�H;��H;X�H;��H;��H;��H;��H;��H;b�H;��H;��H;i�H;��H;��H;W�H;�H;��H;u�H;F�H;!�H;��H;��H;��H;��H;��H;��H;��H;!�H;F�H;u�H;��H;�H;W�H;��H;��H;i�H;��H;��H;b�H;��H;��H;��H;��H;��H;X�H;��H;#�H;�H;��H;&�H;2�H;(�H;��H;L�H;��H;Q�H;Z�H;��H;5�H;      ��H;U�H;7�H;��H;��H;i�H;��H;��H;��H;��H;��H;��H;A�H;��H;��H;!�H;9�H;�H;��H;��H;[�H;��H;��H;e�H; �H;��H;H�H;�H;��H;k�H;7�H;��H;��H;��H;��H;��H;�H;��H;��H;��H;��H;��H;7�H;k�H;��H;�H;H�H;��H; �H;e�H;��H;��H;[�H;��H;��H;�H;9�H;!�H;��H;��H;A�H;��H;��H;��H;��H;��H;��H;i�H;��H;��H;7�H;U�H;      ��H;	�H;�H;w�H;��H;e�H;�H;��H;#�H;��H;��H;!�H;T�H;y�H;k�H;d�H;F�H;�H;��H;z�H;�H;��H;��H;	�H;��H;a�H;�H;��H;k�H;-�H;��H;��H;��H;��H;d�H;K�H;A�H;K�H;d�H;��H;��H;��H;��H;-�H;k�H;��H;�H;a�H;��H;	�H;��H;��H;�H;z�H;��H;�H;F�H;d�H;k�H;y�H;T�H;!�H;��H;��H;#�H;��H;�H;e�H;��H;w�H;�H;	�H;      L�H;p�H;��H;��H;��H;'�H;I�H;w�H;��H;��H;��H;��H;��H;��H;��H;��H;8�H;��H;��H;5�H;��H;��H;�H;��H;r�H;�H;��H;u�H;7�H;��H;��H;��H;w�H;?�H;�H;'�H;(�H;'�H;�H;?�H;w�H;��H;��H;��H;7�H;u�H;��H;�H;r�H;��H;�H;��H;��H;5�H;��H;��H;8�H;��H;��H;��H;��H;��H;��H;��H;��H;w�H;I�H;'�H;��H;��H;��H;p�H;      >�H;B�H;F�H;>�H;V�H;u�H;l�H;��H;��H;v�H;n�H;T�H;%�H;��H;��H;b�H;�H;��H;u�H;�H;��H;B�H;��H;��H;@�H;��H;��H;F�H;��H;��H;��H;_�H;A�H;�H;��H;��H;��H;��H;��H;�H;A�H;_�H;��H;��H;��H;F�H;��H;��H;@�H;��H;��H;B�H;��H;�H;u�H;��H;�H;b�H;��H;��H;%�H;T�H;n�H;v�H;��H;��H;l�H;u�H;V�H;>�H;F�H;B�H;      C�H;6�H;:�H;:�H;3�H;)�H;$�H;�H;��H;��H;��H;n�H;/�H;��H;��H;5�H;��H;��H;P�H;��H;m�H;�H;��H;Y�H;�H;��H;b�H;!�H;��H;��H;w�H;A�H;��H;��H;��H;��H;��H;��H;��H;��H;��H;A�H;w�H;��H;��H;!�H;b�H;��H;�H;Y�H;��H;�H;m�H;��H;P�H;��H;��H;5�H;��H;��H;/�H;n�H;��H;��H;��H;�H;$�H;)�H;3�H;:�H;:�H;6�H;      ��H;��H;��H;��H;��H;h�H;c�H;0�H;�H;��H;��H;Y�H;�H;��H;��H;O�H;��H;]�H;��H;��H;[�H;�H;��H;(�H;��H;��H;D�H;��H;��H;��H;?�H;�H;��H;��H;��H;��H;��H;��H;��H;��H;��H;�H;?�H;��H;��H;��H;D�H;��H;��H;(�H;��H;�H;[�H;��H;��H;]�H;��H;O�H;��H;��H;�H;Y�H;��H;��H;�H;0�H;c�H;h�H;��H;��H;��H;��H;      ��H;��H;��H;��H;��H;��H;s�H;C�H;�H;��H;��H;T�H;�H;��H;h�H;	�H;��H;O�H;��H;��H;*�H;��H;}�H;"�H;��H;o�H;(�H;��H;��H;d�H;�H;��H;��H;��H;��H;��H;��H;��H;��H;��H;��H;��H;�H;d�H;��H;��H;(�H;o�H;��H;"�H;}�H;��H;*�H;��H;��H;O�H;��H;	�H;h�H;��H;�H;T�H;��H;��H;�H;C�H;s�H;��H;��H;��H;��H;��H;      ��H;��H;��H;��H;��H;|�H;X�H;<�H;�H;��H;��H;a�H;�H;��H;K�H;��H;��H;K�H;��H;��H;�H;��H;e�H;�H;��H;\�H;�H;��H;��H;K�H;'�H;��H;��H;��H;��H;��H;��H;��H;��H;��H;��H;��H;'�H;K�H;��H;��H;�H;\�H;��H;�H;e�H;��H;�H;��H;��H;K�H;��H;��H;K�H;��H;�H;a�H;��H;��H;�H;<�H;X�H;|�H;��H;��H;��H;��H;      +�H;$�H;�H;��H;��H;��H;��H;Y�H;$�H;��H;z�H;7�H;��H;��H;m�H;�H;��H;'�H;��H;u�H;�H;��H;L�H;��H;��H;n�H;�H;��H;�H;A�H;(�H;��H;��H;��H;��H;��H;~�H;��H;��H;��H;��H;��H;(�H;A�H;�H;��H;�H;n�H;��H;��H;L�H;��H;�H;u�H;��H;'�H;��H;�H;m�H;��H;��H;7�H;z�H;��H;$�H;Y�H;��H;��H;��H;��H;�H;$�H;      ��H;��H;��H;��H;��H;|�H;X�H;<�H;�H;��H;��H;a�H;�H;��H;K�H;��H;��H;K�H;��H;��H;�H;��H;e�H;�H;��H;\�H;�H;��H;��H;K�H;'�H;��H;��H;��H;��H;��H;��H;��H;��H;��H;��H;��H;'�H;K�H;��H;��H;�H;\�H;��H;�H;e�H;��H;�H;��H;��H;K�H;��H;��H;K�H;��H;�H;a�H;��H;��H;�H;<�H;X�H;|�H;��H;��H;��H;��H;      ��H;��H;��H;��H;��H;��H;s�H;C�H;�H;��H;��H;T�H;�H;��H;h�H;	�H;��H;O�H;��H;��H;*�H;��H;}�H;"�H;��H;o�H;(�H;��H;��H;d�H;�H;��H;��H;��H;��H;��H;��H;��H;��H;��H;��H;��H;�H;d�H;��H;��H;(�H;o�H;��H;"�H;}�H;��H;*�H;��H;��H;O�H;��H;	�H;h�H;��H;�H;T�H;��H;��H;�H;C�H;s�H;��H;��H;��H;��H;��H;      ��H;��H;��H;��H;��H;h�H;c�H;0�H;�H;��H;��H;Y�H;�H;��H;��H;O�H;��H;]�H;��H;��H;[�H;�H;��H;(�H;��H;��H;D�H;��H;��H;��H;?�H;�H;��H;��H;��H;��H;��H;��H;��H;��H;��H;�H;?�H;��H;��H;��H;D�H;��H;��H;(�H;��H;�H;[�H;��H;��H;]�H;��H;O�H;��H;��H;�H;Y�H;��H;��H;�H;0�H;c�H;h�H;��H;��H;��H;��H;      C�H;6�H;:�H;:�H;3�H;)�H;$�H;�H;��H;��H;��H;n�H;/�H;��H;��H;5�H;��H;��H;P�H;��H;m�H;�H;��H;Y�H;�H;��H;b�H;!�H;��H;��H;w�H;A�H;��H;��H;��H;��H;��H;��H;��H;��H;��H;A�H;w�H;��H;��H;!�H;b�H;��H;�H;Y�H;��H;�H;m�H;��H;P�H;��H;��H;5�H;��H;��H;/�H;n�H;��H;��H;��H;�H;$�H;)�H;3�H;:�H;:�H;6�H;      >�H;B�H;F�H;>�H;V�H;u�H;l�H;��H;��H;v�H;n�H;T�H;%�H;��H;��H;b�H;�H;��H;u�H;�H;��H;B�H;��H;��H;@�H;��H;��H;F�H;��H;��H;��H;_�H;A�H;�H;��H;��H;��H;��H;��H;�H;A�H;_�H;��H;��H;��H;F�H;��H;��H;@�H;��H;��H;B�H;��H;�H;u�H;��H;�H;b�H;��H;��H;%�H;T�H;n�H;v�H;��H;��H;l�H;u�H;V�H;>�H;F�H;B�H;      L�H;p�H;��H;��H;��H;'�H;I�H;w�H;��H;��H;��H;��H;��H;��H;��H;��H;8�H;��H;��H;5�H;��H;��H;�H;��H;r�H;�H;��H;u�H;7�H;��H;��H;��H;w�H;?�H;�H;'�H;(�H;'�H;�H;?�H;w�H;��H;��H;��H;7�H;u�H;��H;�H;r�H;��H;�H;��H;��H;5�H;��H;��H;8�H;��H;��H;��H;��H;��H;��H;��H;��H;w�H;I�H;'�H;��H;��H;��H;p�H;      ��H;	�H;�H;w�H;��H;e�H;�H;��H;#�H;��H;��H;!�H;T�H;y�H;k�H;d�H;F�H;�H;��H;z�H;�H;��H;��H;	�H;��H;a�H;�H;��H;k�H;-�H;��H;��H;��H;��H;d�H;K�H;A�H;K�H;d�H;��H;��H;��H;��H;-�H;k�H;��H;�H;a�H;��H;	�H;��H;��H;�H;z�H;��H;�H;F�H;d�H;k�H;y�H;T�H;!�H;��H;��H;#�H;��H;�H;e�H;��H;w�H;�H;	�H;      ��H;U�H;7�H;��H;��H;i�H;��H;��H;��H;��H;��H;��H;A�H;��H;��H;!�H;9�H;�H;��H;��H;[�H;��H;��H;e�H; �H;��H;H�H;�H;��H;k�H;7�H;��H;��H;��H;��H;��H;�H;��H;��H;��H;��H;��H;7�H;k�H;��H;�H;H�H;��H; �H;e�H;��H;��H;[�H;��H;��H;�H;9�H;!�H;��H;��H;A�H;��H;��H;��H;��H;��H;��H;i�H;��H;��H;7�H;U�H;      ��H;5�H;��H;Z�H;Q�H;��H;L�H;��H;(�H;2�H;&�H;��H;�H;#�H;��H;X�H;��H;��H;��H;��H;��H;b�H;��H;��H;i�H;��H;��H;W�H;�H;��H;u�H;F�H;!�H;��H;��H;��H;��H;��H;��H;��H;!�H;F�H;u�H;��H;�H;W�H;��H;��H;i�H;��H;��H;b�H;��H;��H;��H;��H;��H;X�H;��H;#�H;�H;��H;&�H;2�H;(�H;��H;L�H;��H;Q�H;Z�H;��H;5�H;      �H;H;� H;�7H;�SH;KrH;9�H;ժH;��H;��H;|�H;��H;�H;�H;��H;��H;��H;=�H;��H;��H;��H;��H;5�H;��H;��H;_�H;��H;��H;H�H;�H;��H;��H;b�H;D�H;(�H;�H;�H;�H;(�H;D�H;b�H;��H;��H;�H;H�H;��H;��H;_�H;��H;��H;5�H;��H;��H;��H;��H;=�H;��H;��H;��H;�H;�H;��H;|�H;��H;��H;ժH;9�H;KrH;�SH;�7H;� H;H;      nCF;{QF;�yF;�F;�G;�[G;�G;YH;#HH;��H;��H;��H;�H;��H;��H;9�H;��H;7�H;��H;P�H;��H;�H;r�H;D�H;��H;��H;_�H;��H;��H;a�H;�H;��H;��H;��H;o�H;\�H;n�H;\�H;o�H;��H;��H;��H;�H;a�H;��H;��H;_�H;��H;��H;D�H;r�H;�H;��H;P�H;��H;7�H;��H;9�H;��H;��H;�H;��H;��H;��H;#HH;YH;�G;�[G;�G;�F;�yF;{QF;      ��A;B;2oB;�C;��C;|�D;otE;�CF;N�F;��G;�H;eH;�H;��H;[�H;�H;��H;�H;��H;��H;#�H;f�H;��H;j�H;-�H;��H;��H;i�H; �H;��H;r�H;@�H;�H;��H;��H;��H;��H;��H;��H;��H;�H;@�H;r�H;��H; �H;i�H;��H;��H;-�H;j�H;��H;f�H;#�H;��H;��H;�H;��H;�H;[�H;��H;�H;eH;�H;��G;N�F;�CF;otE;|�D;��C;�C;2oB;B;      ~n8;M�8;؎9;��:;��<;
c>;ZQ@;�.B;��C;�OE;�yF;j[G;��G;DhH;8�H;��H;8�H;a�H;-�H;5�H;\�H;��H;b�H;k�H;j�H;D�H;��H;��H;e�H;	�H;��H;��H;Y�H;(�H;"�H;�H;��H;�H;"�H;(�H;Y�H;��H;��H;	�H;e�H;��H;��H;D�H;j�H;k�H;b�H;��H;\�H;5�H;-�H;a�H;8�H;��H;8�H;DhH;��G;j[G;�yF;�OE;��C;�.B;ZQ@;
c>;��<;��:;؎9;M�8;      �R%;i�%;_�';M*;5�-;ʕ1;�5;6�9;�,=;IQ@;�B;��D;9lF;�tG;� H;�H;��H;��H;�H;��H;��H;1�H;�H;b�H;��H;r�H;5�H;��H;��H;��H;�H;��H;��H;��H;}�H;e�H;L�H;e�H;}�H;��H;��H;��H;�H;��H;��H;��H;5�H;r�H;��H;b�H;�H;1�H;��H;��H;�H;��H;��H;�H;� H;�tG;9lF;��D;�B;IQ@;�,=;6�9;�5;ʕ1;5�-;M*;_�';i�%;      �V;�w;1�;Q�
;�;�;)� ;��(;��/;$H6;��;;�?;!C;�OE;�F;�G;�dH;N�H;��H;&�H;P�H;��H;1�H;��H;f�H;�H;��H;b�H;��H;��H;��H;B�H;�H;�H;��H;��H;��H;��H;��H;�H;�H;B�H;��H;��H;��H;b�H;��H;�H;f�H;��H;1�H;��H;P�H;&�H;��H;N�H;�dH;�G;�F;�OE;!C;�?;��;;$H6;��/;��(;)� ;�;�;Q�
;1�;�w;      �:nĆ:pȒ:���:r�:o��:���:��	;v;7�#;��-;#�5;�K<;��@;�'D;3CF;��G;�GH;s�H;�H;��H;P�H;��H;\�H;#�H;��H;��H;��H;[�H;�H;��H;��H;m�H;[�H;*�H;�H;�H;�H;*�H;[�H;m�H;��H;��H;�H;[�H;��H;��H;��H;#�H;\�H;��H;P�H;��H;�H;s�H;�GH;��G;3CF;�'D;��@;�K<;#�5;��-;7�#;v;��	;���:o��:r�:���:pȒ:nĆ:      0.�5��+�깙�K�
9�Z:��k:L�:6��:�x;��;�$;�/;��8;��>;#C;7�E;�[G;]7H;ͤH;�H;&�H;��H;5�H;��H;P�H;��H;��H;��H;z�H;5�H;�H;��H;��H;��H;��H;u�H;��H;��H;��H;��H;�H;5�H;z�H;��H;��H;��H;P�H;��H;5�H;��H;&�H;�H;ͤH;]7H;�[G;7�E;#C;��>;��8;�/;�$;��;�x;6��:L�:��k:�Z:
9��K�+��5��      �Q^��X�UF�\�)��+�+ж���<�jS��k:���:J��:�;}�;M*;	�5;�b=;�oB;��E;�IG;]7H;s�H;��H;�H;-�H;��H;��H;��H;��H;��H;��H;��H;u�H;P�H;��H;��H;��H;��H;��H;��H;��H;P�H;u�H;��H;��H;��H;��H;��H;��H;��H;-�H;�H;��H;s�H;]7H;�IG;��E;�oB;�b=;	�5;M*;}�;�;J��:���:�k:jS���<�+ж��+�\�)�UF��X�      ����o���W��O�ѻf���[ǐ��X��6��
���K�><":gL�:�`�:�h;Z�%;��3;�<;Y/B;��E;�[G;�GH;N�H;��H;a�H;�H;7�H;=�H;��H;�H;�H;��H;��H;��H;]�H;O�H;K�H;'�H;K�H;O�H;]�H;��H;��H;��H;�H;�H;��H;=�H;7�H;�H;a�H;��H;N�H;�GH;�[G;��E;Y/B;�<;��3;Z�%;�h;�`�:gL�:><":�K��
���6��X�[ǐ�f���O�ѻW��o���      ��n��mj���]���J�n�1�L4�k��R���U
x�hX���y�0
9���:ף�:@�;v�#;w�2;�<;�oB;7�E;��G;�dH;��H;8�H;��H;��H;��H;��H;9�H;F�H;8�H;�H;��H;��H;��H;��H;��H;��H;��H;��H;��H;�H;8�H;F�H;9�H;��H;��H;��H;��H;8�H;��H;�dH;��G;7�E;�oB;�<;w�2;v�#;@�;ף�:���:0
9��y�hX�U
x�R���k��L4�n�1���J���]��mj�      B<ͼ��ɼ�����֯�Ҷ��ㄼ��Y�-�*�I���t���X��sѺ�(�N<Q:]��:��
;v�#;��3;�b=;#C;3CF;�G;�H;��H;�H;9�H;��H;X�H;!�H;d�H;��H;b�H;5�H;O�H;	�H;��H;�H;��H;	�H;O�H;5�H;b�H;��H;d�H;!�H;X�H;��H;9�H;�H;��H;�H;�G;3CF;#C;�b=;��3;v�#;��
;]��:N<Q:�(��sѺ�X�t��I���-�*���Y�ㄼҶ���֯�������ɼ      ��'�#�$����y��  ���ۼ����+����]��X!�>ۻ�+��+�c���>:]��:@�;Z�%;	�5;��>;�'D;�F;� H;8�H;[�H;��H;��H;��H;��H;k�H;��H;��H;��H;��H;h�H;K�H;m�H;K�H;h�H;��H;��H;��H;��H;k�H;��H;��H;��H;��H;[�H;8�H;� H;�F;�'D;��>;	�5;Z�%;@�;]��:�>:c��+��+��>ۻ�X!���]��+�������ۼ�  �y����#�$�      �����v����w�]�c��J�Ȅ-�x��;缈沼ㄼ��;�����k��56�c��N<Q:ף�:�h;M*;��8;��@;�OE;�tG;DhH;��H;��H;�H;#�H;��H;y�H;��H;��H;��H;��H;��H;��H;��H;��H;��H;��H;��H;��H;��H;y�H;��H;#�H;�H;��H;��H;DhH;�tG;�OE;��@;��8;M*;�h;ף�:N<Q:c��56�k��������;�ㄼ�沼�;�x�Ȅ-��J�]�c���w��v��      nHͽ̪ɽ�;��"����������[�z0�p��'<ͼо��u�J���k��+��(����:�`�:}�;�/;�K<;!C;9lF;��G;�H;�H;�H;�H;A�H;T�H;��H;%�H;/�H;�H;�H;�H;��H;�H;�H;�H;/�H;%�H;��H;T�H;A�H;�H;�H;�H;�H;��G;9lF;!C;�K<;�/;}�;�`�:���:�(�+�k����u�J�о��'<ͼp��z0���[�������"���;��̪ɽ      ��-�}��|�ű�ƽUP���v���J�D����ۼ��u�J������+���sѺ0
9gL�:�;�$;#�5;�?;��D;j[G;eH;��H;��H;��H;��H;!�H;��H;T�H;n�H;Y�H;T�H;a�H;7�H;a�H;T�H;Y�H;n�H;T�H;��H;!�H;��H;��H;��H;��H;eH;j[G;��D;�?;#�5;�$;�;gL�:0
9�sѺ�+������u�J�����ۼD���J��v��UP��ƽű�|�}��-�       j�Ide�M0X�sD�\{+�z�����k㻽R���IDX������ۼо����;�>ۻ�X���y�><":J��:��;��-;��;;�B;�yF;�H;��H;|�H;&�H;��H;��H;��H;n�H;��H;��H;��H;��H;z�H;��H;��H;��H;��H;n�H;��H;��H;��H;&�H;|�H;��H;�H;�yF;�B;��;;��-;��;J��:><":��y��X�>ۻ��;�о����ۼ���IDX�R���k㻽���z��\{+�sD�M0X�Ide�      ��Fh��b���I���|x���O��C(�y�Īɽ����IDX�D��'<ͼㄼ�X!�t��hX��K����:�x;7�#;$H6;IQ@;�OE;��G;��H;��H;2�H;��H;��H;��H;v�H;��H;��H;��H;��H;��H;��H;��H;��H;��H;v�H;��H;��H;��H;2�H;��H;��H;��G;�OE;IQ@;$H6;7�#;�x;���:�K�hX�t���X!�ㄼ'<ͼD��IDX�����Īɽy��C(���O��|x��I��b��Fh��      /�����������;^ɰ��G����i�.�5��	�ĪɽR����J�p���沼��]�I���U
x��
���k:6��:v;��/;�,=;��C;N�F;#HH;��H;(�H;��H;#�H;��H;��H;��H;�H;�H;�H;$�H;�H;�H;�H;��H;��H;��H;#�H;��H;(�H;��H;#HH;N�F;��C;�,=;��/;v;6��:�k:�
��U
x�I�����]��沼p���J�R���Īɽ�	�.�5���i��G��^ɰ��;��徨���      �2�L�-��"�$E�����4Kɾa��w�s�.�5�y�k㻽�v��z0��;��+��-�*�R����6�jS�L�:��	;��(;6�9;�.B;�CF;YH;ժH;��H;��H;��H;w�H;��H;�H;0�H;C�H;<�H;Y�H;<�H;C�H;0�H;�H;��H;w�H;��H;��H;��H;ժH;YH;�CF;�.B;6�9;��(;��	;L�:jS��6�R���-�*��+���;�z0��v��k㻽y�.�5�w�s�a��4Kɾ����$E��"�L�-�      3s�cm�/�\�]�C�,�%����TҾa����i��C(����UP����[�x������Y�k���X���<���k:���:)� ;�5;ZQ@;otE;�G;9�H;L�H;��H;�H;I�H;l�H;$�H;c�H;s�H;X�H;��H;X�H;s�H;c�H;$�H;l�H;I�H;�H;��H;L�H;9�H;�G;otE;ZQ@;�5;)� ;���:��k:��<��X�k����Y����x���[�UP����콡C(���i�a���TҾ��,�%�]�C�/�\�cm�      �ޞ�������RF�3�W�M�-���4Kɾ�G����O�z��ƽ����Ȅ-���ۼㄼL4�[ǐ�+ж��Z:o��:�;ʕ1;
c>;|�D;�[G;KrH;��H;i�H;e�H;'�H;u�H;)�H;h�H;��H;|�H;��H;|�H;��H;h�H;)�H;u�H;'�H;e�H;i�H;��H;KrH;�[G;|�D;
c>;ʕ1;�;o��:�Z:+ж�[ǐ�L4�ㄼ��ۼȄ-�����ƽz����O��G��4Kɾ��M�-�3�W�RF�������      ��ſ~��Bw���ޞ�|���3�W�,�%�����^ɰ��|x�\{+�ű����J��  �Ҷ��n�1�f����+�
9r�:�;5�-;��<;��C;�G;�SH;Q�H;��H;��H;��H;V�H;3�H;��H;��H;��H;��H;��H;��H;��H;3�H;V�H;��H;��H;��H;Q�H;�SH;�G;��C;��<;5�-;�;r�:
9�+�f���n�1�Ҷ���  ��J���ű�\{+��|x�^ɰ�����,�%�3�W�|����ޞ�Bw��~��      ������Կp���ޞ�RF�]�C�$E��;�I��sD�|�"��]�c�y��֯���J�O�ѻ\�)���K����:Q�
;M*;��:;�C;�F;�7H;Z�H;��H;w�H;��H;>�H;:�H;��H;��H;��H;��H;��H;��H;��H;:�H;>�H;��H;w�H;��H;Z�H;�7H;�F;�C;��:;M*;Q�
;���:��K�\�)�O�ѻ��J��֯�y�]�c�"��|�sD��I���;$E�]�C�RF��ޞ�p���Կ��      ������{���ԿBw�����/�\��"����b��M0X�}���;����w����������]�W��UF�+��pȒ:1�;_�';؎9;2oB;�yF;� H;��H;7�H;�H;��H;F�H;:�H;��H;��H;��H;�H;��H;��H;��H;:�H;F�H;��H;�H;7�H;��H;� H;�yF;2oB;؎9;_�';1�;pȒ:+��UF�W�黼�]����������w��;��}��M0X�b������"�/�\����Bw���Կ{�𿖏�      $��������~�����cm�L�-�����Fh��Ide�-�̪ɽ�v��#�$���ɼ�mj�o����X�5��nĆ:�w;i�%;M�8;B;{QF;H;5�H;U�H;	�H;p�H;B�H;6�H;��H;��H;��H;$�H;��H;��H;��H;6�H;B�H;p�H;	�H;U�H;5�H;H;{QF;B;M�8;i�%;�w;nĆ:5���X�o����mj���ɼ#�$��v��̪ɽ-�Ide�Fh������L�-�cm����~���忖����      Vܿ%�ֿ�aǿ2^��&���Io���7����iþ�(���-=��` ��@����_�&]�&p����I�q�ѻ��)��R�\�:��
;*;D�:;�B;UHF;=�G;�kH;3�H;��H;i�H;��H;��H;p�H;��H;(�H;��H;(�H;��H;p�H;��H;��H;i�H;��H;3�H;�kH;=�G;UHF;�B;D�:;*;��
;\�:�R���)�q�ѻ��I�&p��&]���_��@���` ��-=��(���iþ����7�Io�&���2^���aǿ%�ֿ      %�ֿ5pѿ֊¿������PXi�Õ3��
�GD��;l��1�9�j.���R��\� �\x��1�E��ͻ��$�� ����:��;��*;\�:;.�B;3TF;��G;[mH;ϠH;ݶH;��H;��H;��H;�H;��H;<�H;��H;<�H;��H;�H;��H;��H;��H;ݶH;ϠH;[mH;��G;3TF;.�B;\�:;��*;��;���:� ���$��ͻ1�E�\x�� �\��R��j.��1�9�;l��GD���
�Õ3�PXi�������֊¿5pѿ      �aǿ֊¿���������s"Y��f'�����)o���.}��k/�m��ڟ�<Q�%#�ע��(;�P��������7���:J�;�,;��;;�C;RvF;/�G;�qH;[�H;��H;=�H;�H;�H;��H;��H;j�H;��H;j�H;��H;��H;�H;�H;=�H;��H;[�H;�qH;/�G;RvF;�C;��;;�,;J�;��:��7����P����(;�ע�%#�<Q�ڟ�m���k/��.}�)o�������f'�s"Y����������֊¿      2^������b���Io���@���޾����&ce�"����ڽ绒��f@������R���O*�mG������<^9Ӳ�:[;�c.;'�<;ՏC;G�F;��G;�xH;ĤH;8�H;I�H;��H;��H;��H;�H;��H;6�H;��H;�H;��H;��H;��H;I�H;8�H;ĤH;�xH;��G;G�F;ՏC;'�<;�c.;[;Ӳ�:�<^9���mG���O*��R�������f@�绒���ڽ"��&ce������޾���@�Io�b�������      &����������Io��!J�@�#��\��GD������jPH�����b��C��t +�u�ټ%��������������:���:��;�X1;3>;�/D;��F;�H;r�H;��H;)�H;��H;��H;)�H;��H;p�H;��H;�H;��H;p�H;��H;)�H;��H;��H;)�H;��H;r�H;�H;��F;�/D;3>;�X1;��;���:��:����������%��u�ټt +�C���b�����jPH�����GD���\��@�#��!J�Io��������      Io�PXi�s"Y���@�@�#��
��о�A�� �i���(�i��gr����_��5��ɺ�n�`��<����d�=�\�P�X:PO�:7`;#�4;�?;��D;�7G;�/H;ȊH;��H;��H;.�H;��H;��H;�H;��H;-�H;��H;-�H;��H;�H;��H;��H;.�H;��H;��H;ȊH;�/H;�7G;��D;�?;#�4;7`;PO�:P�X:=�\���d��<��n�`��ɺ��5���_�gr��i����(� �i��A���о�
�@�#���@�s"Y�PXi�      ��7�Õ3��f'���\���о�����.}��-=�o
�y�ĽO��:����������7�?GĻ*�$�	S�����:�z;�C&;E+8;FIA;1�E;��G;�KH;�H;��H;S�H;�H;(�H;��H;��H;@�H;��H;5�H;��H;@�H;��H;��H;(�H;�H;S�H;��H;�H;�KH;��G;1�E;FIA;E+8;�C&;�z;���:	S��*�$�?GĻ�7���������:�O��y�Ľo
��-=��.}������о�\����f'�Õ3�      ���
������޾GD���A���.}��D�[t���ڽ�!��\����P�ļ�
v�F�����Jɺ�N�9���:i';�-;ӊ;;��B;�HF;��G;?eH;ʜH;�H;N�H;��H;��H;��H;{�H;��H;�H;��H;�H;��H;{�H;��H;��H;��H;N�H;�H;ʜH;?eH;��G;�HF;��B;ӊ;;�-;i';���:�N�9�Jɺ��F���
v�P�ļ���\��!����ڽ[t��D��.}��A��GD���޾�����
�      �iþGD��)o���������� �i��-=�[t����R��Tys�m +����s񗼗(;�G�ѻt@�͇!��1j:�O�:4�;�C3;~�>;DED;��F;�H;_{H;��H;��H;W�H;�H;�H;��H;9�H;R�H;��H;�H;��H;R�H;9�H;��H;�H;�H;W�H;��H;��H;_{H;�H;��F;DED;~�>;�C3;4�;�O�:�1j:͇!�t@�G�ѻ�(;�s����m +�Tys��R����[t��-=� �i���������)o��GD��      �(��;l���.}�&ce�jPH���(�o
���ڽ�R����{�4�6�� �$p��\�`�ר�-��JҺ�C^9a��:=�;�}(;t�8;IA;6{E;GiG;�<H;i�H; �H;H�H;��H;N�H;��H;��H;��H;��H;�H;i�H;�H;��H;��H;��H;��H;N�H;��H;H�H; �H;i�H;�<H;GiG;6{E;IA;t�8;�}(;=�;a��:�C^9JҺ-��ר�\�`�$p��� �4�6���{��R����ڽo
���(�jPH�&ce��.}�;l��      �-=�1�9��k/�"�����i��y�Ľ�!��Tys�4�6�#��ɺ��vz����c^��˃$�{����r:���:7�;�X1;?H=;jwC;WvF;R�G;/eH;m�H;��H;��H;��H;v�H;�H;��H;��H;��H;��H;��H;��H;��H;��H;��H;�H;v�H;��H;��H;��H;m�H;/eH;R�G;WvF;jwC;?H=;�X1;7�;���:��r:{��˃$�c^������vz��ɺ�#�4�6�Tys��!��y�Ľi���"���k/�1�9�      �` �j.��m��ڽ�b��gr��O��\�m +�� ��ɺ�<��O*�bͻP6R��ǅ���:���:ڃ;�);6t8;��@;�)E;�7G;t#H;p�H;d�H;�H;J�H;��H;��H;��H;�H;n�H;�H; �H;?�H; �H;�H;n�H;�H;��H;��H;��H;J�H;�H;d�H;p�H;t#H;�7G;�)E;��@;6t8;�);ڃ;���:��:�ǅ�P6R�bͻ�O*�<��ɺ�� �m +�\�O��gr���b����ڽm��j.��      �@���R��ڟ�绒�C����_�:�������$p���vz��O*�5ֻfk������09�:`0;�� ;�C3;��=;�C;kF;��G;�[H;ÖH;o�H;&�H;b�H;��H;��H;��H;�H;'�H;��H;o�H;��H;o�H;��H;'�H;�H;��H;��H;��H;b�H;&�H;o�H;ÖH;�[H;��G;kF;�C;��=;�C3;�� ;`0;�:��09���fk�5ֻ�O*��vz�$p����輙��:���_�C��绒�ڟ��R��      ��_�\�<Q��f@�t +��5�����P�ļs�\�`����bͻfk��Iɺ�	7��:�O�:y�;%d.;��:;Z�A;c{E;�MG;q&H;/�H;�H;��H;��H;J�H;n�H;|�H;S�H;�H;��H;*�H;��H;�H;��H;*�H;��H;�H;S�H;|�H;n�H;J�H;��H;��H;�H;/�H;q&H;�MG;c{E;Z�A;��:;%d.;y�;�O�:�:�	7��Iɺfk�bͻ���\�`�s�P�ļ�����5�t +��f@�<Q�\�      &]� �%#�����u�ټ�ɺ������
v��(;�ר�c^��P6R�����	7����:���:O�;l�*;+8;� @;��D;��F;'�G; eH;��H;��H;žH;��H;�H;��H;B�H;��H;��H;��H;��H;B�H;u�H;B�H;��H;��H;��H;��H;B�H;��H;�H;��H;žH;��H;��H; eH;'�G;��F;��D;� @;+8;l�*;O�;���:���:�	7����P6R�c^��ר��(;��
v������ɺ�u�ټ����%#� �      &p��\x��ע��R��%��n�`��7�F��G�ѻ-��˃$��ǅ���09�:���:�; ~(;�Y6;��>;�C;&HF;�G;DH;s�H;�H;ϸH;3�H;K�H;2�H;�H;��H;��H;��H;,�H;�H;��H;��H;��H;�H;,�H;��H;��H;��H;�H;2�H;K�H;3�H;ϸH;�H;s�H;DH;�G;&HF;�C;��>;�Y6; ~(;�;���:�:��09�ǅ�˃$�-��G�ѻF���7�n�`�%���R��ע�\x��      ��I�1�E��(;��O*�����<��?GĻ��t@�JҺ{��:�:�O�:O�; ~(;S�5;>;qC;k�E;�bG;k#H;"{H;_�H;I�H;��H;��H;Y�H;��H;;�H;x�H;��H;h�H;��H;Y�H;��H;�H;��H;Y�H;��H;h�H;��H;x�H;;�H;��H;Y�H;��H;��H;I�H;_�H;"{H;k#H;�bG;k�E;qC;>;S�5; ~(;O�;�O�:�:��:{��JҺt@���?GĻ�<������O*��(;�1�E�      q�ѻ�ͻP���mG�������d�*�$��Jɺ͇!��C^9��r:���:`0;y�;l�*;�Y6;>;n�B;��E;8G;�H;,mH;A�H;m�H;μH;��H;��H;��H;h�H;�H;��H;��H;�H;�H;��H;�H;<�H;�H;��H;�H;�H;��H;��H;�H;h�H;��H;��H;��H;μH;m�H;A�H;,mH;�H;8G;��E;n�B;>;�Y6;l�*;y�;`0;���:��r:�C^9͇!��Jɺ*�$���d����mG��P����ͻ      ��)���$�����������=�\�	S���N�9�1j:a��:���:ڃ;�� ;%d.;+8;��>;qC;��E;�(G;��G;>cH;��H;��H;��H;��H;T�H;��H;��H;��H;��H;��H;b�H;��H;w�H;�H;I�H;c�H;I�H;�H;w�H;��H;b�H;��H;��H;��H;��H;��H;T�H;��H;��H;��H;��H;>cH;��G;�(G;��E;qC;��>;+8;%d.;�� ;ڃ;���:a��:�1j:�N�9	S��=�\�������������$�      �R�� ���7��<^9��:P�X:���:���:�O�:=�;7�;�);�C3;��:;� @;�C;k�E;8G;��G;�_H;��H;?�H;@�H;��H;d�H;Q�H;i�H;w�H;��H;��H;��H;$�H; �H;��H;@�H;{�H;{�H;{�H;@�H;��H; �H;$�H;��H;��H;��H;w�H;i�H;Q�H;d�H;��H;@�H;?�H;��H;�_H;��G;8G;k�E;�C;� @;��:;�C3;�);7�;=�;�O�:���:���:P�X:��:�<^9��7�� �      \�:���:��:Ӳ�:���:PO�:�z;i';4�;�}(;�X1;6t8;��=;Z�A;��D;&HF;�bG;�H;>cH;��H;m�H;��H;S�H;�H;��H;Y�H;d�H;��H;<�H;��H;��H;��H;m�H;��H;Y�H;��H;��H;��H;Y�H;��H;m�H;��H;��H;��H;<�H;��H;d�H;Y�H;��H;�H;S�H;��H;m�H;��H;>cH;�H;�bG;&HF;��D;Z�A;��=;6t8;�X1;�}(;4�;i';�z;PO�:���:Ӳ�:��:���:      ��
;��;J�;[;��;7`;�C&;�-;�C3;t�8;?H=;��@;�C;c{E;��F;�G;k#H;,mH;��H;?�H;��H;��H;Y�H;:�H;��H;��H;��H;��H;�H;�H;4�H;�H;��H;1�H;r�H;��H;��H;��H;r�H;1�H;��H;�H;4�H;�H;�H;��H;��H;��H;��H;:�H;Y�H;��H;��H;?�H;��H;,mH;k#H;�G;��F;c{E;�C;��@;?H=;t�8;�C3;�-;�C&;7`;��;[;J�;��;      *;��*;�,;�c.;�X1;#�4;E+8;ӊ;;~�>;IA;jwC;�)E;kF;�MG;'�G;DH;"{H;A�H;��H;@�H;S�H;Y�H;��H;�H;�H;w�H;#�H;�H;��H;��H;��H;��H;��H;L�H;��H;��H;��H;��H;��H;L�H;��H;��H;��H;��H;��H;�H;#�H;w�H;�H;�H;��H;Y�H;S�H;@�H;��H;A�H;"{H;DH;'�G;�MG;kF;�)E;jwC;IA;~�>;ӊ;;E+8;#�4;�X1;�c.;�,;��*;      D�:;\�:;��;;'�<;3>;�?;FIA;��B;DED;6{E;WvF;�7G;��G;q&H; eH;s�H;_�H;m�H;��H;��H;�H;:�H;�H;��H;5�H;��H;��H;G�H;��H;~�H;(�H;��H;,�H;l�H;��H;��H;��H;��H;��H;l�H;,�H;��H;(�H;~�H;��H;G�H;��H;��H;5�H;��H;�H;:�H;�H;��H;��H;m�H;_�H;s�H; eH;q&H;��G;�7G;WvF;6{E;DED;��B;FIA;�?;3>;'�<;��;;\�:;      �B;.�B;�C;ՏC;�/D;��D;1�E;�HF;��F;GiG;R�G;t#H;�[H;/�H;��H;�H;I�H;μH;��H;d�H;��H;��H;�H;5�H;��H;��H;�H;T�H;8�H;�H;��H;��H;=�H;��H;��H;��H;��H;��H;��H;��H;=�H;��H;��H;�H;8�H;T�H;�H;��H;��H;5�H;�H;��H;��H;d�H;��H;μH;I�H;�H;��H;/�H;�[H;t#H;R�G;GiG;��F;�HF;1�E;��D;�/D;ՏC;�C;.�B;      UHF;3TF;RvF;G�F;��F;�7G;��G;��G;�H;�<H;/eH;p�H;ÖH;�H;��H;ϸH;��H;��H;T�H;Q�H;Y�H;��H;w�H;��H;��H;	�H;9�H;�H;��H;R�H;��H;.�H;C�H;}�H;��H;��H;��H;��H;��H;}�H;C�H;.�H;��H;R�H;��H;�H;9�H;	�H;��H;��H;w�H;��H;Y�H;Q�H;T�H;��H;��H;ϸH;��H;�H;ÖH;p�H;/eH;�<H;�H;��G;��G;�7G;��F;G�F;RvF;3TF;      =�G;��G;/�G;��G;�H;�/H;�KH;?eH;_{H;i�H;m�H;d�H;o�H;��H;žH;3�H;��H;��H;��H;i�H;d�H;��H;#�H;��H;�H;9�H;�H;��H;[�H;��H;��H;<�H;\�H;�H;��H;��H;��H;��H;��H;�H;\�H;<�H;��H;��H;[�H;��H;�H;9�H;�H;��H;#�H;��H;d�H;i�H;��H;��H;��H;3�H;žH;��H;o�H;d�H;m�H;i�H;_{H;?eH;�KH;�/H;�H;��G;/�G;��G;      �kH;[mH;�qH;�xH;r�H;ȊH;�H;ʜH;��H; �H;��H;�H;&�H;��H;��H;K�H;Y�H;��H;��H;w�H;��H;��H;�H;G�H;T�H;�H;��H;B�H;��H;��H;�H;B�H;k�H;l�H;��H;��H;��H;��H;��H;l�H;k�H;B�H;�H;��H;��H;B�H;��H;�H;T�H;G�H;�H;��H;��H;w�H;��H;��H;Y�H;K�H;��H;��H;&�H;�H;��H; �H;��H;ʜH;�H;ȊH;r�H;�xH;�qH;[mH;      3�H;ϠH;[�H;ĤH;��H;��H;��H;�H;��H;H�H;��H;J�H;b�H;J�H;�H;2�H;��H;h�H;��H;��H;<�H;�H;��H;��H;8�H;��H;[�H;��H;��H;�H;6�H;S�H;j�H;l�H;j�H;u�H;u�H;u�H;j�H;l�H;j�H;S�H;6�H;�H;��H;��H;[�H;��H;8�H;��H;��H;�H;<�H;��H;��H;h�H;��H;2�H;�H;J�H;b�H;J�H;��H;H�H;��H;�H;��H;��H;��H;ĤH;[�H;ϠH;      ��H;ݶH;��H;8�H;)�H;��H;S�H;N�H;W�H;��H;��H;��H;��H;n�H;��H;�H;;�H;�H;��H;��H;��H;�H;��H;~�H;�H;R�H;��H;��H;�H;+�H;J�H;I�H;X�H;h�H;P�H;b�H;{�H;b�H;P�H;h�H;X�H;I�H;J�H;+�H;�H;��H;��H;R�H;�H;~�H;��H;�H;��H;��H;��H;�H;;�H;�H;��H;n�H;��H;��H;��H;��H;W�H;N�H;S�H;��H;)�H;8�H;��H;ݶH;      i�H;��H;=�H;I�H;��H;.�H;�H;��H;�H;N�H;v�H;��H;��H;|�H;B�H;��H;x�H;��H;��H;��H;��H;4�H;��H;(�H;��H;��H;��H;�H;6�H;J�H;a�H;T�H;E�H;E�H;c�H;U�H;6�H;U�H;c�H;E�H;E�H;T�H;a�H;J�H;6�H;�H;��H;��H;��H;(�H;��H;4�H;��H;��H;��H;��H;x�H;��H;B�H;|�H;��H;��H;v�H;N�H;�H;��H;�H;.�H;��H;I�H;=�H;��H;      ��H;��H;�H;��H;��H;��H;(�H;��H;�H;��H;�H;��H;��H;S�H;��H;��H;��H;��H;b�H;$�H;��H;�H;��H;��H;��H;.�H;<�H;B�H;S�H;I�H;T�H;Z�H;C�H;=�H;O�H;4�H;+�H;4�H;O�H;=�H;C�H;Z�H;T�H;I�H;S�H;B�H;<�H;.�H;��H;��H;��H;�H;��H;$�H;b�H;��H;��H;��H;��H;S�H;��H;��H;�H;��H;�H;��H;(�H;��H;��H;��H;�H;��H;      ��H;��H;�H;��H;)�H;��H;��H;��H;��H;��H;��H;�H;�H;�H;��H;��H;h�H;�H;��H; �H;m�H;��H;��H;,�H;=�H;C�H;\�H;k�H;j�H;X�H;E�H;C�H;G�H;C�H;#�H;#�H;S�H;#�H;#�H;C�H;G�H;C�H;E�H;X�H;j�H;k�H;\�H;C�H;=�H;,�H;��H;��H;m�H; �H;��H;�H;h�H;��H;��H;�H;�H;�H;��H;��H;��H;��H;��H;��H;)�H;��H;�H;��H;      p�H;�H;��H;��H;��H;�H;��H;{�H;9�H;��H;��H;n�H;'�H;��H;��H;,�H;��H;�H;w�H;��H;��H;1�H;L�H;l�H;��H;}�H;�H;l�H;l�H;h�H;E�H;=�H;C�H;-�H;�H;$�H;)�H;$�H;�H;-�H;C�H;=�H;E�H;h�H;l�H;l�H;�H;}�H;��H;l�H;L�H;1�H;��H;��H;w�H;�H;��H;,�H;��H;��H;'�H;n�H;��H;��H;9�H;{�H;��H;�H;��H;��H;��H;�H;      ��H;��H;��H;�H;p�H;��H;@�H;��H;R�H;��H;��H;�H;��H;*�H;��H;�H;Y�H;��H;�H;@�H;Y�H;r�H;��H;��H;��H;��H;��H;��H;j�H;P�H;c�H;O�H;#�H;�H;'�H;�H;�H;�H;'�H;�H;#�H;O�H;c�H;P�H;j�H;��H;��H;��H;��H;��H;��H;r�H;Y�H;@�H;�H;��H;Y�H;�H;��H;*�H;��H;�H;��H;��H;R�H;��H;@�H;��H;p�H;�H;��H;��H;      (�H;<�H;j�H;��H;��H;-�H;��H;�H;��H;�H;��H; �H;o�H;��H;B�H;��H;��H;�H;I�H;{�H;��H;��H;��H;��H;��H;��H;��H;��H;u�H;b�H;U�H;4�H;#�H;$�H;�H;�H;�H;�H;�H;$�H;#�H;4�H;U�H;b�H;u�H;��H;��H;��H;��H;��H;��H;��H;��H;{�H;I�H;�H;��H;��H;B�H;��H;o�H; �H;��H;�H;��H;�H;��H;-�H;��H;��H;j�H;<�H;      ��H;��H;��H;6�H;�H;��H;5�H;��H;�H;i�H;��H;?�H;��H;�H;u�H;��H;�H;<�H;c�H;{�H;��H;��H;��H;��H;��H;��H;��H;��H;u�H;{�H;6�H;+�H;S�H;)�H;�H;�H;�H;�H;�H;)�H;S�H;+�H;6�H;{�H;u�H;��H;��H;��H;��H;��H;��H;��H;��H;{�H;c�H;<�H;�H;��H;u�H;�H;��H;?�H;��H;i�H;�H;��H;5�H;��H;�H;6�H;��H;��H;      (�H;<�H;j�H;��H;��H;-�H;��H;�H;��H;�H;��H; �H;o�H;��H;B�H;��H;��H;�H;I�H;{�H;��H;��H;��H;��H;��H;��H;��H;��H;u�H;b�H;U�H;4�H;#�H;$�H;�H;�H;�H;�H;�H;$�H;#�H;4�H;U�H;b�H;u�H;��H;��H;��H;��H;��H;��H;��H;��H;{�H;I�H;�H;��H;��H;B�H;��H;o�H; �H;��H;�H;��H;�H;��H;-�H;��H;��H;j�H;<�H;      ��H;��H;��H;�H;p�H;��H;@�H;��H;R�H;��H;��H;�H;��H;*�H;��H;�H;Y�H;��H;�H;@�H;Y�H;r�H;��H;��H;��H;��H;��H;��H;j�H;P�H;c�H;O�H;#�H;�H;'�H;�H;�H;�H;'�H;�H;#�H;O�H;c�H;P�H;j�H;��H;��H;��H;��H;��H;��H;r�H;Y�H;@�H;�H;��H;Y�H;�H;��H;*�H;��H;�H;��H;��H;R�H;��H;@�H;��H;p�H;�H;��H;��H;      p�H;�H;��H;��H;��H;�H;��H;{�H;9�H;��H;��H;n�H;'�H;��H;��H;,�H;��H;�H;w�H;��H;��H;1�H;L�H;l�H;��H;}�H;�H;l�H;l�H;h�H;E�H;=�H;C�H;-�H;�H;$�H;)�H;$�H;�H;-�H;C�H;=�H;E�H;h�H;l�H;l�H;�H;}�H;��H;l�H;L�H;1�H;��H;��H;w�H;�H;��H;,�H;��H;��H;'�H;n�H;��H;��H;9�H;{�H;��H;�H;��H;��H;��H;�H;      ��H;��H;�H;��H;)�H;��H;��H;��H;��H;��H;��H;�H;�H;�H;��H;��H;h�H;�H;��H; �H;m�H;��H;��H;,�H;=�H;C�H;\�H;k�H;j�H;X�H;E�H;C�H;G�H;C�H;#�H;#�H;S�H;#�H;#�H;C�H;G�H;C�H;E�H;X�H;j�H;k�H;\�H;C�H;=�H;,�H;��H;��H;m�H; �H;��H;�H;h�H;��H;��H;�H;�H;�H;��H;��H;��H;��H;��H;��H;)�H;��H;�H;��H;      ��H;��H;�H;��H;��H;��H;(�H;��H;�H;��H;�H;��H;��H;S�H;��H;��H;��H;��H;b�H;$�H;��H;�H;��H;��H;��H;.�H;<�H;B�H;S�H;I�H;T�H;Z�H;C�H;=�H;O�H;4�H;+�H;4�H;O�H;=�H;C�H;Z�H;T�H;I�H;S�H;B�H;<�H;.�H;��H;��H;��H;�H;��H;$�H;b�H;��H;��H;��H;��H;S�H;��H;��H;�H;��H;�H;��H;(�H;��H;��H;��H;�H;��H;      i�H;��H;=�H;I�H;��H;.�H;�H;��H;�H;N�H;v�H;��H;��H;|�H;B�H;��H;x�H;��H;��H;��H;��H;4�H;��H;(�H;��H;��H;��H;�H;6�H;J�H;a�H;T�H;E�H;E�H;c�H;U�H;6�H;U�H;c�H;E�H;E�H;T�H;a�H;J�H;6�H;�H;��H;��H;��H;(�H;��H;4�H;��H;��H;��H;��H;x�H;��H;B�H;|�H;��H;��H;v�H;N�H;�H;��H;�H;.�H;��H;I�H;=�H;��H;      ��H;ݶH;��H;8�H;)�H;��H;S�H;N�H;W�H;��H;��H;��H;��H;n�H;��H;�H;;�H;�H;��H;��H;��H;�H;��H;~�H;�H;R�H;��H;��H;�H;+�H;J�H;I�H;X�H;h�H;P�H;b�H;{�H;b�H;P�H;h�H;X�H;I�H;J�H;+�H;�H;��H;��H;R�H;�H;~�H;��H;�H;��H;��H;��H;�H;;�H;�H;��H;n�H;��H;��H;��H;��H;W�H;N�H;S�H;��H;)�H;8�H;��H;ݶH;      3�H;ϠH;[�H;ĤH;��H;��H;��H;�H;��H;H�H;��H;J�H;b�H;J�H;�H;2�H;��H;h�H;��H;��H;<�H;�H;��H;��H;8�H;��H;[�H;��H;��H;�H;6�H;S�H;j�H;l�H;j�H;u�H;u�H;u�H;j�H;l�H;j�H;S�H;6�H;�H;��H;��H;[�H;��H;8�H;��H;��H;�H;<�H;��H;��H;h�H;��H;2�H;�H;J�H;b�H;J�H;��H;H�H;��H;�H;��H;��H;��H;ĤH;[�H;ϠH;      �kH;[mH;�qH;�xH;r�H;ȊH;�H;ʜH;��H; �H;��H;�H;&�H;��H;��H;K�H;Y�H;��H;��H;w�H;��H;��H;�H;G�H;T�H;�H;��H;B�H;��H;��H;�H;B�H;k�H;l�H;��H;��H;��H;��H;��H;l�H;k�H;B�H;�H;��H;��H;B�H;��H;�H;T�H;G�H;�H;��H;��H;w�H;��H;��H;Y�H;K�H;��H;��H;&�H;�H;��H; �H;��H;ʜH;�H;ȊH;r�H;�xH;�qH;[mH;      =�G;��G;/�G;��G;�H;�/H;�KH;?eH;_{H;i�H;m�H;d�H;o�H;��H;žH;3�H;��H;��H;��H;i�H;d�H;��H;#�H;��H;�H;9�H;�H;��H;[�H;��H;��H;<�H;\�H;�H;��H;��H;��H;��H;��H;�H;\�H;<�H;��H;��H;[�H;��H;�H;9�H;�H;��H;#�H;��H;d�H;i�H;��H;��H;��H;3�H;žH;��H;o�H;d�H;m�H;i�H;_{H;?eH;�KH;�/H;�H;��G;/�G;��G;      UHF;3TF;RvF;G�F;��F;�7G;��G;��G;�H;�<H;/eH;p�H;ÖH;�H;��H;ϸH;��H;��H;T�H;Q�H;Y�H;��H;w�H;��H;��H;	�H;9�H;�H;��H;R�H;��H;.�H;C�H;}�H;��H;��H;��H;��H;��H;}�H;C�H;.�H;��H;R�H;��H;�H;9�H;	�H;��H;��H;w�H;��H;Y�H;Q�H;T�H;��H;��H;ϸH;��H;�H;ÖH;p�H;/eH;�<H;�H;��G;��G;�7G;��F;G�F;RvF;3TF;      �B;.�B;�C;ՏC;�/D;��D;1�E;�HF;��F;GiG;R�G;t#H;�[H;/�H;��H;�H;I�H;μH;��H;d�H;��H;��H;�H;5�H;��H;��H;�H;T�H;8�H;�H;��H;��H;=�H;��H;��H;��H;��H;��H;��H;��H;=�H;��H;��H;�H;8�H;T�H;�H;��H;��H;5�H;�H;��H;��H;d�H;��H;μH;I�H;�H;��H;/�H;�[H;t#H;R�G;GiG;��F;�HF;1�E;��D;�/D;ՏC;�C;.�B;      D�:;\�:;��;;'�<;3>;�?;FIA;��B;DED;6{E;WvF;�7G;��G;q&H; eH;s�H;_�H;m�H;��H;��H;�H;:�H;�H;��H;5�H;��H;��H;G�H;��H;~�H;(�H;��H;,�H;l�H;��H;��H;��H;��H;��H;l�H;,�H;��H;(�H;~�H;��H;G�H;��H;��H;5�H;��H;�H;:�H;�H;��H;��H;m�H;_�H;s�H; eH;q&H;��G;�7G;WvF;6{E;DED;��B;FIA;�?;3>;'�<;��;;\�:;      *;��*;�,;�c.;�X1;#�4;E+8;ӊ;;~�>;IA;jwC;�)E;kF;�MG;'�G;DH;"{H;A�H;��H;@�H;S�H;Y�H;��H;�H;�H;w�H;#�H;�H;��H;��H;��H;��H;��H;L�H;��H;��H;��H;��H;��H;L�H;��H;��H;��H;��H;��H;�H;#�H;w�H;�H;�H;��H;Y�H;S�H;@�H;��H;A�H;"{H;DH;'�G;�MG;kF;�)E;jwC;IA;~�>;ӊ;;E+8;#�4;�X1;�c.;�,;��*;      ��
;��;J�;[;��;7`;�C&;�-;�C3;t�8;?H=;��@;�C;c{E;��F;�G;k#H;,mH;��H;?�H;��H;��H;Y�H;:�H;��H;��H;��H;��H;�H;�H;4�H;�H;��H;1�H;r�H;��H;��H;��H;r�H;1�H;��H;�H;4�H;�H;�H;��H;��H;��H;��H;:�H;Y�H;��H;��H;?�H;��H;,mH;k#H;�G;��F;c{E;�C;��@;?H=;t�8;�C3;�-;�C&;7`;��;[;J�;��;      \�:���:��:Ӳ�:���:PO�:�z;i';4�;�}(;�X1;6t8;��=;Z�A;��D;&HF;�bG;�H;>cH;��H;m�H;��H;S�H;�H;��H;Y�H;d�H;��H;<�H;��H;��H;��H;m�H;��H;Y�H;��H;��H;��H;Y�H;��H;m�H;��H;��H;��H;<�H;��H;d�H;Y�H;��H;�H;S�H;��H;m�H;��H;>cH;�H;�bG;&HF;��D;Z�A;��=;6t8;�X1;�}(;4�;i';�z;PO�:���:Ӳ�:��:���:      �R�� ���7��<^9��:P�X:���:���:�O�:=�;7�;�);�C3;��:;� @;�C;k�E;8G;��G;�_H;��H;?�H;@�H;��H;d�H;Q�H;i�H;w�H;��H;��H;��H;$�H; �H;��H;@�H;{�H;{�H;{�H;@�H;��H; �H;$�H;��H;��H;��H;w�H;i�H;Q�H;d�H;��H;@�H;?�H;��H;�_H;��G;8G;k�E;�C;� @;��:;�C3;�);7�;=�;�O�:���:���:P�X:��:�<^9��7�� �      ��)���$�����������=�\�	S���N�9�1j:a��:���:ڃ;�� ;%d.;+8;��>;qC;��E;�(G;��G;>cH;��H;��H;��H;��H;T�H;��H;��H;��H;��H;��H;b�H;��H;w�H;�H;I�H;c�H;I�H;�H;w�H;��H;b�H;��H;��H;��H;��H;��H;T�H;��H;��H;��H;��H;>cH;��G;�(G;��E;qC;��>;+8;%d.;�� ;ڃ;���:a��:�1j:�N�9	S��=�\�������������$�      q�ѻ�ͻP���mG�������d�*�$��Jɺ͇!��C^9��r:���:`0;y�;l�*;�Y6;>;n�B;��E;8G;�H;,mH;A�H;m�H;μH;��H;��H;��H;h�H;�H;��H;��H;�H;�H;��H;�H;<�H;�H;��H;�H;�H;��H;��H;�H;h�H;��H;��H;��H;μH;m�H;A�H;,mH;�H;8G;��E;n�B;>;�Y6;l�*;y�;`0;���:��r:�C^9͇!��Jɺ*�$���d����mG��P����ͻ      ��I�1�E��(;��O*�����<��?GĻ��t@�JҺ{��:�:�O�:O�; ~(;S�5;>;qC;k�E;�bG;k#H;"{H;_�H;I�H;��H;��H;Y�H;��H;;�H;x�H;��H;h�H;��H;Y�H;��H;�H;��H;Y�H;��H;h�H;��H;x�H;;�H;��H;Y�H;��H;��H;I�H;_�H;"{H;k#H;�bG;k�E;qC;>;S�5; ~(;O�;�O�:�:��:{��JҺt@���?GĻ�<������O*��(;�1�E�      &p��\x��ע��R��%��n�`��7�F��G�ѻ-��˃$��ǅ���09�:���:�; ~(;�Y6;��>;�C;&HF;�G;DH;s�H;�H;ϸH;3�H;K�H;2�H;�H;��H;��H;��H;,�H;�H;��H;��H;��H;�H;,�H;��H;��H;��H;�H;2�H;K�H;3�H;ϸH;�H;s�H;DH;�G;&HF;�C;��>;�Y6; ~(;�;���:�:��09�ǅ�˃$�-��G�ѻF���7�n�`�%���R��ע�\x��      &]� �%#�����u�ټ�ɺ������
v��(;�ר�c^��P6R�����	7����:���:O�;l�*;+8;� @;��D;��F;'�G; eH;��H;��H;žH;��H;�H;��H;B�H;��H;��H;��H;��H;B�H;u�H;B�H;��H;��H;��H;��H;B�H;��H;�H;��H;žH;��H;��H; eH;'�G;��F;��D;� @;+8;l�*;O�;���:���:�	7����P6R�c^��ר��(;��
v������ɺ�u�ټ����%#� �      ��_�\�<Q��f@�t +��5�����P�ļs�\�`����bͻfk��Iɺ�	7��:�O�:y�;%d.;��:;Z�A;c{E;�MG;q&H;/�H;�H;��H;��H;J�H;n�H;|�H;S�H;�H;��H;*�H;��H;�H;��H;*�H;��H;�H;S�H;|�H;n�H;J�H;��H;��H;�H;/�H;q&H;�MG;c{E;Z�A;��:;%d.;y�;�O�:�:�	7��Iɺfk�bͻ���\�`�s�P�ļ�����5�t +��f@�<Q�\�      �@���R��ڟ�绒�C����_�:�������$p���vz��O*�5ֻfk������09�:`0;�� ;�C3;��=;�C;kF;��G;�[H;ÖH;o�H;&�H;b�H;��H;��H;��H;�H;'�H;��H;o�H;��H;o�H;��H;'�H;�H;��H;��H;��H;b�H;&�H;o�H;ÖH;�[H;��G;kF;�C;��=;�C3;�� ;`0;�:��09���fk�5ֻ�O*��vz�$p����輙��:���_�C��绒�ڟ��R��      �` �j.��m��ڽ�b��gr��O��\�m +�� ��ɺ�<��O*�bͻP6R��ǅ���:���:ڃ;�);6t8;��@;�)E;�7G;t#H;p�H;d�H;�H;J�H;��H;��H;��H;�H;n�H;�H; �H;?�H; �H;�H;n�H;�H;��H;��H;��H;J�H;�H;d�H;p�H;t#H;�7G;�)E;��@;6t8;�);ڃ;���:��:�ǅ�P6R�bͻ�O*�<��ɺ�� �m +�\�O��gr���b����ڽm��j.��      �-=�1�9��k/�"�����i��y�Ľ�!��Tys�4�6�#��ɺ��vz����c^��˃$�{����r:���:7�;�X1;?H=;jwC;WvF;R�G;/eH;m�H;��H;��H;��H;v�H;�H;��H;��H;��H;��H;��H;��H;��H;��H;��H;�H;v�H;��H;��H;��H;m�H;/eH;R�G;WvF;jwC;?H=;�X1;7�;���:��r:{��˃$�c^������vz��ɺ�#�4�6�Tys��!��y�Ľi���"���k/�1�9�      �(��;l���.}�&ce�jPH���(�o
���ڽ�R����{�4�6�� �$p��\�`�ר�-��JҺ�C^9a��:=�;�}(;t�8;IA;6{E;GiG;�<H;i�H; �H;H�H;��H;N�H;��H;��H;��H;��H;�H;i�H;�H;��H;��H;��H;��H;N�H;��H;H�H; �H;i�H;�<H;GiG;6{E;IA;t�8;�}(;=�;a��:�C^9JҺ-��ר�\�`�$p��� �4�6���{��R����ڽo
���(�jPH�&ce��.}�;l��      �iþGD��)o���������� �i��-=�[t����R��Tys�m +����s񗼗(;�G�ѻt@�͇!��1j:�O�:4�;�C3;~�>;DED;��F;�H;_{H;��H;��H;W�H;�H;�H;��H;9�H;R�H;��H;�H;��H;R�H;9�H;��H;�H;�H;W�H;��H;��H;_{H;�H;��F;DED;~�>;�C3;4�;�O�:�1j:͇!�t@�G�ѻ�(;�s����m +�Tys��R����[t��-=� �i���������)o��GD��      ���
������޾GD���A���.}��D�[t���ڽ�!��\����P�ļ�
v�F�����Jɺ�N�9���:i';�-;ӊ;;��B;�HF;��G;?eH;ʜH;�H;N�H;��H;��H;��H;{�H;��H;�H;��H;�H;��H;{�H;��H;��H;��H;N�H;�H;ʜH;?eH;��G;�HF;��B;ӊ;;�-;i';���:�N�9�Jɺ��F���
v�P�ļ���\��!����ڽ[t��D��.}��A��GD���޾�����
�      ��7�Õ3��f'���\���о�����.}��-=�o
�y�ĽO��:����������7�?GĻ*�$�	S�����:�z;�C&;E+8;FIA;1�E;��G;�KH;�H;��H;S�H;�H;(�H;��H;��H;@�H;��H;5�H;��H;@�H;��H;��H;(�H;�H;S�H;��H;�H;�KH;��G;1�E;FIA;E+8;�C&;�z;���:	S��*�$�?GĻ�7���������:�O��y�Ľo
��-=��.}������о�\����f'�Õ3�      Io�PXi�s"Y���@�@�#��
��о�A�� �i���(�i��gr����_��5��ɺ�n�`��<����d�=�\�P�X:PO�:7`;#�4;�?;��D;�7G;�/H;ȊH;��H;��H;.�H;��H;��H;�H;��H;-�H;��H;-�H;��H;�H;��H;��H;.�H;��H;��H;ȊH;�/H;�7G;��D;�?;#�4;7`;PO�:P�X:=�\���d��<��n�`��ɺ��5���_�gr��i����(� �i��A���о�
�@�#���@�s"Y�PXi�      &����������Io��!J�@�#��\��GD������jPH�����b��C��t +�u�ټ%��������������:���:��;�X1;3>;�/D;��F;�H;r�H;��H;)�H;��H;��H;)�H;��H;p�H;��H;�H;��H;p�H;��H;)�H;��H;��H;)�H;��H;r�H;�H;��F;�/D;3>;�X1;��;���:��:����������%��u�ټt +�C���b�����jPH�����GD���\��@�#��!J�Io��������      2^������b���Io���@���޾����&ce�"����ڽ绒��f@������R���O*�mG������<^9Ӳ�:[;�c.;'�<;ՏC;G�F;��G;�xH;ĤH;8�H;I�H;��H;��H;��H;�H;��H;6�H;��H;�H;��H;��H;��H;I�H;8�H;ĤH;�xH;��G;G�F;ՏC;'�<;�c.;[;Ӳ�:�<^9���mG���O*��R�������f@�绒���ڽ"��&ce������޾���@�Io�b�������      �aǿ֊¿���������s"Y��f'�����)o���.}��k/�m��ڟ�<Q�%#�ע��(;�P��������7���:J�;�,;��;;�C;RvF;/�G;�qH;[�H;��H;=�H;�H;�H;��H;��H;j�H;��H;j�H;��H;��H;�H;�H;=�H;��H;[�H;�qH;/�G;RvF;�C;��;;�,;J�;��:��7����P����(;�ע�%#�<Q�ڟ�m���k/��.}�)o�������f'�s"Y����������֊¿      %�ֿ5pѿ֊¿������PXi�Õ3��
�GD��;l��1�9�j.���R��\� �\x��1�E��ͻ��$�� ����:��;��*;\�:;.�B;3TF;��G;[mH;ϠH;ݶH;��H;��H;��H;�H;��H;<�H;��H;<�H;��H;�H;��H;��H;��H;ݶH;ϠH;[mH;��G;3TF;.�B;\�:;��*;��;���:� ���$��ͻ1�E�\x�� �\��R��j.��1�9�;l��GD���
�Õ3�PXi�������֊¿5pѿ      �?��ph��2v��� ��$�X��O/�#y�-�;Ѱ��j+X�����ѽ����Gn;�>�＿����B(�嚩����.�e9��:^;Y.;��<;�VC;@ZF;�G;5/H;tiH;X�H;s�H;��H;E�H;��H;�H;��H;��H;��H;�H;��H;E�H;��H;s�H;X�H;tiH;5/H;�G;@ZF;�VC;��<;Y.;^;��:.�e9���嚩��B(�����>��Gn;�������ѽ��j+X�Ѱ��-�;#y��O/�$�X�� ��2v��ph��      ph��"���V�����y�EvS�aM+��v� 9ɾ�����T�]��[ν����`\8�����x���%�[��������9C,�:��;�.;N�<; nC;�cF;�G;�0H;!jH;ǋH;ңH;��H;��H;��H;��H;��H;��H;��H;��H;��H;��H;��H;ңH;ǋH;!jH;�0H;�G;�cF; nC;N�<;�.;��;C,�:��9���[����%��x�����`\8������[ν]��T����� 9ɾ�v�aM+�EvS���y�V���"���      2v��V���L ��M�h�%E�I��R���i㼾n���nH�È�a�ý�Ȅ��s/��o༼#�����4J���к��9$f�:Nl;�0;P\=; �C;6�F;��G;Q5H;^lH;H�H;ФH;��H;�H;b�H;��H;$�H; �H;$�H;��H;b�H;�H;��H;ФH;H�H;^lH;Q5H;��G;6�F; �C;P\=;�0;Nl;$f�:��9�к4J������#���o��s/��Ȅ�a�ýÈ��nH�n��i㼾R���I��%E�M�h�L ��V���      � ����y�M�h�ބN��O/����-�߾�A���*|�ؕ6�a}��㳽KSt�(�!�Wrμ(F{��_�
Y��f����:���:WZ;2;�N>;�D;��F;��G;J<H;�oH;��H;t�H;��H;��H;��H;��H;��H;�H;��H;��H;��H;��H;��H;t�H;��H;�oH;J<H;��G;��F;�D;�N>;2;WZ;���:�:f���
Y���_�(F{�Wrμ(�!�KSt��㳽a}�ؕ6��*|��A��-�߾����O/�ބN�M�h���y�      $�X�EvS�%E��O/��S�1W����������4S\�� �q�&�����Y�h��������]�|���S�b��Y���Y:�~�:�_;��4;�?;}�D;�F;/�G;5EH;tH;�H;��H;��H;3�H;��H;E�H;7�H;�H;7�H;E�H;��H;3�H;��H;��H;�H;tH;5EH;/�G;�F;}�D;�?;��4;�_;�~�:��Y:�Y�S�b�|�����]�����h����Y�&���q�� �4S\���������1W���S��O/�%E�EvS�      �O/�aM+�I�����1W�� 9ɾ0���Mw�� :�Y��_�ý�L��Dn;�>���bv���E<��˻(�-�����x�:^;%;�7;��@;V4E;�!G;,�G;iOH;1zH;�H;��H;��H;��H;�H;2�H;�H;��H;�H;2�H;�H;��H;��H;��H;�H;1zH;iOH;,�G;�!G;V4E;��@;�7;%;^;�x�:���(�-��˻�E<�bv��>���Dn;��L��_�ýY��� :��Mw�0�� 9ɾ1W�����I��aM+�      #y��v�R���-�߾����0��1����nH���(Ὁu��r�d�O�Prμ<"�����	��1���k89w:�:��;+;�{:;�6B;)�E;FaG;�H;ZH;��H;M�H;ĮH;�H;e�H;e�H;+�H;��H;��H;��H;+�H;e�H;e�H;�H;ĮH;M�H;��H;ZH;�H;FaG;)�E;�6B;�{:;+;��;w:�:�k891��	�����<"��PrμO�r�d��u��(����nH�1���0������-�߾R����v�      -�; 9ɾi㼾�A�������Mw��nH�����Z��㳽����Z\8�O#�������]N�J��-�b�WJx�z5:��:��;8�0;v\=;v�C;�ZF;�G;)H;eH;��H;G�H;g�H;��H;7�H;��H;P�H;��H;��H;��H;P�H;��H;7�H;��H;g�H;G�H;��H;eH;)H;�G;�ZF;v�C;v\=;8�0;��;��:z5:WJx�-�b�J���]N�����O#��Z\8������㳽�Z񽞯��nH��Mw������A��i㼾 9ɾ      Ѱ������n���*|�4S\�� :����Z�U$������K�c���Oļ����������x&�$��P.�:0^;��#;G6;��?;-�D;��F;��G;*?H;�oH;�H;��H;:�H;r�H;J�H;��H;��H;��H;��H;��H;��H;��H;J�H;r�H;:�H;��H;�H;�oH;*?H;��G;��F;-�D;��?;G6;��#;0^;P.�:$��x&������������Oļc���K����U$���Z���� :�4S\��*|�n������      j+X��T��nH�ؕ6�� �Y��(��㳽����mR����ټ�����E<��?ݻad\�a ��%:�c�:8�;z�,;��:;�6B;ͱE;�KG;jH;�RH;�zH;��H;
�H;9�H;`�H;n�H;+�H;��H;�H;��H;�H;��H;+�H;n�H;`�H;9�H;
�H;��H;�zH;�RH;jH;�KG;ͱE;�6B;��:;z�,;8�;�c�:%:a ��ad\��?ݻ�E<������ټ���mR�����㳽(�Y��� �ؕ6��nH��T�      ��]�È�a}�q�_�ý�u�������K����o�Wv���&R���e^�����@���:�A;�";��4;��>;�D;��F;,�G;)H;�cH;��H;5�H;��H;N�H;M�H;��H;��H;<�H;(�H;��H;(�H;<�H;��H;��H;M�H;N�H;��H;5�H;��H;�cH;)H;,�G;��F;�D;��>;��4;�";�A;��:�@���e^�����&R�Wv���o����K������u��_�ýq�a}�È�]�      ��ѽ�[νa�ý�㳽&����L��r�d�Z\8�c���ټWv����Y��_����y��]���Y:@��:�l; r-;Q�:;��A;rnE;�!G;��G;�FH;�rH;�H;��H;�H;J�H;5�H;��H;��H;��H;B�H;�H;B�H;��H;��H;��H;5�H;J�H;�H;��H;�H;�rH;�FH;��G;�!G;rnE;��A;Q�:; r-;�l;@��:��Y:]�y������_���Y�Wv���ټc��Z\8�r�d��L��&����㳽a�ý�[ν      ���������Ȅ�KSt���Y�Dn;�O�O#���Oļ�����&R��_������N3�,�Y�02:�:9�;A?&;)G6;�W?;�D;fwF;�G;c H;�]H;��H;�H;�H;a�H;#�H;�H;��H;(�H;��H;i�H;%�H;i�H;��H;(�H;��H;�H;#�H;a�H;�H;�H;��H;�]H;c H;�G;fwF;�D;�W?;)G6;A?&;9�;�:02:,�Y��N3������_��&R������OļO#��O�Dn;���Y�KSt��Ȅ�����      Gn;�`\8��s/�(�!�h��>���Prμ��������E<�������N3��Ix�f�9��:U^;� ;2;��<;.�B;�E;e4G;2�G;^EH;�pH;��H;h�H;гH;k�H;��H;��H;�H;��H;1�H;��H;�H;��H;1�H;��H;�H;��H;��H;k�H;гH;h�H;��H;�pH;^EH;2�G;e4G;�E;.�B;��<;2;� ;U^;��:f�9�Ix��N3�������E<��������Prμ>���h��(�!��s/�`\8�      >�Ｘ���o�Wrμ����bv��<"���]N�����?ݻe^��y��,�Y�f�9��:���:B�;��.;�{:;2>A;��D;`�F;ߵG;
)H;E`H;5�H;��H;�H;R�H;6�H;R�H;t�H;�H;.�H;k�H;��H;��H;��H;k�H;.�H;�H;t�H;R�H;6�H;R�H;�H;��H;5�H;E`H;
)H;ߵG;`�F;��D;2>A;�{:;��.;B�;���:��:f�9,�Y�y��e^���?ݻ����]N�<"��bv������Wrμ�o༸��      �����x���#��(F{���]��E<����J�뻱���ad\���]�02:��:���:�Z;��,;/�8;a @;0D;�ZF;QzG;
H;jOH;>uH;�H;\�H;�H;C�H;z�H;��H;��H;��H;��H;��H;��H;��H;��H;��H;��H;��H;��H;��H;z�H;C�H;�H;\�H;�H;>uH;jOH;
H;QzG;�ZF;0D;a @;/�8;��,;�Z;���:��:02:]���ad\�����J�뻛���E<���]�(F{��#���x��      �B(��%�����_�|����˻	��-�b�x&�a ���@���Y:�:U^;B�;��,;Z_8;��?;��C;�F;FG;u�G;?H;GjH;#�H; �H;
�H;k�H;��H;�H;��H;/�H;��H;��H;��H;��H;��H;��H;��H;��H;��H;/�H;��H;�H;��H;k�H;
�H; �H;#�H;GjH;?H;u�G;FG;�F;��C;��?;Z_8;��,;B�;U^;�:��Y:�@�a ��x&�-�b�	���˻|����_�����%�      嚩�[���4J��
Y��S�b�(�-�1��WJx�$��%:��:@��:9�;� ;��.;/�8;��?;2�C;�E;f"G;�G;1H;aH;gH;��H;��H;��H;��H;s�H;(�H;I�H;J�H;��H;(�H;��H;H�H;��H;H�H;��H;(�H;��H;J�H;I�H;(�H;s�H;��H;��H;��H;��H;gH;aH;1H;�G;f"G;�E;2�C;��?;/�8;��.;� ;9�;@��:��:%:$��WJx�1��(�-�S�b�
Y��4J��[���      �����뺶кf����Y�����k89z5:P.�:�c�:�A;�l;A?&;2;�{:;a @;��C;�E;�G;�G;}'H;ZH;�yH;W�H;��H;��H;{�H;��H;��H;l�H;��H;�H;[�H;<�H;W�H;
�H;��H;
�H;W�H;<�H;[�H;�H;��H;l�H;��H;��H;{�H;��H;��H;W�H;�yH;ZH;}'H;�G;�G;�E;��C;a @;�{:;2;A?&;�l;�A;�c�:P.�:z5:�k89����Y�f����к���      .�e9��9��9�:��Y:�x�:w:�:��:0^;8�;�"; r-;)G6;��<;2>A;0D;�F;f"G;�G;$H;VH;�uH;��H;Y�H;b�H;��H;!�H;��H;��H;E�H;��H;��H;��H;6�H;�H;��H;�H;��H;�H;6�H;��H;��H;��H;E�H;��H;��H;!�H;��H;b�H;Y�H;��H;�uH;VH;$H;�G;f"G;�F;0D;2>A;��<;)G6; r-;�";8�;0^;��:w:�:�x�:��Y:�:��9��9      ��:C,�:$f�:���:�~�:^;��;��;��#;z�,;��4;Q�:;�W?;.�B;��D;�ZF;FG;�G;}'H;VH;�tH;��H;.�H;�H;<�H;
�H;��H;��H;��H;��H;��H;��H;��H;��H;��H;^�H;b�H;^�H;��H;��H;��H;��H;��H;��H;��H;��H;��H;
�H;<�H;�H;.�H;��H;�tH;VH;}'H;�G;FG;�ZF;��D;.�B;�W?;Q�:;��4;z�,;��#;��;��;^;�~�:���:$f�:C,�:      ^;��;Nl;WZ;�_;%;+;8�0;G6;��:;��>;��A;�D;�E;`�F;QzG;u�G;1H;ZH;�uH;��H;g�H;ܫH;�H;��H;e�H;��H;��H;��H;��H;H�H;G�H;��H;��H;p�H;��H;��H;��H;p�H;��H;��H;G�H;H�H;��H;��H;��H;��H;e�H;��H;�H;ܫH;g�H;��H;�uH;ZH;1H;u�G;QzG;`�F;�E;�D;��A;��>;��:;G6;8�0;+;%;�_;WZ;Nl;��;      Y.;�.;�0;2;��4;�7;�{:;v\=;��?;�6B;�D;rnE;fwF;e4G;ߵG;
H;?H;aH;�yH;��H;.�H;ܫH;`�H;��H;�H;��H;��H;�H;)�H;��H;��H;h�H;c�H;O�H;��H;(�H;P�H;(�H;��H;O�H;c�H;h�H;��H;��H;)�H;�H;��H;��H;�H;��H;`�H;ܫH;.�H;��H;�yH;aH;?H;
H;ߵG;e4G;fwF;rnE;�D;�6B;��?;v\=;�{:;�7;��4;2;�0;�.;      ��<;N�<;P\=;�N>;�?;��@;�6B;v�C;-�D;ͱE;��F;�!G;�G;2�G;
)H;jOH;GjH;gH;W�H;Y�H;�H;�H;��H;H�H;I�H;E�H;W�H;��H;,�H;B�H;�H;�H;�H;��H;I�H;��H;��H;��H;I�H;��H;�H;�H;�H;B�H;,�H;��H;W�H;E�H;I�H;H�H;��H;�H;�H;Y�H;W�H;gH;GjH;jOH;
)H;2�G;�G;�!G;��F;ͱE;-�D;v�C;�6B;��@;�?;�N>;P\=;N�<;      �VC; nC; �C;�D;}�D;V4E;)�E;�ZF;��F;�KG;,�G;��G;c H;^EH;E`H;>uH;#�H;��H;��H;b�H;<�H;��H;�H;I�H;�H;�H;O�H;��H;��H;��H;��H;��H;��H;=�H;��H;��H;��H;��H;��H;=�H;��H;��H;��H;��H;��H;��H;O�H;�H;�H;I�H;�H;��H;<�H;b�H;��H;��H;#�H;>uH;E`H;^EH;c H;��G;,�G;�KG;��F;�ZF;)�E;V4E;}�D;�D; �C; nC;      @ZF;�cF;6�F;��F;�F;�!G;FaG;�G;��G;jH;)H;�FH;�]H;�pH;5�H;�H; �H;��H;��H;��H;
�H;e�H;��H;E�H;�H;5�H;��H;��H;u�H;��H;��H;��H;,�H;~�H;��H;�H;�H;�H;��H;~�H;,�H;��H;��H;��H;u�H;��H;��H;5�H;�H;E�H;��H;e�H;
�H;��H;��H;��H; �H;�H;5�H;�pH;�]H;�FH;)H;jH;��G;�G;FaG;�!G;�F;��F;6�F;�cF;      �G;�G;��G;��G;/�G;,�G;�H;)H;*?H;�RH;�cH;�rH;��H;��H;��H;\�H;
�H;��H;{�H;!�H;��H;��H;��H;W�H;O�H;��H;��H;J�H;��H;��H;j�H; �H;}�H;��H;�H;;�H;Y�H;;�H;�H;��H;}�H; �H;j�H;��H;��H;J�H;��H;��H;O�H;W�H;��H;��H;��H;!�H;{�H;��H;
�H;\�H;��H;��H;��H;�rH;�cH;�RH;*?H;)H;�H;,�G;/�G;��G;��G;�G;      5/H;�0H;Q5H;J<H;5EH;iOH;ZH;eH;�oH;�zH;��H;�H;�H;h�H;�H;�H;k�H;��H;��H;��H;��H;��H;�H;��H;��H;��H;J�H;��H;e�H;S�H;�H;j�H;��H;�H;E�H;[�H;M�H;[�H;E�H;�H;��H;j�H;�H;S�H;e�H;��H;J�H;��H;��H;��H;�H;��H;��H;��H;��H;��H;k�H;�H;�H;h�H;�H;�H;��H;�zH;�oH;eH;ZH;iOH;5EH;J<H;Q5H;�0H;      tiH;!jH;^lH;�oH;tH;1zH;��H;��H;�H;��H;5�H;��H;�H;гH;R�H;C�H;��H;s�H;��H;��H;��H;��H;)�H;,�H;��H;u�H;��H;e�H;[�H;��H;Z�H;��H;��H;5�H;e�H;o�H;b�H;o�H;e�H;5�H;��H;��H;Z�H;��H;[�H;e�H;��H;u�H;��H;,�H;)�H;��H;��H;��H;��H;s�H;��H;C�H;R�H;гH;�H;��H;5�H;��H;�H;��H;��H;1zH;tH;�oH;^lH;!jH;      X�H;ǋH;H�H;��H;�H;�H;M�H;G�H;��H;
�H;��H;�H;a�H;k�H;6�H;z�H;�H;(�H;l�H;E�H;��H;��H;��H;B�H;��H;��H;��H;S�H;��H;K�H;��H;��H;6�H;]�H;h�H;��H;��H;��H;h�H;]�H;6�H;��H;��H;K�H;��H;S�H;��H;��H;��H;B�H;��H;��H;��H;E�H;l�H;(�H;�H;z�H;6�H;k�H;a�H;�H;��H;
�H;��H;G�H;M�H;�H;�H;��H;H�H;ǋH;      s�H;ңH;ФH;t�H;��H;��H;ĮH;g�H;:�H;9�H;N�H;J�H;#�H;��H;R�H;��H;��H;I�H;��H;��H;��H;H�H;��H;�H;��H;��H;j�H;�H;Z�H;��H;��H;)�H;a�H;o�H;��H;��H;��H;��H;��H;o�H;a�H;)�H;��H;��H;Z�H;�H;j�H;��H;��H;�H;��H;H�H;��H;��H;��H;I�H;��H;��H;R�H;��H;#�H;J�H;N�H;9�H;:�H;g�H;ĮH;��H;��H;t�H;ФH;ңH;      ��H;��H;��H;��H;��H;��H;�H;��H;r�H;`�H;M�H;5�H;�H;��H;t�H;��H;/�H;J�H;�H;��H;��H;G�H;h�H;�H;��H;��H; �H;j�H;��H;��H;)�H;A�H;l�H;��H;��H;��H;��H;��H;��H;��H;l�H;A�H;)�H;��H;��H;j�H; �H;��H;��H;�H;h�H;G�H;��H;��H;�H;J�H;/�H;��H;t�H;��H;�H;5�H;M�H;`�H;r�H;��H;�H;��H;��H;��H;��H;��H;      E�H;��H;�H;��H;3�H;��H;e�H;7�H;J�H;n�H;��H;��H;��H;�H;�H;��H;��H;��H;[�H;��H;��H;��H;c�H;�H;��H;,�H;}�H;��H;��H;6�H;a�H;l�H;{�H;��H;��H;��H;��H;��H;��H;��H;{�H;l�H;a�H;6�H;��H;��H;}�H;,�H;��H;�H;c�H;��H;��H;��H;[�H;��H;��H;��H;�H;�H;��H;��H;��H;n�H;J�H;7�H;e�H;��H;3�H;��H;�H;��H;      ��H;��H;b�H;��H;��H;�H;e�H;��H;��H;+�H;��H;��H;(�H;��H;.�H;��H;��H;(�H;<�H;6�H;��H;��H;O�H;��H;=�H;~�H;��H;�H;5�H;]�H;o�H;��H;��H;��H;��H;��H;��H;��H;��H;��H;��H;��H;o�H;]�H;5�H;�H;��H;~�H;=�H;��H;O�H;��H;��H;6�H;<�H;(�H;��H;��H;.�H;��H;(�H;��H;��H;+�H;��H;��H;e�H;�H;��H;��H;b�H;��H;      �H;��H;��H;��H;E�H;2�H;+�H;P�H;��H;��H;<�H;��H;��H;1�H;k�H;��H;��H;��H;W�H;�H;��H;p�H;��H;I�H;��H;��H;�H;E�H;e�H;h�H;��H;��H;��H;��H;��H;��H;��H;��H;��H;��H;��H;��H;��H;h�H;e�H;E�H;�H;��H;��H;I�H;��H;p�H;��H;�H;W�H;��H;��H;��H;k�H;1�H;��H;��H;<�H;��H;��H;P�H;+�H;2�H;E�H;��H;��H;��H;      ��H;��H;$�H;��H;7�H;�H;��H;��H;��H;�H;(�H;B�H;i�H;��H;��H;��H;��H;H�H;
�H;��H;^�H;��H;(�H;��H;��H;�H;;�H;[�H;o�H;��H;��H;��H;��H;��H;��H;��H;��H;��H;��H;��H;��H;��H;��H;��H;o�H;[�H;;�H;�H;��H;��H;(�H;��H;^�H;��H;
�H;H�H;��H;��H;��H;��H;i�H;B�H;(�H;�H;��H;��H;��H;�H;7�H;��H;$�H;��H;      ��H;��H; �H;�H;�H;��H;��H;��H;��H;��H;��H;�H;%�H;�H;��H;��H;��H;��H;��H;�H;b�H;��H;P�H;��H;��H;�H;Y�H;M�H;b�H;��H;��H;��H;��H;��H;��H;��H;��H;��H;��H;��H;��H;��H;��H;��H;b�H;M�H;Y�H;�H;��H;��H;P�H;��H;b�H;�H;��H;��H;��H;��H;��H;�H;%�H;�H;��H;��H;��H;��H;��H;��H;�H;�H; �H;��H;      ��H;��H;$�H;��H;7�H;�H;��H;��H;��H;�H;(�H;B�H;i�H;��H;��H;��H;��H;H�H;
�H;��H;^�H;��H;(�H;��H;��H;�H;;�H;[�H;o�H;��H;��H;��H;��H;��H;��H;��H;��H;��H;��H;��H;��H;��H;��H;��H;o�H;[�H;;�H;�H;��H;��H;(�H;��H;^�H;��H;
�H;H�H;��H;��H;��H;��H;i�H;B�H;(�H;�H;��H;��H;��H;�H;7�H;��H;$�H;��H;      �H;��H;��H;��H;E�H;2�H;+�H;P�H;��H;��H;<�H;��H;��H;1�H;k�H;��H;��H;��H;W�H;�H;��H;p�H;��H;I�H;��H;��H;�H;E�H;e�H;h�H;��H;��H;��H;��H;��H;��H;��H;��H;��H;��H;��H;��H;��H;h�H;e�H;E�H;�H;��H;��H;I�H;��H;p�H;��H;�H;W�H;��H;��H;��H;k�H;1�H;��H;��H;<�H;��H;��H;P�H;+�H;2�H;E�H;��H;��H;��H;      ��H;��H;b�H;��H;��H;�H;e�H;��H;��H;+�H;��H;��H;(�H;��H;.�H;��H;��H;(�H;<�H;6�H;��H;��H;O�H;��H;=�H;~�H;��H;�H;5�H;]�H;o�H;��H;��H;��H;��H;��H;��H;��H;��H;��H;��H;��H;o�H;]�H;5�H;�H;��H;~�H;=�H;��H;O�H;��H;��H;6�H;<�H;(�H;��H;��H;.�H;��H;(�H;��H;��H;+�H;��H;��H;e�H;�H;��H;��H;b�H;��H;      E�H;��H;�H;��H;3�H;��H;e�H;7�H;J�H;n�H;��H;��H;��H;�H;�H;��H;��H;��H;[�H;��H;��H;��H;c�H;�H;��H;,�H;}�H;��H;��H;6�H;a�H;l�H;{�H;��H;��H;��H;��H;��H;��H;��H;{�H;l�H;a�H;6�H;��H;��H;}�H;,�H;��H;�H;c�H;��H;��H;��H;[�H;��H;��H;��H;�H;�H;��H;��H;��H;n�H;J�H;7�H;e�H;��H;3�H;��H;�H;��H;      ��H;��H;��H;��H;��H;��H;�H;��H;r�H;`�H;M�H;5�H;�H;��H;t�H;��H;/�H;J�H;�H;��H;��H;G�H;h�H;�H;��H;��H; �H;j�H;��H;��H;)�H;A�H;l�H;��H;��H;��H;��H;��H;��H;��H;l�H;A�H;)�H;��H;��H;j�H; �H;��H;��H;�H;h�H;G�H;��H;��H;�H;J�H;/�H;��H;t�H;��H;�H;5�H;M�H;`�H;r�H;��H;�H;��H;��H;��H;��H;��H;      s�H;ңH;ФH;t�H;��H;��H;ĮH;g�H;:�H;9�H;N�H;J�H;#�H;��H;R�H;��H;��H;I�H;��H;��H;��H;H�H;��H;�H;��H;��H;j�H;�H;Z�H;��H;��H;)�H;a�H;o�H;��H;��H;��H;��H;��H;o�H;a�H;)�H;��H;��H;Z�H;�H;j�H;��H;��H;�H;��H;H�H;��H;��H;��H;I�H;��H;��H;R�H;��H;#�H;J�H;N�H;9�H;:�H;g�H;ĮH;��H;��H;t�H;ФH;ңH;      X�H;ǋH;H�H;��H;�H;�H;M�H;G�H;��H;
�H;��H;�H;a�H;k�H;6�H;z�H;�H;(�H;l�H;E�H;��H;��H;��H;B�H;��H;��H;��H;S�H;��H;K�H;��H;��H;6�H;]�H;h�H;��H;��H;��H;h�H;]�H;6�H;��H;��H;K�H;��H;S�H;��H;��H;��H;B�H;��H;��H;��H;E�H;l�H;(�H;�H;z�H;6�H;k�H;a�H;�H;��H;
�H;��H;G�H;M�H;�H;�H;��H;H�H;ǋH;      tiH;!jH;^lH;�oH;tH;1zH;��H;��H;�H;��H;5�H;��H;�H;гH;R�H;C�H;��H;s�H;��H;��H;��H;��H;)�H;,�H;��H;u�H;��H;e�H;[�H;��H;Z�H;��H;��H;5�H;e�H;o�H;b�H;o�H;e�H;5�H;��H;��H;Z�H;��H;[�H;e�H;��H;u�H;��H;,�H;)�H;��H;��H;��H;��H;s�H;��H;C�H;R�H;гH;�H;��H;5�H;��H;�H;��H;��H;1zH;tH;�oH;^lH;!jH;      5/H;�0H;Q5H;J<H;5EH;iOH;ZH;eH;�oH;�zH;��H;�H;�H;h�H;�H;�H;k�H;��H;��H;��H;��H;��H;�H;��H;��H;��H;J�H;��H;e�H;S�H;�H;j�H;��H;�H;E�H;[�H;M�H;[�H;E�H;�H;��H;j�H;�H;S�H;e�H;��H;J�H;��H;��H;��H;�H;��H;��H;��H;��H;��H;k�H;�H;�H;h�H;�H;�H;��H;�zH;�oH;eH;ZH;iOH;5EH;J<H;Q5H;�0H;      �G;�G;��G;��G;/�G;,�G;�H;)H;*?H;�RH;�cH;�rH;��H;��H;��H;\�H;
�H;��H;{�H;!�H;��H;��H;��H;W�H;O�H;��H;��H;J�H;��H;��H;j�H; �H;}�H;��H;�H;;�H;Y�H;;�H;�H;��H;}�H; �H;j�H;��H;��H;J�H;��H;��H;O�H;W�H;��H;��H;��H;!�H;{�H;��H;
�H;\�H;��H;��H;��H;�rH;�cH;�RH;*?H;)H;�H;,�G;/�G;��G;��G;�G;      @ZF;�cF;6�F;��F;�F;�!G;FaG;�G;��G;jH;)H;�FH;�]H;�pH;5�H;�H; �H;��H;��H;��H;
�H;e�H;��H;E�H;�H;5�H;��H;��H;u�H;��H;��H;��H;,�H;~�H;��H;�H;�H;�H;��H;~�H;,�H;��H;��H;��H;u�H;��H;��H;5�H;�H;E�H;��H;e�H;
�H;��H;��H;��H; �H;�H;5�H;�pH;�]H;�FH;)H;jH;��G;�G;FaG;�!G;�F;��F;6�F;�cF;      �VC; nC; �C;�D;}�D;V4E;)�E;�ZF;��F;�KG;,�G;��G;c H;^EH;E`H;>uH;#�H;��H;��H;b�H;<�H;��H;�H;I�H;�H;�H;O�H;��H;��H;��H;��H;��H;��H;=�H;��H;��H;��H;��H;��H;=�H;��H;��H;��H;��H;��H;��H;O�H;�H;�H;I�H;�H;��H;<�H;b�H;��H;��H;#�H;>uH;E`H;^EH;c H;��G;,�G;�KG;��F;�ZF;)�E;V4E;}�D;�D; �C; nC;      ��<;N�<;P\=;�N>;�?;��@;�6B;v�C;-�D;ͱE;��F;�!G;�G;2�G;
)H;jOH;GjH;gH;W�H;Y�H;�H;�H;��H;H�H;I�H;E�H;W�H;��H;,�H;B�H;�H;�H;�H;��H;I�H;��H;��H;��H;I�H;��H;�H;�H;�H;B�H;,�H;��H;W�H;E�H;I�H;H�H;��H;�H;�H;Y�H;W�H;gH;GjH;jOH;
)H;2�G;�G;�!G;��F;ͱE;-�D;v�C;�6B;��@;�?;�N>;P\=;N�<;      Y.;�.;�0;2;��4;�7;�{:;v\=;��?;�6B;�D;rnE;fwF;e4G;ߵG;
H;?H;aH;�yH;��H;.�H;ܫH;`�H;��H;�H;��H;��H;�H;)�H;��H;��H;h�H;c�H;O�H;��H;(�H;P�H;(�H;��H;O�H;c�H;h�H;��H;��H;)�H;�H;��H;��H;�H;��H;`�H;ܫH;.�H;��H;�yH;aH;?H;
H;ߵG;e4G;fwF;rnE;�D;�6B;��?;v\=;�{:;�7;��4;2;�0;�.;      ^;��;Nl;WZ;�_;%;+;8�0;G6;��:;��>;��A;�D;�E;`�F;QzG;u�G;1H;ZH;�uH;��H;g�H;ܫH;�H;��H;e�H;��H;��H;��H;��H;H�H;G�H;��H;��H;p�H;��H;��H;��H;p�H;��H;��H;G�H;H�H;��H;��H;��H;��H;e�H;��H;�H;ܫH;g�H;��H;�uH;ZH;1H;u�G;QzG;`�F;�E;�D;��A;��>;��:;G6;8�0;+;%;�_;WZ;Nl;��;      ��:C,�:$f�:���:�~�:^;��;��;��#;z�,;��4;Q�:;�W?;.�B;��D;�ZF;FG;�G;}'H;VH;�tH;��H;.�H;�H;<�H;
�H;��H;��H;��H;��H;��H;��H;��H;��H;��H;^�H;b�H;^�H;��H;��H;��H;��H;��H;��H;��H;��H;��H;
�H;<�H;�H;.�H;��H;�tH;VH;}'H;�G;FG;�ZF;��D;.�B;�W?;Q�:;��4;z�,;��#;��;��;^;�~�:���:$f�:C,�:      .�e9��9��9�:��Y:�x�:w:�:��:0^;8�;�"; r-;)G6;��<;2>A;0D;�F;f"G;�G;$H;VH;�uH;��H;Y�H;b�H;��H;!�H;��H;��H;E�H;��H;��H;��H;6�H;�H;��H;�H;��H;�H;6�H;��H;��H;��H;E�H;��H;��H;!�H;��H;b�H;Y�H;��H;�uH;VH;$H;�G;f"G;�F;0D;2>A;��<;)G6; r-;�";8�;0^;��:w:�:�x�:��Y:�:��9��9      �����뺶кf����Y�����k89z5:P.�:�c�:�A;�l;A?&;2;�{:;a @;��C;�E;�G;�G;}'H;ZH;�yH;W�H;��H;��H;{�H;��H;��H;l�H;��H;�H;[�H;<�H;W�H;
�H;��H;
�H;W�H;<�H;[�H;�H;��H;l�H;��H;��H;{�H;��H;��H;W�H;�yH;ZH;}'H;�G;�G;�E;��C;a @;�{:;2;A?&;�l;�A;�c�:P.�:z5:�k89����Y�f����к���      嚩�[���4J��
Y��S�b�(�-�1��WJx�$��%:��:@��:9�;� ;��.;/�8;��?;2�C;�E;f"G;�G;1H;aH;gH;��H;��H;��H;��H;s�H;(�H;I�H;J�H;��H;(�H;��H;H�H;��H;H�H;��H;(�H;��H;J�H;I�H;(�H;s�H;��H;��H;��H;��H;gH;aH;1H;�G;f"G;�E;2�C;��?;/�8;��.;� ;9�;@��:��:%:$��WJx�1��(�-�S�b�
Y��4J��[���      �B(��%�����_�|����˻	��-�b�x&�a ���@���Y:�:U^;B�;��,;Z_8;��?;��C;�F;FG;u�G;?H;GjH;#�H; �H;
�H;k�H;��H;�H;��H;/�H;��H;��H;��H;��H;��H;��H;��H;��H;��H;/�H;��H;�H;��H;k�H;
�H; �H;#�H;GjH;?H;u�G;FG;�F;��C;��?;Z_8;��,;B�;U^;�:��Y:�@�a ��x&�-�b�	���˻|����_�����%�      �����x���#��(F{���]��E<����J�뻱���ad\���]�02:��:���:�Z;��,;/�8;a @;0D;�ZF;QzG;
H;jOH;>uH;�H;\�H;�H;C�H;z�H;��H;��H;��H;��H;��H;��H;��H;��H;��H;��H;��H;��H;��H;z�H;C�H;�H;\�H;�H;>uH;jOH;
H;QzG;�ZF;0D;a @;/�8;��,;�Z;���:��:02:]���ad\�����J�뻛���E<���]�(F{��#���x��      >�Ｘ���o�Wrμ����bv��<"���]N�����?ݻe^��y��,�Y�f�9��:���:B�;��.;�{:;2>A;��D;`�F;ߵG;
)H;E`H;5�H;��H;�H;R�H;6�H;R�H;t�H;�H;.�H;k�H;��H;��H;��H;k�H;.�H;�H;t�H;R�H;6�H;R�H;�H;��H;5�H;E`H;
)H;ߵG;`�F;��D;2>A;�{:;��.;B�;���:��:f�9,�Y�y��e^���?ݻ����]N�<"��bv������Wrμ�o༸��      Gn;�`\8��s/�(�!�h��>���Prμ��������E<�������N3��Ix�f�9��:U^;� ;2;��<;.�B;�E;e4G;2�G;^EH;�pH;��H;h�H;гH;k�H;��H;��H;�H;��H;1�H;��H;�H;��H;1�H;��H;�H;��H;��H;k�H;гH;h�H;��H;�pH;^EH;2�G;e4G;�E;.�B;��<;2;� ;U^;��:f�9�Ix��N3�������E<��������Prμ>���h��(�!��s/�`\8�      ���������Ȅ�KSt���Y�Dn;�O�O#���Oļ�����&R��_������N3�,�Y�02:�:9�;A?&;)G6;�W?;�D;fwF;�G;c H;�]H;��H;�H;�H;a�H;#�H;�H;��H;(�H;��H;i�H;%�H;i�H;��H;(�H;��H;�H;#�H;a�H;�H;�H;��H;�]H;c H;�G;fwF;�D;�W?;)G6;A?&;9�;�:02:,�Y��N3������_��&R������OļO#��O�Dn;���Y�KSt��Ȅ�����      ��ѽ�[νa�ý�㳽&����L��r�d�Z\8�c���ټWv����Y��_����y��]���Y:@��:�l; r-;Q�:;��A;rnE;�!G;��G;�FH;�rH;�H;��H;�H;J�H;5�H;��H;��H;��H;B�H;�H;B�H;��H;��H;��H;5�H;J�H;�H;��H;�H;�rH;�FH;��G;�!G;rnE;��A;Q�:; r-;�l;@��:��Y:]�y������_���Y�Wv���ټc��Z\8�r�d��L��&����㳽a�ý�[ν      ��]�È�a}�q�_�ý�u�������K����o�Wv���&R���e^�����@���:�A;�";��4;��>;�D;��F;,�G;)H;�cH;��H;5�H;��H;N�H;M�H;��H;��H;<�H;(�H;��H;(�H;<�H;��H;��H;M�H;N�H;��H;5�H;��H;�cH;)H;,�G;��F;�D;��>;��4;�";�A;��:�@���e^�����&R�Wv���o����K������u��_�ýq�a}�È�]�      j+X��T��nH�ؕ6�� �Y��(��㳽����mR����ټ�����E<��?ݻad\�a ��%:�c�:8�;z�,;��:;�6B;ͱE;�KG;jH;�RH;�zH;��H;
�H;9�H;`�H;n�H;+�H;��H;�H;��H;�H;��H;+�H;n�H;`�H;9�H;
�H;��H;�zH;�RH;jH;�KG;ͱE;�6B;��:;z�,;8�;�c�:%:a ��ad\��?ݻ�E<������ټ���mR�����㳽(�Y��� �ؕ6��nH��T�      Ѱ������n���*|�4S\�� :����Z�U$������K�c���Oļ����������x&�$��P.�:0^;��#;G6;��?;-�D;��F;��G;*?H;�oH;�H;��H;:�H;r�H;J�H;��H;��H;��H;��H;��H;��H;��H;J�H;r�H;:�H;��H;�H;�oH;*?H;��G;��F;-�D;��?;G6;��#;0^;P.�:$��x&������������Oļc���K����U$���Z���� :�4S\��*|�n������      -�; 9ɾi㼾�A�������Mw��nH�����Z��㳽����Z\8�O#�������]N�J��-�b�WJx�z5:��:��;8�0;v\=;v�C;�ZF;�G;)H;eH;��H;G�H;g�H;��H;7�H;��H;P�H;��H;��H;��H;P�H;��H;7�H;��H;g�H;G�H;��H;eH;)H;�G;�ZF;v�C;v\=;8�0;��;��:z5:WJx�-�b�J���]N�����O#��Z\8������㳽�Z񽞯��nH��Mw������A��i㼾 9ɾ      #y��v�R���-�߾����0��1����nH���(Ὁu��r�d�O�Prμ<"�����	��1���k89w:�:��;+;�{:;�6B;)�E;FaG;�H;ZH;��H;M�H;ĮH;�H;e�H;e�H;+�H;��H;��H;��H;+�H;e�H;e�H;�H;ĮH;M�H;��H;ZH;�H;FaG;)�E;�6B;�{:;+;��;w:�:�k891��	�����<"��PrμO�r�d��u��(����nH�1���0������-�߾R����v�      �O/�aM+�I�����1W�� 9ɾ0���Mw�� :�Y��_�ý�L��Dn;�>���bv���E<��˻(�-�����x�:^;%;�7;��@;V4E;�!G;,�G;iOH;1zH;�H;��H;��H;��H;�H;2�H;�H;��H;�H;2�H;�H;��H;��H;��H;�H;1zH;iOH;,�G;�!G;V4E;��@;�7;%;^;�x�:���(�-��˻�E<�bv��>���Dn;��L��_�ýY��� :��Mw�0�� 9ɾ1W�����I��aM+�      $�X�EvS�%E��O/��S�1W����������4S\�� �q�&�����Y�h��������]�|���S�b��Y���Y:�~�:�_;��4;�?;}�D;�F;/�G;5EH;tH;�H;��H;��H;3�H;��H;E�H;7�H;�H;7�H;E�H;��H;3�H;��H;��H;�H;tH;5EH;/�G;�F;}�D;�?;��4;�_;�~�:��Y:�Y�S�b�|�����]�����h����Y�&���q�� �4S\���������1W���S��O/�%E�EvS�      � ����y�M�h�ބN��O/����-�߾�A���*|�ؕ6�a}��㳽KSt�(�!�Wrμ(F{��_�
Y��f����:���:WZ;2;�N>;�D;��F;��G;J<H;�oH;��H;t�H;��H;��H;��H;��H;��H;�H;��H;��H;��H;��H;��H;t�H;��H;�oH;J<H;��G;��F;�D;�N>;2;WZ;���:�:f���
Y���_�(F{�Wrμ(�!�KSt��㳽a}�ؕ6��*|��A��-�߾����O/�ބN�M�h���y�      2v��V���L ��M�h�%E�I��R���i㼾n���nH�È�a�ý�Ȅ��s/��o༼#�����4J���к��9$f�:Nl;�0;P\=; �C;6�F;��G;Q5H;^lH;H�H;ФH;��H;�H;b�H;��H;$�H; �H;$�H;��H;b�H;�H;��H;ФH;H�H;^lH;Q5H;��G;6�F; �C;P\=;�0;Nl;$f�:��9�к4J������#���o��s/��Ȅ�a�ýÈ��nH�n��i㼾R���I��%E�M�h�L ��V���      ph��"���V�����y�EvS�aM+��v� 9ɾ�����T�]��[ν����`\8�����x���%�[��������9C,�:��;�.;N�<; nC;�cF;�G;�0H;!jH;ǋH;ңH;��H;��H;��H;��H;��H;��H;��H;��H;��H;��H;��H;ңH;ǋH;!jH;�0H;�G;�cF; nC;N�<;�.;��;C,�:��9���[����%��x�����`\8������[ν]��T����� 9ɾ�v�aM+�EvS���y�V���"���      .Eb�I]�tN�ߛ7����e� �{�˾��	�j��!,�J���0��m���,˼��x�E���1��`���S�:g�:3;��1;n+>;��C;�vF;�G;��G;>H;�gH;Z�H;w�H;9�H;�H;��H;(�H;��H;(�H;��H;�H;9�H;w�H;Z�H;�gH;>H;��G;�G;�vF;��C;n+>;��1;3;g�:S�:`����1��E����x�,˼��m�0��J����!,�	�j���{�˾e� ����ߛ7�tN�I]�      I]�N�W��TI�v3��D�������Ǿb���ȟf� )� ��W;���Fi��k�x�Ǽ�[t�8�	�(Ȅ�sX��џ:���:&�;�I2;�Y>;qD;�~F;\�G;+H;�>H;�hH;�H;�H;r�H;7�H;��H;S�H;��H;S�H;��H;7�H;r�H;�H;�H;�hH;�>H;+H;\�G;�~F;qD;�Y>;�I2;&�;���:џ:sX��(Ȅ�8�	��[t�x�Ǽ�k��Fi�W;�� �� )�ȟf�b�����Ǿ�����D�v3��TI�N�W�      tN��TI���;��'��k���i���f󐾖Z��K ��s�&����&^����"����g����Шu�Q!���1<:��:n
;�f3;-�>;�AD;֕F;�G;�H;UAH;jH;\�H;��H;(�H;ԻH;k�H;��H;B�H;��H;k�H;ԻH;(�H;��H;\�H;jH;UAH;�H;�G;֕F;�AD;-�>;�f3;n
;��:�1<:Q!��Шu������g��"�����&^�&����s潎K ��Z�f�i������k��'���;��TI�      ߛ7�v3��'����e� ��{Ծ
���6���]�F�����ӽ���;�L�1v�x뮼,T�Ƙ��PV�n�=�4(i:`��:!z ;�#5;�?;2�D;�F;�G;�H;�EH;�mH;��H;~�H;j�H;ۼH;4�H;P�H;��H;P�H;4�H;ۼH;j�H;~�H;��H;�mH;�EH;�H;�G;�F;2�D;�?;�#5;!z ;`��:4(i:n�=��PV�Ƙ�,T�x뮼1v�;�L�����ӽ���]�F�6���
����{Ծe� �����'�v3�      ����D��k�e� �<�ݾS���C͓�ȟf��>/�x��~'��n섽/�6�Rt��v��?�:�Tʻ�.�ݷ��s�:2; �$;�X7;��@;	E;:�F;Q�G;�H;EKH;�qH;��H;ɣH;�H;�H;.�H;D�H;��H;D�H;.�H;�H;�H;ɣH;��H;�qH;EKH;�H;Q�G;:�F;	E;��@;�X7; �$;2;�s�:ݷ��.�Tʻ?�:��v��Rt�/�6�n섽~'��x���>/�ȟf�C͓�S���<�ݾe� ��k��D�      e� ������쾻{ԾS���b���9�x�rSC��^�ͻ޽%���Q�e����ѼG������R�����դ8��:�X;��);5�9;.�A;��E;�G;2�G;s H;DRH;�vH;w�H;��H;:�H;��H;r�H;u�H;��H;u�H;r�H;��H;:�H;��H;w�H;�vH;DRH;s H;2�G;�G;��E;.�A;5�9;��);�X;��:դ8����R�����G���Ѽ��Q�e�%���ͻ޽�^�rSC�9�x�b���S����{Ծ�쾃���      {�˾��Ǿi���
���C͓�9�x�ؘJ��K �H��� �������?���t뮼�[�����3|��W��>�:w~�:';�
/;�f<;�C;� F;�MG;��G;:,H;sZH;�|H;ǖH;éH;��H;��H;��H;��H;��H;��H;��H;��H;��H;éH;ǖH;�|H;sZH;:,H;��G;�MG;� F;�C;�f<;�
/;';w~�:>�:�W��3|������[�t뮼����?���� ��H����K �ؘJ�9�x�C͓�
���i�����Ǿ      ��b���f�6���ȟf�rSC��K �Gn����Ž����Z��k��|ռX��Ey-����x.�t���O�:�*�:��;p4;s�>;)D;�vF;I�G;��G;�8H;\cH;x�H;��H;[�H;e�H;��H;��H;K�H;f�H;K�H;��H;��H;e�H;[�H;��H;x�H;\cH;�8H;��G;I�G;�vF;)D;s�>;p4;��;�*�:�O�:t��x.����Ey-�X���|ռ�k��Z������ŽGn���K �rSC�ȟf�6���f�b���      	�j�ȟf��Z�]�F��>/��^�H�����Ž- ���Fi�kQ+�Ot�PT��H�W�����1��hȺ�U�9�O�:	Y;��(;T�8;1A;�E;"�F;|�G;�H;�EH;�lH;��H;��H;8�H;d�H;��H;��H;��H;��H;��H;��H;��H;d�H;8�H;��H;��H;�lH;�EH;�H;|�G;"�F;�E;1A;T�8;��(;	Y;�O�:�U�9hȺ�1�����H�W�PT��Ot�kQ+��Fi�- ����ŽH����^��>/�]�F��Z�ȟf�      �!,� )��K ����x��ͻ޽ ������Fi���0�����跼z�x�����.��b�(�����)i:���:��;�0;��<;�C;��E;)<G;
�G;�#H;kSH;�vH;�H;�H;E�H;t�H;4�H;��H;��H;n�H;��H;��H;4�H;t�H;E�H;�H;�H;�vH;kSH;�#H;
�G;)<G;��E;�C;��<;�0;��;���:�)i:���b�(��.�����z�x��跼�����0��Fi���� ��ͻ޽x������K � )�      J��� ��s��ӽ~'��%�������Z�kQ+�����"��G����0���׻͕b��W���V�9�:�_;�)';0Y7;H#@;S�D;�F;+�G;��G;A7H;aH;��H;Z�H;��H;l�H;��H;��H;{�H;A�H;.�H;A�H;{�H;��H;��H;l�H;��H;Z�H;��H;aH;A7H;��G;+�G;�F;S�D;H#@;0Y7;�)';�_;�:�V�9�W��͕b���׻��0�G���"�����kQ+��Z����%���~'���ӽ�s� ��      0��W;��&������n섽Q�e���?��k�Ot��跼G��ee7�����Ǆ��0��t�_t�: +�:�
;�1;��<;��B;N�E;G;�G;iH;wIH;`nH;��H;��H;�H;��H;��H;�H;��H;�H;��H;�H;��H;�H;��H;��H;�H;��H;��H;`nH;wIH;iH;�G;G;N�E;��B;��<;�1;�
; +�:_t�:�t��0��Ǆ����ee7�G���跼Ot�k���?�Q�e�n섽���&���W;��      m��Fi��&^�;�L�/�6������|ռPT��z�x���0��������0���ڷ�zm`:��:��;��*;~�8;G�@;e�D;��F;}G;��G;�0H;�ZH;n{H;��H;֧H;�H;��H;��H;|�H;��H;��H;d�H;��H;��H;|�H;��H;��H;�H;֧H;��H;n{H;�ZH;�0H;��G;}G;��F;e�D;G�@;~�8;��*;��;��:zm`:�ڷ�0��������껢�0�z�x�PT���|ռ����/�6�;�L��&^��Fi�      ���k���1v�Rt��Ѽt뮼X��H�W������׻�Ǆ�0�����3<:w��:;Y;�s%;=$5;�Y>;.`C;��E;O)G;v�G;#H;GH;lkH;�H;��H;��H;ȻH;��H;��H;��H;g�H;_�H;�H;_�H;g�H;��H;��H;��H;ȻH;��H;��H;�H;lkH;GH;#H;v�G;O)G;��E;.`C;�Y>;=$5;�s%;;Y;w��:�3<:���0���Ǆ���׻���H�W�X��t뮼�ѼRt�1v����k�      ,˼x�Ǽ�"��x뮼�v��G���[�Ey-�����.��͕b��0㺅ڷ��3<:L�:_\;��!;2J2;�f<;/B;RBE;J�F;a�G; �G;�3H;�[H;{H;��H;��H;P�H;��H;6�H;��H;B�H;A�H;��H;��H;��H;A�H;B�H;��H;6�H;��H;P�H;��H;��H;{H;�[H;�3H; �G;a�G;J�F;RBE;/B;�f<;2J2;��!;_\;L�:�3<:�ڷ��0�͕b��.�����Ey-��[�G���v��x뮼�"��x�Ǽ      ��x��[t���g�,T�?�:������������1��b�(��W���t�zm`:w��:_\;pz ;�0;�;;9<A;?�D;�vF;�bG;e�G;� H;�LH;�nH;p�H;~�H;��H;��H;Z�H;��H;H�H;_�H;��H;��H;�H;��H;��H;_�H;H�H;��H;Z�H;��H;��H;~�H;p�H;�nH;�LH;� H;e�G;�bG;�vF;?�D;9<A;�;;�0;pz ;_\;w��:zm`:�t��W��b�(��1������������?�:�,T���g��[t�      E��8�	����Ƙ�Tʻ�R��3|�x.�hȺ����V�9_t�:��:;Y;��!;�0;.�:;�@;5BD;�1F;�7G;��G;�H;k?H;+cH;�H;n�H;;�H;<�H;>�H;��H;��H;��H;[�H;��H;��H;s�H;��H;��H;[�H;��H;��H;��H;>�H;<�H;;�H;n�H;�H;+cH;k?H;�H;��G;�7G;�1F;5BD;�@;.�:;�0;��!;;Y;��:_t�:�V�9���hȺx.�3|��R��TʻƘ����8�	�      �1��(Ȅ�Шu��PV��.�����W��t��U�9�)i:�: +�:��;�s%;2J2;�;;�@;�D;/F;?G;��G;�H;�4H;�YH;5wH;7�H;�H;	�H;�H;I�H;^�H;�H;�H;�H;*�H;E�H;��H;E�H;*�H;�H;�H;�H;^�H;I�H;�H;	�H;�H;7�H;5wH;�YH;�4H;�H;��G;?G;/F;�D;�@;�;;2J2;�s%;��; +�:�:�)i:�U�9t���W������.��PV�Шu�(Ȅ�      `���sX��Q!��n�=�ݷ�դ8>�:�O�:�O�:���:�_;�
;��*;=$5;�f<;9<A;5BD;/F;�G;��G;r�G;�,H;RH;UpH;�H;��H;r�H;�H;)�H;��H;��H;��H;?�H;��H;��H;|�H;��H;|�H;��H;��H;?�H;��H;��H;��H;)�H;�H;r�H;��H;�H;UpH;RH;�,H;r�G;��G;�G;/F;5BD;9<A;�f<;=$5;��*;�
;�_;���:�O�:�O�:>�:դ8ݷ�n�=�Q!��sX��      S�:џ:�1<:4(i:�s�:��:w~�:�*�:	Y;��;�)';�1;~�8;�Y>;/B;?�D;�1F;?G;��G;%�G;�(H;�MH;qkH;C�H;c�H;v�H;��H;�H;t�H;��H;$�H;�H;�H;D�H;��H;��H;��H;��H;��H;D�H;�H;�H;$�H;��H;t�H;�H;��H;v�H;c�H;C�H;qkH;�MH;�(H;%�G;��G;?G;�1F;?�D;/B;�Y>;~�8;�1;�)';��;	Y;�*�:w~�:��:�s�:4(i:�1<:џ:      g�:���:��:`��:2;�X;';��;��(;�0;0Y7;��<;G�@;.`C;RBE;�vF;�7G;��G;r�G;�(H;�KH;�hH;.�H;O�H;��H;��H;��H;O�H;�H;��H;��H;A�H;��H;��H;��H;��H;��H;��H;��H;��H;��H;A�H;��H;��H;�H;O�H;��H;��H;��H;O�H;.�H;�hH;�KH;�(H;r�G;��G;�7G;�vF;RBE;.`C;G�@;��<;0Y7;�0;��(;��;';�X;2;`��:��:���:      3;&�;n
;!z ; �$;��);�
/;p4;T�8;��<;H#@;��B;e�D;��E;J�F;�bG;��G;�H;�,H;�MH;�hH;B�H;��H;��H;ΰH;��H;��H;��H;2�H;��H;^�H;�H;0�H;��H;��H;P�H;��H;P�H;��H;��H;0�H;�H;^�H;��H;2�H;��H;��H;��H;ΰH;��H;��H;B�H;�hH;�MH;�,H;�H;��G;�bG;J�F;��E;e�D;��B;H#@;��<;T�8;p4;�
/;��); �$;!z ;n
;&�;      ��1;�I2;�f3;�#5;�X7;5�9;�f<;s�>;1A;�C;S�D;N�E;��F;O)G;a�G;e�G;�H;�4H;RH;qkH;.�H;��H;�H;ɯH;��H;V�H;L�H; �H;��H;��H;u�H;��H;o�H;��H;��H;�H;\�H;�H;��H;��H;o�H;��H;u�H;��H;��H; �H;L�H;V�H;��H;ɯH;�H;��H;.�H;qkH;RH;�4H;�H;e�G;a�G;O)G;��F;N�E;S�D;�C;1A;s�>;�f<;5�9;�X7;�#5;�f3;�I2;      n+>;�Y>;-�>;�?;��@;.�A;�C;)D;�E;��E;�F;G;}G;v�G; �G;� H;k?H;�YH;UpH;C�H;O�H;��H;ɯH;�H;��H;��H;6�H;��H;��H;��H;O�H; �H;��H;��H;H�H;��H;��H;��H;H�H;��H;��H; �H;O�H;��H;��H;��H;6�H;��H;��H;�H;ɯH;��H;O�H;C�H;UpH;�YH;k?H;� H; �G;v�G;}G;G;�F;��E;�E;)D;�C;.�A;��@;�?;-�>;�Y>;      ��C;qD;�AD;2�D;	E;��E;� F;�vF;"�F;)<G;+�G;�G;��G;#H;�3H;�LH;+cH;5wH;�H;c�H;��H;ΰH;��H;��H;=�H;��H;��H;^�H;c�H;��H;��H;g�H;��H;@�H;��H;D�H;L�H;D�H;��H;@�H;��H;g�H;��H;��H;c�H;^�H;��H;��H;=�H;��H;��H;ΰH;��H;c�H;�H;5wH;+cH;�LH;�3H;#H;��G;�G;+�G;)<G;"�F;�vF;� F;��E;	E;2�D;�AD;qD;      �vF;�~F;֕F;�F;:�F;�G;�MG;I�G;|�G;
�G;��G;iH;�0H;GH;�[H;�nH;�H;7�H;��H;v�H;��H;��H;V�H;��H;��H;W�H;$�H;�H;��H;��H;�H;S�H;6�H;��H;m�H;��H;��H;��H;m�H;��H;6�H;S�H;�H;��H;��H;�H;$�H;W�H;��H;��H;V�H;��H;��H;v�H;��H;7�H;�H;�nH;�[H;GH;�0H;iH;��G;
�G;|�G;I�G;�MG;�G;:�F;�F;֕F;�~F;      �G;\�G;�G;�G;Q�G;2�G;��G;��G;�H;�#H;A7H;wIH;�ZH;lkH;{H;p�H;n�H;�H;r�H;��H;��H;��H;L�H;6�H;��H;$�H;�H;h�H;J�H;��H;7�H;�H;��H;��H;��H;�H;�H;�H;��H;��H;��H;�H;7�H;��H;J�H;h�H;�H;$�H;��H;6�H;L�H;��H;��H;��H;r�H;�H;n�H;p�H;{H;lkH;�ZH;wIH;A7H;�#H;�H;��G;��G;2�G;Q�G;�G;�G;\�G;      ��G;+H;�H;�H;�H;s H;:,H;�8H;�EH;kSH;aH;`nH;n{H;�H;��H;~�H;;�H;	�H;�H;�H;O�H;��H; �H;��H;^�H;�H;h�H;]�H;��H;�H;�H;��H;z�H;��H;�H;^�H;g�H;^�H;�H;��H;z�H;��H;�H;�H;��H;]�H;h�H;�H;^�H;��H; �H;��H;O�H;�H;�H;	�H;;�H;~�H;��H;�H;n{H;`nH;aH;kSH;�EH;�8H;:,H;s H;�H;�H;�H;+H;      >H;�>H;UAH;�EH;EKH;DRH;sZH;\cH;�lH;�vH;��H;��H;��H;��H;��H;��H;<�H;�H;)�H;t�H;�H;2�H;��H;��H;c�H;��H;J�H;��H;$�H;��H;��H;k�H;��H;6�H;p�H;��H;��H;��H;p�H;6�H;��H;k�H;��H;��H;$�H;��H;J�H;��H;c�H;��H;��H;2�H;�H;t�H;)�H;�H;<�H;��H;��H;��H;��H;��H;��H;�vH;�lH;\cH;sZH;DRH;EKH;�EH;UAH;�>H;      �gH;�hH;jH;�mH;�qH;�vH;�|H;x�H;��H;�H;Z�H;��H;֧H;��H;P�H;��H;>�H;I�H;��H;��H;��H;��H;��H;��H;��H;��H;��H;�H;��H;��H;t�H;��H;%�H;y�H;��H;��H;��H;��H;��H;y�H;%�H;��H;t�H;��H;��H;�H;��H;��H;��H;��H;��H;��H;��H;��H;��H;I�H;>�H;��H;P�H;��H;֧H;��H;Z�H;�H;��H;x�H;�|H;�vH;�qH;�mH;jH;�hH;      Z�H;�H;\�H;��H;��H;w�H;ǖH;��H;��H;�H;��H;�H;�H;ȻH;��H;Z�H;��H;^�H;��H;$�H;��H;^�H;u�H;O�H;��H;�H;7�H;�H;��H;t�H;��H;.�H;��H;��H;��H;��H;��H;��H;��H;��H;��H;.�H;��H;t�H;��H;�H;7�H;�H;��H;O�H;u�H;^�H;��H;$�H;��H;^�H;��H;Z�H;��H;ȻH;�H;�H;��H;�H;��H;��H;ǖH;w�H;��H;��H;\�H;�H;      w�H;�H;��H;~�H;ɣH;��H;éH;[�H;8�H;E�H;l�H;��H;��H;��H;6�H;��H;��H;�H;��H;�H;A�H;�H;��H; �H;g�H;S�H;�H;��H;k�H;��H;.�H;{�H;��H;��H;��H;�H;�H;�H;��H;��H;��H;{�H;.�H;��H;k�H;��H;�H;S�H;g�H; �H;��H;�H;A�H;�H;��H;�H;��H;��H;6�H;��H;��H;��H;l�H;E�H;8�H;[�H;éH;��H;ɣH;~�H;��H;�H;      9�H;r�H;(�H;j�H;�H;:�H;��H;e�H;d�H;t�H;��H;��H;��H;��H;��H;H�H;��H;�H;?�H;�H;��H;0�H;o�H;��H;��H;6�H;��H;z�H;��H;%�H;��H;��H;��H;��H;�H;�H;�H;�H;�H;��H;��H;��H;��H;%�H;��H;z�H;��H;6�H;��H;��H;o�H;0�H;��H;�H;?�H;�H;��H;H�H;��H;��H;��H;��H;��H;t�H;d�H;e�H;��H;:�H;�H;j�H;(�H;r�H;      �H;7�H;ԻH;ۼH;�H;��H;��H;��H;��H;4�H;��H;�H;|�H;��H;B�H;_�H;[�H;�H;��H;D�H;��H;��H;��H;��H;@�H;��H;��H;��H;6�H;y�H;��H;��H;��H; �H;.�H;9�H;�H;9�H;.�H; �H;��H;��H;��H;y�H;6�H;��H;��H;��H;@�H;��H;��H;��H;��H;D�H;��H;�H;[�H;_�H;B�H;��H;|�H;�H;��H;4�H;��H;��H;��H;��H;�H;ۼH;ԻH;7�H;      ��H;��H;k�H;4�H;.�H;r�H;��H;��H;��H;��H;{�H;��H;��H;g�H;A�H;��H;��H;*�H;��H;��H;��H;��H;��H;H�H;��H;m�H;��H;�H;p�H;��H;��H;��H;�H;.�H;�H;-�H;J�H;-�H;�H;.�H;�H;��H;��H;��H;p�H;�H;��H;m�H;��H;H�H;��H;��H;��H;��H;��H;*�H;��H;��H;A�H;g�H;��H;��H;{�H;��H;��H;��H;��H;r�H;.�H;4�H;k�H;��H;      (�H;S�H;��H;P�H;D�H;u�H;��H;K�H;��H;��H;A�H;�H;��H;_�H;��H;��H;��H;E�H;|�H;��H;��H;P�H;�H;��H;D�H;��H;�H;^�H;��H;��H;��H;�H;�H;9�H;-�H;$�H;6�H;$�H;-�H;9�H;�H;�H;��H;��H;��H;^�H;�H;��H;D�H;��H;�H;P�H;��H;��H;|�H;E�H;��H;��H;��H;_�H;��H;�H;A�H;��H;��H;K�H;��H;u�H;D�H;P�H;��H;S�H;      ��H;��H;B�H;��H;��H;��H;��H;f�H;��H;n�H;.�H;��H;d�H;�H;��H;�H;s�H;��H;��H;��H;��H;��H;\�H;��H;L�H;��H;�H;g�H;��H;��H;��H;�H;�H;�H;J�H;6�H;#�H;6�H;J�H;�H;�H;�H;��H;��H;��H;g�H;�H;��H;L�H;��H;\�H;��H;��H;��H;��H;��H;s�H;�H;��H;�H;d�H;��H;.�H;n�H;��H;f�H;��H;��H;��H;��H;B�H;��H;      (�H;S�H;��H;P�H;D�H;u�H;��H;K�H;��H;��H;A�H;�H;��H;_�H;��H;��H;��H;E�H;|�H;��H;��H;P�H;�H;��H;D�H;��H;�H;^�H;��H;��H;��H;�H;�H;9�H;-�H;$�H;6�H;$�H;-�H;9�H;�H;�H;��H;��H;��H;^�H;�H;��H;D�H;��H;�H;P�H;��H;��H;|�H;E�H;��H;��H;��H;_�H;��H;�H;A�H;��H;��H;K�H;��H;u�H;D�H;P�H;��H;S�H;      ��H;��H;k�H;4�H;.�H;r�H;��H;��H;��H;��H;{�H;��H;��H;g�H;A�H;��H;��H;*�H;��H;��H;��H;��H;��H;H�H;��H;m�H;��H;�H;p�H;��H;��H;��H;�H;.�H;�H;-�H;J�H;-�H;�H;.�H;�H;��H;��H;��H;p�H;�H;��H;m�H;��H;H�H;��H;��H;��H;��H;��H;*�H;��H;��H;A�H;g�H;��H;��H;{�H;��H;��H;��H;��H;r�H;.�H;4�H;k�H;��H;      �H;7�H;ԻH;ۼH;�H;��H;��H;��H;��H;4�H;��H;�H;|�H;��H;B�H;_�H;[�H;�H;��H;D�H;��H;��H;��H;��H;@�H;��H;��H;��H;6�H;y�H;��H;��H;��H; �H;.�H;9�H;�H;9�H;.�H; �H;��H;��H;��H;y�H;6�H;��H;��H;��H;@�H;��H;��H;��H;��H;D�H;��H;�H;[�H;_�H;B�H;��H;|�H;�H;��H;4�H;��H;��H;��H;��H;�H;ۼH;ԻH;7�H;      9�H;r�H;(�H;j�H;�H;:�H;��H;e�H;d�H;t�H;��H;��H;��H;��H;��H;H�H;��H;�H;?�H;�H;��H;0�H;o�H;��H;��H;6�H;��H;z�H;��H;%�H;��H;��H;��H;��H;�H;�H;�H;�H;�H;��H;��H;��H;��H;%�H;��H;z�H;��H;6�H;��H;��H;o�H;0�H;��H;�H;?�H;�H;��H;H�H;��H;��H;��H;��H;��H;t�H;d�H;e�H;��H;:�H;�H;j�H;(�H;r�H;      w�H;�H;��H;~�H;ɣH;��H;éH;[�H;8�H;E�H;l�H;��H;��H;��H;6�H;��H;��H;�H;��H;�H;A�H;�H;��H; �H;g�H;S�H;�H;��H;k�H;��H;.�H;{�H;��H;��H;��H;�H;�H;�H;��H;��H;��H;{�H;.�H;��H;k�H;��H;�H;S�H;g�H; �H;��H;�H;A�H;�H;��H;�H;��H;��H;6�H;��H;��H;��H;l�H;E�H;8�H;[�H;éH;��H;ɣH;~�H;��H;�H;      Z�H;�H;\�H;��H;��H;w�H;ǖH;��H;��H;�H;��H;�H;�H;ȻH;��H;Z�H;��H;^�H;��H;$�H;��H;^�H;u�H;O�H;��H;�H;7�H;�H;��H;t�H;��H;.�H;��H;��H;��H;��H;��H;��H;��H;��H;��H;.�H;��H;t�H;��H;�H;7�H;�H;��H;O�H;u�H;^�H;��H;$�H;��H;^�H;��H;Z�H;��H;ȻH;�H;�H;��H;�H;��H;��H;ǖH;w�H;��H;��H;\�H;�H;      �gH;�hH;jH;�mH;�qH;�vH;�|H;x�H;��H;�H;Z�H;��H;֧H;��H;P�H;��H;>�H;I�H;��H;��H;��H;��H;��H;��H;��H;��H;��H;�H;��H;��H;t�H;��H;%�H;y�H;��H;��H;��H;��H;��H;y�H;%�H;��H;t�H;��H;��H;�H;��H;��H;��H;��H;��H;��H;��H;��H;��H;I�H;>�H;��H;P�H;��H;֧H;��H;Z�H;�H;��H;x�H;�|H;�vH;�qH;�mH;jH;�hH;      >H;�>H;UAH;�EH;EKH;DRH;sZH;\cH;�lH;�vH;��H;��H;��H;��H;��H;��H;<�H;�H;)�H;t�H;�H;2�H;��H;��H;c�H;��H;J�H;��H;$�H;��H;��H;k�H;��H;6�H;p�H;��H;��H;��H;p�H;6�H;��H;k�H;��H;��H;$�H;��H;J�H;��H;c�H;��H;��H;2�H;�H;t�H;)�H;�H;<�H;��H;��H;��H;��H;��H;��H;�vH;�lH;\cH;sZH;DRH;EKH;�EH;UAH;�>H;      ��G;+H;�H;�H;�H;s H;:,H;�8H;�EH;kSH;aH;`nH;n{H;�H;��H;~�H;;�H;	�H;�H;�H;O�H;��H; �H;��H;^�H;�H;h�H;]�H;��H;�H;�H;��H;z�H;��H;�H;^�H;g�H;^�H;�H;��H;z�H;��H;�H;�H;��H;]�H;h�H;�H;^�H;��H; �H;��H;O�H;�H;�H;	�H;;�H;~�H;��H;�H;n{H;`nH;aH;kSH;�EH;�8H;:,H;s H;�H;�H;�H;+H;      �G;\�G;�G;�G;Q�G;2�G;��G;��G;�H;�#H;A7H;wIH;�ZH;lkH;{H;p�H;n�H;�H;r�H;��H;��H;��H;L�H;6�H;��H;$�H;�H;h�H;J�H;��H;7�H;�H;��H;��H;��H;�H;�H;�H;��H;��H;��H;�H;7�H;��H;J�H;h�H;�H;$�H;��H;6�H;L�H;��H;��H;��H;r�H;�H;n�H;p�H;{H;lkH;�ZH;wIH;A7H;�#H;�H;��G;��G;2�G;Q�G;�G;�G;\�G;      �vF;�~F;֕F;�F;:�F;�G;�MG;I�G;|�G;
�G;��G;iH;�0H;GH;�[H;�nH;�H;7�H;��H;v�H;��H;��H;V�H;��H;��H;W�H;$�H;�H;��H;��H;�H;S�H;6�H;��H;m�H;��H;��H;��H;m�H;��H;6�H;S�H;�H;��H;��H;�H;$�H;W�H;��H;��H;V�H;��H;��H;v�H;��H;7�H;�H;�nH;�[H;GH;�0H;iH;��G;
�G;|�G;I�G;�MG;�G;:�F;�F;֕F;�~F;      ��C;qD;�AD;2�D;	E;��E;� F;�vF;"�F;)<G;+�G;�G;��G;#H;�3H;�LH;+cH;5wH;�H;c�H;��H;ΰH;��H;��H;=�H;��H;��H;^�H;c�H;��H;��H;g�H;��H;@�H;��H;D�H;L�H;D�H;��H;@�H;��H;g�H;��H;��H;c�H;^�H;��H;��H;=�H;��H;��H;ΰH;��H;c�H;�H;5wH;+cH;�LH;�3H;#H;��G;�G;+�G;)<G;"�F;�vF;� F;��E;	E;2�D;�AD;qD;      n+>;�Y>;-�>;�?;��@;.�A;�C;)D;�E;��E;�F;G;}G;v�G; �G;� H;k?H;�YH;UpH;C�H;O�H;��H;ɯH;�H;��H;��H;6�H;��H;��H;��H;O�H; �H;��H;��H;H�H;��H;��H;��H;H�H;��H;��H; �H;O�H;��H;��H;��H;6�H;��H;��H;�H;ɯH;��H;O�H;C�H;UpH;�YH;k?H;� H; �G;v�G;}G;G;�F;��E;�E;)D;�C;.�A;��@;�?;-�>;�Y>;      ��1;�I2;�f3;�#5;�X7;5�9;�f<;s�>;1A;�C;S�D;N�E;��F;O)G;a�G;e�G;�H;�4H;RH;qkH;.�H;��H;�H;ɯH;��H;V�H;L�H; �H;��H;��H;u�H;��H;o�H;��H;��H;�H;\�H;�H;��H;��H;o�H;��H;u�H;��H;��H; �H;L�H;V�H;��H;ɯH;�H;��H;.�H;qkH;RH;�4H;�H;e�G;a�G;O)G;��F;N�E;S�D;�C;1A;s�>;�f<;5�9;�X7;�#5;�f3;�I2;      3;&�;n
;!z ; �$;��);�
/;p4;T�8;��<;H#@;��B;e�D;��E;J�F;�bG;��G;�H;�,H;�MH;�hH;B�H;��H;��H;ΰH;��H;��H;��H;2�H;��H;^�H;�H;0�H;��H;��H;P�H;��H;P�H;��H;��H;0�H;�H;^�H;��H;2�H;��H;��H;��H;ΰH;��H;��H;B�H;�hH;�MH;�,H;�H;��G;�bG;J�F;��E;e�D;��B;H#@;��<;T�8;p4;�
/;��); �$;!z ;n
;&�;      g�:���:��:`��:2;�X;';��;��(;�0;0Y7;��<;G�@;.`C;RBE;�vF;�7G;��G;r�G;�(H;�KH;�hH;.�H;O�H;��H;��H;��H;O�H;�H;��H;��H;A�H;��H;��H;��H;��H;��H;��H;��H;��H;��H;A�H;��H;��H;�H;O�H;��H;��H;��H;O�H;.�H;�hH;�KH;�(H;r�G;��G;�7G;�vF;RBE;.`C;G�@;��<;0Y7;�0;��(;��;';�X;2;`��:��:���:      S�:џ:�1<:4(i:�s�:��:w~�:�*�:	Y;��;�)';�1;~�8;�Y>;/B;?�D;�1F;?G;��G;%�G;�(H;�MH;qkH;C�H;c�H;v�H;��H;�H;t�H;��H;$�H;�H;�H;D�H;��H;��H;��H;��H;��H;D�H;�H;�H;$�H;��H;t�H;�H;��H;v�H;c�H;C�H;qkH;�MH;�(H;%�G;��G;?G;�1F;?�D;/B;�Y>;~�8;�1;�)';��;	Y;�*�:w~�:��:�s�:4(i:�1<:џ:      `���sX��Q!��n�=�ݷ�դ8>�:�O�:�O�:���:�_;�
;��*;=$5;�f<;9<A;5BD;/F;�G;��G;r�G;�,H;RH;UpH;�H;��H;r�H;�H;)�H;��H;��H;��H;?�H;��H;��H;|�H;��H;|�H;��H;��H;?�H;��H;��H;��H;)�H;�H;r�H;��H;�H;UpH;RH;�,H;r�G;��G;�G;/F;5BD;9<A;�f<;=$5;��*;�
;�_;���:�O�:�O�:>�:դ8ݷ�n�=�Q!��sX��      �1��(Ȅ�Шu��PV��.�����W��t��U�9�)i:�: +�:��;�s%;2J2;�;;�@;�D;/F;?G;��G;�H;�4H;�YH;5wH;7�H;�H;	�H;�H;I�H;^�H;�H;�H;�H;*�H;E�H;��H;E�H;*�H;�H;�H;�H;^�H;I�H;�H;	�H;�H;7�H;5wH;�YH;�4H;�H;��G;?G;/F;�D;�@;�;;2J2;�s%;��; +�:�:�)i:�U�9t���W������.��PV�Шu�(Ȅ�      E��8�	����Ƙ�Tʻ�R��3|�x.�hȺ����V�9_t�:��:;Y;��!;�0;.�:;�@;5BD;�1F;�7G;��G;�H;k?H;+cH;�H;n�H;;�H;<�H;>�H;��H;��H;��H;[�H;��H;��H;s�H;��H;��H;[�H;��H;��H;��H;>�H;<�H;;�H;n�H;�H;+cH;k?H;�H;��G;�7G;�1F;5BD;�@;.�:;�0;��!;;Y;��:_t�:�V�9���hȺx.�3|��R��TʻƘ����8�	�      ��x��[t���g�,T�?�:������������1��b�(��W���t�zm`:w��:_\;pz ;�0;�;;9<A;?�D;�vF;�bG;e�G;� H;�LH;�nH;p�H;~�H;��H;��H;Z�H;��H;H�H;_�H;��H;��H;�H;��H;��H;_�H;H�H;��H;Z�H;��H;��H;~�H;p�H;�nH;�LH;� H;e�G;�bG;�vF;?�D;9<A;�;;�0;pz ;_\;w��:zm`:�t��W��b�(��1������������?�:�,T���g��[t�      ,˼x�Ǽ�"��x뮼�v��G���[�Ey-�����.��͕b��0㺅ڷ��3<:L�:_\;��!;2J2;�f<;/B;RBE;J�F;a�G; �G;�3H;�[H;{H;��H;��H;P�H;��H;6�H;��H;B�H;A�H;��H;��H;��H;A�H;B�H;��H;6�H;��H;P�H;��H;��H;{H;�[H;�3H; �G;a�G;J�F;RBE;/B;�f<;2J2;��!;_\;L�:�3<:�ڷ��0�͕b��.�����Ey-��[�G���v��x뮼�"��x�Ǽ      ���k���1v�Rt��Ѽt뮼X��H�W������׻�Ǆ�0�����3<:w��:;Y;�s%;=$5;�Y>;.`C;��E;O)G;v�G;#H;GH;lkH;�H;��H;��H;ȻH;��H;��H;��H;g�H;_�H;�H;_�H;g�H;��H;��H;��H;ȻH;��H;��H;�H;lkH;GH;#H;v�G;O)G;��E;.`C;�Y>;=$5;�s%;;Y;w��:�3<:���0���Ǆ���׻���H�W�X��t뮼�ѼRt�1v����k�      m��Fi��&^�;�L�/�6������|ռPT��z�x���0��������0���ڷ�zm`:��:��;��*;~�8;G�@;e�D;��F;}G;��G;�0H;�ZH;n{H;��H;֧H;�H;��H;��H;|�H;��H;��H;d�H;��H;��H;|�H;��H;��H;�H;֧H;��H;n{H;�ZH;�0H;��G;}G;��F;e�D;G�@;~�8;��*;��;��:zm`:�ڷ�0��������껢�0�z�x�PT���|ռ����/�6�;�L��&^��Fi�      0��W;��&������n섽Q�e���?��k�Ot��跼G��ee7�����Ǆ��0��t�_t�: +�:�
;�1;��<;��B;N�E;G;�G;iH;wIH;`nH;��H;��H;�H;��H;��H;�H;��H;�H;��H;�H;��H;�H;��H;��H;�H;��H;��H;`nH;wIH;iH;�G;G;N�E;��B;��<;�1;�
; +�:_t�:�t��0��Ǆ����ee7�G���跼Ot�k���?�Q�e�n섽���&���W;��      J��� ��s��ӽ~'��%�������Z�kQ+�����"��G����0���׻͕b��W���V�9�:�_;�)';0Y7;H#@;S�D;�F;+�G;��G;A7H;aH;��H;Z�H;��H;l�H;��H;��H;{�H;A�H;.�H;A�H;{�H;��H;��H;l�H;��H;Z�H;��H;aH;A7H;��G;+�G;�F;S�D;H#@;0Y7;�)';�_;�:�V�9�W��͕b���׻��0�G���"�����kQ+��Z����%���~'���ӽ�s� ��      �!,� )��K ����x��ͻ޽ ������Fi���0�����跼z�x�����.��b�(�����)i:���:��;�0;��<;�C;��E;)<G;
�G;�#H;kSH;�vH;�H;�H;E�H;t�H;4�H;��H;��H;n�H;��H;��H;4�H;t�H;E�H;�H;�H;�vH;kSH;�#H;
�G;)<G;��E;�C;��<;�0;��;���:�)i:���b�(��.�����z�x��跼�����0��Fi���� ��ͻ޽x������K � )�      	�j�ȟf��Z�]�F��>/��^�H�����Ž- ���Fi�kQ+�Ot�PT��H�W�����1��hȺ�U�9�O�:	Y;��(;T�8;1A;�E;"�F;|�G;�H;�EH;�lH;��H;��H;8�H;d�H;��H;��H;��H;��H;��H;��H;��H;d�H;8�H;��H;��H;�lH;�EH;�H;|�G;"�F;�E;1A;T�8;��(;	Y;�O�:�U�9hȺ�1�����H�W�PT��Ot�kQ+��Fi�- ����ŽH����^��>/�]�F��Z�ȟf�      ��b���f�6���ȟf�rSC��K �Gn����Ž����Z��k��|ռX��Ey-����x.�t���O�:�*�:��;p4;s�>;)D;�vF;I�G;��G;�8H;\cH;x�H;��H;[�H;e�H;��H;��H;K�H;f�H;K�H;��H;��H;e�H;[�H;��H;x�H;\cH;�8H;��G;I�G;�vF;)D;s�>;p4;��;�*�:�O�:t��x.����Ey-�X���|ռ�k��Z������ŽGn���K �rSC�ȟf�6���f�b���      {�˾��Ǿi���
���C͓�9�x�ؘJ��K �H��� �������?���t뮼�[�����3|��W��>�:w~�:';�
/;�f<;�C;� F;�MG;��G;:,H;sZH;�|H;ǖH;éH;��H;��H;��H;��H;��H;��H;��H;��H;��H;éH;ǖH;�|H;sZH;:,H;��G;�MG;� F;�C;�f<;�
/;';w~�:>�:�W��3|������[�t뮼����?���� ��H����K �ؘJ�9�x�C͓�
���i�����Ǿ      e� ������쾻{ԾS���b���9�x�rSC��^�ͻ޽%���Q�e����ѼG������R�����դ8��:�X;��);5�9;.�A;��E;�G;2�G;s H;DRH;�vH;w�H;��H;:�H;��H;r�H;u�H;��H;u�H;r�H;��H;:�H;��H;w�H;�vH;DRH;s H;2�G;�G;��E;.�A;5�9;��);�X;��:դ8����R�����G���Ѽ��Q�e�%���ͻ޽�^�rSC�9�x�b���S����{Ծ�쾃���      ����D��k�e� �<�ݾS���C͓�ȟf��>/�x��~'��n섽/�6�Rt��v��?�:�Tʻ�.�ݷ��s�:2; �$;�X7;��@;	E;:�F;Q�G;�H;EKH;�qH;��H;ɣH;�H;�H;.�H;D�H;��H;D�H;.�H;�H;�H;ɣH;��H;�qH;EKH;�H;Q�G;:�F;	E;��@;�X7; �$;2;�s�:ݷ��.�Tʻ?�:��v��Rt�/�6�n섽~'��x���>/�ȟf�C͓�S���<�ݾe� ��k��D�      ߛ7�v3��'����e� ��{Ծ
���6���]�F�����ӽ���;�L�1v�x뮼,T�Ƙ��PV�n�=�4(i:`��:!z ;�#5;�?;2�D;�F;�G;�H;�EH;�mH;��H;~�H;j�H;ۼH;4�H;P�H;��H;P�H;4�H;ۼH;j�H;~�H;��H;�mH;�EH;�H;�G;�F;2�D;�?;�#5;!z ;`��:4(i:n�=��PV�Ƙ�,T�x뮼1v�;�L�����ӽ���]�F�6���
����{Ծe� �����'�v3�      tN��TI���;��'��k���i���f󐾖Z��K ��s�&����&^����"����g����Шu�Q!���1<:��:n
;�f3;-�>;�AD;֕F;�G;�H;UAH;jH;\�H;��H;(�H;ԻH;k�H;��H;B�H;��H;k�H;ԻH;(�H;��H;\�H;jH;UAH;�H;�G;֕F;�AD;-�>;�f3;n
;��:�1<:Q!��Шu������g��"�����&^�&����s潎K ��Z�f�i������k��'���;��TI�      I]�N�W��TI�v3��D�������Ǿb���ȟf� )� ��W;���Fi��k�x�Ǽ�[t�8�	�(Ȅ�sX��џ:���:&�;�I2;�Y>;qD;�~F;\�G;+H;�>H;�hH;�H;�H;r�H;7�H;��H;S�H;��H;S�H;��H;7�H;r�H;�H;�H;�hH;�>H;+H;\�G;�~F;qD;�Y>;�I2;&�;���:џ:sX��(Ȅ�8�	��[t�x�Ǽ�k��Fi�W;�� �� )�ȟf�b�����Ǿ�����D�v3��TI�N�W�      �$��� ���������þ�*��
Dx�}�=����\Pν鰒��&K�xc����;�V�s���D^���S��v[:���:�d;��4;�_?;�lD;��F;puG;M�G;�H;�NH;�rH;�H;��H;��H;�H;q�H;E�H;q�H;�H;��H;��H;�H;�rH;�NH;�H;M�G;puG;��F;�lD;�_?;��4;�d;���:�v[:��S��D^�s��;�V����xc��&K�鰒�\Pν���}�=�
Dx��*���þ��������� �      �� �k��>��=���������0���s���:�N9���ʽZ����G��8��-��z5S�v���/X���D��Ad:�A�:� ;y�4;	�?;#~D;q�F;3xG;��G;�H;NOH;IsH;:�H;�H;�H;W�H;��H;U�H;��H;W�H;�H;�H;:�H;IsH;NOH;�H;��G;3xG;q�F;#~D;	�?;y�4;� ;�A�:�Ad:��D��/X�v��z5S��-���8���G�Z����ʽN9���:��s��0��������=��>��k��      ���>��&�
�����fYؾ���ȥ����f���0�C[�*8������ȟ>�|���#Ȥ�Y6H�,�ܻ�qF�.��6�}:���:�";��5;6�?;��D;��F;/�G;��G;s"H;�QH;�tH;z�H;�H;��H;�H;�H;��H;�H;�H;��H;�H;z�H;�tH;�QH;s"H;��G;/�G;��F;��D;6�?;��5;�";���:6�}:.���qF�,�ܻY6H�#Ȥ�|���ȟ>�����*8��C[���0���f�ȥ�����fYؾ����&�
�>��      ��=������I��þ�R��&���QS��Q"��s�����}��0���d���x�6��ƻ'}*����_�:�w;�%;Rl7;�@;�D;�F;��G;��G;3'H;UH;�wH;�H;f�H;ñH;ۺH;�H;��H;�H;ۺH;ñH;f�H;�H;�wH;UH;3'H;��G;��G;�F;�D;�@;Rl7;�%;�w;_�:���'}*��ƻx�6�d����켟0���}�����s��Q"�QS�&����R���þIᾁ���=��      ����fYؾ�þ�ê�f쏾jk���:�e�R�ؽ�����c�:y���Ҽݫ��� �B�'����'7��:�
;d�(;�^9;��A;�[E;��F;�G;��G;�-H;�YH;{H;�H;i�H;u�H;6�H;�H;��H;�H;6�H;u�H;i�H;�H;{H;�YH;�-H;��G;�G;��F;�[E;��A;�^9;d�(;�
;��:��'7'��B�� �ݫ����Ҽ:y��c�����R�ؽe���:�jk�f쏾�ê��þfYؾ��      �þ��������R��f쏾�s��H����������������D�vc�g����f�3,�����P����90��:6;�i-;��;;��B;+�E;�G;��G;��G;�5H;�_H;�H;{�H;��H;r�H;ɽH;r�H;��H;r�H;ɽH;r�H;��H;{�H;�H;�_H;�5H;��G;��G;�G;+�E;��B;��;;�i-;6;0��:��9�P�����3,��f�g���vc���D���������������H��s�f쏾�R���������      �*���0��ȥ��&���jk��H��#%�B[�ZPν�s��0�f�/%�d��`���G�=�n?ػgFL��D�c�R:C�:��;�2;�=;��C;�/F;�FG;�G;WH;?H;�fH;��H;V�H;ͫH;��H;��H;�H;��H;�H;��H;��H;ͫH;V�H;��H;�fH;?H;WH;�G;�FG;�/F;��C;�=;�2;��;C�:c�R:�D�gFL�n?ػG�=�`���d��/%�0�f��s��ZPνB[��#%��H�jk�&���ȥ���0��      
Dx��s���f�QS���:����B[��7ս�榽��}�u�;��8�)�����r����G������Ҭ����:��;}$;,�6;f�?;3�D;�F; pG;��G;H;XIH;dnH;i�H;��H;�H;[�H;��H;��H;G�H;��H;��H;[�H;�H;��H;i�H;dnH;XIH;H;��G; pG;�F;3�D;f�?;,�6;}$;��;���:�Ҭ����G�������r�)����8�u�;���}��榽�7սB[������:�QS���f��s�      }�=���:���0��Q"�e�����ZPν�榽%����G�����Ҽ���E:�	�ܻ�D^�θ��kh:���:P;�{,;�:;��A;~hE;��F;]�G;��G;�'H;eTH;�vH;��H;L�H;��H;�H;��H;��H;4�H;��H;��H;�H;��H;L�H;��H;�vH;eTH;�'H;��G;]�G;��F;~hE;��A;�:;�{,;P;���:kh:θ���D^�	�ܻE:������Ҽ����G�%���榽ZPν����e��Q"���0���:�      ���N9�C[��s�R�ؽ���s����}���G��K��	c��!�V�$,��*�����"����:@��:� ;ǂ3;0>;�C;#F;$8G;l�G;�H;7H;�_H;,H;�H; �H;g�H;�H;m�H;��H;3�H;��H;m�H;�H;g�H; �H;�H;,H;�_H;7H;�H;l�G;$8G;#F;�C;0>;ǂ3;� ;@��:��:"������*��$,�!�V�	c��K�����G���}��s����R�ؽ�s�C[�N9�      \Pν��ʽ*8�������������0�f�u�;���K��Ȥ���f���#ߵ�>o5�2�D�N�-:���:X>;H+;_9;�A;��D;[�F;�uG;�G;IH;�FH;�kH;�H;��H;�H;H�H;�H;��H;"�H;F�H;"�H;��H;�H;H�H;�H;��H;�H;�kH;�FH;IH;�G;�uG;[�F;��D;�A;_9;H+;X>;���:N�-:2�D�>o5�#ߵ�����f�Ȥ�K����u�;�0�f������������*8����ʽ      鰒�Z��������}��c���D�/%��8���Ҽ	c����f�����ƻY/X�t������9g�:ȏ;G";�3;�>;�XC;��E;G;'�G;��G;�+H;/VH;9wH;��H;W�H;�H;.�H;�H;Q�H;`�H;O�H;`�H;Q�H;�H;.�H;�H;W�H;��H;9wH;/VH;�+H;��G;'�G;G;��E;�XC;�>;�3;G";ȏ;g�:���9t���Y/X��ƻ�����f�	c����Ҽ�8�/%���D��c���}�����Z��      �&K���G�ȟ>��0�:y�vc�d��)������!�V����ƻfod���º>Q(7�3�:���: �;^P.;:�:;ayA;y�D;�F;�mG;u�G;!H;�?H;MeH;��H;R�H;ժH;��H;�H;
�H;��H;��H;V�H;��H;��H;
�H;�H;��H;ժH;R�H;��H;MeH;�?H;!H;u�G;�mG;�F;y�D;ayA;:�:;^P.; �;���:�3�:>Q(7��ºfod��ƻ��!�V����)���d��vc�:y��0�ȟ>���G�      xc��8�|����켔�Ҽg���`�����r�E:�$,�#ߵ�Y/X���º�ˬ�G�}:? �:v;��);�l7;i�?;�C;KF;�(G;F�G;��G;2)H;�RH;�sH;��H;��H;�H;ͼH;��H;��H;,�H;��H;l�H;��H;,�H;��H;��H;ͼH;�H;��H;��H;�sH;�RH;2)H;��G;F�G;�(G;KF;�C;i�?;�l7;��);v;? �:G�}:�ˬ���ºY/X�#ߵ�$,�E:���r�`���g�����Ҽ��|����8�      ����-��#Ȥ�d���ݫ���f�G�=����	�ܻ�*��>o5�t���>Q(7G�}:�m�:��;>&;��4;C�=;�B;,�E;S�F;ˀG;$�G;cH;�@H;�dH;d�H;��H;x�H;��H;��H;;�H;��H;��H;��H;l�H;��H;��H;��H;;�H;��H;��H;x�H;��H;d�H;�dH;�@H;cH;$�G;ˀG;S�F;,�E;�B;C�=;��4;>&;��;�m�:G�}:>Q(7t���>o5��*��	�ܻ���G�=��f�ݫ��d���#Ȥ��-��      ;�V�z5S�Y6H�x�6�� �3,�n?ػG���D^����2�D����9�3�:? �:��;^%;��3;p�<;�B;�
E;?�F;�WG;8�G;t�G;�/H;xVH;�uH;�H;��H;ܰH;��H;��H;��H;k�H;��H;��H;Q�H;��H;��H;k�H;��H;��H;��H;ܰH;��H;�H;�uH;xVH;�/H;t�G;8�G;�WG;?�F;�
E;�B;p�<;��3;^%;��;? �:�3�:���92�D�����D^�G��n?ػ3,�� �x�6�Y6H�z5S�      s��v��,�ܻ�ƻB󩻜��gFL����θ��"��N�-:g�:���:v;>&;��3;�8<;`�A;%�D;�YF;Z4G;3�G;�G;� H;aIH;VjH;ńH;ٙH;��H;��H;�H;��H;��H;��H;��H;v�H;�H;v�H;��H;��H;��H;��H;�H;��H;��H;ٙH;ńH;VjH;aIH;� H;�G;3�G;Z4G;�YF;%�D;`�A;�8<;��3;>&;v;���:g�:N�-:"��θ�����gFL����B��ƻ,�ܻv��      �D^��/X��qF�'}*�'���P���D��Ҭ�kh:��:���:ȏ; �;��);��4;p�<;`�A;f�D;�8F;
G;��G;w�G;jH;C>H;�`H;5|H;��H;��H;��H;��H;��H;}�H;��H;4�H;��H;8�H;��H;8�H;��H;4�H;��H;}�H;��H;��H;��H;��H;��H;5|H;�`H;C>H;jH;w�G;��G;
G;�8F;f�D;`�A;p�<;��4;��); �;ȏ;���:��:kh:�Ҭ��D��P��'��'}*��qF��/X�      ��S���D�.�������'7��9c�R:���:���:@��:X>;G";^P.;�l7;C�=;�B;%�D;�8F;YG;R�G;��G;�H;�5H;�XH;	uH;=�H;�H;�H;�H;��H;9�H;��H;-�H;M�H;r�H;��H;�H;��H;r�H;M�H;-�H;��H;9�H;��H;�H;�H;�H;=�H;	uH;�XH;�5H;�H;��G;R�G;YG;�8F;%�D;�B;C�=;�l7;^P.;G";X>;@��:���:���:c�R:��9��'7���.����D�      �v[:�Ad:6�}:_�:��:0��:C�:��;P;� ;H+;�3;:�:;i�?;�B;�
E;�YF;
G;R�G;��G;nH;�0H;�RH;�oH;�H;f�H;�H;��H;��H;��H;�H;��H;��H;5�H;�H;(�H;q�H;(�H;�H;5�H;��H;��H;�H;��H;��H;��H;�H;f�H;�H;�oH;�RH;�0H;nH;��G;R�G;
G;�YF;�
E;�B;i�?;:�:;�3;H+;� ;P;��;C�:0��:��:_�:6�}:�Ad:      ���:�A�:���:�w;�
;6;��;}$;�{,;ǂ3;_9;�>;ayA;�C;,�E;?�F;Z4G;��G;��G;nH;�.H;PH;'lH;i�H;��H;��H;��H;�H;��H;)�H;r�H;��H;��H;��H;z�H;W�H;��H;W�H;z�H;��H;��H;��H;r�H;)�H;��H;�H;��H;��H;��H;i�H;'lH;PH;�.H;nH;��G;��G;Z4G;?�F;,�E;�C;ayA;�>;_9;ǂ3;�{,;}$;��;6;�
;�w;���:�A�:      �d;� ;�";�%;d�(;�i-;�2;,�6;�:;0>;�A;�XC;y�D;KF;S�F;�WG;3�G;w�G;�H;�0H;PH;�jH;��H;��H;V�H;E�H;�H;��H;��H;�H;��H;��H;��H;�H;��H;j�H;��H;j�H;��H;�H;��H;��H;��H;�H;��H;��H;�H;E�H;V�H;��H;��H;�jH;PH;�0H;�H;w�G;3�G;�WG;S�F;KF;y�D;�XC;�A;0>;�:;,�6;�2;�i-;d�(;�%;�";� ;      ��4;y�4;��5;Rl7;�^9;��;;�=;f�?;��A;�C;��D;��E;�F;�(G;ˀG;8�G;�G;jH;�5H;�RH;'lH;��H;˓H;#�H;گH;g�H;<�H;H�H;��H;��H;(�H;��H;C�H;��H;��H;m�H;��H;m�H;��H;��H;C�H;��H;(�H;��H;��H;H�H;<�H;g�H;گH;#�H;˓H;��H;'lH;�RH;�5H;jH;�G;8�G;ˀG;�(G;�F;��E;��D;�C;��A;f�?;�=;��;;�^9;Rl7;��5;y�4;      �_?;	�?;6�?;�@;��A;��B;��C;3�D;~hE;#F;[�F;G;�mG;F�G;$�G;t�G;� H;C>H;�XH;�oH;i�H;��H;#�H;\�H;��H;;�H;Y�H;�H;��H;��H;g�H;��H;��H;��H;��H;E�H;^�H;E�H;��H;��H;��H;��H;g�H;��H;��H;�H;Y�H;;�H;��H;\�H;#�H;��H;i�H;�oH;�XH;C>H;� H;t�G;$�G;F�G;�mG;G;[�F;#F;~hE;3�D;��C;��B;��A;�@;6�?;	�?;      �lD;#~D;��D;�D;�[E;+�E;�/F;�F;��F;$8G;�uG;'�G;u�G;��G;cH;�/H;aIH;�`H;	uH;�H;��H;V�H;گH;��H;�H;��H;}�H;#�H;��H;�H;n�H;N�H;��H;��H;��H;��H;6�H;��H;��H;��H;��H;N�H;n�H;�H;��H;#�H;}�H;��H;�H;��H;گH;V�H;��H;�H;	uH;�`H;aIH;�/H;cH;��G;u�G;'�G;�uG;$8G;��F;�F;�/F;+�E;�[E;�D;��D;#~D;      ��F;q�F;��F;�F;��F;�G;�FG; pG;]�G;l�G;�G;��G;!H;2)H;�@H;xVH;VjH;5|H;=�H;f�H;��H;E�H;g�H;;�H;��H;E�H;��H;��H;��H;�H;�H;��H;��H;��H;B�H;��H;��H;��H;B�H;��H;��H;��H;�H;�H;��H;��H;��H;E�H;��H;;�H;g�H;E�H;��H;f�H;=�H;5|H;VjH;xVH;�@H;2)H;!H;��G;�G;l�G;]�G; pG;�FG;�G;��F;�F;��F;q�F;      puG;3xG;/�G;��G;�G;��G;�G;��G;��G;�H;IH;�+H;�?H;�RH;�dH;�uH;ńH;��H;�H;�H;��H;�H;<�H;Y�H;}�H;��H;t�H;m�H;��H;��H;n�H;��H;��H;L�H;��H;-�H;.�H;-�H;��H;L�H;��H;��H;n�H;��H;��H;m�H;t�H;��H;}�H;Y�H;<�H;�H;��H;�H;�H;��H;ńH;�uH;�dH;�RH;�?H;�+H;IH;�H;��G;��G;�G;��G;�G;��G;/�G;3xG;      M�G;��G;��G;��G;��G;��G;WH;H;�'H;7H;�FH;/VH;MeH;�sH;d�H;�H;ٙH;��H;�H;��H;�H;��H;H�H;�H;#�H;��H;m�H;��H;��H;p�H;��H;��H;c�H;��H;V�H;��H;��H;��H;V�H;��H;c�H;��H;��H;p�H;��H;��H;m�H;��H;#�H;�H;H�H;��H;�H;��H;�H;��H;ٙH;�H;d�H;�sH;MeH;/VH;�FH;7H;�'H;H;WH;��G;��G;��G;��G;��G;      �H;�H;s"H;3'H;�-H;�5H;?H;XIH;eTH;�_H;�kH;9wH;��H;��H;��H;��H;��H;��H;�H;��H;��H;��H;��H;��H;��H;��H;��H;��H;>�H;��H;��H;X�H;��H;y�H;��H;��H;��H;��H;��H;y�H;��H;X�H;��H;��H;>�H;��H;��H;��H;��H;��H;��H;��H;��H;��H;�H;��H;��H;��H;��H;��H;��H;9wH;�kH;�_H;eTH;XIH;?H;�5H;�-H;3'H;s"H;�H;      �NH;NOH;�QH;UH;�YH;�_H;�fH;dnH;�vH;,H;�H;��H;R�H;��H;x�H;ܰH;��H;��H;��H;��H;)�H;�H;��H;��H;�H;�H;��H;p�H;��H;��H;V�H;��H;q�H;��H;�H;%�H;?�H;%�H;�H;��H;q�H;��H;V�H;��H;��H;p�H;��H;�H;�H;��H;��H;�H;)�H;��H;��H;��H;��H;ܰH;x�H;��H;R�H;��H;�H;,H;�vH;dnH;�fH;�_H;�YH;UH;�QH;NOH;      �rH;IsH;�tH;�wH;{H;�H;��H;i�H;��H;�H;��H;W�H;ժH;�H;��H;��H;�H;��H;9�H;�H;r�H;��H;(�H;g�H;n�H;�H;n�H;��H;��H;V�H;��H;q�H;��H;�H;_�H;l�H;d�H;l�H;_�H;�H;��H;q�H;��H;V�H;��H;��H;n�H;�H;n�H;g�H;(�H;��H;r�H;�H;9�H;��H;�H;��H;��H;�H;ժH;W�H;��H;�H;��H;i�H;��H;�H;{H;�wH;�tH;IsH;      �H;:�H;z�H;�H;�H;{�H;V�H;��H;L�H; �H;�H;�H;��H;ͼH;��H;��H;��H;}�H;��H;��H;��H;��H;��H;��H;N�H;��H;��H;��H;X�H;��H;q�H;��H;�H;_�H;��H;��H;��H;��H;��H;_�H;�H;��H;q�H;��H;X�H;��H;��H;��H;N�H;��H;��H;��H;��H;��H;��H;}�H;��H;��H;��H;ͼH;��H;�H;�H; �H;L�H;��H;V�H;{�H;�H;�H;z�H;:�H;      ��H;�H;�H;f�H;i�H;��H;ͫH;�H;��H;g�H;H�H;.�H;�H;��H;;�H;��H;��H;��H;-�H;��H;��H;��H;C�H;��H;��H;��H;��H;c�H;��H;q�H;��H;�H;X�H;��H;��H;��H;��H;��H;��H;��H;X�H;�H;��H;q�H;��H;c�H;��H;��H;��H;��H;C�H;��H;��H;��H;-�H;��H;��H;��H;;�H;��H;�H;.�H;H�H;g�H;��H;�H;ͫH;��H;i�H;f�H;�H;�H;      ��H;�H;��H;ñH;u�H;r�H;��H;[�H;�H;�H;�H;�H;
�H;��H;��H;k�H;��H;4�H;M�H;5�H;��H;�H;��H;��H;��H;��H;L�H;��H;y�H;��H;�H;_�H;��H;��H;��H;��H;��H;��H;��H;��H;��H;_�H;�H;��H;y�H;��H;L�H;��H;��H;��H;��H;�H;��H;5�H;M�H;4�H;��H;k�H;��H;��H;
�H;�H;�H;�H;�H;[�H;��H;r�H;u�H;ñH;��H;�H;      �H;W�H;�H;ۺH;6�H;ɽH;��H;��H;��H;m�H;��H;Q�H;��H;,�H;��H;��H;��H;��H;r�H;�H;z�H;��H;��H;��H;��H;B�H;��H;V�H;��H;�H;_�H;��H;��H;��H;��H;��H;��H;��H;��H;��H;��H;��H;_�H;�H;��H;V�H;��H;B�H;��H;��H;��H;��H;z�H;�H;r�H;��H;��H;��H;��H;,�H;��H;Q�H;��H;m�H;��H;��H;��H;ɽH;6�H;ۺH;�H;W�H;      q�H;��H;�H;�H;�H;r�H;�H;��H;��H;��H;"�H;`�H;��H;��H;��H;��H;v�H;8�H;��H;(�H;W�H;j�H;m�H;E�H;��H;��H;-�H;��H;��H;%�H;l�H;��H;��H;��H;��H;��H;��H;��H;��H;��H;��H;��H;l�H;%�H;��H;��H;-�H;��H;��H;E�H;m�H;j�H;W�H;(�H;��H;8�H;v�H;��H;��H;��H;��H;`�H;"�H;��H;��H;��H;�H;r�H;�H;�H;�H;��H;      E�H;U�H;��H;��H;��H;��H;��H;G�H;4�H;3�H;F�H;O�H;V�H;l�H;l�H;Q�H;�H;��H;�H;q�H;��H;��H;��H;^�H;6�H;��H;.�H;��H;��H;?�H;d�H;��H;��H;��H;��H;��H;��H;��H;��H;��H;��H;��H;d�H;?�H;��H;��H;.�H;��H;6�H;^�H;��H;��H;��H;q�H;�H;��H;�H;Q�H;l�H;l�H;V�H;O�H;F�H;3�H;4�H;G�H;��H;��H;��H;��H;��H;U�H;      q�H;��H;�H;�H;�H;r�H;�H;��H;��H;��H;"�H;`�H;��H;��H;��H;��H;v�H;8�H;��H;(�H;W�H;j�H;m�H;E�H;��H;��H;-�H;��H;��H;%�H;l�H;��H;��H;��H;��H;��H;��H;��H;��H;��H;��H;��H;l�H;%�H;��H;��H;-�H;��H;��H;E�H;m�H;j�H;W�H;(�H;��H;8�H;v�H;��H;��H;��H;��H;`�H;"�H;��H;��H;��H;�H;r�H;�H;�H;�H;��H;      �H;W�H;�H;ۺH;6�H;ɽH;��H;��H;��H;m�H;��H;Q�H;��H;,�H;��H;��H;��H;��H;r�H;�H;z�H;��H;��H;��H;��H;B�H;��H;V�H;��H;�H;_�H;��H;��H;��H;��H;��H;��H;��H;��H;��H;��H;��H;_�H;�H;��H;V�H;��H;B�H;��H;��H;��H;��H;z�H;�H;r�H;��H;��H;��H;��H;,�H;��H;Q�H;��H;m�H;��H;��H;��H;ɽH;6�H;ۺH;�H;W�H;      ��H;�H;��H;ñH;u�H;r�H;��H;[�H;�H;�H;�H;�H;
�H;��H;��H;k�H;��H;4�H;M�H;5�H;��H;�H;��H;��H;��H;��H;L�H;��H;y�H;��H;�H;_�H;��H;��H;��H;��H;��H;��H;��H;��H;��H;_�H;�H;��H;y�H;��H;L�H;��H;��H;��H;��H;�H;��H;5�H;M�H;4�H;��H;k�H;��H;��H;
�H;�H;�H;�H;�H;[�H;��H;r�H;u�H;ñH;��H;�H;      ��H;�H;�H;f�H;i�H;��H;ͫH;�H;��H;g�H;H�H;.�H;�H;��H;;�H;��H;��H;��H;-�H;��H;��H;��H;C�H;��H;��H;��H;��H;c�H;��H;q�H;��H;�H;X�H;��H;��H;��H;��H;��H;��H;��H;X�H;�H;��H;q�H;��H;c�H;��H;��H;��H;��H;C�H;��H;��H;��H;-�H;��H;��H;��H;;�H;��H;�H;.�H;H�H;g�H;��H;�H;ͫH;��H;i�H;f�H;�H;�H;      �H;:�H;z�H;�H;�H;{�H;V�H;��H;L�H; �H;�H;�H;��H;ͼH;��H;��H;��H;}�H;��H;��H;��H;��H;��H;��H;N�H;��H;��H;��H;X�H;��H;q�H;��H;�H;_�H;��H;��H;��H;��H;��H;_�H;�H;��H;q�H;��H;X�H;��H;��H;��H;N�H;��H;��H;��H;��H;��H;��H;}�H;��H;��H;��H;ͼH;��H;�H;�H; �H;L�H;��H;V�H;{�H;�H;�H;z�H;:�H;      �rH;IsH;�tH;�wH;{H;�H;��H;i�H;��H;�H;��H;W�H;ժH;�H;��H;��H;�H;��H;9�H;�H;r�H;��H;(�H;g�H;n�H;�H;n�H;��H;��H;V�H;��H;q�H;��H;�H;_�H;l�H;d�H;l�H;_�H;�H;��H;q�H;��H;V�H;��H;��H;n�H;�H;n�H;g�H;(�H;��H;r�H;�H;9�H;��H;�H;��H;��H;�H;ժH;W�H;��H;�H;��H;i�H;��H;�H;{H;�wH;�tH;IsH;      �NH;NOH;�QH;UH;�YH;�_H;�fH;dnH;�vH;,H;�H;��H;R�H;��H;x�H;ܰH;��H;��H;��H;��H;)�H;�H;��H;��H;�H;�H;��H;p�H;��H;��H;V�H;��H;q�H;��H;�H;%�H;?�H;%�H;�H;��H;q�H;��H;V�H;��H;��H;p�H;��H;�H;�H;��H;��H;�H;)�H;��H;��H;��H;��H;ܰH;x�H;��H;R�H;��H;�H;,H;�vH;dnH;�fH;�_H;�YH;UH;�QH;NOH;      �H;�H;s"H;3'H;�-H;�5H;?H;XIH;eTH;�_H;�kH;9wH;��H;��H;��H;��H;��H;��H;�H;��H;��H;��H;��H;��H;��H;��H;��H;��H;>�H;��H;��H;X�H;��H;y�H;��H;��H;��H;��H;��H;y�H;��H;X�H;��H;��H;>�H;��H;��H;��H;��H;��H;��H;��H;��H;��H;�H;��H;��H;��H;��H;��H;��H;9wH;�kH;�_H;eTH;XIH;?H;�5H;�-H;3'H;s"H;�H;      M�G;��G;��G;��G;��G;��G;WH;H;�'H;7H;�FH;/VH;MeH;�sH;d�H;�H;ٙH;��H;�H;��H;�H;��H;H�H;�H;#�H;��H;m�H;��H;��H;p�H;��H;��H;c�H;��H;V�H;��H;��H;��H;V�H;��H;c�H;��H;��H;p�H;��H;��H;m�H;��H;#�H;�H;H�H;��H;�H;��H;�H;��H;ٙH;�H;d�H;�sH;MeH;/VH;�FH;7H;�'H;H;WH;��G;��G;��G;��G;��G;      puG;3xG;/�G;��G;�G;��G;�G;��G;��G;�H;IH;�+H;�?H;�RH;�dH;�uH;ńH;��H;�H;�H;��H;�H;<�H;Y�H;}�H;��H;t�H;m�H;��H;��H;n�H;��H;��H;L�H;��H;-�H;.�H;-�H;��H;L�H;��H;��H;n�H;��H;��H;m�H;t�H;��H;}�H;Y�H;<�H;�H;��H;�H;�H;��H;ńH;�uH;�dH;�RH;�?H;�+H;IH;�H;��G;��G;�G;��G;�G;��G;/�G;3xG;      ��F;q�F;��F;�F;��F;�G;�FG; pG;]�G;l�G;�G;��G;!H;2)H;�@H;xVH;VjH;5|H;=�H;f�H;��H;E�H;g�H;;�H;��H;E�H;��H;��H;��H;�H;�H;��H;��H;��H;B�H;��H;��H;��H;B�H;��H;��H;��H;�H;�H;��H;��H;��H;E�H;��H;;�H;g�H;E�H;��H;f�H;=�H;5|H;VjH;xVH;�@H;2)H;!H;��G;�G;l�G;]�G; pG;�FG;�G;��F;�F;��F;q�F;      �lD;#~D;��D;�D;�[E;+�E;�/F;�F;��F;$8G;�uG;'�G;u�G;��G;cH;�/H;aIH;�`H;	uH;�H;��H;V�H;گH;��H;�H;��H;}�H;#�H;��H;�H;n�H;N�H;��H;��H;��H;��H;6�H;��H;��H;��H;��H;N�H;n�H;�H;��H;#�H;}�H;��H;�H;��H;گH;V�H;��H;�H;	uH;�`H;aIH;�/H;cH;��G;u�G;'�G;�uG;$8G;��F;�F;�/F;+�E;�[E;�D;��D;#~D;      �_?;	�?;6�?;�@;��A;��B;��C;3�D;~hE;#F;[�F;G;�mG;F�G;$�G;t�G;� H;C>H;�XH;�oH;i�H;��H;#�H;\�H;��H;;�H;Y�H;�H;��H;��H;g�H;��H;��H;��H;��H;E�H;^�H;E�H;��H;��H;��H;��H;g�H;��H;��H;�H;Y�H;;�H;��H;\�H;#�H;��H;i�H;�oH;�XH;C>H;� H;t�G;$�G;F�G;�mG;G;[�F;#F;~hE;3�D;��C;��B;��A;�@;6�?;	�?;      ��4;y�4;��5;Rl7;�^9;��;;�=;f�?;��A;�C;��D;��E;�F;�(G;ˀG;8�G;�G;jH;�5H;�RH;'lH;��H;˓H;#�H;گH;g�H;<�H;H�H;��H;��H;(�H;��H;C�H;��H;��H;m�H;��H;m�H;��H;��H;C�H;��H;(�H;��H;��H;H�H;<�H;g�H;گH;#�H;˓H;��H;'lH;�RH;�5H;jH;�G;8�G;ˀG;�(G;�F;��E;��D;�C;��A;f�?;�=;��;;�^9;Rl7;��5;y�4;      �d;� ;�";�%;d�(;�i-;�2;,�6;�:;0>;�A;�XC;y�D;KF;S�F;�WG;3�G;w�G;�H;�0H;PH;�jH;��H;��H;V�H;E�H;�H;��H;��H;�H;��H;��H;��H;�H;��H;j�H;��H;j�H;��H;�H;��H;��H;��H;�H;��H;��H;�H;E�H;V�H;��H;��H;�jH;PH;�0H;�H;w�G;3�G;�WG;S�F;KF;y�D;�XC;�A;0>;�:;,�6;�2;�i-;d�(;�%;�";� ;      ���:�A�:���:�w;�
;6;��;}$;�{,;ǂ3;_9;�>;ayA;�C;,�E;?�F;Z4G;��G;��G;nH;�.H;PH;'lH;i�H;��H;��H;��H;�H;��H;)�H;r�H;��H;��H;��H;z�H;W�H;��H;W�H;z�H;��H;��H;��H;r�H;)�H;��H;�H;��H;��H;��H;i�H;'lH;PH;�.H;nH;��G;��G;Z4G;?�F;,�E;�C;ayA;�>;_9;ǂ3;�{,;}$;��;6;�
;�w;���:�A�:      �v[:�Ad:6�}:_�:��:0��:C�:��;P;� ;H+;�3;:�:;i�?;�B;�
E;�YF;
G;R�G;��G;nH;�0H;�RH;�oH;�H;f�H;�H;��H;��H;��H;�H;��H;��H;5�H;�H;(�H;q�H;(�H;�H;5�H;��H;��H;�H;��H;��H;��H;�H;f�H;�H;�oH;�RH;�0H;nH;��G;R�G;
G;�YF;�
E;�B;i�?;:�:;�3;H+;� ;P;��;C�:0��:��:_�:6�}:�Ad:      ��S���D�.�������'7��9c�R:���:���:@��:X>;G";^P.;�l7;C�=;�B;%�D;�8F;YG;R�G;��G;�H;�5H;�XH;	uH;=�H;�H;�H;�H;��H;9�H;��H;-�H;M�H;r�H;��H;�H;��H;r�H;M�H;-�H;��H;9�H;��H;�H;�H;�H;=�H;	uH;�XH;�5H;�H;��G;R�G;YG;�8F;%�D;�B;C�=;�l7;^P.;G";X>;@��:���:���:c�R:��9��'7���.����D�      �D^��/X��qF�'}*�'���P���D��Ҭ�kh:��:���:ȏ; �;��);��4;p�<;`�A;f�D;�8F;
G;��G;w�G;jH;C>H;�`H;5|H;��H;��H;��H;��H;��H;}�H;��H;4�H;��H;8�H;��H;8�H;��H;4�H;��H;}�H;��H;��H;��H;��H;��H;5|H;�`H;C>H;jH;w�G;��G;
G;�8F;f�D;`�A;p�<;��4;��); �;ȏ;���:��:kh:�Ҭ��D��P��'��'}*��qF��/X�      s��v��,�ܻ�ƻB󩻜��gFL����θ��"��N�-:g�:���:v;>&;��3;�8<;`�A;%�D;�YF;Z4G;3�G;�G;� H;aIH;VjH;ńH;ٙH;��H;��H;�H;��H;��H;��H;��H;v�H;�H;v�H;��H;��H;��H;��H;�H;��H;��H;ٙH;ńH;VjH;aIH;� H;�G;3�G;Z4G;�YF;%�D;`�A;�8<;��3;>&;v;���:g�:N�-:"��θ�����gFL����B��ƻ,�ܻv��      ;�V�z5S�Y6H�x�6�� �3,�n?ػG���D^����2�D����9�3�:? �:��;^%;��3;p�<;�B;�
E;?�F;�WG;8�G;t�G;�/H;xVH;�uH;�H;��H;ܰH;��H;��H;��H;k�H;��H;��H;Q�H;��H;��H;k�H;��H;��H;��H;ܰH;��H;�H;�uH;xVH;�/H;t�G;8�G;�WG;?�F;�
E;�B;p�<;��3;^%;��;? �:�3�:���92�D�����D^�G��n?ػ3,�� �x�6�Y6H�z5S�      ����-��#Ȥ�d���ݫ���f�G�=����	�ܻ�*��>o5�t���>Q(7G�}:�m�:��;>&;��4;C�=;�B;,�E;S�F;ˀG;$�G;cH;�@H;�dH;d�H;��H;x�H;��H;��H;;�H;��H;��H;��H;l�H;��H;��H;��H;;�H;��H;��H;x�H;��H;d�H;�dH;�@H;cH;$�G;ˀG;S�F;,�E;�B;C�=;��4;>&;��;�m�:G�}:>Q(7t���>o5��*��	�ܻ���G�=��f�ݫ��d���#Ȥ��-��      xc��8�|����켔�Ҽg���`�����r�E:�$,�#ߵ�Y/X���º�ˬ�G�}:? �:v;��);�l7;i�?;�C;KF;�(G;F�G;��G;2)H;�RH;�sH;��H;��H;�H;ͼH;��H;��H;,�H;��H;l�H;��H;,�H;��H;��H;ͼH;�H;��H;��H;�sH;�RH;2)H;��G;F�G;�(G;KF;�C;i�?;�l7;��);v;? �:G�}:�ˬ���ºY/X�#ߵ�$,�E:���r�`���g�����Ҽ��|����8�      �&K���G�ȟ>��0�:y�vc�d��)������!�V����ƻfod���º>Q(7�3�:���: �;^P.;:�:;ayA;y�D;�F;�mG;u�G;!H;�?H;MeH;��H;R�H;ժH;��H;�H;
�H;��H;��H;V�H;��H;��H;
�H;�H;��H;ժH;R�H;��H;MeH;�?H;!H;u�G;�mG;�F;y�D;ayA;:�:;^P.; �;���:�3�:>Q(7��ºfod��ƻ��!�V����)���d��vc�:y��0�ȟ>���G�      鰒�Z��������}��c���D�/%��8���Ҽ	c����f�����ƻY/X�t������9g�:ȏ;G";�3;�>;�XC;��E;G;'�G;��G;�+H;/VH;9wH;��H;W�H;�H;.�H;�H;Q�H;`�H;O�H;`�H;Q�H;�H;.�H;�H;W�H;��H;9wH;/VH;�+H;��G;'�G;G;��E;�XC;�>;�3;G";ȏ;g�:���9t���Y/X��ƻ�����f�	c����Ҽ�8�/%���D��c���}�����Z��      \Pν��ʽ*8�������������0�f�u�;���K��Ȥ���f���#ߵ�>o5�2�D�N�-:���:X>;H+;_9;�A;��D;[�F;�uG;�G;IH;�FH;�kH;�H;��H;�H;H�H;�H;��H;"�H;F�H;"�H;��H;�H;H�H;�H;��H;�H;�kH;�FH;IH;�G;�uG;[�F;��D;�A;_9;H+;X>;���:N�-:2�D�>o5�#ߵ�����f�Ȥ�K����u�;�0�f������������*8����ʽ      ���N9�C[��s�R�ؽ���s����}���G��K��	c��!�V�$,��*�����"����:@��:� ;ǂ3;0>;�C;#F;$8G;l�G;�H;7H;�_H;,H;�H; �H;g�H;�H;m�H;��H;3�H;��H;m�H;�H;g�H; �H;�H;,H;�_H;7H;�H;l�G;$8G;#F;�C;0>;ǂ3;� ;@��:��:"������*��$,�!�V�	c��K�����G���}��s����R�ؽ�s�C[�N9�      }�=���:���0��Q"�e�����ZPν�榽%����G�����Ҽ���E:�	�ܻ�D^�θ��kh:���:P;�{,;�:;��A;~hE;��F;]�G;��G;�'H;eTH;�vH;��H;L�H;��H;�H;��H;��H;4�H;��H;��H;�H;��H;L�H;��H;�vH;eTH;�'H;��G;]�G;��F;~hE;��A;�:;�{,;P;���:kh:θ���D^�	�ܻE:������Ҽ����G�%���榽ZPν����e��Q"���0���:�      
Dx��s���f�QS���:����B[��7ս�榽��}�u�;��8�)�����r����G������Ҭ����:��;}$;,�6;f�?;3�D;�F; pG;��G;H;XIH;dnH;i�H;��H;�H;[�H;��H;��H;G�H;��H;��H;[�H;�H;��H;i�H;dnH;XIH;H;��G; pG;�F;3�D;f�?;,�6;}$;��;���:�Ҭ����G�������r�)����8�u�;���}��榽�7սB[������:�QS���f��s�      �*���0��ȥ��&���jk��H��#%�B[�ZPν�s��0�f�/%�d��`���G�=�n?ػgFL��D�c�R:C�:��;�2;�=;��C;�/F;�FG;�G;WH;?H;�fH;��H;V�H;ͫH;��H;��H;�H;��H;�H;��H;��H;ͫH;V�H;��H;�fH;?H;WH;�G;�FG;�/F;��C;�=;�2;��;C�:c�R:�D�gFL�n?ػG�=�`���d��/%�0�f��s��ZPνB[��#%��H�jk�&���ȥ���0��      �þ��������R��f쏾�s��H����������������D�vc�g����f�3,�����P����90��:6;�i-;��;;��B;+�E;�G;��G;��G;�5H;�_H;�H;{�H;��H;r�H;ɽH;r�H;��H;r�H;ɽH;r�H;��H;{�H;�H;�_H;�5H;��G;��G;�G;+�E;��B;��;;�i-;6;0��:��9�P�����3,��f�g���vc���D���������������H��s�f쏾�R���������      ����fYؾ�þ�ê�f쏾jk���:�e�R�ؽ�����c�:y���Ҽݫ��� �B�'����'7��:�
;d�(;�^9;��A;�[E;��F;�G;��G;�-H;�YH;{H;�H;i�H;u�H;6�H;�H;��H;�H;6�H;u�H;i�H;�H;{H;�YH;�-H;��G;�G;��F;�[E;��A;�^9;d�(;�
;��:��'7'��B�� �ݫ����Ҽ:y��c�����R�ؽe���:�jk�f쏾�ê��þfYؾ��      ��=������I��þ�R��&���QS��Q"��s�����}��0���d���x�6��ƻ'}*����_�:�w;�%;Rl7;�@;�D;�F;��G;��G;3'H;UH;�wH;�H;f�H;ñH;ۺH;�H;��H;�H;ۺH;ñH;f�H;�H;�wH;UH;3'H;��G;��G;�F;�D;�@;Rl7;�%;�w;_�:���'}*��ƻx�6�d����켟0���}�����s��Q"�QS�&����R���þIᾁ���=��      ���>��&�
�����fYؾ���ȥ����f���0�C[�*8������ȟ>�|���#Ȥ�Y6H�,�ܻ�qF�.��6�}:���:�";��5;6�?;��D;��F;/�G;��G;s"H;�QH;�tH;z�H;�H;��H;�H;�H;��H;�H;�H;��H;�H;z�H;�tH;�QH;s"H;��G;/�G;��F;��D;6�?;��5;�";���:6�}:.���qF�,�ܻY6H�#Ȥ�|���ȟ>�����*8��C[���0���f�ȥ�����fYؾ����&�
�>��      �� �k��>��=���������0���s���:�N9���ʽZ����G��8��-��z5S�v���/X���D��Ad:�A�:� ;y�4;	�?;#~D;q�F;3xG;��G;�H;NOH;IsH;:�H;�H;�H;W�H;��H;U�H;��H;W�H;�H;�H;:�H;IsH;NOH;�H;��G;3xG;q�F;#~D;	�?;y�4;� ;�A�:�Ad:��D��/X�v��z5S��-���8���G�Z����ʽN9���:��s��0��������=��>��k��      3F�/h��ǰ�3Vھ�������~���S��#��o��S��R₽�6�-���<y��FB��Eֻ_A?��	�Y�:���:�";�36;�@;��D;�F;�mG;&�G;>H;9?H;fH;w�H;P�H;��H;��H;�H;�H;�H;��H;��H;P�H;w�H;fH;9?H;>H;&�G;�mG;�F;��D;�@;�36;�";���:Y�:�	�_A?��EֻFB�<y��-����6�R₽S���o���#��S��~��������3Vھǰ�/h��      /h���b���쾅*־�v������)�� �O�6� ��r�r���؀��3����ݜ��>��ѻ��9�����n�:�$ ;�L#;˃6;�@@;C�D;�F;<pG;��G;TH;@H;�fH;�H;��H;�H;>�H;�H;��H;�H;>�H;�H;��H;�H;�fH;@H;TH;��G;<pG;�F;C�D;�@@;˃6;�L#;�$ ;�n�:�����9��ѻ�>�ݜ�����3��؀��r���r�6� � �O��)������v���*־�쾼b��      ǰ�쾐�޾5ʾ/;���:����v��E�A'���L����u�X�+�aW缨A��r�4�n�Ļ�8)��j��W�:�;�%;kk7;g�@;B�D;4�F;wG;��G;vH;cBH;YhH;B�H;��H;ƩH;�H;��H;��H;��H;�H;ƩH;��H;B�H;YhH;cBH;vH;��G;wG;4�F;B�D;g�@;kk7;�%;�;W�:�j���8)�n�Ļr�4��A��aW�X�+���u�L����A'��E���v��:��/;��5ʾ��޾��      3Vھ�*־5ʾT��������M���9b��5���}�սn���Xc�ݟ���ռ�I��$�$�4T���Z�_����:��;��';��8;]QA;�8E;��F;�G;%�G;�H;-FH;@kH;u�H;Z�H;�H;�H;��H;t�H;��H;�H;�H;Z�H;u�H;@kH;-FH;�H;%�G;�G;��F;�8E;]QA;��8;��';��;��:_���Z�4T��$�$��I����ռݟ��Xc�n��}�ս���5��9b��M������T���5ʾ�*־      ���v��/;������:P���r�U�H�6� ��~��@������Q�K�<��վ���s�F��_�~ܺ3u9�%�:��;��+;��:;"B;��E;,�F;��G;�G;nH;[KH;(oH;k�H;��H;ƬH;_�H;��H;��H;��H;_�H;ƬH;��H;k�H;(oH;[KH;nH;�G;��G;,�F;��E;"B;��:;��+;��;�%�:3u9~ܺ_�F����s��վ�<�Q�K�����@���~��6� �U�H��r�:P������/;���v��      ��������:���M���r� �O��",�<�
��gٽKĥ�|�u�K1�(����Τ�m�P��Z�q.o�kp���:Դ�:{P;��/;��<;F
C;f�E;� G;^�G;5�G;�$H;�QH;�sH;%�H;f�H;��H;*�H;{�H;&�H;{�H;*�H;��H;f�H;%�H;�sH;�QH;�$H;5�G;^�G;� G;f�E;F
C;��<;��/;{P;Դ�:�:kp��q.o��Z�m�P��Τ�(���K1�|�u�Kĥ��gٽ<�
��",� �O��r��M���:�����      �~���)����v��9b�U�H��",�0Z���S��X^��e�N�{����μ�I���%+�ۚ����.������i~:���:�l;@�3;��>;�C;�OF;�EG;|�G;"�G;�.H;'YH;�yH;p�H;��H;��H;F�H;K�H;��H;K�H;F�H;��H;��H;p�H;�yH;'YH;�.H;"�G;|�G;�EG;�OF;�C;��>;@�3;�l;���:�i~:������.�ۚ���%+��I����μ{��e�N�X^��S����0Z��",�U�H��9b���v��)��      �S� �O��E��5�6� �<�
���|9��l���Xc���(����߈��Z�[����nݎ�ܺH99���:��	;�c';��7;��@;��D;.�F;biG;��G;�H;�9H;faH;�H;/�H;P�H;g�H;��H;Y�H;��H;Y�H;��H;g�H;P�H;/�H;�H;faH;�9H;�H;��G;biG;.�F;��D;��@;��7;�c';��	;���:H99ܺnݎ����Z�[�߈�������(��Xc�l��|9����<�
�6� ��5��E� �O�      �#�6� �A'����~���gٽS��l���j��3�ji��վ�T����(�P�Ļ+A?���B�6�@:[�:�P;w�.;Q�;;�sB;\�E;��F;l�G;'�G;H;�EH;KjH;��H;H�H;.�H;��H;0�H;��H;�H;��H;0�H;��H;.�H;H�H;��H;KjH;�EH;H;'�G;l�G;��F;\�E;�sB;Q�;;w�.;�P;[�:6�@:��B�+A?�P�Ļ�(�T����վ�ji��3��j�l��S���gٽ�~����A'�6� �      �o���r���}�ս@��Kĥ�X^���Xc��3���	���˼t]��FB��Z򻆜��DӺ8��8�:z�;RM#;�<5;x?;��C;�?F;J9G;,�G;M�G;c&H;�QH;�sH;ۍH;��H;H�H;кH;��H;��H;a�H;��H;��H;кH;H�H;��H;ۍH;�sH;�QH;c&H;M�G;,�G;J9G;�?F;��C;x?;�<5;RM#;z�;�:8��8DӺ�����Z�FB�t]����˼��	��3��Xc�X^��Kĥ�@��}�ս���r�      S���r��L��n������|�u�e�N���(�ji���˼�A��b�P�=s��|������\:�:�;�m-;F�:;N�A;�+E;��F;mnG;,�G;�H;�6H;k^H;0}H;�H;&�H;��H;/�H;��H;Z�H;��H;Z�H;��H;/�H;��H;&�H;�H;0}H;k^H;�6H;�H;,�G;mnG;��F;�+E;N�A;F�:;�m-;�;�:�\:����|��=s�b�P��A����˼ji���(�e�N�|�u�����n��L���r��      R₽�؀���u��Xc�Q�K�K1�{�����վ�t]��b�P�l��	T��g�9��o�k2�9�%�:��	;�%;��5;�>;��C;	F;� G;ݙG;�G;pH;�GH;�jH;ʆH;s�H;��H;̸H;��H;l�H;��H;��H;��H;l�H;��H;̸H;��H;s�H;ʆH;�jH;�GH;pH;�G;ݙG;� G;	F;��C;�>;��5;�%;��	;�%�:k2�9�o�g�9�	T��l��b�P�t]���վ����{��K1�Q�K��Xc���u��؀�      �6��3�X�+�ݟ�<�(�����μ߈��T���FB�=s�	T����D��{���8u91q�:���:�X;at0;T�;;1B;C9E;/�F;:gG;�G;<�G;�/H;�WH;SwH;G�H;��H;$�H;�H; �H;2�H;I�H;S�H;I�H;2�H; �H;�H;$�H;��H;G�H;SwH;�WH;�/H;<�G;�G;:gG;/�F;C9E;1B;T�;;at0;�X;���:1q�:�8u9�{����D�	T��=s�FB�T���߈����μ(���<�ݟ�X�+��3�      -������aW缑�ռ�վ��Τ��I��Z�[��(��Z�g�9��{���99�W�:�W�:�P;�,;�8;�@@;ZAD;�?F;�+G;ÛG;��G;�H;�CH;HgH;W�H;y�H;��H;�H;>�H;:�H;��H;��H;��H;��H;��H;:�H;>�H;�H;��H;y�H;W�H;HgH;�CH;�H;��G;ÛG;�+G;�?F;ZAD;�@@;�8;�,;�P;�W�:�W�:�99�{��g�9���Z��(�Z�[��I���Τ��վ���ռaW缧��      <y��ݜ��A���I����s�m�P��%+����P�Ļ����|��o��8u9�W�:9+�:�;]);8�6;ذ>;�OC;��E;:�F;�wG;a�G;� H;�0H;@WH;)vH;ԎH;8�H;#�H;��H;4�H;^�H;��H;�H;��H;�H;��H;^�H;4�H;��H;#�H;8�H;ԎH;)vH;@WH;�0H;� H;a�G;�wG;:�F;��E;�OC;ذ>;8�6;]);�;9+�:�W�:�8u9�o�|�����P�Ļ����%+�m�P���s��I���A��ݜ�      FB��>�r�4�$�$�F���Z�ۚ��nݎ�+A?�DӺ����k2�91q�:�W�:�;D�';�<5;֜=;Z�B;jFE;��F;�TG;Y�G;�G;�H;�GH;9iH;�H;��H;g�H;T�H;f�H;��H;[�H;(�H;5�H;��H;5�H;(�H;[�H;��H;f�H;T�H;g�H;��H;�H;9iH;�GH;�H;�G;Y�G;�TG;��F;jFE;Z�B;֜=;�<5;D�';�;�W�:1q�:k2�9����DӺ+A?�nݎ�ۚ���Z�F��$�$�r�4��>�      �Eֻ�ѻn�Ļ4T��_�q.o���.�ܺ��B�8��8�\:�%�:���:�P;]);�<5;K:=;x"B;��D;!uF;,6G;��G;��G;�H;�9H;:]H;�yH;�H;��H;�H;'�H;��H;u�H;6�H;��H;B�H;��H;B�H;��H;6�H;u�H;��H;'�H;�H;��H;�H;�yH;:]H;�9H;�H;��G;��G;,6G;!uF;��D;x"B;K:=;�<5;]);�P;���:�%�:�\:8��8��B�ܺ��.�q.o�_�4T��n�Ļ�ѻ      _A?���9��8)��Z�~ܺkp������H996�@:�:�:��	;�X;�,;8�6;֜=;x"B; �D;�WF;!G;��G;T�G;�H; .H;�RH;�pH;�H;ԜH;��H;׸H;��H;��H;��H;��H;��H;0�H;��H;0�H;��H;��H;��H;��H;��H;׸H;��H;ԜH;�H;�pH;�RH; .H;�H;T�G;��G;!G;�WF; �D;x"B;֜=;8�6;�,;�X;��	;�:�:6�@:H99����kp��~ܺ�Z��8)���9�      �	�����j��_��3u9�:�i~:���:[�:z�;�;�%;at0;�8;ذ>;Z�B;��D;�WF;sG;��G;��G;��G;%H;.JH;�hH;�H;��H;T�H;��H;�H;x�H;��H;��H;H�H;��H;��H;i�H;��H;��H;H�H;��H;��H;x�H;�H;��H;T�H;��H;�H;�hH;.JH;%H;��G;��G;��G;sG;�WF;��D;Z�B;ذ>;�8;at0;�%;�;z�;[�:���:�i~:�:3u9_���j�����      Y�:�n�:W�:��:�%�:Դ�:���:��	;�P;RM#;�m-;��5;T�;;�@@;�OC;jFE;!uF;!G;��G;�G;F�G;wH;7DH;�bH;e|H;��H;ԢH;��H;ۻH;��H;��H;B�H;i�H;e�H;^�H;��H;��H;��H;^�H;e�H;i�H;B�H;��H;��H;ۻH;��H;ԢH;��H;e|H;�bH;7DH;wH;F�G;�G;��G;!G;!uF;jFE;�OC;�@@;T�;;��5;�m-;RM#;�P;��	;���:Դ�:�%�:��:W�:�n�:      ���:�$ ;�;��;��;{P;�l;�c';w�.;�<5;F�:;�>;1B;ZAD;��E;��F;,6G;��G;��G;F�G;�H;AH;/_H;mxH;��H;<�H;m�H;��H;b�H;��H;��H;F�H;��H;S�H;�H;��H;Z�H;��H;�H;S�H;��H;F�H;��H;��H;b�H;��H;m�H;<�H;��H;mxH;/_H;AH;�H;F�G;��G;��G;,6G;��F;��E;ZAD;1B;�>;F�:;�<5;w�.;�c';�l;{P;��;��;�;�$ ;      �";�L#;�%;��';��+;��/;@�3;��7;Q�;;x?;N�A;��C;C9E;�?F;:�F;�TG;��G;T�G;��G;wH;AH;�]H;hvH;9�H;��H;��H;��H;E�H;�H;7�H;1�H;��H;��H;��H;x�H;U�H;��H;U�H;x�H;��H;��H;��H;1�H;7�H;�H;E�H;��H;��H;��H;9�H;hvH;�]H;AH;wH;��G;T�G;��G;�TG;:�F;�?F;C9E;��C;N�A;x?;Q�;;��7;@�3;��/;��+;��';�%;�L#;      �36;˃6;kk7;��8;��:;��<;��>;��@;�sB;��C;�+E;	F;/�F;�+G;�wG;Y�G;��G;�H;%H;7DH;/_H;hvH;O�H;P�H;h�H;��H;��H;��H;��H;�H;=�H;Q�H;��H;m�H;��H;{�H;��H;{�H;��H;m�H;��H;Q�H;=�H;�H;��H;��H;��H;��H;h�H;P�H;O�H;hvH;/_H;7DH;%H;�H;��G;Y�G;�wG;�+G;/�F;	F;�+E;��C;�sB;��@;��>;��<;��:;��8;kk7;˃6;      �@;�@@;g�@;]QA;"B;F
C;�C;��D;\�E;�?F;��F;� G;:gG;ÛG;a�G;�G;�H; .H;.JH;�bH;mxH;9�H;P�H;ܨH;#�H;��H;��H;��H;"�H;[�H;��H;[�H;K�H;��H;��H;i�H;��H;i�H;��H;��H;K�H;[�H;��H;[�H;"�H;��H;��H;��H;#�H;ܨH;P�H;9�H;mxH;�bH;.JH; .H;�H;�G;a�G;ÛG;:gG;� G;��F;�?F;\�E;��D;�C;F
C;"B;]QA;g�@;�@@;      ��D;C�D;B�D;�8E;��E;f�E;�OF;.�F;��F;J9G;mnG;ݙG;�G;��G;� H;�H;�9H;�RH;�hH;e|H;��H;��H;h�H;#�H;U�H;��H;@�H;}�H;��H;9�H;��H;�H;��H;��H;��H;-�H;q�H;-�H;��H;��H;��H;�H;��H;9�H;��H;}�H;@�H;��H;U�H;#�H;h�H;��H;��H;e|H;�hH;�RH;�9H;�H;� H;��G;�G;ݙG;mnG;J9G;��F;.�F;�OF;f�E;��E;�8E;B�D;C�D;      �F;�F;4�F;��F;,�F;� G;�EG;biG;l�G;,�G;,�G;�G;<�G;�H;�0H;�GH;:]H;�pH;�H;��H;<�H;��H;��H;��H;��H;�H;/�H;k�H;��H;��H;��H;��H;��H;��H;��H;��H;�H;��H;��H;��H;��H;��H;��H;��H;��H;k�H;/�H;�H;��H;��H;��H;��H;<�H;��H;�H;�pH;:]H;�GH;�0H;�H;<�G;�G;,�G;,�G;l�G;biG;�EG;� G;,�F;��F;4�F;�F;      �mG;<pG;wG;�G;��G;^�G;|�G;��G;'�G;M�G;�H;pH;�/H;�CH;@WH;9iH;�yH;�H;��H;ԢH;m�H;��H;��H;��H;@�H;/�H;N�H;��H;h�H;��H;X�H;��H;��H;��H;;�H;��H;��H;��H;;�H;��H;��H;��H;X�H;��H;h�H;��H;N�H;/�H;@�H;��H;��H;��H;m�H;ԢH;��H;�H;�yH;9iH;@WH;�CH;�/H;pH;�H;M�G;'�G;��G;|�G;^�G;��G;�G;wG;<pG;      &�G;��G;��G;%�G;�G;5�G;"�G;�H;H;c&H;�6H;�GH;�WH;HgH;)vH;�H;�H;ԜH;T�H;��H;��H;E�H;��H;��H;}�H;k�H;��H;G�H;��H;L�H;��H;��H;��H;k�H;��H;�H; �H;�H;��H;k�H;��H;��H;��H;L�H;��H;G�H;��H;k�H;}�H;��H;��H;E�H;��H;��H;T�H;ԜH;�H;�H;)vH;HgH;�WH;�GH;�6H;c&H;H;�H;"�G;5�G;�G;%�G;��G;��G;      >H;TH;vH;�H;nH;�$H;�.H;�9H;�EH;�QH;k^H;�jH;SwH;W�H;ԎH;��H;��H;��H;��H;ۻH;b�H;�H;��H;"�H;��H;��H;h�H;��H;,�H;��H;��H;��H;b�H;��H;L�H;�H;��H;�H;L�H;��H;b�H;��H;��H;��H;,�H;��H;h�H;��H;��H;"�H;��H;�H;b�H;ۻH;��H;��H;��H;��H;ԎH;W�H;SwH;�jH;k^H;�QH;�EH;�9H;�.H;�$H;nH;�H;vH;TH;      9?H;@H;cBH;-FH;[KH;�QH;'YH;faH;KjH;�sH;0}H;ʆH;G�H;y�H;8�H;g�H;�H;׸H;�H;��H;��H;7�H;�H;[�H;9�H;��H;��H;L�H;��H;��H;��H;m�H;�H;T�H;��H;��H;��H;��H;��H;T�H;�H;m�H;��H;��H;��H;L�H;��H;��H;9�H;[�H;�H;7�H;��H;��H;�H;׸H;�H;g�H;8�H;y�H;G�H;ʆH;0}H;�sH;KjH;faH;'YH;�QH;[KH;-FH;cBH;@H;      fH;�fH;YhH;@kH;(oH;�sH;�yH;�H;��H;ۍH;�H;s�H;��H;��H;#�H;T�H;'�H;��H;x�H;��H;��H;1�H;=�H;��H;��H;��H;X�H;��H;��H;��H;t�H;�H;h�H;��H;��H;�H;0�H;�H;��H;��H;h�H;�H;t�H;��H;��H;��H;X�H;��H;��H;��H;=�H;1�H;��H;��H;x�H;��H;'�H;T�H;#�H;��H;��H;s�H;�H;ۍH;��H;�H;�yH;�sH;(oH;@kH;YhH;�fH;      w�H;�H;B�H;u�H;k�H;%�H;p�H;/�H;H�H;��H;&�H;��H;$�H;�H;��H;f�H;��H;��H;��H;B�H;F�H;��H;Q�H;[�H;�H;��H;��H;��H;��H;m�H;�H;z�H;��H; �H;,�H;J�H;I�H;J�H;,�H; �H;��H;z�H;�H;m�H;��H;��H;��H;��H;�H;[�H;Q�H;��H;F�H;B�H;��H;��H;��H;f�H;��H;�H;$�H;��H;&�H;��H;H�H;/�H;p�H;%�H;k�H;u�H;B�H;�H;      P�H;��H;��H;Z�H;��H;f�H;��H;P�H;.�H;H�H;��H;̸H;�H;>�H;4�H;��H;u�H;��H;��H;i�H;��H;��H;��H;K�H;��H;��H;��H;��H;b�H;�H;h�H;��H;	�H;9�H;X�H;��H;��H;��H;X�H;9�H;	�H;��H;h�H;�H;b�H;��H;��H;��H;��H;K�H;��H;��H;��H;i�H;��H;��H;u�H;��H;4�H;>�H;�H;̸H;��H;H�H;.�H;P�H;��H;f�H;��H;Z�H;��H;��H;      ��H;�H;ƩH;�H;ƬH;��H;��H;g�H;��H;кH;/�H;��H; �H;:�H;^�H;[�H;6�H;��H;H�H;e�H;S�H;��H;m�H;��H;��H;��H;��H;k�H;��H;T�H;��H; �H;9�H;u�H;��H;��H;��H;��H;��H;u�H;9�H; �H;��H;T�H;��H;k�H;��H;��H;��H;��H;m�H;��H;S�H;e�H;H�H;��H;6�H;[�H;^�H;:�H; �H;��H;/�H;кH;��H;g�H;��H;��H;ƬH;�H;ƩH;�H;      ��H;>�H;�H;�H;_�H;*�H;F�H;��H;0�H;��H;��H;l�H;2�H;��H;��H;(�H;��H;��H;��H;^�H;�H;x�H;��H;��H;��H;��H;;�H;��H;L�H;��H;��H;,�H;X�H;��H;��H;��H;��H;��H;��H;��H;X�H;,�H;��H;��H;L�H;��H;;�H;��H;��H;��H;��H;x�H;�H;^�H;��H;��H;��H;(�H;��H;��H;2�H;l�H;��H;��H;0�H;��H;F�H;*�H;_�H;�H;�H;>�H;      �H;�H;��H;��H;��H;{�H;K�H;Y�H;��H;��H;Z�H;��H;I�H;��H;�H;5�H;B�H;0�H;��H;��H;��H;U�H;{�H;i�H;-�H;��H;��H;�H;�H;��H;�H;J�H;��H;��H;��H;��H;��H;��H;��H;��H;��H;J�H;�H;��H;�H;�H;��H;��H;-�H;i�H;{�H;U�H;��H;��H;��H;0�H;B�H;5�H;�H;��H;I�H;��H;Z�H;��H;��H;Y�H;K�H;{�H;��H;��H;��H;�H;      �H;��H;��H;t�H;��H;&�H;��H;��H;�H;a�H;��H;��H;S�H;��H;��H;��H;��H;��H;i�H;��H;Z�H;��H;��H;��H;q�H;�H;��H; �H;��H;��H;0�H;I�H;��H;��H;��H;��H;��H;��H;��H;��H;��H;I�H;0�H;��H;��H; �H;��H;�H;q�H;��H;��H;��H;Z�H;��H;i�H;��H;��H;��H;��H;��H;S�H;��H;��H;a�H;�H;��H;��H;&�H;��H;t�H;��H;��H;      �H;�H;��H;��H;��H;{�H;K�H;Y�H;��H;��H;Z�H;��H;I�H;��H;�H;5�H;B�H;0�H;��H;��H;��H;U�H;{�H;i�H;-�H;��H;��H;�H;�H;��H;�H;J�H;��H;��H;��H;��H;��H;��H;��H;��H;��H;J�H;�H;��H;�H;�H;��H;��H;-�H;i�H;{�H;U�H;��H;��H;��H;0�H;B�H;5�H;�H;��H;I�H;��H;Z�H;��H;��H;Y�H;K�H;{�H;��H;��H;��H;�H;      ��H;>�H;�H;�H;_�H;*�H;F�H;��H;0�H;��H;��H;l�H;2�H;��H;��H;(�H;��H;��H;��H;^�H;�H;x�H;��H;��H;��H;��H;;�H;��H;L�H;��H;��H;,�H;X�H;��H;��H;��H;��H;��H;��H;��H;X�H;,�H;��H;��H;L�H;��H;;�H;��H;��H;��H;��H;x�H;�H;^�H;��H;��H;��H;(�H;��H;��H;2�H;l�H;��H;��H;0�H;��H;F�H;*�H;_�H;�H;�H;>�H;      ��H;�H;ƩH;�H;ƬH;��H;��H;g�H;��H;кH;/�H;��H; �H;:�H;^�H;[�H;6�H;��H;H�H;e�H;S�H;��H;m�H;��H;��H;��H;��H;k�H;��H;T�H;��H; �H;9�H;u�H;��H;��H;��H;��H;��H;u�H;9�H; �H;��H;T�H;��H;k�H;��H;��H;��H;��H;m�H;��H;S�H;e�H;H�H;��H;6�H;[�H;^�H;:�H; �H;��H;/�H;кH;��H;g�H;��H;��H;ƬH;�H;ƩH;�H;      P�H;��H;��H;Z�H;��H;f�H;��H;P�H;.�H;H�H;��H;̸H;�H;>�H;4�H;��H;u�H;��H;��H;i�H;��H;��H;��H;K�H;��H;��H;��H;��H;b�H;�H;h�H;��H;	�H;9�H;X�H;��H;��H;��H;X�H;9�H;	�H;��H;h�H;�H;b�H;��H;��H;��H;��H;K�H;��H;��H;��H;i�H;��H;��H;u�H;��H;4�H;>�H;�H;̸H;��H;H�H;.�H;P�H;��H;f�H;��H;Z�H;��H;��H;      w�H;�H;B�H;u�H;k�H;%�H;p�H;/�H;H�H;��H;&�H;��H;$�H;�H;��H;f�H;��H;��H;��H;B�H;F�H;��H;Q�H;[�H;�H;��H;��H;��H;��H;m�H;�H;z�H;��H; �H;,�H;J�H;I�H;J�H;,�H; �H;��H;z�H;�H;m�H;��H;��H;��H;��H;�H;[�H;Q�H;��H;F�H;B�H;��H;��H;��H;f�H;��H;�H;$�H;��H;&�H;��H;H�H;/�H;p�H;%�H;k�H;u�H;B�H;�H;      fH;�fH;YhH;@kH;(oH;�sH;�yH;�H;��H;ۍH;�H;s�H;��H;��H;#�H;T�H;'�H;��H;x�H;��H;��H;1�H;=�H;��H;��H;��H;X�H;��H;��H;��H;t�H;�H;h�H;��H;��H;�H;0�H;�H;��H;��H;h�H;�H;t�H;��H;��H;��H;X�H;��H;��H;��H;=�H;1�H;��H;��H;x�H;��H;'�H;T�H;#�H;��H;��H;s�H;�H;ۍH;��H;�H;�yH;�sH;(oH;@kH;YhH;�fH;      9?H;@H;cBH;-FH;[KH;�QH;'YH;faH;KjH;�sH;0}H;ʆH;G�H;y�H;8�H;g�H;�H;׸H;�H;��H;��H;7�H;�H;[�H;9�H;��H;��H;L�H;��H;��H;��H;m�H;�H;T�H;��H;��H;��H;��H;��H;T�H;�H;m�H;��H;��H;��H;L�H;��H;��H;9�H;[�H;�H;7�H;��H;��H;�H;׸H;�H;g�H;8�H;y�H;G�H;ʆH;0}H;�sH;KjH;faH;'YH;�QH;[KH;-FH;cBH;@H;      >H;TH;vH;�H;nH;�$H;�.H;�9H;�EH;�QH;k^H;�jH;SwH;W�H;ԎH;��H;��H;��H;��H;ۻH;b�H;�H;��H;"�H;��H;��H;h�H;��H;,�H;��H;��H;��H;b�H;��H;L�H;�H;��H;�H;L�H;��H;b�H;��H;��H;��H;,�H;��H;h�H;��H;��H;"�H;��H;�H;b�H;ۻH;��H;��H;��H;��H;ԎH;W�H;SwH;�jH;k^H;�QH;�EH;�9H;�.H;�$H;nH;�H;vH;TH;      &�G;��G;��G;%�G;�G;5�G;"�G;�H;H;c&H;�6H;�GH;�WH;HgH;)vH;�H;�H;ԜH;T�H;��H;��H;E�H;��H;��H;}�H;k�H;��H;G�H;��H;L�H;��H;��H;��H;k�H;��H;�H; �H;�H;��H;k�H;��H;��H;��H;L�H;��H;G�H;��H;k�H;}�H;��H;��H;E�H;��H;��H;T�H;ԜH;�H;�H;)vH;HgH;�WH;�GH;�6H;c&H;H;�H;"�G;5�G;�G;%�G;��G;��G;      �mG;<pG;wG;�G;��G;^�G;|�G;��G;'�G;M�G;�H;pH;�/H;�CH;@WH;9iH;�yH;�H;��H;ԢH;m�H;��H;��H;��H;@�H;/�H;N�H;��H;h�H;��H;X�H;��H;��H;��H;;�H;��H;��H;��H;;�H;��H;��H;��H;X�H;��H;h�H;��H;N�H;/�H;@�H;��H;��H;��H;m�H;ԢH;��H;�H;�yH;9iH;@WH;�CH;�/H;pH;�H;M�G;'�G;��G;|�G;^�G;��G;�G;wG;<pG;      �F;�F;4�F;��F;,�F;� G;�EG;biG;l�G;,�G;,�G;�G;<�G;�H;�0H;�GH;:]H;�pH;�H;��H;<�H;��H;��H;��H;��H;�H;/�H;k�H;��H;��H;��H;��H;��H;��H;��H;��H;�H;��H;��H;��H;��H;��H;��H;��H;��H;k�H;/�H;�H;��H;��H;��H;��H;<�H;��H;�H;�pH;:]H;�GH;�0H;�H;<�G;�G;,�G;,�G;l�G;biG;�EG;� G;,�F;��F;4�F;�F;      ��D;C�D;B�D;�8E;��E;f�E;�OF;.�F;��F;J9G;mnG;ݙG;�G;��G;� H;�H;�9H;�RH;�hH;e|H;��H;��H;h�H;#�H;U�H;��H;@�H;}�H;��H;9�H;��H;�H;��H;��H;��H;-�H;q�H;-�H;��H;��H;��H;�H;��H;9�H;��H;}�H;@�H;��H;U�H;#�H;h�H;��H;��H;e|H;�hH;�RH;�9H;�H;� H;��G;�G;ݙG;mnG;J9G;��F;.�F;�OF;f�E;��E;�8E;B�D;C�D;      �@;�@@;g�@;]QA;"B;F
C;�C;��D;\�E;�?F;��F;� G;:gG;ÛG;a�G;�G;�H; .H;.JH;�bH;mxH;9�H;P�H;ܨH;#�H;��H;��H;��H;"�H;[�H;��H;[�H;K�H;��H;��H;i�H;��H;i�H;��H;��H;K�H;[�H;��H;[�H;"�H;��H;��H;��H;#�H;ܨH;P�H;9�H;mxH;�bH;.JH; .H;�H;�G;a�G;ÛG;:gG;� G;��F;�?F;\�E;��D;�C;F
C;"B;]QA;g�@;�@@;      �36;˃6;kk7;��8;��:;��<;��>;��@;�sB;��C;�+E;	F;/�F;�+G;�wG;Y�G;��G;�H;%H;7DH;/_H;hvH;O�H;P�H;h�H;��H;��H;��H;��H;�H;=�H;Q�H;��H;m�H;��H;{�H;��H;{�H;��H;m�H;��H;Q�H;=�H;�H;��H;��H;��H;��H;h�H;P�H;O�H;hvH;/_H;7DH;%H;�H;��G;Y�G;�wG;�+G;/�F;	F;�+E;��C;�sB;��@;��>;��<;��:;��8;kk7;˃6;      �";�L#;�%;��';��+;��/;@�3;��7;Q�;;x?;N�A;��C;C9E;�?F;:�F;�TG;��G;T�G;��G;wH;AH;�]H;hvH;9�H;��H;��H;��H;E�H;�H;7�H;1�H;��H;��H;��H;x�H;U�H;��H;U�H;x�H;��H;��H;��H;1�H;7�H;�H;E�H;��H;��H;��H;9�H;hvH;�]H;AH;wH;��G;T�G;��G;�TG;:�F;�?F;C9E;��C;N�A;x?;Q�;;��7;@�3;��/;��+;��';�%;�L#;      ���:�$ ;�;��;��;{P;�l;�c';w�.;�<5;F�:;�>;1B;ZAD;��E;��F;,6G;��G;��G;F�G;�H;AH;/_H;mxH;��H;<�H;m�H;��H;b�H;��H;��H;F�H;��H;S�H;�H;��H;Z�H;��H;�H;S�H;��H;F�H;��H;��H;b�H;��H;m�H;<�H;��H;mxH;/_H;AH;�H;F�G;��G;��G;,6G;��F;��E;ZAD;1B;�>;F�:;�<5;w�.;�c';�l;{P;��;��;�;�$ ;      Y�:�n�:W�:��:�%�:Դ�:���:��	;�P;RM#;�m-;��5;T�;;�@@;�OC;jFE;!uF;!G;��G;�G;F�G;wH;7DH;�bH;e|H;��H;ԢH;��H;ۻH;��H;��H;B�H;i�H;e�H;^�H;��H;��H;��H;^�H;e�H;i�H;B�H;��H;��H;ۻH;��H;ԢH;��H;e|H;�bH;7DH;wH;F�G;�G;��G;!G;!uF;jFE;�OC;�@@;T�;;��5;�m-;RM#;�P;��	;���:Դ�:�%�:��:W�:�n�:      �	�����j��_��3u9�:�i~:���:[�:z�;�;�%;at0;�8;ذ>;Z�B;��D;�WF;sG;��G;��G;��G;%H;.JH;�hH;�H;��H;T�H;��H;�H;x�H;��H;��H;H�H;��H;��H;i�H;��H;��H;H�H;��H;��H;x�H;�H;��H;T�H;��H;�H;�hH;.JH;%H;��G;��G;��G;sG;�WF;��D;Z�B;ذ>;�8;at0;�%;�;z�;[�:���:�i~:�:3u9_���j�����      _A?���9��8)��Z�~ܺkp������H996�@:�:�:��	;�X;�,;8�6;֜=;x"B; �D;�WF;!G;��G;T�G;�H; .H;�RH;�pH;�H;ԜH;��H;׸H;��H;��H;��H;��H;��H;0�H;��H;0�H;��H;��H;��H;��H;��H;׸H;��H;ԜH;�H;�pH;�RH; .H;�H;T�G;��G;!G;�WF; �D;x"B;֜=;8�6;�,;�X;��	;�:�:6�@:H99����kp��~ܺ�Z��8)���9�      �Eֻ�ѻn�Ļ4T��_�q.o���.�ܺ��B�8��8�\:�%�:���:�P;]);�<5;K:=;x"B;��D;!uF;,6G;��G;��G;�H;�9H;:]H;�yH;�H;��H;�H;'�H;��H;u�H;6�H;��H;B�H;��H;B�H;��H;6�H;u�H;��H;'�H;�H;��H;�H;�yH;:]H;�9H;�H;��G;��G;,6G;!uF;��D;x"B;K:=;�<5;]);�P;���:�%�:�\:8��8��B�ܺ��.�q.o�_�4T��n�Ļ�ѻ      FB��>�r�4�$�$�F���Z�ۚ��nݎ�+A?�DӺ����k2�91q�:�W�:�;D�';�<5;֜=;Z�B;jFE;��F;�TG;Y�G;�G;�H;�GH;9iH;�H;��H;g�H;T�H;f�H;��H;[�H;(�H;5�H;��H;5�H;(�H;[�H;��H;f�H;T�H;g�H;��H;�H;9iH;�GH;�H;�G;Y�G;�TG;��F;jFE;Z�B;֜=;�<5;D�';�;�W�:1q�:k2�9����DӺ+A?�nݎ�ۚ���Z�F��$�$�r�4��>�      <y��ݜ��A���I����s�m�P��%+����P�Ļ����|��o��8u9�W�:9+�:�;]);8�6;ذ>;�OC;��E;:�F;�wG;a�G;� H;�0H;@WH;)vH;ԎH;8�H;#�H;��H;4�H;^�H;��H;�H;��H;�H;��H;^�H;4�H;��H;#�H;8�H;ԎH;)vH;@WH;�0H;� H;a�G;�wG;:�F;��E;�OC;ذ>;8�6;]);�;9+�:�W�:�8u9�o�|�����P�Ļ����%+�m�P���s��I���A��ݜ�      -������aW缑�ռ�վ��Τ��I��Z�[��(��Z�g�9��{���99�W�:�W�:�P;�,;�8;�@@;ZAD;�?F;�+G;ÛG;��G;�H;�CH;HgH;W�H;y�H;��H;�H;>�H;:�H;��H;��H;��H;��H;��H;:�H;>�H;�H;��H;y�H;W�H;HgH;�CH;�H;��G;ÛG;�+G;�?F;ZAD;�@@;�8;�,;�P;�W�:�W�:�99�{��g�9���Z��(�Z�[��I���Τ��վ���ռaW缧��      �6��3�X�+�ݟ�<�(�����μ߈��T���FB�=s�	T����D��{���8u91q�:���:�X;at0;T�;;1B;C9E;/�F;:gG;�G;<�G;�/H;�WH;SwH;G�H;��H;$�H;�H; �H;2�H;I�H;S�H;I�H;2�H; �H;�H;$�H;��H;G�H;SwH;�WH;�/H;<�G;�G;:gG;/�F;C9E;1B;T�;;at0;�X;���:1q�:�8u9�{����D�	T��=s�FB�T���߈����μ(���<�ݟ�X�+��3�      R₽�؀���u��Xc�Q�K�K1�{�����վ�t]��b�P�l��	T��g�9��o�k2�9�%�:��	;�%;��5;�>;��C;	F;� G;ݙG;�G;pH;�GH;�jH;ʆH;s�H;��H;̸H;��H;l�H;��H;��H;��H;l�H;��H;̸H;��H;s�H;ʆH;�jH;�GH;pH;�G;ݙG;� G;	F;��C;�>;��5;�%;��	;�%�:k2�9�o�g�9�	T��l��b�P�t]���վ����{��K1�Q�K��Xc���u��؀�      S���r��L��n������|�u�e�N���(�ji���˼�A��b�P�=s��|������\:�:�;�m-;F�:;N�A;�+E;��F;mnG;,�G;�H;�6H;k^H;0}H;�H;&�H;��H;/�H;��H;Z�H;��H;Z�H;��H;/�H;��H;&�H;�H;0}H;k^H;�6H;�H;,�G;mnG;��F;�+E;N�A;F�:;�m-;�;�:�\:����|��=s�b�P��A����˼ji���(�e�N�|�u�����n��L���r��      �o���r���}�ս@��Kĥ�X^���Xc��3���	���˼t]��FB��Z򻆜��DӺ8��8�:z�;RM#;�<5;x?;��C;�?F;J9G;,�G;M�G;c&H;�QH;�sH;ۍH;��H;H�H;кH;��H;��H;a�H;��H;��H;кH;H�H;��H;ۍH;�sH;�QH;c&H;M�G;,�G;J9G;�?F;��C;x?;�<5;RM#;z�;�:8��8DӺ�����Z�FB�t]����˼��	��3��Xc�X^��Kĥ�@��}�ս���r�      �#�6� �A'����~���gٽS��l���j��3�ji��վ�T����(�P�Ļ+A?���B�6�@:[�:�P;w�.;Q�;;�sB;\�E;��F;l�G;'�G;H;�EH;KjH;��H;H�H;.�H;��H;0�H;��H;�H;��H;0�H;��H;.�H;H�H;��H;KjH;�EH;H;'�G;l�G;��F;\�E;�sB;Q�;;w�.;�P;[�:6�@:��B�+A?�P�Ļ�(�T����վ�ji��3��j�l��S���gٽ�~����A'�6� �      �S� �O��E��5�6� �<�
���|9��l���Xc���(����߈��Z�[����nݎ�ܺH99���:��	;�c';��7;��@;��D;.�F;biG;��G;�H;�9H;faH;�H;/�H;P�H;g�H;��H;Y�H;��H;Y�H;��H;g�H;P�H;/�H;�H;faH;�9H;�H;��G;biG;.�F;��D;��@;��7;�c';��	;���:H99ܺnݎ����Z�[�߈�������(��Xc�l��|9����<�
�6� ��5��E� �O�      �~���)����v��9b�U�H��",�0Z���S��X^��e�N�{����μ�I���%+�ۚ����.������i~:���:�l;@�3;��>;�C;�OF;�EG;|�G;"�G;�.H;'YH;�yH;p�H;��H;��H;F�H;K�H;��H;K�H;F�H;��H;��H;p�H;�yH;'YH;�.H;"�G;|�G;�EG;�OF;�C;��>;@�3;�l;���:�i~:������.�ۚ���%+��I����μ{��e�N�X^��S����0Z��",�U�H��9b���v��)��      ��������:���M���r� �O��",�<�
��gٽKĥ�|�u�K1�(����Τ�m�P��Z�q.o�kp���:Դ�:{P;��/;��<;F
C;f�E;� G;^�G;5�G;�$H;�QH;�sH;%�H;f�H;��H;*�H;{�H;&�H;{�H;*�H;��H;f�H;%�H;�sH;�QH;�$H;5�G;^�G;� G;f�E;F
C;��<;��/;{P;Դ�:�:kp��q.o��Z�m�P��Τ�(���K1�|�u�Kĥ��gٽ<�
��",� �O��r��M���:�����      ���v��/;������:P���r�U�H�6� ��~��@������Q�K�<��վ���s�F��_�~ܺ3u9�%�:��;��+;��:;"B;��E;,�F;��G;�G;nH;[KH;(oH;k�H;��H;ƬH;_�H;��H;��H;��H;_�H;ƬH;��H;k�H;(oH;[KH;nH;�G;��G;,�F;��E;"B;��:;��+;��;�%�:3u9~ܺ_�F����s��վ�<�Q�K�����@���~��6� �U�H��r�:P������/;���v��      3Vھ�*־5ʾT��������M���9b��5���}�սn���Xc�ݟ���ռ�I��$�$�4T���Z�_����:��;��';��8;]QA;�8E;��F;�G;%�G;�H;-FH;@kH;u�H;Z�H;�H;�H;��H;t�H;��H;�H;�H;Z�H;u�H;@kH;-FH;�H;%�G;�G;��F;�8E;]QA;��8;��';��;��:_���Z�4T��$�$��I����ռݟ��Xc�n��}�ս���5��9b��M������T���5ʾ�*־      ǰ�쾐�޾5ʾ/;���:����v��E�A'���L����u�X�+�aW缨A��r�4�n�Ļ�8)��j��W�:�;�%;kk7;g�@;B�D;4�F;wG;��G;vH;cBH;YhH;B�H;��H;ƩH;�H;��H;��H;��H;�H;ƩH;��H;B�H;YhH;cBH;vH;��G;wG;4�F;B�D;g�@;kk7;�%;�;W�:�j���8)�n�Ļr�4��A��aW�X�+���u�L����A'��E���v��:��/;��5ʾ��޾��      /h���b���쾅*־�v������)�� �O�6� ��r�r���؀��3����ݜ��>��ѻ��9�����n�:�$ ;�L#;˃6;�@@;C�D;�F;<pG;��G;TH;@H;�fH;�H;��H;�H;>�H;�H;��H;�H;>�H;�H;��H;�H;�fH;@H;TH;��G;<pG;�F;C�D;�@@;˃6;�L#;�$ ;�n�:�����9��ѻ�>�ݜ�����3��؀��r���r�6� � �O��)������v���*־�쾼b��      ����]�0_ݾ��ɾK*��Ы���zx��G�0,�U�뽘b�� @{�|�/�\���䙼�J;��ͻ��4�)Wṻ��:�;]�#;��6;UZ@;��D;��F;�kG;��G;{H;�9H;�aH;�H;M�H;V�H;�H;�H;��H;�H;�H;V�H;M�H;�H;�aH;�9H;{H;��G;�kG;��F;��D;UZ@;��6;]�#;�;���:)Wṫ�4��ͻ�J;��䙼\��|�/� @{��b��U��0,��G��zx�Ы��K*����ɾ0_ݾ�]�      �]����:پZ�žI�������8t�I�C�����罽���`w�-�l���_����7��Rɻ�K/�yƹc��:P/;f$;)7;~@;��D;��F;nG;-�G;gH;�:H;�bH;��H;��H;��H;5�H;M�H;B�H;M�H;5�H;��H;��H;��H;�bH;�:H;gH;-�G;nG;��F;��D;~@;)7;f$;P/;c��:yƹ�K/��Rɻ��7��_��l��-�`w����������I�C��8t����I���Z�ž�:پ��      0_ݾ�:پ�V;�*���Ƥ�3a����g�g$:��Z�?ݽkƣ�Al�:.%��߼=��n9.�����#V�2p��@�:�w;�'&;��7;~�@;P
E;F�F;�tG;Z�G;�
H;=H;|dH;��H;��H;t�H;ֱH;ݷH;عH;ݷH;ֱH;t�H;��H;��H;|dH;=H;�
H;Z�G;�tG;F�F;P
E;~�@;��7;�'&;�w;�@�:2p�#V�����n9.�=���߼:.%�Al�kƣ�?ݽ�Z�g$:���g�3a���Ƥ��*���V;�:پ      ��ɾZ�ž�*��Sת�Ы��	�����T��J+��a2̽ss���yZ����μ>y�����!Ϩ�+,�u��6���:��
;��(;�M9;C�A;�ME;��F;�~G;�G;�H;�@H;agH;�H;`�H;��H;��H;ǸH;��H;ǸH;��H;��H;`�H;�H;agH;�@H;�H;�G;�~G;��F;�ME;C�A;�M9;��(;��
;���:u��6+,�!Ϩ����>y��μ����yZ�ss��a2̽��J+���T�	���Ы��Sת��*��Z�ž      K*��I����Ƥ�Ы���/���c��G=����z�gж��ɇ� �C�����!��);k�z&�|-��F�˺PX�9	��:�8;hh,;8	;;@PB;��E; G;�G;�G;�H;2FH;}kH;/�H;��H;��H;e�H;&�H;��H;&�H;e�H;��H;��H;/�H;}kH;2FH;�H;�G;�G; G;��E;@PB;8	;;hh,;�8;	��:PX�9F�˺|-��z&�);k��!����� �C��ɇ�gж��z����G=��c��/��Ы���Ƥ�I���      Ы�����3a��	����c�J�C�Z#���$vϽ����Al�8g*�T��v
���I�W��p\c��쀺2t,:h��:u�;D_0;��<;�0C;2�E;�"G;}�G;B�G;GH;�LH;fpH;׊H;��H;�H;T�H;��H;��H;��H;T�H;�H;��H;׊H;fpH;�LH;GH;B�G;}�G;�"G;2�E;�0C;��<;D_0;u�;h��:2t,:�쀺p\c�W�軞I�v
��T��8g*�Al�����$vϽ��Z#�J�C��c�	���3a�����      �zx��8t���g���T��G=�Z#��5�?ݽ�b������G������Ǽ>y���$�'����$�!vƹ磆:7&�:2� ;�~4;��>;�D;[F;�EG;��G;:�G;7)H;�TH;%vH;&�H;�H;��H;��H;��H;M�H;��H;��H;��H;�H;&�H;%vH;�TH;7)H;:�G;��G;�EG;[F;�D;��>;�~4;2� ;7&�:磆:!vƹ�$�'����$�>y����Ǽ���G������b��?ݽ�5�Z#��G=���T���g��8t�      �G�I�C�g$:��J+�����?ݽ4���I���yZ�Ơ"�k�鼢���T�Y� ��L��i�˺�m9�ض:�;�_(;}8;��@;��D;'�F;�gG;��G;� H;e4H; ]H;�|H;�H;ۥH;y�H;�H;ʿH;X�H;ʿH;�H;y�H;ۥH;�H;�|H; ]H;e4H;� H;��G;�gG;'�F;��D;��@;}8;�_(;�;�ض:�m9i�˺�L��Y� �T�����k��Ơ"��yZ�I��4���?ݽ�����J+�g$:�I�C�      0,����Z���z�$vϽ�b��I��.]a�-�D� ��!��)�{��!�f���h�4��P(�=nQ:L�:��;H�/;:'<;A�B;=�E;)�F;φG;��G;hH;o@H;=fH;y�H;]�H;�H;��H;��H;�H;u�H;�H;��H;��H;�H;]�H;y�H;=fH;o@H;hH;��G;φG;)�F;=�E;A�B;:'<;H�/;��;L�:=nQ:�P(�h�4�f����!�)�{��!��D� �-�.]a�I���b��$vϽ�z���Z���      U�뽱��?ݽa2̽gж����������yZ�-�����`ļ-O���J;�5��&�|�^�ºHM@9<��:��;Tf$;��5;)N?;�D;�KF;@:G;�G;$�G;� H;MH;�oH;��H;��H;K�H;�H;f�H;��H;��H;��H;f�H;�H;K�H;��H;��H;�oH;MH;� H;$�G;�G;@:G;�KF;�D;)N?;��5;Tf$;��;<��:HM@9^�º&�|�5�軃J;�-O���`ļ���-��yZ���������gж�a2̽?ݽ���      �b������kƣ�ss���ɇ�Al�G�Ơ"�D� ��`ļ6���I��C��ۙ��Suƹ��k:��:��;�=.;|	;;*�A;.AE;��F;OlG;��G;��G;�1H;ZH;�yH;�H;��H;��H;|�H;O�H;�H;3�H;�H;O�H;|�H;��H;��H;�H;�yH;ZH;�1H;��G;��G;OlG;��F;.AE;*�A;|	;;�=.;��;��:��k:Suƹ��ۙ��C��I�6���`ļD� �Ơ"�G�Al��ɇ�ss��kƣ�����       @{�`w�Al��yZ� �C�8g*����k���!��-O���I�|��Ψ�3K/�`$T��P:���:3�;6(&;]#6;%?;��C;�"F;9#G;^�G;��G;�H;XBH;gH;��H;��H;��H;�H;�H;?�H;��H;��H;��H;?�H;�H;�H;��H;��H;��H;gH;XBH;�H;��G;^�G;9#G;�"F;��C;%?;]#6;6(&;3�;���:�P:`$T�3K/��Ψ�|��I�-O���!��k�鼇��8g*� �C��yZ�Al�`w�      |�/�-�:.%�������T���Ǽ����)�{��J;��C��Ψ�
O:�����zZ�9M��:;�;�-1;k'<;$5B;%NE;Z�F;jeG;�G;h�G;"*H;
SH;�sH;F�H;�H;@�H;i�H;��H;�H;�H;=�H;�H;�H;��H;i�H;@�H;�H;F�H;�sH;
SH;"*H;h�G;�G;jeG;Z�F;%NE;$5B;k'<;�-1;�;;M��:zZ�9����
O:��Ψ��C��J;�)�{�������ǼT��������:.%�-�      \��l�鼟߼μ�!��v
��>y��T��!�5�軉ۙ�3K/�����pm9pA�:���:ƽ;��,;,N9;�~@;^D;
LF;�-G;�G;��G;�H;�>H;CcH;<�H;��H;+�H;��H;��H;��H;��H;��H;��H;��H;��H;��H;��H;��H;+�H;��H;<�H;CcH;�>H;�H;��G;�G;�-G;
LF;^D;�~@;,N9;��,;ƽ;���:pA�:pm9����3K/��ۙ�5���!�T�>y��v
���!��μ�߼l��      �䙼�_��=��>y��);k��I��$�Y� �f���&�|��`$T�zZ�9pA�:���:��;��);�7;=�>; tC;_�E;1�F;%uG;O�G;��G;/+H;�RH;�rH;��H;��H;0�H;�H;��H;S�H;��H;�H;��H;�H;��H;S�H;��H;�H;0�H;��H;��H;�rH;�RH;/+H;��G;O�G;%uG;1�F;_�E; tC;=�>;�7;��);��;���:pA�:zZ�9`$T��&�|�f���Y� ��$��I�);k�>y��=���_��      �J;���7�n9.����z&�W��'����L��h�4�^�ºSuƹ�P:M��:���:��;-�(;-�5;#�=;�B;�ZE;��F;TG;�G;��G;�H;�BH;9eH;�H;��H;�H;��H;�H;��H;p�H;�H;R�H;9�H;R�H;�H;p�H;��H;�H;��H;�H;��H;�H;9eH;�BH;�H;��G;�G;TG;��F;�ZE;�B;#�=;-�5;-�(;��;���:M��:�P:Suƹ^�ºh�4��L��'���W��z&����n9.���7�      �ͻ�Rɻ����!Ϩ�|-��p\c��$�i�˺�P(�HM@9��k:���:;ƽ;��);-�5;��=;vPB;�
E;5F;d7G;z�G;|�G;�H;�4H;�XH;gvH;��H;ѠH;�H;��H;��H;l�H;<�H;��H;��H;9�H;��H;��H;<�H;l�H;��H;��H;�H;ѠH;��H;gvH;�XH;�4H;�H;|�G;z�G;d7G;5F;�
E;vPB;��=;-�5;��);ƽ;;���:��k:HM@9�P(�i�˺�$�p\c�|-��!Ϩ������Rɻ      ��4��K/�#V�+,�F�˺�쀺!vƹ�m9=nQ:<��:��:3�;�;��,;�7;#�=;vPB;�D;�bF;]#G;�G;�G;�G;�(H;�MH;�lH;��H;�H;E�H;-�H;-�H;��H;��H;��H;��H;��H;'�H;��H;��H;��H;��H;��H;-�H;-�H;E�H;�H;��H;�lH;�MH;�(H;�G;�G;�G;]#G;�bF;�D;vPB;#�=;�7;��,;�;3�;��:<��:=nQ:�m9!vƹ�쀺F�˺+,�#V��K/�      )W�yƹ2p�u��6PX�92t,:磆:�ض:L�:��;��;6(&;�-1;,N9;=�>;�B;�
E;�bF;+G;eG;�G;��G;�H;EH;�dH;�~H;ړH;�H;ҲH;��H;(�H;��H;��H;g�H;�H;Z�H;��H;Z�H;�H;g�H;��H;��H;(�H;��H;ҲH;�H;ړH;�~H;�dH;EH;�H;��G;�G;eG;+G;�bF;�
E;�B;=�>;,N9;�-1;6(&;��;��;L�:�ض:磆:2t,:PX�9u��62p�yƹ      ���:c��:�@�:���:	��:h��:7&�:�;��;Tf$;�=.;]#6;k'<;�~@; tC;�ZE;5F;]#G;eG;�G;L�G;�H;?H;�^H;yH;y�H;<�H;ѮH;J�H;��H;��H;d�H;��H;��H;��H;�H;|�H;�H;��H;��H;��H;d�H;��H;��H;J�H;ѮH;<�H;y�H;yH;�^H;?H;�H;L�G;�G;eG;]#G;5F;�ZE; tC;�~@;k'<;]#6;�=.;Tf$;��;�;7&�:h��:	��:���:�@�:c��:      �;P/;�w;��
;�8;u�;2� ;�_(;H�/;��5;|	;;%?;$5B;^D;_�E;��F;d7G;�G;�G;L�G;�H;�;H;�ZH;
uH;��H;p�H;U�H;U�H;��H;��H;��H;~�H;�H;��H;��H;��H;��H;��H;��H;��H;�H;~�H;��H;��H;��H;U�H;U�H;p�H;��H;
uH;�ZH;�;H;�H;L�G;�G;�G;d7G;��F;_�E;^D;$5B;%?;|	;;��5;H�/;�_(;2� ;u�;�8;��
;�w;P/;      ]�#;f$;�'&;��(;hh,;D_0;�~4;}8;:'<;)N?;*�A;��C;%NE;
LF;1�F;TG;z�G;�G;��G;�H;�;H;�YH;sH;�H;��H;��H;�H;�H;��H;)�H;Q�H;F�H;e�H;��H;��H;��H;%�H;��H;��H;��H;e�H;F�H;Q�H;)�H;��H;�H;�H;��H;��H;�H;sH;�YH;�;H;�H;��G;�G;z�G;TG;1�F;
LF;%NE;��C;*�A;)N?;:'<;}8;�~4;D_0;hh,;��(;�'&;f$;      ��6;)7;��7;�M9;8	;;��<;��>;��@;A�B;�D;.AE;�"F;Z�F;�-G;%uG;�G;|�G;�G;�H;?H;�ZH;sH;V�H;r�H;�H;?�H;�H;;�H;�H;4�H;d�H;��H;U�H;>�H;G�H;�H;@�H;�H;G�H;>�H;U�H;��H;d�H;4�H;�H;;�H;�H;?�H;�H;r�H;V�H;sH;�ZH;?H;�H;�G;|�G;�G;%uG;�-G;Z�F;�"F;.AE;�D;A�B;��@;��>;��<;8	;;�M9;��7;)7;      UZ@;~@;~�@;C�A;@PB;�0C;�D;��D;=�E;�KF;��F;9#G;jeG;�G;O�G;��G;�H;�(H;EH;�^H;
uH;�H;r�H;}�H;W�H;/�H;@�H;��H;c�H;��H;�H;��H;��H;x�H;t�H;
�H;Q�H;
�H;t�H;x�H;��H;��H;�H;��H;c�H;��H;@�H;/�H;W�H;}�H;r�H;�H;
uH;�^H;EH;�(H;�H;��G;O�G;�G;jeG;9#G;��F;�KF;=�E;��D;�D;�0C;@PB;C�A;~�@;~@;      ��D;��D;P
E;�ME;��E;2�E;[F;'�F;)�F;@:G;OlG;^�G;�G;��G;��G;�H;�4H;�MH;�dH;yH;��H;��H;�H;W�H;��H;��H;=�H;��H;�H;��H;c�H;��H;b�H;��H;��H;��H;�H;��H;��H;��H;b�H;��H;c�H;��H;�H;��H;=�H;��H;��H;W�H;�H;��H;��H;yH;�dH;�MH;�4H;�H;��G;��G;�G;^�G;OlG;@:G;)�F;'�F;[F;2�E;��E;�ME;P
E;��D;      ��F;��F;F�F;��F; G;�"G;�EG;�gG;φG;�G;��G;��G;h�G;�H;/+H;�BH;�XH;�lH;�~H;y�H;p�H;��H;?�H;/�H;��H;�H;H�H;��H;#�H;)�H;k�H;�H;��H;��H;f�H;��H;��H;��H;f�H;��H;��H;�H;k�H;)�H;#�H;��H;H�H;�H;��H;/�H;?�H;��H;p�H;y�H;�~H;�lH;�XH;�BH;/+H;�H;h�G;��G;��G;�G;φG;�gG;�EG;�"G; G;��F;F�F;��F;      �kG;nG;�tG;�~G;�G;}�G;��G;��G;��G;$�G;��G;�H;"*H;�>H;�RH;9eH;gvH;��H;ړH;<�H;U�H;�H;�H;@�H;=�H;H�H;e�H;��H;��H;5�H;*�H;t�H;��H;x�H;�H;d�H;��H;d�H;�H;x�H;��H;t�H;*�H;5�H;��H;��H;e�H;H�H;=�H;@�H;�H;�H;U�H;<�H;ړH;��H;gvH;9eH;�RH;�>H;"*H;�H;��G;$�G;��G;��G;��G;}�G;�G;�~G;�tG;nG;      ��G;-�G;Z�G;�G;�G;B�G;:�G;� H;hH;� H;�1H;XBH;
SH;CcH;�rH;�H;��H;�H;�H;ѮH;U�H;�H;;�H;��H;��H;��H;��H;��H;�H;��H;q�H;��H;��H;B�H;��H;��H;#�H;��H;��H;B�H;��H;��H;q�H;��H;�H;��H;��H;��H;��H;��H;;�H;�H;U�H;ѮH;�H;�H;��H;�H;�rH;CcH;
SH;XBH;�1H;� H;hH;� H;:�G;B�G;�G;�G;Z�G;-�G;      {H;gH;�
H;�H;�H;GH;7)H;e4H;o@H;MH;ZH;gH;�sH;<�H;��H;��H;ѠH;E�H;ҲH;J�H;��H;��H;�H;c�H;�H;#�H;��H;�H;��H;V�H;�H;��H;A�H;��H;�H;V�H;b�H;V�H;�H;��H;A�H;��H;�H;V�H;��H;�H;��H;#�H;�H;c�H;�H;��H;��H;J�H;ҲH;E�H;ѠH;��H;��H;<�H;�sH;gH;ZH;MH;o@H;e4H;7)H;GH;�H;�H;�
H;gH;      �9H;�:H;=H;�@H;2FH;�LH;�TH; ]H;=fH;�oH;�yH;��H;F�H;��H;��H;�H;�H;-�H;��H;��H;��H;)�H;4�H;��H;��H;)�H;5�H;��H;V�H;��H;w�H;1�H;��H;8�H;��H;��H;��H;��H;��H;8�H;��H;1�H;w�H;��H;V�H;��H;5�H;)�H;��H;��H;4�H;)�H;��H;��H;��H;-�H;�H;�H;��H;��H;F�H;��H;�yH;�oH;=fH; ]H;�TH;�LH;2FH;�@H;=H;�:H;      �aH;�bH;|dH;agH;}kH;fpH;%vH;�|H;y�H;��H;�H;��H;�H;+�H;0�H;��H;��H;-�H;(�H;��H;��H;Q�H;d�H;�H;c�H;k�H;*�H;q�H;�H;w�H;H�H;��H;2�H;��H;��H;��H;�H;��H;��H;��H;2�H;��H;H�H;w�H;�H;q�H;*�H;k�H;c�H;�H;d�H;Q�H;��H;��H;(�H;-�H;��H;��H;0�H;+�H;�H;��H;�H;��H;y�H;�|H;%vH;fpH;}kH;agH;|dH;�bH;      �H;��H;��H;�H;/�H;׊H;&�H;�H;]�H;��H;��H;��H;@�H;��H;�H;�H;��H;��H;��H;d�H;~�H;F�H;��H;��H;��H;�H;t�H;��H;��H;1�H;��H;B�H;��H;��H;�H;C�H;5�H;C�H;�H;��H;��H;B�H;��H;1�H;��H;��H;t�H;�H;��H;��H;��H;F�H;~�H;d�H;��H;��H;��H;�H;�H;��H;@�H;��H;��H;��H;]�H;�H;&�H;׊H;/�H;�H;��H;��H;      M�H;��H;��H;`�H;��H;��H;�H;ۥH;�H;K�H;��H;�H;i�H;��H;��H;��H;l�H;��H;��H;��H;�H;e�H;U�H;��H;b�H;��H;��H;��H;A�H;��H;2�H;��H;�H;�H;V�H;l�H;7�H;l�H;V�H;�H;�H;��H;2�H;��H;A�H;��H;��H;��H;b�H;��H;U�H;e�H;�H;��H;��H;��H;l�H;��H;��H;��H;i�H;�H;��H;K�H;�H;ۥH;�H;��H;��H;`�H;��H;��H;      V�H;��H;t�H;��H;��H;�H;��H;y�H;��H;�H;|�H;�H;��H;��H;S�H;p�H;<�H;��H;g�H;��H;��H;��H;>�H;x�H;��H;��H;x�H;B�H;��H;8�H;��H;��H;�H;M�H;m�H;y�H;��H;y�H;m�H;M�H;�H;��H;��H;8�H;��H;B�H;x�H;��H;��H;x�H;>�H;��H;��H;��H;g�H;��H;<�H;p�H;S�H;��H;��H;�H;|�H;�H;��H;y�H;��H;�H;��H;��H;t�H;��H;      �H;5�H;ֱH;��H;e�H;T�H;��H;�H;��H;f�H;O�H;?�H;�H;��H;��H;�H;��H;��H;�H;��H;��H;��H;G�H;t�H;��H;f�H;�H;��H;�H;��H;��H;�H;V�H;m�H;u�H;��H;��H;��H;u�H;m�H;V�H;�H;��H;��H;�H;��H;�H;f�H;��H;t�H;G�H;��H;��H;��H;�H;��H;��H;�H;��H;��H;�H;?�H;O�H;f�H;��H;�H;��H;T�H;e�H;��H;ֱH;5�H;      �H;M�H;ݷH;ǸH;&�H;��H;��H;ʿH;�H;��H;�H;��H;�H;��H;�H;R�H;��H;��H;Z�H;�H;��H;��H;�H;
�H;��H;��H;d�H;��H;V�H;��H;��H;C�H;l�H;y�H;��H;��H;��H;��H;��H;y�H;l�H;C�H;��H;��H;V�H;��H;d�H;��H;��H;
�H;�H;��H;��H;�H;Z�H;��H;��H;R�H;�H;��H;�H;��H;�H;��H;�H;ʿH;��H;��H;&�H;ǸH;ݷH;M�H;      ��H;B�H;عH;��H;��H;��H;M�H;X�H;u�H;��H;3�H;��H;=�H;��H;��H;9�H;9�H;'�H;��H;|�H;��H;%�H;@�H;Q�H;�H;��H;��H;#�H;b�H;��H;�H;5�H;7�H;��H;��H;��H;��H;��H;��H;��H;7�H;5�H;�H;��H;b�H;#�H;��H;��H;�H;Q�H;@�H;%�H;��H;|�H;��H;'�H;9�H;9�H;��H;��H;=�H;��H;3�H;��H;u�H;X�H;M�H;��H;��H;��H;عH;B�H;      �H;M�H;ݷH;ǸH;&�H;��H;��H;ʿH;�H;��H;�H;��H;�H;��H;�H;R�H;��H;��H;Z�H;�H;��H;��H;�H;
�H;��H;��H;d�H;��H;V�H;��H;��H;C�H;l�H;y�H;��H;��H;��H;��H;��H;y�H;l�H;C�H;��H;��H;V�H;��H;d�H;��H;��H;
�H;�H;��H;��H;�H;Z�H;��H;��H;R�H;�H;��H;�H;��H;�H;��H;�H;ʿH;��H;��H;&�H;ǸH;ݷH;M�H;      �H;5�H;ֱH;��H;e�H;T�H;��H;�H;��H;f�H;O�H;?�H;�H;��H;��H;�H;��H;��H;�H;��H;��H;��H;G�H;t�H;��H;f�H;�H;��H;�H;��H;��H;�H;V�H;m�H;u�H;��H;��H;��H;u�H;m�H;V�H;�H;��H;��H;�H;��H;�H;f�H;��H;t�H;G�H;��H;��H;��H;�H;��H;��H;�H;��H;��H;�H;?�H;O�H;f�H;��H;�H;��H;T�H;e�H;��H;ֱH;5�H;      V�H;��H;t�H;��H;��H;�H;��H;y�H;��H;�H;|�H;�H;��H;��H;S�H;p�H;<�H;��H;g�H;��H;��H;��H;>�H;x�H;��H;��H;x�H;B�H;��H;8�H;��H;��H;�H;M�H;m�H;y�H;��H;y�H;m�H;M�H;�H;��H;��H;8�H;��H;B�H;x�H;��H;��H;x�H;>�H;��H;��H;��H;g�H;��H;<�H;p�H;S�H;��H;��H;�H;|�H;�H;��H;y�H;��H;�H;��H;��H;t�H;��H;      M�H;��H;��H;`�H;��H;��H;�H;ۥH;�H;K�H;��H;�H;i�H;��H;��H;��H;l�H;��H;��H;��H;�H;e�H;U�H;��H;b�H;��H;��H;��H;A�H;��H;2�H;��H;�H;�H;V�H;l�H;7�H;l�H;V�H;�H;�H;��H;2�H;��H;A�H;��H;��H;��H;b�H;��H;U�H;e�H;�H;��H;��H;��H;l�H;��H;��H;��H;i�H;�H;��H;K�H;�H;ۥH;�H;��H;��H;`�H;��H;��H;      �H;��H;��H;�H;/�H;׊H;&�H;�H;]�H;��H;��H;��H;@�H;��H;�H;�H;��H;��H;��H;d�H;~�H;F�H;��H;��H;��H;�H;t�H;��H;��H;1�H;��H;B�H;��H;��H;�H;C�H;5�H;C�H;�H;��H;��H;B�H;��H;1�H;��H;��H;t�H;�H;��H;��H;��H;F�H;~�H;d�H;��H;��H;��H;�H;�H;��H;@�H;��H;��H;��H;]�H;�H;&�H;׊H;/�H;�H;��H;��H;      �aH;�bH;|dH;agH;}kH;fpH;%vH;�|H;y�H;��H;�H;��H;�H;+�H;0�H;��H;��H;-�H;(�H;��H;��H;Q�H;d�H;�H;c�H;k�H;*�H;q�H;�H;w�H;H�H;��H;2�H;��H;��H;��H;�H;��H;��H;��H;2�H;��H;H�H;w�H;�H;q�H;*�H;k�H;c�H;�H;d�H;Q�H;��H;��H;(�H;-�H;��H;��H;0�H;+�H;�H;��H;�H;��H;y�H;�|H;%vH;fpH;}kH;agH;|dH;�bH;      �9H;�:H;=H;�@H;2FH;�LH;�TH; ]H;=fH;�oH;�yH;��H;F�H;��H;��H;�H;�H;-�H;��H;��H;��H;)�H;4�H;��H;��H;)�H;5�H;��H;V�H;��H;w�H;1�H;��H;8�H;��H;��H;��H;��H;��H;8�H;��H;1�H;w�H;��H;V�H;��H;5�H;)�H;��H;��H;4�H;)�H;��H;��H;��H;-�H;�H;�H;��H;��H;F�H;��H;�yH;�oH;=fH; ]H;�TH;�LH;2FH;�@H;=H;�:H;      {H;gH;�
H;�H;�H;GH;7)H;e4H;o@H;MH;ZH;gH;�sH;<�H;��H;��H;ѠH;E�H;ҲH;J�H;��H;��H;�H;c�H;�H;#�H;��H;�H;��H;V�H;�H;��H;A�H;��H;�H;V�H;b�H;V�H;�H;��H;A�H;��H;�H;V�H;��H;�H;��H;#�H;�H;c�H;�H;��H;��H;J�H;ҲH;E�H;ѠH;��H;��H;<�H;�sH;gH;ZH;MH;o@H;e4H;7)H;GH;�H;�H;�
H;gH;      ��G;-�G;Z�G;�G;�G;B�G;:�G;� H;hH;� H;�1H;XBH;
SH;CcH;�rH;�H;��H;�H;�H;ѮH;U�H;�H;;�H;��H;��H;��H;��H;��H;�H;��H;q�H;��H;��H;B�H;��H;��H;#�H;��H;��H;B�H;��H;��H;q�H;��H;�H;��H;��H;��H;��H;��H;;�H;�H;U�H;ѮH;�H;�H;��H;�H;�rH;CcH;
SH;XBH;�1H;� H;hH;� H;:�G;B�G;�G;�G;Z�G;-�G;      �kG;nG;�tG;�~G;�G;}�G;��G;��G;��G;$�G;��G;�H;"*H;�>H;�RH;9eH;gvH;��H;ړH;<�H;U�H;�H;�H;@�H;=�H;H�H;e�H;��H;��H;5�H;*�H;t�H;��H;x�H;�H;d�H;��H;d�H;�H;x�H;��H;t�H;*�H;5�H;��H;��H;e�H;H�H;=�H;@�H;�H;�H;U�H;<�H;ړH;��H;gvH;9eH;�RH;�>H;"*H;�H;��G;$�G;��G;��G;��G;}�G;�G;�~G;�tG;nG;      ��F;��F;F�F;��F; G;�"G;�EG;�gG;φG;�G;��G;��G;h�G;�H;/+H;�BH;�XH;�lH;�~H;y�H;p�H;��H;?�H;/�H;��H;�H;H�H;��H;#�H;)�H;k�H;�H;��H;��H;f�H;��H;��H;��H;f�H;��H;��H;�H;k�H;)�H;#�H;��H;H�H;�H;��H;/�H;?�H;��H;p�H;y�H;�~H;�lH;�XH;�BH;/+H;�H;h�G;��G;��G;�G;φG;�gG;�EG;�"G; G;��F;F�F;��F;      ��D;��D;P
E;�ME;��E;2�E;[F;'�F;)�F;@:G;OlG;^�G;�G;��G;��G;�H;�4H;�MH;�dH;yH;��H;��H;�H;W�H;��H;��H;=�H;��H;�H;��H;c�H;��H;b�H;��H;��H;��H;�H;��H;��H;��H;b�H;��H;c�H;��H;�H;��H;=�H;��H;��H;W�H;�H;��H;��H;yH;�dH;�MH;�4H;�H;��G;��G;�G;^�G;OlG;@:G;)�F;'�F;[F;2�E;��E;�ME;P
E;��D;      UZ@;~@;~�@;C�A;@PB;�0C;�D;��D;=�E;�KF;��F;9#G;jeG;�G;O�G;��G;�H;�(H;EH;�^H;
uH;�H;r�H;}�H;W�H;/�H;@�H;��H;c�H;��H;�H;��H;��H;x�H;t�H;
�H;Q�H;
�H;t�H;x�H;��H;��H;�H;��H;c�H;��H;@�H;/�H;W�H;}�H;r�H;�H;
uH;�^H;EH;�(H;�H;��G;O�G;�G;jeG;9#G;��F;�KF;=�E;��D;�D;�0C;@PB;C�A;~�@;~@;      ��6;)7;��7;�M9;8	;;��<;��>;��@;A�B;�D;.AE;�"F;Z�F;�-G;%uG;�G;|�G;�G;�H;?H;�ZH;sH;V�H;r�H;�H;?�H;�H;;�H;�H;4�H;d�H;��H;U�H;>�H;G�H;�H;@�H;�H;G�H;>�H;U�H;��H;d�H;4�H;�H;;�H;�H;?�H;�H;r�H;V�H;sH;�ZH;?H;�H;�G;|�G;�G;%uG;�-G;Z�F;�"F;.AE;�D;A�B;��@;��>;��<;8	;;�M9;��7;)7;      ]�#;f$;�'&;��(;hh,;D_0;�~4;}8;:'<;)N?;*�A;��C;%NE;
LF;1�F;TG;z�G;�G;��G;�H;�;H;�YH;sH;�H;��H;��H;�H;�H;��H;)�H;Q�H;F�H;e�H;��H;��H;��H;%�H;��H;��H;��H;e�H;F�H;Q�H;)�H;��H;�H;�H;��H;��H;�H;sH;�YH;�;H;�H;��G;�G;z�G;TG;1�F;
LF;%NE;��C;*�A;)N?;:'<;}8;�~4;D_0;hh,;��(;�'&;f$;      �;P/;�w;��
;�8;u�;2� ;�_(;H�/;��5;|	;;%?;$5B;^D;_�E;��F;d7G;�G;�G;L�G;�H;�;H;�ZH;
uH;��H;p�H;U�H;U�H;��H;��H;��H;~�H;�H;��H;��H;��H;��H;��H;��H;��H;�H;~�H;��H;��H;��H;U�H;U�H;p�H;��H;
uH;�ZH;�;H;�H;L�G;�G;�G;d7G;��F;_�E;^D;$5B;%?;|	;;��5;H�/;�_(;2� ;u�;�8;��
;�w;P/;      ���:c��:�@�:���:	��:h��:7&�:�;��;Tf$;�=.;]#6;k'<;�~@; tC;�ZE;5F;]#G;eG;�G;L�G;�H;?H;�^H;yH;y�H;<�H;ѮH;J�H;��H;��H;d�H;��H;��H;��H;�H;|�H;�H;��H;��H;��H;d�H;��H;��H;J�H;ѮH;<�H;y�H;yH;�^H;?H;�H;L�G;�G;eG;]#G;5F;�ZE; tC;�~@;k'<;]#6;�=.;Tf$;��;�;7&�:h��:	��:���:�@�:c��:      )W�yƹ2p�u��6PX�92t,:磆:�ض:L�:��;��;6(&;�-1;,N9;=�>;�B;�
E;�bF;+G;eG;�G;��G;�H;EH;�dH;�~H;ړH;�H;ҲH;��H;(�H;��H;��H;g�H;�H;Z�H;��H;Z�H;�H;g�H;��H;��H;(�H;��H;ҲH;�H;ړH;�~H;�dH;EH;�H;��G;�G;eG;+G;�bF;�
E;�B;=�>;,N9;�-1;6(&;��;��;L�:�ض:磆:2t,:PX�9u��62p�yƹ      ��4��K/�#V�+,�F�˺�쀺!vƹ�m9=nQ:<��:��:3�;�;��,;�7;#�=;vPB;�D;�bF;]#G;�G;�G;�G;�(H;�MH;�lH;��H;�H;E�H;-�H;-�H;��H;��H;��H;��H;��H;'�H;��H;��H;��H;��H;��H;-�H;-�H;E�H;�H;��H;�lH;�MH;�(H;�G;�G;�G;]#G;�bF;�D;vPB;#�=;�7;��,;�;3�;��:<��:=nQ:�m9!vƹ�쀺F�˺+,�#V��K/�      �ͻ�Rɻ����!Ϩ�|-��p\c��$�i�˺�P(�HM@9��k:���:;ƽ;��);-�5;��=;vPB;�
E;5F;d7G;z�G;|�G;�H;�4H;�XH;gvH;��H;ѠH;�H;��H;��H;l�H;<�H;��H;��H;9�H;��H;��H;<�H;l�H;��H;��H;�H;ѠH;��H;gvH;�XH;�4H;�H;|�G;z�G;d7G;5F;�
E;vPB;��=;-�5;��);ƽ;;���:��k:HM@9�P(�i�˺�$�p\c�|-��!Ϩ������Rɻ      �J;���7�n9.����z&�W��'����L��h�4�^�ºSuƹ�P:M��:���:��;-�(;-�5;#�=;�B;�ZE;��F;TG;�G;��G;�H;�BH;9eH;�H;��H;�H;��H;�H;��H;p�H;�H;R�H;9�H;R�H;�H;p�H;��H;�H;��H;�H;��H;�H;9eH;�BH;�H;��G;�G;TG;��F;�ZE;�B;#�=;-�5;-�(;��;���:M��:�P:Suƹ^�ºh�4��L��'���W��z&����n9.���7�      �䙼�_��=��>y��);k��I��$�Y� �f���&�|��`$T�zZ�9pA�:���:��;��);�7;=�>; tC;_�E;1�F;%uG;O�G;��G;/+H;�RH;�rH;��H;��H;0�H;�H;��H;S�H;��H;�H;��H;�H;��H;S�H;��H;�H;0�H;��H;��H;�rH;�RH;/+H;��G;O�G;%uG;1�F;_�E; tC;=�>;�7;��);��;���:pA�:zZ�9`$T��&�|�f���Y� ��$��I�);k�>y��=���_��      \��l�鼟߼μ�!��v
��>y��T��!�5�軉ۙ�3K/�����pm9pA�:���:ƽ;��,;,N9;�~@;^D;
LF;�-G;�G;��G;�H;�>H;CcH;<�H;��H;+�H;��H;��H;��H;��H;��H;��H;��H;��H;��H;��H;��H;+�H;��H;<�H;CcH;�>H;�H;��G;�G;�-G;
LF;^D;�~@;,N9;��,;ƽ;���:pA�:pm9����3K/��ۙ�5���!�T�>y��v
���!��μ�߼l��      |�/�-�:.%�������T���Ǽ����)�{��J;��C��Ψ�
O:�����zZ�9M��:;�;�-1;k'<;$5B;%NE;Z�F;jeG;�G;h�G;"*H;
SH;�sH;F�H;�H;@�H;i�H;��H;�H;�H;=�H;�H;�H;��H;i�H;@�H;�H;F�H;�sH;
SH;"*H;h�G;�G;jeG;Z�F;%NE;$5B;k'<;�-1;�;;M��:zZ�9����
O:��Ψ��C��J;�)�{�������ǼT��������:.%�-�       @{�`w�Al��yZ� �C�8g*����k���!��-O���I�|��Ψ�3K/�`$T��P:���:3�;6(&;]#6;%?;��C;�"F;9#G;^�G;��G;�H;XBH;gH;��H;��H;��H;�H;�H;?�H;��H;��H;��H;?�H;�H;�H;��H;��H;��H;gH;XBH;�H;��G;^�G;9#G;�"F;��C;%?;]#6;6(&;3�;���:�P:`$T�3K/��Ψ�|��I�-O���!��k�鼇��8g*� �C��yZ�Al�`w�      �b������kƣ�ss���ɇ�Al�G�Ơ"�D� ��`ļ6���I��C��ۙ��Suƹ��k:��:��;�=.;|	;;*�A;.AE;��F;OlG;��G;��G;�1H;ZH;�yH;�H;��H;��H;|�H;O�H;�H;3�H;�H;O�H;|�H;��H;��H;�H;�yH;ZH;�1H;��G;��G;OlG;��F;.AE;*�A;|	;;�=.;��;��:��k:Suƹ��ۙ��C��I�6���`ļD� �Ơ"�G�Al��ɇ�ss��kƣ�����      U�뽱��?ݽa2̽gж����������yZ�-�����`ļ-O���J;�5��&�|�^�ºHM@9<��:��;Tf$;��5;)N?;�D;�KF;@:G;�G;$�G;� H;MH;�oH;��H;��H;K�H;�H;f�H;��H;��H;��H;f�H;�H;K�H;��H;��H;�oH;MH;� H;$�G;�G;@:G;�KF;�D;)N?;��5;Tf$;��;<��:HM@9^�º&�|�5�軃J;�-O���`ļ���-��yZ���������gж�a2̽?ݽ���      0,����Z���z�$vϽ�b��I��.]a�-�D� ��!��)�{��!�f���h�4��P(�=nQ:L�:��;H�/;:'<;A�B;=�E;)�F;φG;��G;hH;o@H;=fH;y�H;]�H;�H;��H;��H;�H;u�H;�H;��H;��H;�H;]�H;y�H;=fH;o@H;hH;��G;φG;)�F;=�E;A�B;:'<;H�/;��;L�:=nQ:�P(�h�4�f����!�)�{��!��D� �-�.]a�I���b��$vϽ�z���Z���      �G�I�C�g$:��J+�����?ݽ4���I���yZ�Ơ"�k�鼢���T�Y� ��L��i�˺�m9�ض:�;�_(;}8;��@;��D;'�F;�gG;��G;� H;e4H; ]H;�|H;�H;ۥH;y�H;�H;ʿH;X�H;ʿH;�H;y�H;ۥH;�H;�|H; ]H;e4H;� H;��G;�gG;'�F;��D;��@;}8;�_(;�;�ض:�m9i�˺�L��Y� �T�����k��Ơ"��yZ�I��4���?ݽ�����J+�g$:�I�C�      �zx��8t���g���T��G=�Z#��5�?ݽ�b������G������Ǽ>y���$�'����$�!vƹ磆:7&�:2� ;�~4;��>;�D;[F;�EG;��G;:�G;7)H;�TH;%vH;&�H;�H;��H;��H;��H;M�H;��H;��H;��H;�H;&�H;%vH;�TH;7)H;:�G;��G;�EG;[F;�D;��>;�~4;2� ;7&�:磆:!vƹ�$�'����$�>y����Ǽ���G������b��?ݽ�5�Z#��G=���T���g��8t�      Ы�����3a��	����c�J�C�Z#���$vϽ����Al�8g*�T��v
���I�W��p\c��쀺2t,:h��:u�;D_0;��<;�0C;2�E;�"G;}�G;B�G;GH;�LH;fpH;׊H;��H;�H;T�H;��H;��H;��H;T�H;�H;��H;׊H;fpH;�LH;GH;B�G;}�G;�"G;2�E;�0C;��<;D_0;u�;h��:2t,:�쀺p\c�W�軞I�v
��T��8g*�Al�����$vϽ��Z#�J�C��c�	���3a�����      K*��I����Ƥ�Ы���/���c��G=����z�gж��ɇ� �C�����!��);k�z&�|-��F�˺PX�9	��:�8;hh,;8	;;@PB;��E; G;�G;�G;�H;2FH;}kH;/�H;��H;��H;e�H;&�H;��H;&�H;e�H;��H;��H;/�H;}kH;2FH;�H;�G;�G; G;��E;@PB;8	;;hh,;�8;	��:PX�9F�˺|-��z&�);k��!����� �C��ɇ�gж��z����G=��c��/��Ы���Ƥ�I���      ��ɾZ�ž�*��Sת�Ы��	�����T��J+��a2̽ss���yZ����μ>y�����!Ϩ�+,�u��6���:��
;��(;�M9;C�A;�ME;��F;�~G;�G;�H;�@H;agH;�H;`�H;��H;��H;ǸH;��H;ǸH;��H;��H;`�H;�H;agH;�@H;�H;�G;�~G;��F;�ME;C�A;�M9;��(;��
;���:u��6+,�!Ϩ����>y��μ����yZ�ss��a2̽��J+���T�	���Ы��Sת��*��Z�ž      0_ݾ�:پ�V;�*���Ƥ�3a����g�g$:��Z�?ݽkƣ�Al�:.%��߼=��n9.�����#V�2p��@�:�w;�'&;��7;~�@;P
E;F�F;�tG;Z�G;�
H;=H;|dH;��H;��H;t�H;ֱH;ݷH;عH;ݷH;ֱH;t�H;��H;��H;|dH;=H;�
H;Z�G;�tG;F�F;P
E;~�@;��7;�'&;�w;�@�:2p�#V�����n9.�=���߼:.%�Al�kƣ�?ݽ�Z�g$:���g�3a���Ƥ��*���V;�:پ      �]����:پZ�žI�������8t�I�C�����罽���`w�-�l���_����7��Rɻ�K/�yƹc��:P/;f$;)7;~@;��D;��F;nG;-�G;gH;�:H;�bH;��H;��H;��H;5�H;M�H;B�H;M�H;5�H;��H;��H;��H;�bH;�:H;gH;-�G;nG;��F;��D;~@;)7;f$;P/;c��:yƹ�K/��Rɻ��7��_��l��-�`w����������I�C��8t����I���Z�ž�:پ��      3F�/h��ǰ�3Vھ�������~���S��#��o��S��R₽�6�-���<y��FB��Eֻ_A?��	�Y�:���:�";�36;�@;��D;�F;�mG;&�G;>H;9?H;fH;w�H;P�H;��H;��H;�H;�H;�H;��H;��H;P�H;w�H;fH;9?H;>H;&�G;�mG;�F;��D;�@;�36;�";���:Y�:�	�_A?��EֻFB�<y��-����6�R₽S���o���#��S��~��������3Vھǰ�/h��      /h���b���쾅*־�v������)�� �O�6� ��r�r���؀��3����ݜ��>��ѻ��9�����n�:�$ ;�L#;˃6;�@@;B�D;�F;<pG;��G;TH;@H;�fH;�H;��H;�H;=�H;�H;��H;�H;=�H;�H;��H;�H;�fH;@H;TH;��G;<pG;�F;B�D;�@@;˃6;�L#;�$ ;�n�:�����9��ѻ�>�ݜ�����3��؀��r���r�6� � �O��)������v���*־�쾼b��      ǰ�쾐�޾5ʾ/;���:����v��E�A'���L����u�X�+�bW缨A��s�4�n�Ļ�8)��j��W�:�;�%;kk7;g�@;B�D;4�F;wG;��G;vH;cBH;YhH;B�H;��H;ƩH;�H;��H;��H;��H;�H;ƩH;��H;B�H;YhH;cBH;vH;��G;wG;4�F;B�D;g�@;kk7;�%;�;W�:�j���8)�n�Ļs�4��A��bW�X�+���u�L����A'��E���v��:��/;��5ʾ��޾��      3Vھ�*־5ʾT��������M���9b��5���}�սn���Xc�ݟ���ռ�I��$�$�4T���Z�_����:��;��';��8;]QA;�8E;��F;�G;%�G;�H;-FH;@kH;u�H;Z�H;�H;�H;��H;t�H;��H;�H;�H;Z�H;u�H;@kH;-FH;�H;%�G;�G;��F;�8E;]QA;��8;��';��;��:_���Z�4T��$�$��I����ռݟ��Xc�n��}�ս���5��9b��M������T���5ʾ�*־      ���v��/;������:P���r�U�H�6� ��~��@������Q�K�<��վ���s�F��_�ܺ3u9�%�:��;��+;��:;"B;��E;,�F;��G;�G;nH;[KH;'oH;k�H;��H;ƬH;_�H;��H;��H;��H;_�H;ƬH;��H;k�H;'oH;[KH;nH;�G;��G;,�F;��E;"B;��:;��+;��;�%�:3u9ܺ_�F����s��վ�<�Q�K�����@���~��6� �U�H��r�:P������/;���v��      ��������:���M���r� �O��",�<�
��gٽKĥ�|�u�K1�(����Τ�m�P��Z�q.o�kp���:Դ�:{P;��/;��<;F
C;e�E;� G;^�G;5�G;�$H;�QH;�sH;%�H;f�H;��H;*�H;{�H;&�H;{�H;*�H;��H;f�H;%�H;�sH;�QH;�$H;5�G;^�G;� G;e�E;F
C;��<;��/;{P;Դ�:�:kp��q.o��Z�m�P��Τ�(���K1�|�u�Kĥ��gٽ<�
��",� �O��r��M���:�����      �~���)����v��9b�U�H��",�0Z���S��X^��e�N�{����μ�I���%+�ۚ����.������i~:���:�l;@�3;��>;�C;�OF;�EG;{�G;"�G;�.H;'YH;�yH;p�H;��H;��H;E�H;K�H;��H;K�H;E�H;��H;��H;p�H;�yH;'YH;�.H;"�G;{�G;�EG;�OF;�C;��>;@�3;�l;���:�i~:������.�ۚ���%+��I����μ{��e�N�X^��S����0Z��",�U�H��9b���v��)��      �S� �O��E��5�6� �<�
���|9��l���Xc���(����߈��Z�[����oݎ�ܺF99���:��	;�c';��7;��@;��D;.�F;biG;��G;�H;�9H;faH;�H;/�H;P�H;g�H;��H;Y�H;��H;Y�H;��H;g�H;P�H;/�H;�H;faH;�9H;�H;��G;biG;.�F;��D;��@;��7;�c';��	;���:F99ܺoݎ����Z�[�߈�������(��Xc�l��|9����<�
�6� ��5��E� �O�      �#�6� �A'����~���gٽS��l���j��3�ji��վ�T����(�P�Ļ,A?���B�6�@:[�:�P;w�.;Q�;;�sB;\�E;��F;l�G;'�G;H;�EH;JjH;��H;H�H;.�H;��H;0�H;��H;�H;��H;0�H;��H;.�H;H�H;��H;JjH;�EH;H;'�G;l�G;��F;\�E;�sB;Q�;;w�.;�P;[�:6�@:��B�,A?�P�Ļ�(�T����վ�ji��3��j�l��S���gٽ�~����A'�6� �      �o���r���}�ս@��Kĥ�X^���Xc��3���	���˼t]��FB��Z򻆜��DӺ3��8�:z�;RM#;�<5;x?;��C;�?F;J9G;,�G;M�G;c&H;�QH;�sH;ۍH;��H;H�H;кH;��H;��H;a�H;��H;��H;кH;H�H;��H;ۍH;�sH;�QH;c&H;M�G;,�G;J9G;�?F;��C;x?;�<5;RM#;z�;�:3��8DӺ�����Z�FB�t]����˼��	��3��Xc�X^��Kĥ�@��}�ս���r�      S���r��L��n������|�u�e�N���(�ji���˼�A��b�P�=s��|������\:�:�;�m-;E�:;N�A;�+E;��F;mnG;,�G;�H;�6H;k^H;0}H;�H;&�H;��H;/�H;��H;Z�H;��H;Z�H;��H;/�H;��H;&�H;�H;0}H;k^H;�6H;�H;,�G;mnG;��F;�+E;N�A;E�:;�m-;�;�:�\:����|��=s�b�P��A����˼ji���(�e�N�|�u�����n��L���r��      R₽�؀���u��Xc�Q�K�K1�{�����վ�t]��b�P�m��	T��g�9��o�j2�9�%�:��	;�%;��5;�>;��C;	F;� G;ݙG;�G;pH;�GH;�jH;ʆH;s�H;��H;̸H;��H;l�H;��H;��H;��H;l�H;��H;̸H;��H;s�H;ʆH;�jH;�GH;pH;�G;ݙG;� G;	F;��C;�>;��5;�%;��	;�%�:j2�9�o�g�9�	T��m��b�P�t]���վ����{��K1�Q�K��Xc���u��؀�      �6��3�X�+�ݟ�<�(�����μ߈��T���FB�=s�	T����D��{���8u91q�:���:�X;at0;T�;;1B;C9E;/�F;:gG;�G;<�G;�/H;�WH;SwH;G�H;��H;#�H;�H; �H;2�H;I�H;S�H;I�H;2�H; �H;�H;#�H;��H;G�H;SwH;�WH;�/H;<�G;�G;:gG;/�F;C9E;1B;T�;;at0;�X;���:1q�:�8u9�{����D�	T��=s�FB�T���߈����μ(���<�ݟ�X�+��3�      -������bW缑�ռ�վ��Τ��I��Z�[��(��Z�g�9��{���99�W�:�W�:�P;�,;�8;�@@;ZAD;�?F;�+G;ÛG;��G;�H;�CH;HgH;W�H;y�H;��H;�H;>�H;:�H;��H;��H;��H;��H;��H;:�H;>�H;�H;��H;y�H;W�H;HgH;�CH;�H;��G;ÛG;�+G;�?F;ZAD;�@@;�8;�,;�P;�W�:�W�:�99�{��g�9���Z��(�Z�[��I���Τ��վ���ռbW缧��      <y��ݜ��A���I����s�m�P��%+����P�Ļ����|��o��8u9�W�:9+�:�;]);8�6;ذ>;�OC;��E;9�F;�wG;a�G;� H;�0H;@WH;)vH;ԎH;8�H;#�H;��H;4�H;^�H;��H;�H;��H;�H;��H;^�H;4�H;��H;#�H;8�H;ԎH;)vH;@WH;�0H;� H;a�G;�wG;9�F;��E;�OC;ذ>;8�6;]);�;9+�:�W�:�8u9�o�|�����P�Ļ����%+�m�P���s��I���A��ݜ�      FB��>�s�4�$�$�F���Z�ۚ��oݎ�,A?�DӺ����j2�91q�:�W�:�;D�';�<5;֜=;Z�B;jFE;��F;�TG;Y�G;�G;�H;�GH;9iH;�H;��H;f�H;T�H;f�H;��H;[�H;(�H;5�H;��H;5�H;(�H;[�H;��H;f�H;T�H;f�H;��H;�H;9iH;�GH;�H;�G;Y�G;�TG;��F;jFE;Z�B;֜=;�<5;D�';�;�W�:1q�:j2�9����DӺ,A?�oݎ�ۚ���Z�F��$�$�s�4��>�      �Eֻ�ѻn�Ļ4T��_�q.o���.�ܺ��B�3��8�\:�%�:���:�P;]);�<5;K:=;x"B;��D;!uF;,6G;��G;��G;�H;�9H;:]H;�yH;�H;��H;�H;'�H;��H;u�H;6�H;��H;B�H;��H;B�H;��H;6�H;u�H;��H;'�H;�H;��H;�H;�yH;:]H;�9H;�H;��G;��G;,6G;!uF;��D;x"B;K:=;�<5;]);�P;���:�%�:�\:3��8��B�ܺ��.�q.o�_�4T��n�Ļ�ѻ      _A?���9��8)��Z�ܺkp������F996�@:�:�:��	;�X;�,;8�6;֜=;x"B; �D;�WF;!G;��G;S�G;�H; .H;�RH;�pH;�H;ԜH;��H;׸H;��H;��H;��H;��H;��H;0�H;��H;0�H;��H;��H;��H;��H;��H;׸H;��H;ԜH;�H;�pH;�RH; .H;�H;S�G;��G;!G;�WF; �D;x"B;֜=;8�6;�,;�X;��	;�:�:6�@:F99����kp��ܺ�Z��8)���9�      �	�����j��_��3u9�:�i~:���:[�:z�;�;�%;at0;�8;ذ>;Z�B;��D;�WF;sG;��G;��G;��G;%H;.JH;�hH;�H;��H;T�H;��H;�H;x�H;��H;��H;H�H;��H;��H;i�H;��H;��H;H�H;��H;��H;x�H;�H;��H;T�H;��H;�H;�hH;.JH;%H;��G;��G;��G;sG;�WF;��D;Z�B;ذ>;�8;at0;�%;�;z�;[�:���:�i~:�:3u9_���j�����      Y�:�n�:W�:��:�%�:Դ�:���:��	;�P;RM#;�m-;��5;T�;;�@@;�OC;jFE;!uF;!G;��G;�G;F�G;wH;7DH;�bH;e|H;��H;ԢH;��H;ۻH;��H;��H;B�H;i�H;e�H;^�H;��H;��H;��H;^�H;e�H;i�H;B�H;��H;��H;ۻH;��H;ԢH;��H;e|H;�bH;7DH;wH;F�G;�G;��G;!G;!uF;jFE;�OC;�@@;T�;;��5;�m-;RM#;�P;��	;���:Դ�:�%�:��:W�:�n�:      ���:�$ ;�;��;��;{P;�l;�c';w�.;�<5;E�:;�>;1B;ZAD;��E;��F;,6G;��G;��G;F�G;�H;AH;/_H;mxH;��H;<�H;m�H;��H;b�H;��H;��H;F�H;��H;S�H;�H;��H;Z�H;��H;�H;S�H;��H;F�H;��H;��H;b�H;��H;m�H;<�H;��H;mxH;/_H;AH;�H;F�G;��G;��G;,6G;��F;��E;ZAD;1B;�>;E�:;�<5;w�.;�c';�l;{P;��;��;�;�$ ;      �";�L#;�%;��';��+;��/;@�3;��7;Q�;;x?;N�A;��C;C9E;�?F;9�F;�TG;��G;S�G;��G;wH;AH;�]H;hvH;9�H;��H;��H;��H;E�H;�H;7�H;1�H;��H;��H;��H;x�H;U�H;��H;U�H;x�H;��H;��H;��H;1�H;7�H;�H;E�H;��H;��H;��H;9�H;hvH;�]H;AH;wH;��G;S�G;��G;�TG;9�F;�?F;C9E;��C;N�A;x?;Q�;;��7;@�3;��/;��+;��';�%;�L#;      �36;˃6;kk7;��8;��:;��<;��>;��@;�sB;��C;�+E;	F;/�F;�+G;�wG;Y�G;��G;�H;%H;7DH;/_H;hvH;O�H;P�H;h�H;��H;��H;��H;��H;�H;=�H;Q�H;��H;m�H;��H;{�H;��H;{�H;��H;m�H;��H;Q�H;=�H;�H;��H;��H;��H;��H;h�H;P�H;O�H;hvH;/_H;7DH;%H;�H;��G;Y�G;�wG;�+G;/�F;	F;�+E;��C;�sB;��@;��>;��<;��:;��8;kk7;˃6;      �@;�@@;g�@;]QA;"B;F
C;�C;��D;\�E;�?F;��F;� G;:gG;ÛG;a�G;�G;�H; .H;.JH;�bH;mxH;9�H;P�H;ܨH;#�H;��H;��H;��H;"�H;[�H;��H;[�H;K�H;��H;��H;i�H;��H;i�H;��H;��H;K�H;[�H;��H;[�H;"�H;��H;��H;��H;#�H;ܨH;P�H;9�H;mxH;�bH;.JH; .H;�H;�G;a�G;ÛG;:gG;� G;��F;�?F;\�E;��D;�C;F
C;"B;]QA;g�@;�@@;      ��D;B�D;B�D;�8E;��E;e�E;�OF;.�F;��F;J9G;mnG;ݙG;�G;��G;� H;�H;�9H;�RH;�hH;e|H;��H;��H;h�H;#�H;U�H;��H;@�H;}�H;��H;9�H;��H;�H;��H;��H;��H;-�H;q�H;-�H;��H;��H;��H;�H;��H;9�H;��H;}�H;@�H;��H;U�H;#�H;h�H;��H;��H;e|H;�hH;�RH;�9H;�H;� H;��G;�G;ݙG;mnG;J9G;��F;.�F;�OF;e�E;��E;�8E;B�D;B�D;      �F;�F;4�F;��F;,�F;� G;�EG;biG;l�G;,�G;,�G;�G;<�G;�H;�0H;�GH;:]H;�pH;�H;��H;<�H;��H;��H;��H;��H;�H;/�H;k�H;��H;��H;��H;��H;��H;��H;��H;��H;�H;��H;��H;��H;��H;��H;��H;��H;��H;k�H;/�H;�H;��H;��H;��H;��H;<�H;��H;�H;�pH;:]H;�GH;�0H;�H;<�G;�G;,�G;,�G;l�G;biG;�EG;� G;,�F;��F;4�F;�F;      �mG;<pG;wG;�G;��G;^�G;{�G;��G;'�G;M�G;�H;pH;�/H;�CH;@WH;9iH;�yH;�H;��H;ԢH;m�H;��H;��H;��H;@�H;/�H;N�H;��H;h�H;��H;X�H;��H;��H;��H;;�H;��H;��H;��H;;�H;��H;��H;��H;X�H;��H;h�H;��H;N�H;/�H;@�H;��H;��H;��H;m�H;ԢH;��H;�H;�yH;9iH;@WH;�CH;�/H;pH;�H;M�G;'�G;��G;{�G;^�G;��G;�G;wG;<pG;      &�G;��G;��G;%�G;�G;5�G;"�G;�H;H;c&H;�6H;�GH;�WH;HgH;)vH;�H;�H;ԜH;T�H;��H;��H;E�H;��H;��H;}�H;k�H;��H;G�H;��H;K�H;��H;��H;��H;k�H;��H;�H; �H;�H;��H;k�H;��H;��H;��H;K�H;��H;G�H;��H;k�H;}�H;��H;��H;E�H;��H;��H;T�H;ԜH;�H;�H;)vH;HgH;�WH;�GH;�6H;c&H;H;�H;"�G;5�G;�G;%�G;��G;��G;      >H;TH;vH;�H;nH;�$H;�.H;�9H;�EH;�QH;k^H;�jH;SwH;W�H;ԎH;��H;��H;��H;��H;ۻH;b�H;�H;��H;"�H;��H;��H;h�H;��H;,�H;��H;��H;��H;b�H;��H;L�H;�H;��H;�H;L�H;��H;b�H;��H;��H;��H;,�H;��H;h�H;��H;��H;"�H;��H;�H;b�H;ۻH;��H;��H;��H;��H;ԎH;W�H;SwH;�jH;k^H;�QH;�EH;�9H;�.H;�$H;nH;�H;vH;TH;      9?H;@H;cBH;-FH;[KH;�QH;'YH;faH;JjH;�sH;0}H;ʆH;G�H;y�H;8�H;f�H;�H;׸H;�H;��H;��H;7�H;�H;[�H;9�H;��H;��H;K�H;��H;��H;��H;m�H;�H;T�H;��H;��H;��H;��H;��H;T�H;�H;m�H;��H;��H;��H;K�H;��H;��H;9�H;[�H;�H;7�H;��H;��H;�H;׸H;�H;f�H;8�H;y�H;G�H;ʆH;0}H;�sH;JjH;faH;'YH;�QH;[KH;-FH;cBH;@H;      fH;�fH;YhH;@kH;'oH;�sH;�yH;�H;��H;ۍH;�H;s�H;��H;��H;#�H;T�H;'�H;��H;x�H;��H;��H;1�H;=�H;��H;��H;��H;X�H;��H;��H;��H;t�H;�H;h�H;��H;��H;�H;0�H;�H;��H;��H;h�H;�H;t�H;��H;��H;��H;X�H;��H;��H;��H;=�H;1�H;��H;��H;x�H;��H;'�H;T�H;#�H;��H;��H;s�H;�H;ۍH;��H;�H;�yH;�sH;'oH;@kH;YhH;�fH;      w�H;�H;B�H;u�H;k�H;%�H;p�H;/�H;H�H;��H;&�H;��H;#�H;�H;��H;f�H;��H;��H;��H;B�H;F�H;��H;Q�H;[�H;�H;��H;��H;��H;��H;m�H;�H;z�H;��H; �H;,�H;J�H;I�H;J�H;,�H; �H;��H;z�H;�H;m�H;��H;��H;��H;��H;�H;[�H;Q�H;��H;F�H;B�H;��H;��H;��H;f�H;��H;�H;#�H;��H;&�H;��H;H�H;/�H;p�H;%�H;k�H;u�H;B�H;�H;      P�H;��H;��H;Z�H;��H;f�H;��H;P�H;.�H;H�H;��H;̸H;�H;>�H;4�H;��H;u�H;��H;��H;i�H;��H;��H;��H;K�H;��H;��H;��H;��H;b�H;�H;h�H;��H;	�H;9�H;X�H;��H;��H;��H;X�H;9�H;	�H;��H;h�H;�H;b�H;��H;��H;��H;��H;K�H;��H;��H;��H;i�H;��H;��H;u�H;��H;4�H;>�H;�H;̸H;��H;H�H;.�H;P�H;��H;f�H;��H;Z�H;��H;��H;      ��H;�H;ƩH;�H;ƬH;��H;��H;g�H;��H;кH;/�H;��H; �H;:�H;^�H;[�H;6�H;��H;H�H;e�H;S�H;��H;m�H;��H;��H;��H;��H;k�H;��H;T�H;��H; �H;9�H;u�H;��H;��H;��H;��H;��H;u�H;9�H; �H;��H;T�H;��H;k�H;��H;��H;��H;��H;m�H;��H;S�H;e�H;H�H;��H;6�H;[�H;^�H;:�H; �H;��H;/�H;кH;��H;g�H;��H;��H;ƬH;�H;ƩH;�H;      ��H;=�H;�H;�H;_�H;*�H;E�H;��H;0�H;��H;��H;l�H;2�H;��H;��H;(�H;��H;��H;��H;^�H;�H;x�H;��H;��H;��H;��H;;�H;��H;L�H;��H;��H;,�H;X�H;��H;��H;��H;��H;��H;��H;��H;X�H;,�H;��H;��H;L�H;��H;;�H;��H;��H;��H;��H;x�H;�H;^�H;��H;��H;��H;(�H;��H;��H;2�H;l�H;��H;��H;0�H;��H;E�H;*�H;_�H;�H;�H;=�H;      �H;�H;��H;��H;��H;{�H;K�H;Y�H;��H;��H;Z�H;��H;I�H;��H;�H;5�H;B�H;0�H;��H;��H;��H;U�H;{�H;i�H;-�H;��H;��H;�H;�H;��H;�H;J�H;��H;��H;��H;��H;��H;��H;��H;��H;��H;J�H;�H;��H;�H;�H;��H;��H;-�H;i�H;{�H;U�H;��H;��H;��H;0�H;B�H;5�H;�H;��H;I�H;��H;Z�H;��H;��H;Y�H;K�H;{�H;��H;��H;��H;�H;      �H;��H;��H;t�H;��H;&�H;��H;��H;�H;a�H;��H;��H;S�H;��H;��H;��H;��H;��H;i�H;��H;Z�H;��H;��H;��H;q�H;�H;��H; �H;��H;��H;0�H;I�H;��H;��H;��H;��H;��H;��H;��H;��H;��H;I�H;0�H;��H;��H; �H;��H;�H;q�H;��H;��H;��H;Z�H;��H;i�H;��H;��H;��H;��H;��H;S�H;��H;��H;a�H;�H;��H;��H;&�H;��H;t�H;��H;��H;      �H;�H;��H;��H;��H;{�H;K�H;Y�H;��H;��H;Z�H;��H;I�H;��H;�H;5�H;B�H;0�H;��H;��H;��H;U�H;{�H;i�H;-�H;��H;��H;�H;�H;��H;�H;J�H;��H;��H;��H;��H;��H;��H;��H;��H;��H;J�H;�H;��H;�H;�H;��H;��H;-�H;i�H;{�H;U�H;��H;��H;��H;0�H;B�H;5�H;�H;��H;I�H;��H;Z�H;��H;��H;Y�H;K�H;{�H;��H;��H;��H;�H;      ��H;=�H;�H;�H;_�H;*�H;E�H;��H;0�H;��H;��H;l�H;2�H;��H;��H;(�H;��H;��H;��H;^�H;�H;x�H;��H;��H;��H;��H;;�H;��H;L�H;��H;��H;,�H;X�H;��H;��H;��H;��H;��H;��H;��H;X�H;,�H;��H;��H;L�H;��H;;�H;��H;��H;��H;��H;x�H;�H;^�H;��H;��H;��H;(�H;��H;��H;2�H;l�H;��H;��H;0�H;��H;E�H;*�H;_�H;�H;�H;=�H;      ��H;�H;ƩH;�H;ƬH;��H;��H;g�H;��H;кH;/�H;��H; �H;:�H;^�H;[�H;6�H;��H;H�H;e�H;S�H;��H;m�H;��H;��H;��H;��H;k�H;��H;T�H;��H; �H;9�H;u�H;��H;��H;��H;��H;��H;u�H;9�H; �H;��H;T�H;��H;k�H;��H;��H;��H;��H;m�H;��H;S�H;e�H;H�H;��H;6�H;[�H;^�H;:�H; �H;��H;/�H;кH;��H;g�H;��H;��H;ƬH;�H;ƩH;�H;      P�H;��H;��H;Z�H;��H;f�H;��H;P�H;.�H;H�H;��H;̸H;�H;>�H;4�H;��H;u�H;��H;��H;i�H;��H;��H;��H;K�H;��H;��H;��H;��H;b�H;�H;h�H;��H;	�H;9�H;X�H;��H;��H;��H;X�H;9�H;	�H;��H;h�H;�H;b�H;��H;��H;��H;��H;K�H;��H;��H;��H;i�H;��H;��H;u�H;��H;4�H;>�H;�H;̸H;��H;H�H;.�H;P�H;��H;f�H;��H;Z�H;��H;��H;      w�H;�H;B�H;u�H;k�H;%�H;p�H;/�H;H�H;��H;&�H;��H;#�H;�H;��H;f�H;��H;��H;��H;B�H;F�H;��H;Q�H;[�H;�H;��H;��H;��H;��H;m�H;�H;z�H;��H; �H;,�H;J�H;I�H;J�H;,�H; �H;��H;z�H;�H;m�H;��H;��H;��H;��H;�H;[�H;Q�H;��H;F�H;B�H;��H;��H;��H;f�H;��H;�H;#�H;��H;&�H;��H;H�H;/�H;p�H;%�H;k�H;u�H;B�H;�H;      fH;�fH;YhH;@kH;'oH;�sH;�yH;�H;��H;ۍH;�H;s�H;��H;��H;#�H;T�H;'�H;��H;x�H;��H;��H;1�H;=�H;��H;��H;��H;X�H;��H;��H;��H;t�H;�H;h�H;��H;��H;�H;0�H;�H;��H;��H;h�H;�H;t�H;��H;��H;��H;X�H;��H;��H;��H;=�H;1�H;��H;��H;x�H;��H;'�H;T�H;#�H;��H;��H;s�H;�H;ۍH;��H;�H;�yH;�sH;'oH;@kH;YhH;�fH;      9?H;@H;cBH;-FH;[KH;�QH;'YH;faH;JjH;�sH;0}H;ʆH;G�H;y�H;8�H;f�H;�H;׸H;�H;��H;��H;7�H;�H;[�H;9�H;��H;��H;K�H;��H;��H;��H;m�H;�H;T�H;��H;��H;��H;��H;��H;T�H;�H;m�H;��H;��H;��H;K�H;��H;��H;9�H;[�H;�H;7�H;��H;��H;�H;׸H;�H;f�H;8�H;y�H;G�H;ʆH;0}H;�sH;JjH;faH;'YH;�QH;[KH;-FH;cBH;@H;      >H;TH;vH;�H;nH;�$H;�.H;�9H;�EH;�QH;k^H;�jH;SwH;W�H;ԎH;��H;��H;��H;��H;ۻH;b�H;�H;��H;"�H;��H;��H;h�H;��H;,�H;��H;��H;��H;b�H;��H;L�H;�H;��H;�H;L�H;��H;b�H;��H;��H;��H;,�H;��H;h�H;��H;��H;"�H;��H;�H;b�H;ۻH;��H;��H;��H;��H;ԎH;W�H;SwH;�jH;k^H;�QH;�EH;�9H;�.H;�$H;nH;�H;vH;TH;      &�G;��G;��G;%�G;�G;5�G;"�G;�H;H;c&H;�6H;�GH;�WH;HgH;)vH;�H;�H;ԜH;T�H;��H;��H;E�H;��H;��H;}�H;k�H;��H;G�H;��H;K�H;��H;��H;��H;k�H;��H;�H; �H;�H;��H;k�H;��H;��H;��H;K�H;��H;G�H;��H;k�H;}�H;��H;��H;E�H;��H;��H;T�H;ԜH;�H;�H;)vH;HgH;�WH;�GH;�6H;c&H;H;�H;"�G;5�G;�G;%�G;��G;��G;      �mG;<pG;wG;�G;��G;^�G;{�G;��G;'�G;M�G;�H;pH;�/H;�CH;@WH;9iH;�yH;�H;��H;ԢH;m�H;��H;��H;��H;@�H;/�H;N�H;��H;h�H;��H;X�H;��H;��H;��H;;�H;��H;��H;��H;;�H;��H;��H;��H;X�H;��H;h�H;��H;N�H;/�H;@�H;��H;��H;��H;m�H;ԢH;��H;�H;�yH;9iH;@WH;�CH;�/H;pH;�H;M�G;'�G;��G;{�G;^�G;��G;�G;wG;<pG;      �F;�F;4�F;��F;,�F;� G;�EG;biG;l�G;,�G;,�G;�G;<�G;�H;�0H;�GH;:]H;�pH;�H;��H;<�H;��H;��H;��H;��H;�H;/�H;k�H;��H;��H;��H;��H;��H;��H;��H;��H;�H;��H;��H;��H;��H;��H;��H;��H;��H;k�H;/�H;�H;��H;��H;��H;��H;<�H;��H;�H;�pH;:]H;�GH;�0H;�H;<�G;�G;,�G;,�G;l�G;biG;�EG;� G;,�F;��F;4�F;�F;      ��D;B�D;B�D;�8E;��E;e�E;�OF;.�F;��F;J9G;mnG;ݙG;�G;��G;� H;�H;�9H;�RH;�hH;e|H;��H;��H;h�H;#�H;U�H;��H;@�H;}�H;��H;9�H;��H;�H;��H;��H;��H;-�H;q�H;-�H;��H;��H;��H;�H;��H;9�H;��H;}�H;@�H;��H;U�H;#�H;h�H;��H;��H;e|H;�hH;�RH;�9H;�H;� H;��G;�G;ݙG;mnG;J9G;��F;.�F;�OF;e�E;��E;�8E;B�D;B�D;      �@;�@@;g�@;]QA;"B;F
C;�C;��D;\�E;�?F;��F;� G;:gG;ÛG;a�G;�G;�H; .H;.JH;�bH;mxH;9�H;P�H;ܨH;#�H;��H;��H;��H;"�H;[�H;��H;[�H;K�H;��H;��H;i�H;��H;i�H;��H;��H;K�H;[�H;��H;[�H;"�H;��H;��H;��H;#�H;ܨH;P�H;9�H;mxH;�bH;.JH; .H;�H;�G;a�G;ÛG;:gG;� G;��F;�?F;\�E;��D;�C;F
C;"B;]QA;g�@;�@@;      �36;˃6;kk7;��8;��:;��<;��>;��@;�sB;��C;�+E;	F;/�F;�+G;�wG;Y�G;��G;�H;%H;7DH;/_H;hvH;O�H;P�H;h�H;��H;��H;��H;��H;�H;=�H;Q�H;��H;m�H;��H;{�H;��H;{�H;��H;m�H;��H;Q�H;=�H;�H;��H;��H;��H;��H;h�H;P�H;O�H;hvH;/_H;7DH;%H;�H;��G;Y�G;�wG;�+G;/�F;	F;�+E;��C;�sB;��@;��>;��<;��:;��8;kk7;˃6;      �";�L#;�%;��';��+;��/;@�3;��7;Q�;;x?;N�A;��C;C9E;�?F;9�F;�TG;��G;S�G;��G;wH;AH;�]H;hvH;9�H;��H;��H;��H;E�H;�H;7�H;1�H;��H;��H;��H;x�H;U�H;��H;U�H;x�H;��H;��H;��H;1�H;7�H;�H;E�H;��H;��H;��H;9�H;hvH;�]H;AH;wH;��G;S�G;��G;�TG;9�F;�?F;C9E;��C;N�A;x?;Q�;;��7;@�3;��/;��+;��';�%;�L#;      ���:�$ ;�;��;��;{P;�l;�c';w�.;�<5;E�:;�>;1B;ZAD;��E;��F;,6G;��G;��G;F�G;�H;AH;/_H;mxH;��H;<�H;m�H;��H;b�H;��H;��H;F�H;��H;S�H;�H;��H;Z�H;��H;�H;S�H;��H;F�H;��H;��H;b�H;��H;m�H;<�H;��H;mxH;/_H;AH;�H;F�G;��G;��G;,6G;��F;��E;ZAD;1B;�>;E�:;�<5;w�.;�c';�l;{P;��;��;�;�$ ;      Y�:�n�:W�:��:�%�:Դ�:���:��	;�P;RM#;�m-;��5;T�;;�@@;�OC;jFE;!uF;!G;��G;�G;F�G;wH;7DH;�bH;e|H;��H;ԢH;��H;ۻH;��H;��H;B�H;i�H;e�H;^�H;��H;��H;��H;^�H;e�H;i�H;B�H;��H;��H;ۻH;��H;ԢH;��H;e|H;�bH;7DH;wH;F�G;�G;��G;!G;!uF;jFE;�OC;�@@;T�;;��5;�m-;RM#;�P;��	;���:Դ�:�%�:��:W�:�n�:      �	�����j��_��3u9�:�i~:���:[�:z�;�;�%;at0;�8;ذ>;Z�B;��D;�WF;sG;��G;��G;��G;%H;.JH;�hH;�H;��H;T�H;��H;�H;x�H;��H;��H;H�H;��H;��H;i�H;��H;��H;H�H;��H;��H;x�H;�H;��H;T�H;��H;�H;�hH;.JH;%H;��G;��G;��G;sG;�WF;��D;Z�B;ذ>;�8;at0;�%;�;z�;[�:���:�i~:�:3u9_���j�����      _A?���9��8)��Z�ܺkp������F996�@:�:�:��	;�X;�,;8�6;֜=;x"B; �D;�WF;!G;��G;S�G;�H; .H;�RH;�pH;�H;ԜH;��H;׸H;��H;��H;��H;��H;��H;0�H;��H;0�H;��H;��H;��H;��H;��H;׸H;��H;ԜH;�H;�pH;�RH; .H;�H;S�G;��G;!G;�WF; �D;x"B;֜=;8�6;�,;�X;��	;�:�:6�@:F99����kp��ܺ�Z��8)���9�      �Eֻ�ѻn�Ļ4T��_�q.o���.�ܺ��B�3��8�\:�%�:���:�P;]);�<5;K:=;x"B;��D;!uF;,6G;��G;��G;�H;�9H;:]H;�yH;�H;��H;�H;'�H;��H;u�H;6�H;��H;B�H;��H;B�H;��H;6�H;u�H;��H;'�H;�H;��H;�H;�yH;:]H;�9H;�H;��G;��G;,6G;!uF;��D;x"B;K:=;�<5;]);�P;���:�%�:�\:3��8��B�ܺ��.�q.o�_�4T��n�Ļ�ѻ      FB��>�s�4�$�$�F���Z�ۚ��oݎ�,A?�DӺ����j2�91q�:�W�:�;D�';�<5;֜=;Z�B;jFE;��F;�TG;Y�G;�G;�H;�GH;9iH;�H;��H;f�H;T�H;f�H;��H;[�H;(�H;5�H;��H;5�H;(�H;[�H;��H;f�H;T�H;f�H;��H;�H;9iH;�GH;�H;�G;Y�G;�TG;��F;jFE;Z�B;֜=;�<5;D�';�;�W�:1q�:j2�9����DӺ,A?�oݎ�ۚ���Z�F��$�$�s�4��>�      <y��ݜ��A���I����s�m�P��%+����P�Ļ����|��o��8u9�W�:9+�:�;]);8�6;ذ>;�OC;��E;9�F;�wG;a�G;� H;�0H;@WH;)vH;ԎH;8�H;#�H;��H;4�H;^�H;��H;�H;��H;�H;��H;^�H;4�H;��H;#�H;8�H;ԎH;)vH;@WH;�0H;� H;a�G;�wG;9�F;��E;�OC;ذ>;8�6;]);�;9+�:�W�:�8u9�o�|�����P�Ļ����%+�m�P���s��I���A��ݜ�      -������bW缑�ռ�վ��Τ��I��Z�[��(��Z�g�9��{���99�W�:�W�:�P;�,;�8;�@@;ZAD;�?F;�+G;ÛG;��G;�H;�CH;HgH;W�H;y�H;��H;�H;>�H;:�H;��H;��H;��H;��H;��H;:�H;>�H;�H;��H;y�H;W�H;HgH;�CH;�H;��G;ÛG;�+G;�?F;ZAD;�@@;�8;�,;�P;�W�:�W�:�99�{��g�9���Z��(�Z�[��I���Τ��վ���ռbW缧��      �6��3�X�+�ݟ�<�(�����μ߈��T���FB�=s�	T����D��{���8u91q�:���:�X;at0;T�;;1B;C9E;/�F;:gG;�G;<�G;�/H;�WH;SwH;G�H;��H;#�H;�H; �H;2�H;I�H;S�H;I�H;2�H; �H;�H;#�H;��H;G�H;SwH;�WH;�/H;<�G;�G;:gG;/�F;C9E;1B;T�;;at0;�X;���:1q�:�8u9�{����D�	T��=s�FB�T���߈����μ(���<�ݟ�X�+��3�      R₽�؀���u��Xc�Q�K�K1�{�����վ�t]��b�P�m��	T��g�9��o�j2�9�%�:��	;�%;��5;�>;��C;	F;� G;ݙG;�G;pH;�GH;�jH;ʆH;s�H;��H;̸H;��H;l�H;��H;��H;��H;l�H;��H;̸H;��H;s�H;ʆH;�jH;�GH;pH;�G;ݙG;� G;	F;��C;�>;��5;�%;��	;�%�:j2�9�o�g�9�	T��m��b�P�t]���վ����{��K1�Q�K��Xc���u��؀�      S���r��L��n������|�u�e�N���(�ji���˼�A��b�P�=s��|������\:�:�;�m-;E�:;N�A;�+E;��F;mnG;,�G;�H;�6H;k^H;0}H;�H;&�H;��H;/�H;��H;Z�H;��H;Z�H;��H;/�H;��H;&�H;�H;0}H;k^H;�6H;�H;,�G;mnG;��F;�+E;N�A;E�:;�m-;�;�:�\:����|��=s�b�P��A����˼ji���(�e�N�|�u�����n��L���r��      �o���r���}�ս@��Kĥ�X^���Xc��3���	���˼t]��FB��Z򻆜��DӺ3��8�:z�;RM#;�<5;x?;��C;�?F;J9G;,�G;M�G;c&H;�QH;�sH;ۍH;��H;H�H;кH;��H;��H;a�H;��H;��H;кH;H�H;��H;ۍH;�sH;�QH;c&H;M�G;,�G;J9G;�?F;��C;x?;�<5;RM#;z�;�:3��8DӺ�����Z�FB�t]����˼��	��3��Xc�X^��Kĥ�@��}�ս���r�      �#�6� �A'����~���gٽS��l���j��3�ji��վ�T����(�P�Ļ,A?���B�6�@:[�:�P;w�.;Q�;;�sB;\�E;��F;l�G;'�G;H;�EH;JjH;��H;H�H;.�H;��H;0�H;��H;�H;��H;0�H;��H;.�H;H�H;��H;JjH;�EH;H;'�G;l�G;��F;\�E;�sB;Q�;;w�.;�P;[�:6�@:��B�,A?�P�Ļ�(�T����վ�ji��3��j�l��S���gٽ�~����A'�6� �      �S� �O��E��5�6� �<�
���|9��l���Xc���(����߈��Z�[����oݎ�ܺF99���:��	;�c';��7;��@;��D;.�F;biG;��G;�H;�9H;faH;�H;/�H;P�H;g�H;��H;Y�H;��H;Y�H;��H;g�H;P�H;/�H;�H;faH;�9H;�H;��G;biG;.�F;��D;��@;��7;�c';��	;���:F99ܺoݎ����Z�[�߈�������(��Xc�l��|9����<�
�6� ��5��E� �O�      �~���)����v��9b�U�H��",�0Z���S��X^��e�N�{����μ�I���%+�ۚ����.������i~:���:�l;@�3;��>;�C;�OF;�EG;{�G;"�G;�.H;'YH;�yH;p�H;��H;��H;E�H;K�H;��H;K�H;E�H;��H;��H;p�H;�yH;'YH;�.H;"�G;{�G;�EG;�OF;�C;��>;@�3;�l;���:�i~:������.�ۚ���%+��I����μ{��e�N�X^��S����0Z��",�U�H��9b���v��)��      ��������:���M���r� �O��",�<�
��gٽKĥ�|�u�K1�(����Τ�m�P��Z�q.o�kp���:Դ�:{P;��/;��<;F
C;e�E;� G;^�G;5�G;�$H;�QH;�sH;%�H;f�H;��H;*�H;{�H;&�H;{�H;*�H;��H;f�H;%�H;�sH;�QH;�$H;5�G;^�G;� G;e�E;F
C;��<;��/;{P;Դ�:�:kp��q.o��Z�m�P��Τ�(���K1�|�u�Kĥ��gٽ<�
��",� �O��r��M���:�����      ���v��/;������:P���r�U�H�6� ��~��@������Q�K�<��վ���s�F��_�ܺ3u9�%�:��;��+;��:;"B;��E;,�F;��G;�G;nH;[KH;'oH;k�H;��H;ƬH;_�H;��H;��H;��H;_�H;ƬH;��H;k�H;'oH;[KH;nH;�G;��G;,�F;��E;"B;��:;��+;��;�%�:3u9ܺ_�F����s��վ�<�Q�K�����@���~��6� �U�H��r�:P������/;���v��      3Vھ�*־5ʾT��������M���9b��5���}�սn���Xc�ݟ���ռ�I��$�$�4T���Z�_����:��;��';��8;]QA;�8E;��F;�G;%�G;�H;-FH;@kH;u�H;Z�H;�H;�H;��H;t�H;��H;�H;�H;Z�H;u�H;@kH;-FH;�H;%�G;�G;��F;�8E;]QA;��8;��';��;��:_���Z�4T��$�$��I����ռݟ��Xc�n��}�ս���5��9b��M������T���5ʾ�*־      ǰ�쾐�޾5ʾ/;���:����v��E�A'���L����u�X�+�bW缨A��s�4�n�Ļ�8)��j��W�:�;�%;kk7;g�@;B�D;4�F;wG;��G;vH;cBH;YhH;B�H;��H;ƩH;�H;��H;��H;��H;�H;ƩH;��H;B�H;YhH;cBH;vH;��G;wG;4�F;B�D;g�@;kk7;�%;�;W�:�j���8)�n�Ļs�4��A��bW�X�+���u�L����A'��E���v��:��/;��5ʾ��޾��      /h���b���쾅*־�v������)�� �O�6� ��r�r���؀��3����ݜ��>��ѻ��9�����n�:�$ ;�L#;˃6;�@@;B�D;�F;<pG;��G;TH;@H;�fH;�H;��H;�H;=�H;�H;��H;�H;=�H;�H;��H;�H;�fH;@H;TH;��G;<pG;�F;B�D;�@@;˃6;�L#;�$ ;�n�:�����9��ѻ�>�ݜ�����3��؀��r���r�6� � �O��)������v���*־�쾼b��      �$��� ���������þ�*��
Dx�}�=����\Pν鰒��&K�xc����;�V�s���D^���S��v[:���:�d;��4;�_?;�lD;��F;puG;M�G;�H;�NH;�rH;�H;��H;��H;�H;q�H;E�H;q�H;�H;��H;��H;�H;�rH;�NH;�H;M�G;puG;��F;�lD;�_?;��4;�d;���:�v[:��S��D^�s��;�V����xc��&K�鰒�\Pν���}�=�
Dx��*���þ��������� �      �� �k��>��=���������0���s���:�N9���ʽZ����G��8��-��z5S�v���/X���D��Ad:�A�:� ;x�4;	�?;#~D;q�F;3xG;��G;�H;NOH;HsH;:�H;�H;�H;W�H;��H;U�H;��H;W�H;�H;�H;:�H;HsH;NOH;�H;��G;3xG;q�F;#~D;	�?;x�4;� ;�A�:�Ad:��D��/X�v��z5S��-���8���G�Z����ʽN9���:��s��0��������=��>��k��      ���>��&�
�����fYؾ���ȥ����f���0�C[�*8������ȟ>�|���#Ȥ�Y6H�,�ܻ�qF�/��5�}:���:�";��5;6�?;��D;��F;/�G;��G;s"H;�QH;�tH;z�H;�H;��H;�H;�H;��H;�H;�H;��H;�H;z�H;�tH;�QH;s"H;��G;/�G;��F;��D;6�?;��5;�";���:5�}:/���qF�,�ܻY6H�#Ȥ�|���ȟ>�����*8��C[���0���f�ȥ�����fYؾ����&�
�>��      ��=������I��þ�R��&���QS��Q"��s�����}��0���d���x�6��ƻ(}*����^�:�w;�%;Rl7;�@;�D;�F;��G;��G;3'H;UH;�wH;�H;f�H;ñH;ۺH;�H;��H;�H;ۺH;ñH;f�H;�H;�wH;UH;3'H;��G;��G;�F;�D;�@;Rl7;�%;�w;^�:���(}*��ƻx�6�d����켟0���}�����s��Q"�QS�&����R���þIᾁ���=��      ����fYؾ�þ�ê�f쏾jk���:�e�R�ؽ�����c�:y���Ҽݫ��� �B�'��E�'7��:�
;d�(;�^9;��A;�[E;��F;�G;��G;�-H;�YH;{H;�H;i�H;u�H;6�H;�H;��H;�H;6�H;u�H;i�H;�H;{H;�YH;�-H;��G;�G;��F;�[E;��A;�^9;d�(;�
;��:E�'7'��B�� �ݫ����Ҽ:y��c�����R�ؽe���:�jk�f쏾�ê��þfYؾ��      �þ��������R��f쏾�s��H����������������D�vc�g����f�3,�����P����9/��:5;�i-;��;;��B;+�E;�G;��G;��G;�5H;�_H;�H;{�H;�H;r�H;ɽH;r�H;��H;r�H;ɽH;r�H;�H;{�H;�H;�_H;�5H;��G;��G;�G;+�E;��B;��;;�i-;5;/��:��9�P�����3,��f�g���vc���D���������������H��s�f쏾�R���������      �*���0��ȥ��&���jk��H��#%�B[�ZPν�s��0�f�/%�d��`���G�=�n?ػgFL��D�a�R:C�:��;�2;�=;��C;�/F;�FG;�G;WH;?H;�fH;��H;V�H;ͫH;��H;��H;�H;��H;�H;��H;��H;ͫH;V�H;��H;�fH;?H;WH;�G;�FG;�/F;��C;�=;�2;��;C�:a�R:�D�gFL�n?ػG�=�`���d��/%�0�f��s��ZPνB[��#%��H�jk�&���ȥ���0��      
Dx��s���f�QS���:����B[��7ս�榽��}�u�;��8�)�����r����G������Ҭ����:��;}$;,�6;f�?;3�D;�F; pG;��G;H;XIH;dnH;i�H;��H;�H;[�H;��H;��H;G�H;��H;��H;[�H;�H;��H;i�H;dnH;XIH;H;��G; pG;�F;3�D;f�?;,�6;}$;��;���:�Ҭ����G�������r�)����8�u�;���}��榽�7սB[������:�QS���f��s�      }�=���:���0��Q"�e�����ZPν�榽%����G�����Ҽ���E:�	�ܻ�D^�θ��jh:���:P;�{,;�:;��A;~hE;��F;\�G;��G;�'H;eTH;�vH;��H;L�H;��H;�H;��H;��H;4�H;��H;��H;�H;��H;L�H;��H;�vH;eTH;�'H;��G;\�G;��F;~hE;��A;�:;�{,;P;���:jh:θ���D^�	�ܻE:������Ҽ����G�%���榽ZPν����e��Q"���0���:�      ���N9�C[��s�R�ؽ���s����}���G��K��	c��!�V�%,��*�����&����:@��:� ;ǂ3;0>;�C;#F;$8G;l�G;�H;7H;�_H;,H;�H; �H;g�H;�H;m�H;��H;3�H;��H;m�H;�H;g�H; �H;�H;,H;�_H;7H;�H;l�G;$8G;#F;�C;0>;ǂ3;� ;@��:��:&������*��%,�!�V�	c��K�����G���}��s����R�ؽ�s�C[�N9�      \Pν��ʽ*8�������������0�f�u�;���K��Ȥ���f���#ߵ�>o5�4�D�M�-:���:X>;G+;_9;�A;��D;[�F;�uG;�G;IH;�FH;�kH;�H;��H;�H;H�H;�H;��H;"�H;F�H;"�H;��H;�H;H�H;�H;��H;�H;�kH;�FH;IH;�G;�uG;[�F;��D;�A;_9;G+;X>;���:M�-:4�D�>o5�#ߵ�����f�Ȥ�K����u�;�0�f������������*8����ʽ      鰒�Z��������}��c���D�/%��8���Ҽ	c����f�����ƻY/X�u����9g�:ȏ;G";�3;�>;�XC;��E;G;'�G;��G;�+H;/VH;9wH;��H;W�H;�H;.�H;�H;Q�H;`�H;O�H;`�H;Q�H;�H;.�H;�H;W�H;��H;9wH;/VH;�+H;��G;'�G;G;��E;�XC;�>;�3;G";ȏ;g�:�9u���Y/X��ƻ�����f�	c����Ҽ�8�/%���D��c���}�����Z��      �&K���G�ȟ>��0�:y�vc�d��)������!�V����ƻfod���º�P(7�3�:���: �;]P.;:�:;ayA;y�D;�F;�mG;t�G;!H;�?H;MeH;��H;R�H;ժH;��H;�H;
�H;��H;��H;V�H;��H;��H;
�H;�H;��H;ժH;R�H;��H;MeH;�?H;!H;t�G;�mG;�F;y�D;ayA;:�:;]P.; �;���:�3�:�P(7��ºfod��ƻ��!�V����)���d��vc�:y��0�ȟ>���G�      xc��8�|����켔�Ҽg���`�����r�E:�%,�#ߵ�Y/X���º̬�F�}:> �:v;��);�l7;i�?;�C;KF;�(G;E�G;��G;2)H;�RH;�sH;��H;��H;�H;ͼH;��H;��H;,�H;��H;l�H;��H;,�H;��H;��H;ͼH;�H;��H;��H;�sH;�RH;2)H;��G;E�G;�(G;KF;�C;i�?;�l7;��);v;> �:F�}:̬���ºY/X�#ߵ�%,�E:���r�`���g�����Ҽ��|����8�      ����-��#Ȥ�d���ݫ���f�G�=����	�ܻ�*��>o5�u����P(7F�}:�m�:��;>&;��4;B�=;�B;,�E;S�F;ˀG;$�G;cH;�@H;�dH;d�H;��H;x�H;��H;��H;;�H;��H;��H;��H;l�H;��H;��H;��H;;�H;��H;��H;x�H;��H;d�H;�dH;�@H;cH;$�G;ˀG;S�F;,�E;�B;B�=;��4;>&;��;�m�:F�}:�P(7u���>o5��*��	�ܻ���G�=��f�ݫ��d���#Ȥ��-��      ;�V�z5S�Y6H�x�6�� �3,�n?ػG���D^����4�D��9�3�:> �:��;]%;��3;p�<;�B;�
E;>�F;�WG;8�G;t�G;�/H;xVH;�uH;�H;��H;ܰH;��H;��H;��H;k�H;��H;��H;Q�H;��H;��H;k�H;��H;��H;��H;ܰH;��H;�H;�uH;xVH;�/H;t�G;8�G;�WG;>�F;�
E;�B;p�<;��3;]%;��;> �:�3�:�94�D�����D^�G��n?ػ3,�� �x�6�Y6H�z5S�      s��v��,�ܻ�ƻB󩻜��gFL����θ��&��M�-:g�:���:v;>&;��3;�8<;`�A;%�D;�YF;Z4G;3�G;�G;� H;aIH;VjH;ńH;ٙH;��H;��H;�H;��H;��H;��H;��H;v�H;�H;v�H;��H;��H;��H;��H;�H;��H;��H;ٙH;ńH;VjH;aIH;� H;�G;3�G;Z4G;�YF;%�D;`�A;�8<;��3;>&;v;���:g�:M�-:&��θ�����gFL����B��ƻ,�ܻv��      �D^��/X��qF�(}*�'���P���D��Ҭ�jh:��:���:ȏ; �;��);��4;p�<;`�A;f�D;�8F;
G;��G;w�G;jH;C>H;�`H;5|H;��H;��H;��H;��H;��H;|�H;��H;4�H;��H;8�H;��H;8�H;��H;4�H;��H;|�H;��H;��H;��H;��H;��H;5|H;�`H;C>H;jH;w�G;��G;
G;�8F;f�D;`�A;p�<;��4;��); �;ȏ;���:��:jh:�Ҭ��D��P��'��(}*��qF��/X�      ��S���D�/�����E�'7��9a�R:���:���:@��:X>;G";]P.;�l7;B�=;�B;%�D;�8F;XG;R�G;��G;�H;�5H;�XH;uH;=�H;�H;�H;�H;��H;9�H;��H;-�H;M�H;r�H;��H;�H;��H;r�H;M�H;-�H;��H;9�H;��H;�H;�H;�H;=�H;uH;�XH;�5H;�H;��G;R�G;XG;�8F;%�D;�B;B�=;�l7;]P.;G";X>;@��:���:���:a�R:��9E�'7���/����D�      �v[:�Ad:5�}:^�:��:/��:C�:��;P;� ;G+;�3;:�:;i�?;�B;�
E;�YF;
G;R�G;��G;nH;�0H;�RH;�oH;�H;f�H;�H;��H;��H;��H;�H;��H;��H;5�H;�H;(�H;q�H;(�H;�H;5�H;��H;��H;�H;��H;��H;��H;�H;f�H;�H;�oH;�RH;�0H;nH;��G;R�G;
G;�YF;�
E;�B;i�?;:�:;�3;G+;� ;P;��;C�:/��:��:^�:5�}:�Ad:      ���:�A�:���:�w;�
;5;��;}$;�{,;ǂ3;_9;�>;ayA;�C;,�E;>�F;Z4G;��G;��G;nH;�.H;PH;&lH;i�H;��H;��H;��H;�H;��H;)�H;r�H;��H;��H;��H;z�H;W�H;��H;W�H;z�H;��H;��H;��H;r�H;)�H;��H;�H;��H;��H;��H;i�H;&lH;PH;�.H;nH;��G;��G;Z4G;>�F;,�E;�C;ayA;�>;_9;ǂ3;�{,;}$;��;5;�
;�w;���:�A�:      �d;� ;�";�%;d�(;�i-;�2;,�6;�:;0>;�A;�XC;y�D;KF;S�F;�WG;3�G;w�G;�H;�0H;PH;�jH;��H;��H;V�H;E�H;�H;��H;��H;�H;��H;��H;��H;�H;��H;j�H;��H;j�H;��H;�H;��H;��H;��H;�H;��H;��H;�H;E�H;V�H;��H;��H;�jH;PH;�0H;�H;w�G;3�G;�WG;S�F;KF;y�D;�XC;�A;0>;�:;,�6;�2;�i-;d�(;�%;�";� ;      ��4;x�4;��5;Rl7;�^9;��;;�=;f�?;��A;�C;��D;��E;�F;�(G;ˀG;8�G;�G;jH;�5H;�RH;&lH;��H;˓H;#�H;گH;g�H;<�H;H�H;��H;��H;(�H;��H;C�H;��H;��H;m�H;��H;m�H;��H;��H;C�H;��H;(�H;��H;��H;H�H;<�H;g�H;گH;#�H;˓H;��H;&lH;�RH;�5H;jH;�G;8�G;ˀG;�(G;�F;��E;��D;�C;��A;f�?;�=;��;;�^9;Rl7;��5;x�4;      �_?;	�?;6�?;�@;��A;��B;��C;3�D;~hE;#F;[�F;G;�mG;E�G;$�G;t�G;� H;C>H;�XH;�oH;i�H;��H;#�H;\�H;��H;;�H;Y�H;�H;��H;��H;g�H;��H;��H;��H;��H;E�H;^�H;E�H;��H;��H;��H;��H;g�H;��H;��H;�H;Y�H;;�H;��H;\�H;#�H;��H;i�H;�oH;�XH;C>H;� H;t�G;$�G;E�G;�mG;G;[�F;#F;~hE;3�D;��C;��B;��A;�@;6�?;	�?;      �lD;#~D;��D;�D;�[E;+�E;�/F;�F;��F;$8G;�uG;'�G;t�G;��G;cH;�/H;aIH;�`H;uH;�H;��H;V�H;گH;��H;�H;��H;}�H;#�H;��H;�H;n�H;N�H;��H;��H;��H;��H;6�H;��H;��H;��H;��H;N�H;n�H;�H;��H;#�H;}�H;��H;�H;��H;گH;V�H;��H;�H;uH;�`H;aIH;�/H;cH;��G;t�G;'�G;�uG;$8G;��F;�F;�/F;+�E;�[E;�D;��D;#~D;      ��F;q�F;��F;�F;��F;�G;�FG; pG;\�G;l�G;�G;��G;!H;2)H;�@H;xVH;VjH;5|H;=�H;f�H;��H;E�H;g�H;;�H;��H;E�H;��H;��H;��H;�H;�H;��H;��H;��H;B�H;��H;��H;��H;B�H;��H;��H;��H;�H;�H;��H;��H;��H;E�H;��H;;�H;g�H;E�H;��H;f�H;=�H;5|H;VjH;xVH;�@H;2)H;!H;��G;�G;l�G;\�G; pG;�FG;�G;��F;�F;��F;q�F;      puG;3xG;/�G;��G;�G;��G;�G;��G;��G;�H;IH;�+H;�?H;�RH;�dH;�uH;ńH;��H;�H;�H;��H;�H;<�H;Y�H;}�H;��H;t�H;m�H;��H;��H;n�H;��H;��H;L�H;��H;-�H;.�H;-�H;��H;L�H;��H;��H;n�H;��H;��H;m�H;t�H;��H;}�H;Y�H;<�H;�H;��H;�H;�H;��H;ńH;�uH;�dH;�RH;�?H;�+H;IH;�H;��G;��G;�G;��G;�G;��G;/�G;3xG;      M�G;��G;��G;��G;��G;��G;WH;H;�'H;7H;�FH;/VH;MeH;�sH;d�H;�H;ٙH;��H;�H;��H;�H;��H;H�H;�H;#�H;��H;m�H;��H;��H;p�H;��H;��H;c�H;��H;V�H;��H;��H;��H;V�H;��H;c�H;��H;��H;p�H;��H;��H;m�H;��H;#�H;�H;H�H;��H;�H;��H;�H;��H;ٙH;�H;d�H;�sH;MeH;/VH;�FH;7H;�'H;H;WH;��G;��G;��G;��G;��G;      �H;�H;s"H;3'H;�-H;�5H;?H;XIH;eTH;�_H;�kH;9wH;��H;��H;��H;��H;��H;��H;�H;��H;��H;��H;��H;��H;��H;��H;��H;��H;>�H;��H;��H;X�H;��H;y�H;��H;��H;��H;��H;��H;y�H;��H;X�H;��H;��H;>�H;��H;��H;��H;��H;��H;��H;��H;��H;��H;�H;��H;��H;��H;��H;��H;��H;9wH;�kH;�_H;eTH;XIH;?H;�5H;�-H;3'H;s"H;�H;      �NH;NOH;�QH;UH;�YH;�_H;�fH;dnH;�vH;,H;�H;��H;R�H;��H;x�H;ܰH;��H;��H;��H;��H;)�H;�H;��H;��H;�H;�H;��H;p�H;��H;��H;V�H;��H;q�H;��H;�H;%�H;?�H;%�H;�H;��H;q�H;��H;V�H;��H;��H;p�H;��H;�H;�H;��H;��H;�H;)�H;��H;��H;��H;��H;ܰH;x�H;��H;R�H;��H;�H;,H;�vH;dnH;�fH;�_H;�YH;UH;�QH;NOH;      �rH;HsH;�tH;�wH;{H;�H;��H;i�H;��H;�H;��H;W�H;ժH;�H;��H;��H;�H;��H;9�H;�H;r�H;��H;(�H;g�H;n�H;�H;n�H;��H;��H;V�H;��H;q�H;��H;�H;_�H;l�H;d�H;l�H;_�H;�H;��H;q�H;��H;V�H;��H;��H;n�H;�H;n�H;g�H;(�H;��H;r�H;�H;9�H;��H;�H;��H;��H;�H;ժH;W�H;��H;�H;��H;i�H;��H;�H;{H;�wH;�tH;HsH;      �H;:�H;z�H;�H;�H;{�H;V�H;��H;L�H; �H;�H;�H;��H;ͼH;��H;��H;��H;|�H;��H;��H;��H;��H;��H;��H;N�H;��H;��H;��H;X�H;��H;q�H;��H;�H;_�H;��H;��H;��H;��H;��H;_�H;�H;��H;q�H;��H;X�H;��H;��H;��H;N�H;��H;��H;��H;��H;��H;��H;|�H;��H;��H;��H;ͼH;��H;�H;�H; �H;L�H;��H;V�H;{�H;�H;�H;z�H;:�H;      ��H;�H;�H;f�H;i�H;�H;ͫH;�H;��H;g�H;H�H;.�H;�H;��H;;�H;��H;��H;��H;-�H;��H;��H;��H;C�H;��H;��H;��H;��H;c�H;��H;q�H;��H;�H;X�H;��H;��H;��H;��H;��H;��H;��H;X�H;�H;��H;q�H;��H;c�H;��H;��H;��H;��H;C�H;��H;��H;��H;-�H;��H;��H;��H;;�H;��H;�H;.�H;H�H;g�H;��H;�H;ͫH;�H;i�H;f�H;�H;�H;      ��H;�H;��H;ñH;u�H;r�H;��H;[�H;�H;�H;�H;�H;
�H;��H;��H;k�H;��H;4�H;M�H;5�H;��H;�H;��H;��H;��H;��H;L�H;��H;y�H;��H;�H;_�H;��H;��H;��H;��H;��H;��H;��H;��H;��H;_�H;�H;��H;y�H;��H;L�H;��H;��H;��H;��H;�H;��H;5�H;M�H;4�H;��H;k�H;��H;��H;
�H;�H;�H;�H;�H;[�H;��H;r�H;u�H;ñH;��H;�H;      �H;W�H;�H;ۺH;6�H;ɽH;��H;��H;��H;m�H;��H;Q�H;��H;,�H;��H;��H;��H;��H;r�H;�H;z�H;��H;��H;��H;��H;B�H;��H;V�H;��H;�H;_�H;��H;��H;��H;��H;��H;��H;��H;��H;��H;��H;��H;_�H;�H;��H;V�H;��H;B�H;��H;��H;��H;��H;z�H;�H;r�H;��H;��H;��H;��H;,�H;��H;Q�H;��H;m�H;��H;��H;��H;ɽH;6�H;ۺH;�H;W�H;      q�H;��H;�H;�H;�H;r�H;�H;��H;��H;��H;"�H;`�H;��H;��H;��H;��H;v�H;8�H;��H;(�H;W�H;j�H;m�H;E�H;��H;��H;-�H;��H;��H;%�H;l�H;��H;��H;��H;��H;��H;��H;��H;��H;��H;��H;��H;l�H;%�H;��H;��H;-�H;��H;��H;E�H;m�H;j�H;W�H;(�H;��H;8�H;v�H;��H;��H;��H;��H;`�H;"�H;��H;��H;��H;�H;r�H;�H;�H;�H;��H;      E�H;U�H;��H;��H;��H;��H;��H;G�H;4�H;3�H;F�H;O�H;V�H;l�H;l�H;Q�H;�H;��H;�H;q�H;��H;��H;��H;^�H;6�H;��H;.�H;��H;��H;?�H;d�H;��H;��H;��H;��H;��H;��H;��H;��H;��H;��H;��H;d�H;?�H;��H;��H;.�H;��H;6�H;^�H;��H;��H;��H;q�H;�H;��H;�H;Q�H;l�H;l�H;V�H;O�H;F�H;3�H;4�H;G�H;��H;��H;��H;��H;��H;U�H;      q�H;��H;�H;�H;�H;r�H;�H;��H;��H;��H;"�H;`�H;��H;��H;��H;��H;v�H;8�H;��H;(�H;W�H;j�H;m�H;E�H;��H;��H;-�H;��H;��H;%�H;l�H;��H;��H;��H;��H;��H;��H;��H;��H;��H;��H;��H;l�H;%�H;��H;��H;-�H;��H;��H;E�H;m�H;j�H;W�H;(�H;��H;8�H;v�H;��H;��H;��H;��H;`�H;"�H;��H;��H;��H;�H;r�H;�H;�H;�H;��H;      �H;W�H;�H;ۺH;6�H;ɽH;��H;��H;��H;m�H;��H;Q�H;��H;,�H;��H;��H;��H;��H;r�H;�H;z�H;��H;��H;��H;��H;B�H;��H;V�H;��H;�H;_�H;��H;��H;��H;��H;��H;��H;��H;��H;��H;��H;��H;_�H;�H;��H;V�H;��H;B�H;��H;��H;��H;��H;z�H;�H;r�H;��H;��H;��H;��H;,�H;��H;Q�H;��H;m�H;��H;��H;��H;ɽH;6�H;ۺH;�H;W�H;      ��H;�H;��H;ñH;u�H;r�H;��H;[�H;�H;�H;�H;�H;
�H;��H;��H;k�H;��H;4�H;M�H;5�H;��H;�H;��H;��H;��H;��H;L�H;��H;y�H;��H;�H;_�H;��H;��H;��H;��H;��H;��H;��H;��H;��H;_�H;�H;��H;y�H;��H;L�H;��H;��H;��H;��H;�H;��H;5�H;M�H;4�H;��H;k�H;��H;��H;
�H;�H;�H;�H;�H;[�H;��H;r�H;u�H;ñH;��H;�H;      ��H;�H;�H;f�H;i�H;�H;ͫH;�H;��H;g�H;H�H;.�H;�H;��H;;�H;��H;��H;��H;-�H;��H;��H;��H;C�H;��H;��H;��H;��H;c�H;��H;q�H;��H;�H;X�H;��H;��H;��H;��H;��H;��H;��H;X�H;�H;��H;q�H;��H;c�H;��H;��H;��H;��H;C�H;��H;��H;��H;-�H;��H;��H;��H;;�H;��H;�H;.�H;H�H;g�H;��H;�H;ͫH;�H;i�H;f�H;�H;�H;      �H;:�H;z�H;�H;�H;{�H;V�H;��H;L�H; �H;�H;�H;��H;ͼH;��H;��H;��H;|�H;��H;��H;��H;��H;��H;��H;N�H;��H;��H;��H;X�H;��H;q�H;��H;�H;_�H;��H;��H;��H;��H;��H;_�H;�H;��H;q�H;��H;X�H;��H;��H;��H;N�H;��H;��H;��H;��H;��H;��H;|�H;��H;��H;��H;ͼH;��H;�H;�H; �H;L�H;��H;V�H;{�H;�H;�H;z�H;:�H;      �rH;HsH;�tH;�wH;{H;�H;��H;i�H;��H;�H;��H;W�H;ժH;�H;��H;��H;�H;��H;9�H;�H;r�H;��H;(�H;g�H;n�H;�H;n�H;��H;��H;V�H;��H;q�H;��H;�H;_�H;l�H;d�H;l�H;_�H;�H;��H;q�H;��H;V�H;��H;��H;n�H;�H;n�H;g�H;(�H;��H;r�H;�H;9�H;��H;�H;��H;��H;�H;ժH;W�H;��H;�H;��H;i�H;��H;�H;{H;�wH;�tH;HsH;      �NH;NOH;�QH;UH;�YH;�_H;�fH;dnH;�vH;,H;�H;��H;R�H;��H;x�H;ܰH;��H;��H;��H;��H;)�H;�H;��H;��H;�H;�H;��H;p�H;��H;��H;V�H;��H;q�H;��H;�H;%�H;?�H;%�H;�H;��H;q�H;��H;V�H;��H;��H;p�H;��H;�H;�H;��H;��H;�H;)�H;��H;��H;��H;��H;ܰH;x�H;��H;R�H;��H;�H;,H;�vH;dnH;�fH;�_H;�YH;UH;�QH;NOH;      �H;�H;s"H;3'H;�-H;�5H;?H;XIH;eTH;�_H;�kH;9wH;��H;��H;��H;��H;��H;��H;�H;��H;��H;��H;��H;��H;��H;��H;��H;��H;>�H;��H;��H;X�H;��H;y�H;��H;��H;��H;��H;��H;y�H;��H;X�H;��H;��H;>�H;��H;��H;��H;��H;��H;��H;��H;��H;��H;�H;��H;��H;��H;��H;��H;��H;9wH;�kH;�_H;eTH;XIH;?H;�5H;�-H;3'H;s"H;�H;      M�G;��G;��G;��G;��G;��G;WH;H;�'H;7H;�FH;/VH;MeH;�sH;d�H;�H;ٙH;��H;�H;��H;�H;��H;H�H;�H;#�H;��H;m�H;��H;��H;p�H;��H;��H;c�H;��H;V�H;��H;��H;��H;V�H;��H;c�H;��H;��H;p�H;��H;��H;m�H;��H;#�H;�H;H�H;��H;�H;��H;�H;��H;ٙH;�H;d�H;�sH;MeH;/VH;�FH;7H;�'H;H;WH;��G;��G;��G;��G;��G;      puG;3xG;/�G;��G;�G;��G;�G;��G;��G;�H;IH;�+H;�?H;�RH;�dH;�uH;ńH;��H;�H;�H;��H;�H;<�H;Y�H;}�H;��H;t�H;m�H;��H;��H;n�H;��H;��H;L�H;��H;-�H;.�H;-�H;��H;L�H;��H;��H;n�H;��H;��H;m�H;t�H;��H;}�H;Y�H;<�H;�H;��H;�H;�H;��H;ńH;�uH;�dH;�RH;�?H;�+H;IH;�H;��G;��G;�G;��G;�G;��G;/�G;3xG;      ��F;q�F;��F;�F;��F;�G;�FG; pG;\�G;l�G;�G;��G;!H;2)H;�@H;xVH;VjH;5|H;=�H;f�H;��H;E�H;g�H;;�H;��H;E�H;��H;��H;��H;�H;�H;��H;��H;��H;B�H;��H;��H;��H;B�H;��H;��H;��H;�H;�H;��H;��H;��H;E�H;��H;;�H;g�H;E�H;��H;f�H;=�H;5|H;VjH;xVH;�@H;2)H;!H;��G;�G;l�G;\�G; pG;�FG;�G;��F;�F;��F;q�F;      �lD;#~D;��D;�D;�[E;+�E;�/F;�F;��F;$8G;�uG;'�G;t�G;��G;cH;�/H;aIH;�`H;uH;�H;��H;V�H;گH;��H;�H;��H;}�H;#�H;��H;�H;n�H;N�H;��H;��H;��H;��H;6�H;��H;��H;��H;��H;N�H;n�H;�H;��H;#�H;}�H;��H;�H;��H;گH;V�H;��H;�H;uH;�`H;aIH;�/H;cH;��G;t�G;'�G;�uG;$8G;��F;�F;�/F;+�E;�[E;�D;��D;#~D;      �_?;	�?;6�?;�@;��A;��B;��C;3�D;~hE;#F;[�F;G;�mG;E�G;$�G;t�G;� H;C>H;�XH;�oH;i�H;��H;#�H;\�H;��H;;�H;Y�H;�H;��H;��H;g�H;��H;��H;��H;��H;E�H;^�H;E�H;��H;��H;��H;��H;g�H;��H;��H;�H;Y�H;;�H;��H;\�H;#�H;��H;i�H;�oH;�XH;C>H;� H;t�G;$�G;E�G;�mG;G;[�F;#F;~hE;3�D;��C;��B;��A;�@;6�?;	�?;      ��4;x�4;��5;Rl7;�^9;��;;�=;f�?;��A;�C;��D;��E;�F;�(G;ˀG;8�G;�G;jH;�5H;�RH;&lH;��H;˓H;#�H;گH;g�H;<�H;H�H;��H;��H;(�H;��H;C�H;��H;��H;m�H;��H;m�H;��H;��H;C�H;��H;(�H;��H;��H;H�H;<�H;g�H;گH;#�H;˓H;��H;&lH;�RH;�5H;jH;�G;8�G;ˀG;�(G;�F;��E;��D;�C;��A;f�?;�=;��;;�^9;Rl7;��5;x�4;      �d;� ;�";�%;d�(;�i-;�2;,�6;�:;0>;�A;�XC;y�D;KF;S�F;�WG;3�G;w�G;�H;�0H;PH;�jH;��H;��H;V�H;E�H;�H;��H;��H;�H;��H;��H;��H;�H;��H;j�H;��H;j�H;��H;�H;��H;��H;��H;�H;��H;��H;�H;E�H;V�H;��H;��H;�jH;PH;�0H;�H;w�G;3�G;�WG;S�F;KF;y�D;�XC;�A;0>;�:;,�6;�2;�i-;d�(;�%;�";� ;      ���:�A�:���:�w;�
;5;��;}$;�{,;ǂ3;_9;�>;ayA;�C;,�E;>�F;Z4G;��G;��G;nH;�.H;PH;&lH;i�H;��H;��H;��H;�H;��H;)�H;r�H;��H;��H;��H;z�H;W�H;��H;W�H;z�H;��H;��H;��H;r�H;)�H;��H;�H;��H;��H;��H;i�H;&lH;PH;�.H;nH;��G;��G;Z4G;>�F;,�E;�C;ayA;�>;_9;ǂ3;�{,;}$;��;5;�
;�w;���:�A�:      �v[:�Ad:5�}:^�:��:/��:C�:��;P;� ;G+;�3;:�:;i�?;�B;�
E;�YF;
G;R�G;��G;nH;�0H;�RH;�oH;�H;f�H;�H;��H;��H;��H;�H;��H;��H;5�H;�H;(�H;q�H;(�H;�H;5�H;��H;��H;�H;��H;��H;��H;�H;f�H;�H;�oH;�RH;�0H;nH;��G;R�G;
G;�YF;�
E;�B;i�?;:�:;�3;G+;� ;P;��;C�:/��:��:^�:5�}:�Ad:      ��S���D�/�����E�'7��9a�R:���:���:@��:X>;G";]P.;�l7;B�=;�B;%�D;�8F;XG;R�G;��G;�H;�5H;�XH;uH;=�H;�H;�H;�H;��H;9�H;��H;-�H;M�H;r�H;��H;�H;��H;r�H;M�H;-�H;��H;9�H;��H;�H;�H;�H;=�H;uH;�XH;�5H;�H;��G;R�G;XG;�8F;%�D;�B;B�=;�l7;]P.;G";X>;@��:���:���:a�R:��9E�'7���/����D�      �D^��/X��qF�(}*�'���P���D��Ҭ�jh:��:���:ȏ; �;��);��4;p�<;`�A;f�D;�8F;
G;��G;w�G;jH;C>H;�`H;5|H;��H;��H;��H;��H;��H;|�H;��H;4�H;��H;8�H;��H;8�H;��H;4�H;��H;|�H;��H;��H;��H;��H;��H;5|H;�`H;C>H;jH;w�G;��G;
G;�8F;f�D;`�A;p�<;��4;��); �;ȏ;���:��:jh:�Ҭ��D��P��'��(}*��qF��/X�      s��v��,�ܻ�ƻB󩻜��gFL����θ��&��M�-:g�:���:v;>&;��3;�8<;`�A;%�D;�YF;Z4G;3�G;�G;� H;aIH;VjH;ńH;ٙH;��H;��H;�H;��H;��H;��H;��H;v�H;�H;v�H;��H;��H;��H;��H;�H;��H;��H;ٙH;ńH;VjH;aIH;� H;�G;3�G;Z4G;�YF;%�D;`�A;�8<;��3;>&;v;���:g�:M�-:&��θ�����gFL����B��ƻ,�ܻv��      ;�V�z5S�Y6H�x�6�� �3,�n?ػG���D^����4�D��9�3�:> �:��;]%;��3;p�<;�B;�
E;>�F;�WG;8�G;t�G;�/H;xVH;�uH;�H;��H;ܰH;��H;��H;��H;k�H;��H;��H;Q�H;��H;��H;k�H;��H;��H;��H;ܰH;��H;�H;�uH;xVH;�/H;t�G;8�G;�WG;>�F;�
E;�B;p�<;��3;]%;��;> �:�3�:�94�D�����D^�G��n?ػ3,�� �x�6�Y6H�z5S�      ����-��#Ȥ�d���ݫ���f�G�=����	�ܻ�*��>o5�u����P(7F�}:�m�:��;>&;��4;B�=;�B;,�E;S�F;ˀG;$�G;cH;�@H;�dH;d�H;��H;x�H;��H;��H;;�H;��H;��H;��H;l�H;��H;��H;��H;;�H;��H;��H;x�H;��H;d�H;�dH;�@H;cH;$�G;ˀG;S�F;,�E;�B;B�=;��4;>&;��;�m�:F�}:�P(7u���>o5��*��	�ܻ���G�=��f�ݫ��d���#Ȥ��-��      xc��8�|����켔�Ҽg���`�����r�E:�%,�#ߵ�Y/X���º̬�F�}:> �:v;��);�l7;i�?;�C;KF;�(G;E�G;��G;2)H;�RH;�sH;��H;��H;�H;ͼH;��H;��H;,�H;��H;l�H;��H;,�H;��H;��H;ͼH;�H;��H;��H;�sH;�RH;2)H;��G;E�G;�(G;KF;�C;i�?;�l7;��);v;> �:F�}:̬���ºY/X�#ߵ�%,�E:���r�`���g�����Ҽ��|����8�      �&K���G�ȟ>��0�:y�vc�d��)������!�V����ƻfod���º�P(7�3�:���: �;]P.;:�:;ayA;y�D;�F;�mG;t�G;!H;�?H;MeH;��H;R�H;ժH;��H;�H;
�H;��H;��H;V�H;��H;��H;
�H;�H;��H;ժH;R�H;��H;MeH;�?H;!H;t�G;�mG;�F;y�D;ayA;:�:;]P.; �;���:�3�:�P(7��ºfod��ƻ��!�V����)���d��vc�:y��0�ȟ>���G�      鰒�Z��������}��c���D�/%��8���Ҽ	c����f�����ƻY/X�u����9g�:ȏ;G";�3;�>;�XC;��E;G;'�G;��G;�+H;/VH;9wH;��H;W�H;�H;.�H;�H;Q�H;`�H;O�H;`�H;Q�H;�H;.�H;�H;W�H;��H;9wH;/VH;�+H;��G;'�G;G;��E;�XC;�>;�3;G";ȏ;g�:�9u���Y/X��ƻ�����f�	c����Ҽ�8�/%���D��c���}�����Z��      \Pν��ʽ*8�������������0�f�u�;���K��Ȥ���f���#ߵ�>o5�4�D�M�-:���:X>;G+;_9;�A;��D;[�F;�uG;�G;IH;�FH;�kH;�H;��H;�H;H�H;�H;��H;"�H;F�H;"�H;��H;�H;H�H;�H;��H;�H;�kH;�FH;IH;�G;�uG;[�F;��D;�A;_9;G+;X>;���:M�-:4�D�>o5�#ߵ�����f�Ȥ�K����u�;�0�f������������*8����ʽ      ���N9�C[��s�R�ؽ���s����}���G��K��	c��!�V�%,��*�����&����:@��:� ;ǂ3;0>;�C;#F;$8G;l�G;�H;7H;�_H;,H;�H; �H;g�H;�H;m�H;��H;3�H;��H;m�H;�H;g�H; �H;�H;,H;�_H;7H;�H;l�G;$8G;#F;�C;0>;ǂ3;� ;@��:��:&������*��%,�!�V�	c��K�����G���}��s����R�ؽ�s�C[�N9�      }�=���:���0��Q"�e�����ZPν�榽%����G�����Ҽ���E:�	�ܻ�D^�θ��jh:���:P;�{,;�:;��A;~hE;��F;\�G;��G;�'H;eTH;�vH;��H;L�H;��H;�H;��H;��H;4�H;��H;��H;�H;��H;L�H;��H;�vH;eTH;�'H;��G;\�G;��F;~hE;��A;�:;�{,;P;���:jh:θ���D^�	�ܻE:������Ҽ����G�%���榽ZPν����e��Q"���0���:�      
Dx��s���f�QS���:����B[��7ս�榽��}�u�;��8�)�����r����G������Ҭ����:��;}$;,�6;f�?;3�D;�F; pG;��G;H;XIH;dnH;i�H;��H;�H;[�H;��H;��H;G�H;��H;��H;[�H;�H;��H;i�H;dnH;XIH;H;��G; pG;�F;3�D;f�?;,�6;}$;��;���:�Ҭ����G�������r�)����8�u�;���}��榽�7սB[������:�QS���f��s�      �*���0��ȥ��&���jk��H��#%�B[�ZPν�s��0�f�/%�d��`���G�=�n?ػgFL��D�a�R:C�:��;�2;�=;��C;�/F;�FG;�G;WH;?H;�fH;��H;V�H;ͫH;��H;��H;�H;��H;�H;��H;��H;ͫH;V�H;��H;�fH;?H;WH;�G;�FG;�/F;��C;�=;�2;��;C�:a�R:�D�gFL�n?ػG�=�`���d��/%�0�f��s��ZPνB[��#%��H�jk�&���ȥ���0��      �þ��������R��f쏾�s��H����������������D�vc�g����f�3,�����P����9/��:5;�i-;��;;��B;+�E;�G;��G;��G;�5H;�_H;�H;{�H;�H;r�H;ɽH;r�H;��H;r�H;ɽH;r�H;�H;{�H;�H;�_H;�5H;��G;��G;�G;+�E;��B;��;;�i-;5;/��:��9�P�����3,��f�g���vc���D���������������H��s�f쏾�R���������      ����fYؾ�þ�ê�f쏾jk���:�e�R�ؽ�����c�:y���Ҽݫ��� �B�'��E�'7��:�
;d�(;�^9;��A;�[E;��F;�G;��G;�-H;�YH;{H;�H;i�H;u�H;6�H;�H;��H;�H;6�H;u�H;i�H;�H;{H;�YH;�-H;��G;�G;��F;�[E;��A;�^9;d�(;�
;��:E�'7'��B�� �ݫ����Ҽ:y��c�����R�ؽe���:�jk�f쏾�ê��þfYؾ��      ��=������I��þ�R��&���QS��Q"��s�����}��0���d���x�6��ƻ(}*����^�:�w;�%;Rl7;�@;�D;�F;��G;��G;3'H;UH;�wH;�H;f�H;ñH;ۺH;�H;��H;�H;ۺH;ñH;f�H;�H;�wH;UH;3'H;��G;��G;�F;�D;�@;Rl7;�%;�w;^�:���(}*��ƻx�6�d����켟0���}�����s��Q"�QS�&����R���þIᾁ���=��      ���>��&�
�����fYؾ���ȥ����f���0�C[�*8������ȟ>�|���#Ȥ�Y6H�,�ܻ�qF�/��5�}:���:�";��5;6�?;��D;��F;/�G;��G;s"H;�QH;�tH;z�H;�H;��H;�H;�H;��H;�H;�H;��H;�H;z�H;�tH;�QH;s"H;��G;/�G;��F;��D;6�?;��5;�";���:5�}:/���qF�,�ܻY6H�#Ȥ�|���ȟ>�����*8��C[���0���f�ȥ�����fYؾ����&�
�>��      �� �k��>��=���������0���s���:�N9���ʽZ����G��8��-��z5S�v���/X���D��Ad:�A�:� ;x�4;	�?;#~D;q�F;3xG;��G;�H;NOH;HsH;:�H;�H;�H;W�H;��H;U�H;��H;W�H;�H;�H;:�H;HsH;NOH;�H;��G;3xG;q�F;#~D;	�?;x�4;� ;�A�:�Ad:��D��/X�v��z5S��-���8���G�Z����ʽN9���:��s��0��������=��>��k��      .Eb�I]�tN�ߛ7����e� �{�˾��	�j��!,�J���0��m���,˼��x�E���1��a���R�:f�:2;��1;n+>;��C;�vF;�G;��G;>H;�gH;Z�H;v�H;8�H;�H;��H;(�H;��H;(�H;��H;�H;8�H;v�H;Z�H;�gH;>H;��G;�G;�vF;��C;n+>;��1;2;f�:R�:a����1��E����x�,˼��m�0��J����!,�	�j���{�˾e� ����ߛ7�tN�I]�      I]�N�W��TI�v3��D�������Ǿb���ȟf� )� ��W;���Fi��k�x�Ǽ�[t�8�	�(Ȅ�sX��ϟ:���:%�;�I2;�Y>;qD;�~F;\�G;+H;�>H;�hH;�H;�H;r�H;7�H;��H;S�H;��H;S�H;��H;7�H;r�H;�H;�H;�hH;�>H;+H;\�G;�~F;qD;�Y>;�I2;%�;���:ϟ:sX��(Ȅ�8�	��[t�x�Ǽ�k��Fi�W;�� �� )�ȟf�b�����Ǿ�����D�v3��TI�N�W�      tN��TI���;��'��k���i���f󐾖Z��K ��s�&����&^����"����g����Ѩu�R!���1<:��:n
;�f3;-�>;�AD;ՕF;�G;�H;UAH;jH;\�H;ߟH;(�H;ԻH;k�H;��H;B�H;��H;k�H;ԻH;(�H;ߟH;\�H;jH;UAH;�H;�G;ՕF;�AD;-�>;�f3;n
;��:�1<:R!��Ѩu������g��"�����&^�&����s潎K ��Z�f�i������k��'���;��TI�      ߛ7�v3��'����e� ��{Ծ
���6���]�F�����ӽ���;�L�1v�x뮼,T�ǘ��PV�p�=�2(i:`��:!z ;�#5;�?;2�D;�F;�G;�H;�EH;�mH;��H;}�H;j�H;ۼH;4�H;O�H;��H;O�H;4�H;ۼH;j�H;}�H;��H;�mH;�EH;�H;�G;�F;2�D;�?;�#5;!z ;`��:2(i:p�=��PV�ǘ�,T�x뮼1v�;�L�����ӽ���]�F�6���
����{Ծe� �����'�v3�      ����D��k�e� �<�ݾS���C͓�ȟf��>/�x��~'��n섽/�6�Rt��v��?�:�Tʻ�.�ݷ��s�:2; �$;�X7;��@;	E;:�F;P�G;�H;EKH;�qH;��H;ɣH;�H;�H;.�H;D�H;��H;D�H;.�H;�H;�H;ɣH;��H;�qH;EKH;�H;P�G;:�F;	E;��@;�X7; �$;2;�s�:ݷ��.�Tʻ?�:��v��Rt�/�6�n섽~'��x���>/�ȟf�C͓�S���<�ݾe� ��k��D�      e� ������쾻{ԾS���b���9�x�rSC��^�ͻ޽%���Q�e����ѼG������R�����դ8��:�X;��);5�9;-�A;��E;�G;2�G;s H;DRH;�vH;v�H;��H;:�H;��H;r�H;u�H;��H;u�H;r�H;��H;:�H;��H;v�H;�vH;DRH;s H;2�G;�G;��E;-�A;5�9;��);�X;��:դ8����R�����G���Ѽ��Q�e�%���ͻ޽�^�rSC�9�x�b���S����{Ծ�쾃���      {�˾��Ǿi���
���C͓�9�x�ؘJ��K �H��� �������?���t뮼�[�����3|��W��<�:v~�:';�
/;�f<;�C;� F;�MG;��G;9,H;sZH;�|H;ǖH;©H;��H;��H;��H;��H;��H;��H;��H;��H;��H;©H;ǖH;�|H;sZH;9,H;��G;�MG;� F;�C;�f<;�
/;';v~�:<�:�W��3|������[�t뮼����?���� ��H����K �ؘJ�9�x�C͓�
���i�����Ǿ      ��b���f�6���ȟf�rSC��K �Gn����Ž����Z��k��|ռX��Ey-����x.�w���O�:�*�:��;o4;s�>;)D;�vF;I�G;��G;�8H;\cH;x�H;��H;[�H;e�H;��H;��H;K�H;f�H;K�H;��H;��H;e�H;[�H;��H;x�H;\cH;�8H;��G;I�G;�vF;)D;s�>;o4;��;�*�:�O�:w��x.����Ey-�X���|ռ�k��Z������ŽGn���K �rSC�ȟf�6���f�b���      	�j�ȟf��Z�]�F��>/��^�H�����Ž- ���Fi�kQ+�Ot�PT��H�W�����1��iȺ�U�9�O�:	Y;��(;T�8;1A;�E;!�F;|�G;�H;�EH;�lH;��H;��H;8�H;d�H;��H;��H;��H;��H;��H;��H;��H;d�H;8�H;��H;��H;�lH;�EH;�H;|�G;!�F;�E;1A;T�8;��(;	Y;�O�:�U�9iȺ�1�����H�W�PT��Ot�kQ+��Fi�- ����ŽH����^��>/�]�F��Z�ȟf�      �!,� )��K ����x��ͻ޽ ������Fi���0�����跼z�x�����.��b�(�����)i:���:��;�0;��<;�C;��E;)<G;
�G;�#H;kSH;�vH;�H;�H;E�H;t�H;4�H;��H;��H;n�H;��H;��H;4�H;t�H;E�H;�H;�H;�vH;kSH;�#H;
�G;)<G;��E;�C;��<;�0;��;���:�)i:���b�(��.�����z�x��跼�����0��Fi���� ��ͻ޽x������K � )�      J��� ��s��ӽ~'��%�������Z�kQ+�����"��G����0���׻͕b��W���V�9�:�_;�)';/Y7;G#@;S�D;�F;+�G;��G;A7H;aH;��H;Z�H;��H;l�H;��H;��H;{�H;A�H;.�H;A�H;{�H;��H;��H;l�H;��H;Z�H;��H;aH;A7H;��G;+�G;�F;S�D;G#@;/Y7;�)';�_;�:�V�9�W��͕b���׻��0�G���"�����kQ+��Z����%���~'���ӽ�s� ��      0��W;��&������n섽Q�e���?��k�Ot��跼G��ee7�����Ǆ��0�6�t�^t�:�*�:�
;�1;��<;��B;N�E;G;�G;iH;wIH;`nH;��H;��H;�H;��H;��H;�H;��H;�H;��H;�H;��H;�H;��H;��H;�H;��H;��H;`nH;wIH;iH;�G;G;N�E;��B;��<;�1;�
;�*�:^t�:6�t��0��Ǆ����ee7�G���跼Ot�k���?�Q�e�n섽���&���W;��      m��Fi��&^�;�L�/�6������|ռPT��z�x���0��������0���ڷ�xm`:��:��;��*;}�8;G�@;d�D;��F;}G;��G;�0H;�ZH;m{H;��H;֧H;�H;��H;��H;|�H;��H;��H;d�H;��H;��H;|�H;��H;��H;�H;֧H;��H;m{H;�ZH;�0H;��G;}G;��F;d�D;G�@;}�8;��*;��;��:xm`:�ڷ�0��������껣�0�z�x�PT���|ռ����/�6�;�L��&^��Fi�      ���k���1v�Rt��Ѽt뮼X��H�W������׻�Ǆ�0�����3<:v��:;Y;�s%;=$5;�Y>;-`C;��E;O)G;u�G;"H;GH;lkH;�H;��H;��H;ȻH;��H;��H;��H;g�H;_�H;�H;_�H;g�H;��H;��H;��H;ȻH;��H;��H;�H;lkH;GH;"H;u�G;O)G;��E;-`C;�Y>;=$5;�s%;;Y;v��:�3<:���0���Ǆ���׻���H�W�X��t뮼�ѼRt�1v����k�      ,˼x�Ǽ�"��x뮼�v��G���[�Ey-�����.��͕b��0㺈ڷ��3<:L�:_\;��!;1J2;�f<;/B;QBE;J�F;a�G; �G;�3H;�[H;{H;��H;��H;P�H;��H;6�H;��H;B�H;A�H;��H;��H;��H;A�H;B�H;��H;6�H;��H;P�H;��H;��H;{H;�[H;�3H; �G;a�G;J�F;QBE;/B;�f<;1J2;��!;_\;L�:�3<:�ڷ��0�͕b��.�����Ey-��[�G���v��x뮼�"��x�Ǽ      ��x��[t���g�,T�?�:������������1��b�(��W��6�t�xm`:v��:_\;pz ;�0;�;;9<A;?�D;�vF;�bG;d�G;� H;�LH;�nH;p�H;~�H;��H;��H;Z�H;��H;H�H;_�H;��H;��H;�H;��H;��H;_�H;H�H;��H;Z�H;��H;��H;~�H;p�H;�nH;�LH;� H;d�G;�bG;�vF;?�D;9<A;�;;�0;pz ;_\;v��:xm`:6�t��W��b�(��1������������?�:�,T���g��[t�      E��8�	����ǘ�Tʻ�R��3|�x.�iȺ����V�9^t�:��:;Y;��!;�0;-�:;�@;4BD;�1F;�7G;��G;�H;k?H;*cH;�H;m�H;:�H;<�H;>�H;��H;��H;��H;[�H;��H;��H;s�H;��H;��H;[�H;��H;��H;��H;>�H;<�H;:�H;m�H;�H;*cH;k?H;�H;��G;�7G;�1F;4BD;�@;-�:;�0;��!;;Y;��:^t�:�V�9���iȺx.�3|��R��Tʻǘ����8�	�      �1��(Ȅ�Ѩu��PV��.�����W��w��U�9�)i:�:�*�:��;�s%;1J2;�;;�@;�D;/F;>G;��G;�H;�4H;�YH;5wH;7�H;�H;	�H;�H;I�H;^�H;�H;�H;�H;*�H;E�H;��H;E�H;*�H;�H;�H;�H;^�H;I�H;�H;	�H;�H;7�H;5wH;�YH;�4H;�H;��G;>G;/F;�D;�@;�;;1J2;�s%;��;�*�:�:�)i:�U�9w���W������.��PV�Ѩu�(Ȅ�      a���sX��R!��p�=�ݷ�դ8<�:�O�:�O�:���:�_;�
;��*;=$5;�f<;9<A;4BD;/F;�G;��G;r�G;�,H;RH;UpH;�H;��H;r�H;�H;)�H;��H;��H;��H;?�H;��H;��H;|�H;��H;|�H;��H;��H;?�H;��H;��H;��H;)�H;�H;r�H;��H;�H;UpH;RH;�,H;r�G;��G;�G;/F;4BD;9<A;�f<;=$5;��*;�
;�_;���:�O�:�O�:<�:դ8ݷ�p�=�R!��sX��      R�:ϟ:�1<:2(i:�s�:��:v~�:�*�:	Y;��;�)';�1;}�8;�Y>;/B;?�D;�1F;>G;��G;%�G;�(H;�MH;qkH;C�H;c�H;v�H;��H;�H;t�H;��H;$�H;�H;�H;D�H;��H;��H;��H;��H;��H;D�H;�H;�H;$�H;��H;t�H;�H;��H;v�H;c�H;C�H;qkH;�MH;�(H;%�G;��G;>G;�1F;?�D;/B;�Y>;}�8;�1;�)';��;	Y;�*�:v~�:��:�s�:2(i:�1<:ϟ:      f�:���:��:`��:2;�X;';��;��(;�0;/Y7;��<;G�@;-`C;QBE;�vF;�7G;��G;r�G;�(H;�KH;�hH;.�H;O�H;��H;��H;��H;O�H;�H;��H;��H;A�H;��H;��H;��H;��H;��H;��H;��H;��H;��H;A�H;��H;��H;�H;O�H;��H;��H;��H;O�H;.�H;�hH;�KH;�(H;r�G;��G;�7G;�vF;QBE;-`C;G�@;��<;/Y7;�0;��(;��;';�X;2;`��:��:���:      2;%�;n
;!z ; �$;��);�
/;o4;T�8;��<;G#@;��B;d�D;��E;J�F;�bG;��G;�H;�,H;�MH;�hH;B�H;��H;��H;ΰH;��H;��H;��H;2�H;��H;^�H;�H;0�H;��H;��H;P�H;��H;P�H;��H;��H;0�H;�H;^�H;��H;2�H;��H;��H;��H;ΰH;��H;��H;B�H;�hH;�MH;�,H;�H;��G;�bG;J�F;��E;d�D;��B;G#@;��<;T�8;o4;�
/;��); �$;!z ;n
;%�;      ��1;�I2;�f3;�#5;�X7;5�9;�f<;s�>;1A;�C;S�D;N�E;��F;O)G;a�G;d�G;�H;�4H;RH;qkH;.�H;��H;�H;ɯH;�H;V�H;L�H; �H;��H;��H;u�H;��H;o�H;��H;��H;�H;\�H;�H;��H;��H;o�H;��H;u�H;��H;��H; �H;L�H;V�H;�H;ɯH;�H;��H;.�H;qkH;RH;�4H;�H;d�G;a�G;O)G;��F;N�E;S�D;�C;1A;s�>;�f<;5�9;�X7;�#5;�f3;�I2;      n+>;�Y>;-�>;�?;��@;-�A;�C;)D;�E;��E;�F;G;}G;u�G; �G;� H;k?H;�YH;UpH;C�H;O�H;��H;ɯH;�H;��H;��H;6�H;��H;��H;��H;O�H; �H;��H;��H;H�H;��H;��H;��H;H�H;��H;��H; �H;O�H;��H;��H;��H;6�H;��H;��H;�H;ɯH;��H;O�H;C�H;UpH;�YH;k?H;� H; �G;u�G;}G;G;�F;��E;�E;)D;�C;-�A;��@;�?;-�>;�Y>;      ��C;qD;�AD;2�D;	E;��E;� F;�vF;!�F;)<G;+�G;�G;��G;"H;�3H;�LH;*cH;5wH;�H;c�H;��H;ΰH;�H;��H;=�H;��H;��H;^�H;c�H;��H;��H;f�H;��H;@�H;��H;C�H;L�H;C�H;��H;@�H;��H;f�H;��H;��H;c�H;^�H;��H;��H;=�H;��H;�H;ΰH;��H;c�H;�H;5wH;*cH;�LH;�3H;"H;��G;�G;+�G;)<G;!�F;�vF;� F;��E;	E;2�D;�AD;qD;      �vF;�~F;ՕF;�F;:�F;�G;�MG;I�G;|�G;
�G;��G;iH;�0H;GH;�[H;�nH;�H;7�H;��H;v�H;��H;��H;V�H;��H;��H;W�H;$�H;�H;��H;��H;�H;S�H;6�H;��H;m�H;��H;��H;��H;m�H;��H;6�H;S�H;�H;��H;��H;�H;$�H;W�H;��H;��H;V�H;��H;��H;v�H;��H;7�H;�H;�nH;�[H;GH;�0H;iH;��G;
�G;|�G;I�G;�MG;�G;:�F;�F;ՕF;�~F;      �G;\�G;�G;�G;P�G;2�G;��G;��G;�H;�#H;A7H;wIH;�ZH;lkH;{H;p�H;m�H;�H;r�H;��H;��H;��H;L�H;6�H;��H;$�H;�H;h�H;J�H;��H;7�H;�H;��H;��H;��H;�H;�H;�H;��H;��H;��H;�H;7�H;��H;J�H;h�H;�H;$�H;��H;6�H;L�H;��H;��H;��H;r�H;�H;m�H;p�H;{H;lkH;�ZH;wIH;A7H;�#H;�H;��G;��G;2�G;P�G;�G;�G;\�G;      ��G;+H;�H;�H;�H;s H;9,H;�8H;�EH;kSH;aH;`nH;m{H;�H;��H;~�H;:�H;	�H;�H;�H;O�H;��H; �H;��H;^�H;�H;h�H;]�H;��H;�H;�H;��H;z�H;��H;�H;^�H;g�H;^�H;�H;��H;z�H;��H;�H;�H;��H;]�H;h�H;�H;^�H;��H; �H;��H;O�H;�H;�H;	�H;:�H;~�H;��H;�H;m{H;`nH;aH;kSH;�EH;�8H;9,H;s H;�H;�H;�H;+H;      >H;�>H;UAH;�EH;EKH;DRH;sZH;\cH;�lH;�vH;��H;��H;��H;��H;��H;��H;<�H;�H;)�H;t�H;�H;2�H;��H;��H;c�H;��H;J�H;��H;$�H;��H;��H;k�H;��H;5�H;p�H;��H;��H;��H;p�H;5�H;��H;k�H;��H;��H;$�H;��H;J�H;��H;c�H;��H;��H;2�H;�H;t�H;)�H;�H;<�H;��H;��H;��H;��H;��H;��H;�vH;�lH;\cH;sZH;DRH;EKH;�EH;UAH;�>H;      �gH;�hH;jH;�mH;�qH;�vH;�|H;x�H;��H;�H;Z�H;��H;֧H;��H;P�H;��H;>�H;I�H;��H;��H;��H;��H;��H;��H;��H;��H;��H;�H;��H;��H;t�H;��H;%�H;y�H;��H;��H;��H;��H;��H;y�H;%�H;��H;t�H;��H;��H;�H;��H;��H;��H;��H;��H;��H;��H;��H;��H;I�H;>�H;��H;P�H;��H;֧H;��H;Z�H;�H;��H;x�H;�|H;�vH;�qH;�mH;jH;�hH;      Z�H;�H;\�H;��H;��H;v�H;ǖH;��H;��H;�H;��H;�H;�H;ȻH;��H;Z�H;��H;^�H;��H;$�H;��H;^�H;u�H;O�H;��H;�H;7�H;�H;��H;t�H;��H;.�H;��H;��H;��H;��H;��H;��H;��H;��H;��H;.�H;��H;t�H;��H;�H;7�H;�H;��H;O�H;u�H;^�H;��H;$�H;��H;^�H;��H;Z�H;��H;ȻH;�H;�H;��H;�H;��H;��H;ǖH;v�H;��H;��H;\�H;�H;      v�H;�H;ߟH;}�H;ɣH;��H;©H;[�H;8�H;E�H;l�H;��H;��H;��H;6�H;��H;��H;�H;��H;�H;A�H;�H;��H; �H;f�H;S�H;�H;��H;k�H;��H;.�H;z�H;��H;��H;��H;�H;�H;�H;��H;��H;��H;z�H;.�H;��H;k�H;��H;�H;S�H;f�H; �H;��H;�H;A�H;�H;��H;�H;��H;��H;6�H;��H;��H;��H;l�H;E�H;8�H;[�H;©H;��H;ɣH;}�H;ߟH;�H;      8�H;r�H;(�H;j�H;�H;:�H;��H;e�H;d�H;t�H;��H;��H;��H;��H;��H;H�H;��H;�H;?�H;�H;��H;0�H;o�H;��H;��H;6�H;��H;z�H;��H;%�H;��H;��H;��H;��H;�H;�H;�H;�H;�H;��H;��H;��H;��H;%�H;��H;z�H;��H;6�H;��H;��H;o�H;0�H;��H;�H;?�H;�H;��H;H�H;��H;��H;��H;��H;��H;t�H;d�H;e�H;��H;:�H;�H;j�H;(�H;r�H;      �H;7�H;ԻH;ۼH;�H;��H;��H;��H;��H;4�H;��H;�H;|�H;��H;B�H;_�H;[�H;�H;��H;D�H;��H;��H;��H;��H;@�H;��H;��H;��H;5�H;y�H;��H;��H;��H; �H;.�H;9�H;�H;9�H;.�H; �H;��H;��H;��H;y�H;5�H;��H;��H;��H;@�H;��H;��H;��H;��H;D�H;��H;�H;[�H;_�H;B�H;��H;|�H;�H;��H;4�H;��H;��H;��H;��H;�H;ۼH;ԻH;7�H;      ��H;��H;k�H;4�H;.�H;r�H;��H;��H;��H;��H;{�H;��H;��H;g�H;A�H;��H;��H;*�H;��H;��H;��H;��H;��H;H�H;��H;m�H;��H;�H;p�H;��H;��H;��H;�H;.�H;�H;-�H;J�H;-�H;�H;.�H;�H;��H;��H;��H;p�H;�H;��H;m�H;��H;H�H;��H;��H;��H;��H;��H;*�H;��H;��H;A�H;g�H;��H;��H;{�H;��H;��H;��H;��H;r�H;.�H;4�H;k�H;��H;      (�H;S�H;��H;O�H;D�H;u�H;��H;K�H;��H;��H;A�H;�H;��H;_�H;��H;��H;��H;E�H;|�H;��H;��H;P�H;�H;��H;C�H;��H;�H;^�H;��H;��H;��H;�H;�H;9�H;-�H;$�H;6�H;$�H;-�H;9�H;�H;�H;��H;��H;��H;^�H;�H;��H;C�H;��H;�H;P�H;��H;��H;|�H;E�H;��H;��H;��H;_�H;��H;�H;A�H;��H;��H;K�H;��H;u�H;D�H;O�H;��H;S�H;      ��H;��H;B�H;��H;��H;��H;��H;f�H;��H;n�H;.�H;��H;d�H;�H;��H;�H;s�H;��H;��H;��H;��H;��H;\�H;��H;L�H;��H;�H;g�H;��H;��H;��H;�H;�H;�H;J�H;6�H;#�H;6�H;J�H;�H;�H;�H;��H;��H;��H;g�H;�H;��H;L�H;��H;\�H;��H;��H;��H;��H;��H;s�H;�H;��H;�H;d�H;��H;.�H;n�H;��H;f�H;��H;��H;��H;��H;B�H;��H;      (�H;S�H;��H;O�H;D�H;u�H;��H;K�H;��H;��H;A�H;�H;��H;_�H;��H;��H;��H;E�H;|�H;��H;��H;P�H;�H;��H;C�H;��H;�H;^�H;��H;��H;��H;�H;�H;9�H;-�H;$�H;6�H;$�H;-�H;9�H;�H;�H;��H;��H;��H;^�H;�H;��H;C�H;��H;�H;P�H;��H;��H;|�H;E�H;��H;��H;��H;_�H;��H;�H;A�H;��H;��H;K�H;��H;u�H;D�H;O�H;��H;S�H;      ��H;��H;k�H;4�H;.�H;r�H;��H;��H;��H;��H;{�H;��H;��H;g�H;A�H;��H;��H;*�H;��H;��H;��H;��H;��H;H�H;��H;m�H;��H;�H;p�H;��H;��H;��H;�H;.�H;�H;-�H;J�H;-�H;�H;.�H;�H;��H;��H;��H;p�H;�H;��H;m�H;��H;H�H;��H;��H;��H;��H;��H;*�H;��H;��H;A�H;g�H;��H;��H;{�H;��H;��H;��H;��H;r�H;.�H;4�H;k�H;��H;      �H;7�H;ԻH;ۼH;�H;��H;��H;��H;��H;4�H;��H;�H;|�H;��H;B�H;_�H;[�H;�H;��H;D�H;��H;��H;��H;��H;@�H;��H;��H;��H;5�H;y�H;��H;��H;��H; �H;.�H;9�H;�H;9�H;.�H; �H;��H;��H;��H;y�H;5�H;��H;��H;��H;@�H;��H;��H;��H;��H;D�H;��H;�H;[�H;_�H;B�H;��H;|�H;�H;��H;4�H;��H;��H;��H;��H;�H;ۼH;ԻH;7�H;      8�H;r�H;(�H;j�H;�H;:�H;��H;e�H;d�H;t�H;��H;��H;��H;��H;��H;H�H;��H;�H;?�H;�H;��H;0�H;o�H;��H;��H;6�H;��H;z�H;��H;%�H;��H;��H;��H;��H;�H;�H;�H;�H;�H;��H;��H;��H;��H;%�H;��H;z�H;��H;6�H;��H;��H;o�H;0�H;��H;�H;?�H;�H;��H;H�H;��H;��H;��H;��H;��H;t�H;d�H;e�H;��H;:�H;�H;j�H;(�H;r�H;      v�H;�H;ߟH;}�H;ɣH;��H;©H;[�H;8�H;E�H;l�H;��H;��H;��H;6�H;��H;��H;�H;��H;�H;A�H;�H;��H; �H;f�H;S�H;�H;��H;k�H;��H;.�H;z�H;��H;��H;��H;�H;�H;�H;��H;��H;��H;z�H;.�H;��H;k�H;��H;�H;S�H;f�H; �H;��H;�H;A�H;�H;��H;�H;��H;��H;6�H;��H;��H;��H;l�H;E�H;8�H;[�H;©H;��H;ɣH;}�H;ߟH;�H;      Z�H;�H;\�H;��H;��H;v�H;ǖH;��H;��H;�H;��H;�H;�H;ȻH;��H;Z�H;��H;^�H;��H;$�H;��H;^�H;u�H;O�H;��H;�H;7�H;�H;��H;t�H;��H;.�H;��H;��H;��H;��H;��H;��H;��H;��H;��H;.�H;��H;t�H;��H;�H;7�H;�H;��H;O�H;u�H;^�H;��H;$�H;��H;^�H;��H;Z�H;��H;ȻH;�H;�H;��H;�H;��H;��H;ǖH;v�H;��H;��H;\�H;�H;      �gH;�hH;jH;�mH;�qH;�vH;�|H;x�H;��H;�H;Z�H;��H;֧H;��H;P�H;��H;>�H;I�H;��H;��H;��H;��H;��H;��H;��H;��H;��H;�H;��H;��H;t�H;��H;%�H;y�H;��H;��H;��H;��H;��H;y�H;%�H;��H;t�H;��H;��H;�H;��H;��H;��H;��H;��H;��H;��H;��H;��H;I�H;>�H;��H;P�H;��H;֧H;��H;Z�H;�H;��H;x�H;�|H;�vH;�qH;�mH;jH;�hH;      >H;�>H;UAH;�EH;EKH;DRH;sZH;\cH;�lH;�vH;��H;��H;��H;��H;��H;��H;<�H;�H;)�H;t�H;�H;2�H;��H;��H;c�H;��H;J�H;��H;$�H;��H;��H;k�H;��H;5�H;p�H;��H;��H;��H;p�H;5�H;��H;k�H;��H;��H;$�H;��H;J�H;��H;c�H;��H;��H;2�H;�H;t�H;)�H;�H;<�H;��H;��H;��H;��H;��H;��H;�vH;�lH;\cH;sZH;DRH;EKH;�EH;UAH;�>H;      ��G;+H;�H;�H;�H;s H;9,H;�8H;�EH;kSH;aH;`nH;m{H;�H;��H;~�H;:�H;	�H;�H;�H;O�H;��H; �H;��H;^�H;�H;h�H;]�H;��H;�H;�H;��H;z�H;��H;�H;^�H;g�H;^�H;�H;��H;z�H;��H;�H;�H;��H;]�H;h�H;�H;^�H;��H; �H;��H;O�H;�H;�H;	�H;:�H;~�H;��H;�H;m{H;`nH;aH;kSH;�EH;�8H;9,H;s H;�H;�H;�H;+H;      �G;\�G;�G;�G;P�G;2�G;��G;��G;�H;�#H;A7H;wIH;�ZH;lkH;{H;p�H;m�H;�H;r�H;��H;��H;��H;L�H;6�H;��H;$�H;�H;h�H;J�H;��H;7�H;�H;��H;��H;��H;�H;�H;�H;��H;��H;��H;�H;7�H;��H;J�H;h�H;�H;$�H;��H;6�H;L�H;��H;��H;��H;r�H;�H;m�H;p�H;{H;lkH;�ZH;wIH;A7H;�#H;�H;��G;��G;2�G;P�G;�G;�G;\�G;      �vF;�~F;ՕF;�F;:�F;�G;�MG;I�G;|�G;
�G;��G;iH;�0H;GH;�[H;�nH;�H;7�H;��H;v�H;��H;��H;V�H;��H;��H;W�H;$�H;�H;��H;��H;�H;S�H;6�H;��H;m�H;��H;��H;��H;m�H;��H;6�H;S�H;�H;��H;��H;�H;$�H;W�H;��H;��H;V�H;��H;��H;v�H;��H;7�H;�H;�nH;�[H;GH;�0H;iH;��G;
�G;|�G;I�G;�MG;�G;:�F;�F;ՕF;�~F;      ��C;qD;�AD;2�D;	E;��E;� F;�vF;!�F;)<G;+�G;�G;��G;"H;�3H;�LH;*cH;5wH;�H;c�H;��H;ΰH;�H;��H;=�H;��H;��H;^�H;c�H;��H;��H;f�H;��H;@�H;��H;C�H;L�H;C�H;��H;@�H;��H;f�H;��H;��H;c�H;^�H;��H;��H;=�H;��H;�H;ΰH;��H;c�H;�H;5wH;*cH;�LH;�3H;"H;��G;�G;+�G;)<G;!�F;�vF;� F;��E;	E;2�D;�AD;qD;      n+>;�Y>;-�>;�?;��@;-�A;�C;)D;�E;��E;�F;G;}G;u�G; �G;� H;k?H;�YH;UpH;C�H;O�H;��H;ɯH;�H;��H;��H;6�H;��H;��H;��H;O�H; �H;��H;��H;H�H;��H;��H;��H;H�H;��H;��H; �H;O�H;��H;��H;��H;6�H;��H;��H;�H;ɯH;��H;O�H;C�H;UpH;�YH;k?H;� H; �G;u�G;}G;G;�F;��E;�E;)D;�C;-�A;��@;�?;-�>;�Y>;      ��1;�I2;�f3;�#5;�X7;5�9;�f<;s�>;1A;�C;S�D;N�E;��F;O)G;a�G;d�G;�H;�4H;RH;qkH;.�H;��H;�H;ɯH;�H;V�H;L�H; �H;��H;��H;u�H;��H;o�H;��H;��H;�H;\�H;�H;��H;��H;o�H;��H;u�H;��H;��H; �H;L�H;V�H;�H;ɯH;�H;��H;.�H;qkH;RH;�4H;�H;d�G;a�G;O)G;��F;N�E;S�D;�C;1A;s�>;�f<;5�9;�X7;�#5;�f3;�I2;      2;%�;n
;!z ; �$;��);�
/;o4;T�8;��<;G#@;��B;d�D;��E;J�F;�bG;��G;�H;�,H;�MH;�hH;B�H;��H;��H;ΰH;��H;��H;��H;2�H;��H;^�H;�H;0�H;��H;��H;P�H;��H;P�H;��H;��H;0�H;�H;^�H;��H;2�H;��H;��H;��H;ΰH;��H;��H;B�H;�hH;�MH;�,H;�H;��G;�bG;J�F;��E;d�D;��B;G#@;��<;T�8;o4;�
/;��); �$;!z ;n
;%�;      f�:���:��:`��:2;�X;';��;��(;�0;/Y7;��<;G�@;-`C;QBE;�vF;�7G;��G;r�G;�(H;�KH;�hH;.�H;O�H;��H;��H;��H;O�H;�H;��H;��H;A�H;��H;��H;��H;��H;��H;��H;��H;��H;��H;A�H;��H;��H;�H;O�H;��H;��H;��H;O�H;.�H;�hH;�KH;�(H;r�G;��G;�7G;�vF;QBE;-`C;G�@;��<;/Y7;�0;��(;��;';�X;2;`��:��:���:      R�:ϟ:�1<:2(i:�s�:��:v~�:�*�:	Y;��;�)';�1;}�8;�Y>;/B;?�D;�1F;>G;��G;%�G;�(H;�MH;qkH;C�H;c�H;v�H;��H;�H;t�H;��H;$�H;�H;�H;D�H;��H;��H;��H;��H;��H;D�H;�H;�H;$�H;��H;t�H;�H;��H;v�H;c�H;C�H;qkH;�MH;�(H;%�G;��G;>G;�1F;?�D;/B;�Y>;}�8;�1;�)';��;	Y;�*�:v~�:��:�s�:2(i:�1<:ϟ:      a���sX��R!��p�=�ݷ�դ8<�:�O�:�O�:���:�_;�
;��*;=$5;�f<;9<A;4BD;/F;�G;��G;r�G;�,H;RH;UpH;�H;��H;r�H;�H;)�H;��H;��H;��H;?�H;��H;��H;|�H;��H;|�H;��H;��H;?�H;��H;��H;��H;)�H;�H;r�H;��H;�H;UpH;RH;�,H;r�G;��G;�G;/F;4BD;9<A;�f<;=$5;��*;�
;�_;���:�O�:�O�:<�:դ8ݷ�p�=�R!��sX��      �1��(Ȅ�Ѩu��PV��.�����W��w��U�9�)i:�:�*�:��;�s%;1J2;�;;�@;�D;/F;>G;��G;�H;�4H;�YH;5wH;7�H;�H;	�H;�H;I�H;^�H;�H;�H;�H;*�H;E�H;��H;E�H;*�H;�H;�H;�H;^�H;I�H;�H;	�H;�H;7�H;5wH;�YH;�4H;�H;��G;>G;/F;�D;�@;�;;1J2;�s%;��;�*�:�:�)i:�U�9w���W������.��PV�Ѩu�(Ȅ�      E��8�	����ǘ�Tʻ�R��3|�x.�iȺ����V�9^t�:��:;Y;��!;�0;-�:;�@;4BD;�1F;�7G;��G;�H;k?H;*cH;�H;m�H;:�H;<�H;>�H;��H;��H;��H;[�H;��H;��H;s�H;��H;��H;[�H;��H;��H;��H;>�H;<�H;:�H;m�H;�H;*cH;k?H;�H;��G;�7G;�1F;4BD;�@;-�:;�0;��!;;Y;��:^t�:�V�9���iȺx.�3|��R��Tʻǘ����8�	�      ��x��[t���g�,T�?�:������������1��b�(��W��6�t�xm`:v��:_\;pz ;�0;�;;9<A;?�D;�vF;�bG;d�G;� H;�LH;�nH;p�H;~�H;��H;��H;Z�H;��H;H�H;_�H;��H;��H;�H;��H;��H;_�H;H�H;��H;Z�H;��H;��H;~�H;p�H;�nH;�LH;� H;d�G;�bG;�vF;?�D;9<A;�;;�0;pz ;_\;v��:xm`:6�t��W��b�(��1������������?�:�,T���g��[t�      ,˼x�Ǽ�"��x뮼�v��G���[�Ey-�����.��͕b��0㺈ڷ��3<:L�:_\;��!;1J2;�f<;/B;QBE;J�F;a�G; �G;�3H;�[H;{H;��H;��H;P�H;��H;6�H;��H;B�H;A�H;��H;��H;��H;A�H;B�H;��H;6�H;��H;P�H;��H;��H;{H;�[H;�3H; �G;a�G;J�F;QBE;/B;�f<;1J2;��!;_\;L�:�3<:�ڷ��0�͕b��.�����Ey-��[�G���v��x뮼�"��x�Ǽ      ���k���1v�Rt��Ѽt뮼X��H�W������׻�Ǆ�0�����3<:v��:;Y;�s%;=$5;�Y>;-`C;��E;O)G;u�G;"H;GH;lkH;�H;��H;��H;ȻH;��H;��H;��H;g�H;_�H;�H;_�H;g�H;��H;��H;��H;ȻH;��H;��H;�H;lkH;GH;"H;u�G;O)G;��E;-`C;�Y>;=$5;�s%;;Y;v��:�3<:���0���Ǆ���׻���H�W�X��t뮼�ѼRt�1v����k�      m��Fi��&^�;�L�/�6������|ռPT��z�x���0��������0���ڷ�xm`:��:��;��*;}�8;G�@;d�D;��F;}G;��G;�0H;�ZH;m{H;��H;֧H;�H;��H;��H;|�H;��H;��H;d�H;��H;��H;|�H;��H;��H;�H;֧H;��H;m{H;�ZH;�0H;��G;}G;��F;d�D;G�@;}�8;��*;��;��:xm`:�ڷ�0��������껣�0�z�x�PT���|ռ����/�6�;�L��&^��Fi�      0��W;��&������n섽Q�e���?��k�Ot��跼G��ee7�����Ǆ��0�6�t�^t�:�*�:�
;�1;��<;��B;N�E;G;�G;iH;wIH;`nH;��H;��H;�H;��H;��H;�H;��H;�H;��H;�H;��H;�H;��H;��H;�H;��H;��H;`nH;wIH;iH;�G;G;N�E;��B;��<;�1;�
;�*�:^t�:6�t��0��Ǆ����ee7�G���跼Ot�k���?�Q�e�n섽���&���W;��      J��� ��s��ӽ~'��%�������Z�kQ+�����"��G����0���׻͕b��W���V�9�:�_;�)';/Y7;G#@;S�D;�F;+�G;��G;A7H;aH;��H;Z�H;��H;l�H;��H;��H;{�H;A�H;.�H;A�H;{�H;��H;��H;l�H;��H;Z�H;��H;aH;A7H;��G;+�G;�F;S�D;G#@;/Y7;�)';�_;�:�V�9�W��͕b���׻��0�G���"�����kQ+��Z����%���~'���ӽ�s� ��      �!,� )��K ����x��ͻ޽ ������Fi���0�����跼z�x�����.��b�(�����)i:���:��;�0;��<;�C;��E;)<G;
�G;�#H;kSH;�vH;�H;�H;E�H;t�H;4�H;��H;��H;n�H;��H;��H;4�H;t�H;E�H;�H;�H;�vH;kSH;�#H;
�G;)<G;��E;�C;��<;�0;��;���:�)i:���b�(��.�����z�x��跼�����0��Fi���� ��ͻ޽x������K � )�      	�j�ȟf��Z�]�F��>/��^�H�����Ž- ���Fi�kQ+�Ot�PT��H�W�����1��iȺ�U�9�O�:	Y;��(;T�8;1A;�E;!�F;|�G;�H;�EH;�lH;��H;��H;8�H;d�H;��H;��H;��H;��H;��H;��H;��H;d�H;8�H;��H;��H;�lH;�EH;�H;|�G;!�F;�E;1A;T�8;��(;	Y;�O�:�U�9iȺ�1�����H�W�PT��Ot�kQ+��Fi�- ����ŽH����^��>/�]�F��Z�ȟf�      ��b���f�6���ȟf�rSC��K �Gn����Ž����Z��k��|ռX��Ey-����x.�w���O�:�*�:��;o4;s�>;)D;�vF;I�G;��G;�8H;\cH;x�H;��H;[�H;e�H;��H;��H;K�H;f�H;K�H;��H;��H;e�H;[�H;��H;x�H;\cH;�8H;��G;I�G;�vF;)D;s�>;o4;��;�*�:�O�:w��x.����Ey-�X���|ռ�k��Z������ŽGn���K �rSC�ȟf�6���f�b���      {�˾��Ǿi���
���C͓�9�x�ؘJ��K �H��� �������?���t뮼�[�����3|��W��<�:v~�:';�
/;�f<;�C;� F;�MG;��G;9,H;sZH;�|H;ǖH;©H;��H;��H;��H;��H;��H;��H;��H;��H;��H;©H;ǖH;�|H;sZH;9,H;��G;�MG;� F;�C;�f<;�
/;';v~�:<�:�W��3|������[�t뮼����?���� ��H����K �ؘJ�9�x�C͓�
���i�����Ǿ      e� ������쾻{ԾS���b���9�x�rSC��^�ͻ޽%���Q�e����ѼG������R�����դ8��:�X;��);5�9;-�A;��E;�G;2�G;s H;DRH;�vH;v�H;��H;:�H;��H;r�H;u�H;��H;u�H;r�H;��H;:�H;��H;v�H;�vH;DRH;s H;2�G;�G;��E;-�A;5�9;��);�X;��:դ8����R�����G���Ѽ��Q�e�%���ͻ޽�^�rSC�9�x�b���S����{Ծ�쾃���      ����D��k�e� �<�ݾS���C͓�ȟf��>/�x��~'��n섽/�6�Rt��v��?�:�Tʻ�.�ݷ��s�:2; �$;�X7;��@;	E;:�F;P�G;�H;EKH;�qH;��H;ɣH;�H;�H;.�H;D�H;��H;D�H;.�H;�H;�H;ɣH;��H;�qH;EKH;�H;P�G;:�F;	E;��@;�X7; �$;2;�s�:ݷ��.�Tʻ?�:��v��Rt�/�6�n섽~'��x���>/�ȟf�C͓�S���<�ݾe� ��k��D�      ߛ7�v3��'����e� ��{Ծ
���6���]�F�����ӽ���;�L�1v�x뮼,T�ǘ��PV�p�=�2(i:`��:!z ;�#5;�?;2�D;�F;�G;�H;�EH;�mH;��H;}�H;j�H;ۼH;4�H;O�H;��H;O�H;4�H;ۼH;j�H;}�H;��H;�mH;�EH;�H;�G;�F;2�D;�?;�#5;!z ;`��:2(i:p�=��PV�ǘ�,T�x뮼1v�;�L�����ӽ���]�F�6���
����{Ծe� �����'�v3�      tN��TI���;��'��k���i���f󐾖Z��K ��s�&����&^����"����g����Ѩu�R!���1<:��:n
;�f3;-�>;�AD;ՕF;�G;�H;UAH;jH;\�H;ߟH;(�H;ԻH;k�H;��H;B�H;��H;k�H;ԻH;(�H;ߟH;\�H;jH;UAH;�H;�G;ՕF;�AD;-�>;�f3;n
;��:�1<:R!��Ѩu������g��"�����&^�&����s潎K ��Z�f�i������k��'���;��TI�      I]�N�W��TI�v3��D�������Ǿb���ȟf� )� ��W;���Fi��k�x�Ǽ�[t�8�	�(Ȅ�sX��ϟ:���:%�;�I2;�Y>;qD;�~F;\�G;+H;�>H;�hH;�H;�H;r�H;7�H;��H;S�H;��H;S�H;��H;7�H;r�H;�H;�H;�hH;�>H;+H;\�G;�~F;qD;�Y>;�I2;%�;���:ϟ:sX��(Ȅ�8�	��[t�x�Ǽ�k��Fi�W;�� �� )�ȟf�b�����Ǿ�����D�v3��TI�N�W�      �?��ph��1v��� ��$�X��O/�#y�-�;Ѱ��j+X�����ѽ����Gn;�>�＿����B(�暩����%�e9��:^;Y.;��<;�VC;?ZF;�G;5/H;tiH;X�H;s�H;��H;E�H;��H;�H;��H;��H;��H;�H;��H;E�H;��H;s�H;X�H;tiH;5/H;�G;?ZF;�VC;��<;Y.;^;��:%�e9���暩��B(�����>��Gn;�������ѽ��j+X�Ѱ��-�;#y��O/�$�X�� ��1v��ph��      ph��"���V�����y�EvS�aM+��v� 9ɾ�����T�]��[ν����`\8�����x���%�\��������9B,�:��;�.;M�<; nC;�cF;�G;�0H;!jH;ǋH;ѣH;��H;��H;��H;��H;��H;��H;��H;��H;��H;��H;��H;ѣH;ǋH;!jH;�0H;�G;�cF; nC;M�<;�.;��;B,�:��9���\����%��x�����`\8������[ν]��T����� 9ɾ�v�aM+�EvS���y�V���"���      1v��V���L ��M�h�%E�I��R���i㼾n���nH�È�a�ý�Ȅ��s/��o༼#�����4J���к��9#f�:Ml;�0;P\=; �C;5�F;��G;Q5H;^lH;H�H;ϤH;��H;�H;b�H;��H;#�H; �H;#�H;��H;b�H;�H;��H;ϤH;H�H;^lH;Q5H;��G;5�F; �C;P\=;�0;Ml;#f�:��9�к4J������#���o��s/��Ȅ�a�ýÈ��nH�n��i㼾R���I��%E�M�h�L ��V���      � ����y�M�h�ބN��O/����-�߾�A���*|�ؕ6�a}��㳽KSt�(�!�Wrμ(F{��_�Y��h����:���:VZ;2;�N>;�D;��F;��G;J<H;�oH;��H;t�H;��H;��H;��H;��H;��H;�H;��H;��H;��H;��H;��H;t�H;��H;�oH;J<H;��G;��F;�D;�N>;2;VZ;���:�:h���Y���_�(F{�Wrμ(�!�KSt��㳽a}�ؕ6��*|��A��-�߾����O/�ބN�M�h���y�      $�X�EvS�%E��O/��S�1W����������4S\�� �q�&�����Y�h��������]�}���T�b��Y���Y:~�:�_;��4;�?;|�D;�F;/�G;5EH;tH;�H;��H;��H;3�H;��H;E�H;7�H;�H;7�H;E�H;��H;3�H;��H;��H;�H;tH;5EH;/�G;�F;|�D;�?;��4;�_;~�:��Y:�Y�T�b�}�����]�����h����Y�&���q�� �4S\���������1W���S��O/�%E�EvS�      �O/�aM+�I�����1W�� 9ɾ0���Mw�� :�Y��_�ý�L��Dn;�>���bv���E<��˻)�-����x�:^;%;�7;��@;V4E;�!G;,�G;hOH;1zH;��H;��H;��H;��H;�H;2�H;�H;��H;�H;2�H;�H;��H;��H;��H;��H;1zH;hOH;,�G;�!G;V4E;��@;�7;%;^;�x�:��)�-��˻�E<�bv��>���Dn;��L��_�ýY��� :��Mw�0�� 9ɾ1W�����I��aM+�      #y��v�R���-�߾����0��1����nH���(Ὁu��r�d�O�Prμ="�����	��3���k89v:�:��;+;�{:;�6B;)�E;EaG;�H;ZH;��H;M�H;ĮH;�H;e�H;e�H;*�H;��H;��H;��H;*�H;e�H;e�H;�H;ĮH;M�H;��H;ZH;�H;EaG;)�E;�6B;�{:;+;��;v:�:�k893��	�����="��PrμO�r�d��u��(����nH�1���0������-�߾R����v�      -�; 9ɾi㼾�A�������Mw��nH�����Z��㳽����Z\8�P#�������]N�J��.�b�YJx�w5:��:��;8�0;v\=;u�C;�ZF;�G;)H;eH;��H;F�H;g�H;��H;7�H;��H;P�H;��H;��H;��H;P�H;��H;7�H;��H;g�H;F�H;��H;eH;)H;�G;�ZF;u�C;v\=;8�0;��;��:w5:YJx�.�b�J���]N�����P#��Z\8������㳽�Z񽞯��nH��Mw������A��i㼾 9ɾ      Ѱ������n���*|�4S\�� :����Z�U$������K�c���Oļ����������x&�-��O.�:0^;��#;G6;��?;-�D;��F;��G;)?H;�oH;�H;��H;:�H;q�H;J�H;��H;��H;��H;��H;��H;��H;��H;J�H;q�H;:�H;��H;�H;�oH;)?H;��G;��F;-�D;��?;G6;��#;0^;O.�:-��x&������������Oļc���K����U$���Z���� :�4S\��*|�n������      j+X��T��nH�ؕ6�� �Y��(��㳽����mR����ټ�����E<��?ݻbd\�c ��#:�c�:8�;y�,;��:;�6B;ͱE;�KG;iH;�RH;�zH;��H;
�H;9�H;`�H;n�H;+�H;��H;�H;��H;�H;��H;+�H;n�H;`�H;9�H;
�H;��H;�zH;�RH;iH;�KG;ͱE;�6B;��:;y�,;8�;�c�:#:c ��bd\��?ݻ�E<������ټ���mR�����㳽(�Y��� �ؕ6��nH��T�      ��]�È�a}�q�_�ý�u�������K����o�Wv���&R���f^����@���:�A;�";��4;��>;�D;��F;,�G; )H;�cH;��H;5�H;��H;N�H;M�H;��H;��H;<�H;(�H;��H;(�H;<�H;��H;��H;M�H;N�H;��H;5�H;��H;�cH; )H;,�G;��F;�D;��>;��4;�";�A;��:@���f^�����&R�Wv���o����K������u��_�ýq�a}�È�]�      ��ѽ�[νa�ý�㳽&����L��r�d�Z\8�c���ټWv����Y��_����z��]���Y:?��:�l;r-;Q�:;��A;rnE;�!G;��G;�FH;�rH;�H;��H;�H;J�H;5�H;��H;��H;��H;B�H;�H;B�H;��H;��H;��H;5�H;J�H;�H;��H;�H;�rH;�FH;��G;�!G;rnE;��A;Q�:;r-;�l;?��:��Y:]�z������_���Y�Wv���ټc��Z\8�r�d��L��&����㳽a�ý�[ν      ���������Ȅ�KSt���Y�Dn;�O�P#���Oļ�����&R��_������N3�.�Y�-2:�:9�;@?&;(G6;�W?;�D;fwF;�G;c H;�]H;��H;�H;�H;a�H;#�H;�H;��H;(�H;��H;i�H;%�H;i�H;��H;(�H;��H;�H;#�H;a�H;�H;�H;��H;�]H;c H;�G;fwF;�D;�W?;(G6;@?&;9�;�:-2:.�Y��N3������_��&R������OļP#��O�Dn;���Y�KSt��Ȅ�����      Gn;�`\8��s/�(�!�h��>���Prμ��������E<�������N3��Ix�a�9��:T^;� ;~2;��<;.�B;�E;e4G;1�G;^EH;�pH;��H;h�H;ϳH;k�H;��H;��H;�H;��H;1�H;��H;�H;��H;1�H;��H;�H;��H;��H;k�H;ϳH;h�H;��H;�pH;^EH;1�G;e4G;�E;.�B;��<;~2;� ;T^;��:a�9�Ix��N3�������E<��������Prμ>���h��(�!��s/�`\8�      >�Ｘ���o�Wrμ����bv��="���]N�����?ݻf^��z��.�Y�a�9��:���:B�;��.;�{:;2>A;��D;`�F;ߵG;
)H;D`H;5�H;��H;�H;R�H;6�H;R�H;t�H;�H;.�H;k�H;��H;��H;��H;k�H;.�H;�H;t�H;R�H;6�H;R�H;�H;��H;5�H;D`H;
)H;ߵG;`�F;��D;2>A;�{:;��.;B�;���:��:a�9.�Y�z��f^���?ݻ����]N�="��bv������Wrμ�o༸��      �����x���#��(F{���]��E<����J�뻲���bd\���]�-2:��:���:�Z;��,;/�8;` @;0D;�ZF;PzG;
H;iOH;=uH;�H;[�H;�H;C�H;z�H;��H;��H;��H;��H;��H;��H;��H;��H;��H;��H;��H;��H;��H;z�H;C�H;�H;[�H;�H;=uH;iOH;
H;PzG;�ZF;0D;` @;/�8;��,;�Z;���:��:-2:]���bd\�����J�뻛���E<���]�(F{��#���x��      �B(��%�����_�}����˻	��.�b�x&�c ��@���Y:�:T^;B�;��,;Z_8;��?;��C;�F;FG;t�G;?H;FjH;#�H; �H;
�H;k�H;��H;~�H;��H;/�H;��H;��H;��H;��H;��H;��H;��H;��H;��H;/�H;��H;~�H;��H;k�H;
�H; �H;#�H;FjH;?H;t�G;FG;�F;��C;��?;Z_8;��,;B�;T^;�:��Y:@�c ��x&�.�b�	���˻}����_�����%�      暩�\���4J��Y��T�b�)�-�3��YJx�-��#:��:?��:9�;� ;��.;/�8;��?;2�C;�E;f"G;�G;1H;aH;gH;��H;��H;��H;��H;s�H;(�H;I�H;J�H;��H;(�H;��H;G�H;��H;G�H;��H;(�H;��H;J�H;I�H;(�H;s�H;��H;��H;��H;��H;gH;aH;1H;�G;f"G;�E;2�C;��?;/�8;��.;� ;9�;?��:��:#:-��YJx�3��)�-�T�b�Y��4J��\���      �����뺸кh����Y����k89w5:O.�:�c�:�A;�l;@?&;~2;�{:;` @;��C;�E;�G;�G;}'H;ZH;�yH;W�H;��H;��H;{�H;��H;��H;l�H;��H;
�H;[�H;<�H;W�H;
�H;��H;
�H;W�H;<�H;[�H;
�H;��H;l�H;��H;��H;{�H;��H;��H;W�H;�yH;ZH;}'H;�G;�G;�E;��C;` @;�{:;~2;@?&;�l;�A;�c�:O.�:w5:�k89���Y�h����к���      %�e9��9��9�:��Y:�x�:v:�:��:0^;8�;�";r-;(G6;��<;2>A;0D;�F;f"G;�G;$H;VH;�uH;��H;Y�H;b�H;��H;!�H;��H;��H;E�H;��H;��H;��H;6�H;�H;��H;�H;��H;�H;6�H;��H;��H;��H;E�H;��H;��H;!�H;��H;b�H;Y�H;��H;�uH;VH;$H;�G;f"G;�F;0D;2>A;��<;(G6;r-;�";8�;0^;��:v:�:�x�:��Y:�:��9��9      ��:B,�:#f�:���:~�:^;��;��;��#;y�,;��4;Q�:;�W?;.�B;��D;�ZF;FG;�G;}'H;VH;�tH;��H;.�H;�H;<�H;	�H;��H;��H;��H;��H;��H;��H;��H;��H;��H;^�H;b�H;^�H;��H;��H;��H;��H;��H;��H;��H;��H;��H;	�H;<�H;�H;.�H;��H;�tH;VH;}'H;�G;FG;�ZF;��D;.�B;�W?;Q�:;��4;y�,;��#;��;��;^;~�:���:#f�:B,�:      ^;��;Ml;VZ;�_;%;+;8�0;G6;��:;��>;��A;�D;�E;`�F;PzG;t�G;1H;ZH;�uH;��H;g�H;ܫH;߷H;��H;e�H;��H;��H;��H;��H;H�H;G�H;��H;��H;p�H;��H;��H;��H;p�H;��H;��H;G�H;H�H;��H;��H;��H;��H;e�H;��H;߷H;ܫH;g�H;��H;�uH;ZH;1H;t�G;PzG;`�F;�E;�D;��A;��>;��:;G6;8�0;+;%;�_;VZ;Ml;��;      Y.;�.;�0;2;��4;�7;�{:;v\=;��?;�6B;�D;rnE;fwF;e4G;ߵG;
H;?H;aH;�yH;��H;.�H;ܫH;`�H;��H;�H;��H;��H;�H;)�H;��H;��H;h�H;c�H;O�H;��H;(�H;P�H;(�H;��H;O�H;c�H;h�H;��H;��H;)�H;�H;��H;��H;�H;��H;`�H;ܫH;.�H;��H;�yH;aH;?H;
H;ߵG;e4G;fwF;rnE;�D;�6B;��?;v\=;�{:;�7;��4;2;�0;�.;      ��<;M�<;P\=;�N>;�?;��@;�6B;u�C;-�D;ͱE;��F;�!G;�G;1�G;
)H;iOH;FjH;gH;W�H;Y�H;�H;߷H;��H;H�H;I�H;E�H;W�H;��H;,�H;B�H;�H;�H;�H;��H;H�H;��H;��H;��H;H�H;��H;�H;�H;�H;B�H;,�H;��H;W�H;E�H;I�H;H�H;��H;߷H;�H;Y�H;W�H;gH;FjH;iOH;
)H;1�G;�G;�!G;��F;ͱE;-�D;u�C;�6B;��@;�?;�N>;P\=;M�<;      �VC; nC; �C;�D;|�D;V4E;)�E;�ZF;��F;�KG;,�G;��G;c H;^EH;D`H;=uH;#�H;��H;��H;b�H;<�H;��H;�H;I�H;�H;�H;O�H;��H;��H;��H;��H;��H;��H;=�H;��H;��H;��H;��H;��H;=�H;��H;��H;��H;��H;��H;��H;O�H;�H;�H;I�H;�H;��H;<�H;b�H;��H;��H;#�H;=uH;D`H;^EH;c H;��G;,�G;�KG;��F;�ZF;)�E;V4E;|�D;�D; �C; nC;      ?ZF;�cF;5�F;��F;�F;�!G;EaG;�G;��G;iH; )H;�FH;�]H;�pH;5�H;�H; �H;��H;��H;��H;	�H;e�H;��H;E�H;�H;5�H;��H;��H;u�H;��H;��H;��H;,�H;~�H;��H;�H;�H;�H;��H;~�H;,�H;��H;��H;��H;u�H;��H;��H;5�H;�H;E�H;��H;e�H;	�H;��H;��H;��H; �H;�H;5�H;�pH;�]H;�FH; )H;iH;��G;�G;EaG;�!G;�F;��F;5�F;�cF;      �G;�G;��G;��G;/�G;,�G;�H;)H;)?H;�RH;�cH;�rH;��H;��H;��H;[�H;
�H;��H;{�H;!�H;��H;��H;��H;W�H;O�H;��H;��H;J�H;��H;��H;j�H; �H;}�H;��H;�H;;�H;Y�H;;�H;�H;��H;}�H; �H;j�H;��H;��H;J�H;��H;��H;O�H;W�H;��H;��H;��H;!�H;{�H;��H;
�H;[�H;��H;��H;��H;�rH;�cH;�RH;)?H;)H;�H;,�G;/�G;��G;��G;�G;      5/H;�0H;Q5H;J<H;5EH;hOH;ZH;eH;�oH;�zH;��H;�H;�H;h�H;�H;�H;k�H;��H;��H;��H;��H;��H;�H;��H;��H;��H;J�H;��H;e�H;S�H;�H;i�H;��H;�H;E�H;[�H;M�H;[�H;E�H;�H;��H;i�H;�H;S�H;e�H;��H;J�H;��H;��H;��H;�H;��H;��H;��H;��H;��H;k�H;�H;�H;h�H;�H;�H;��H;�zH;�oH;eH;ZH;hOH;5EH;J<H;Q5H;�0H;      tiH;!jH;^lH;�oH;tH;1zH;��H;��H;�H;��H;5�H;��H;�H;ϳH;R�H;C�H;��H;s�H;��H;��H;��H;��H;)�H;,�H;��H;u�H;��H;e�H;[�H;��H;Y�H;��H;��H;5�H;e�H;o�H;b�H;o�H;e�H;5�H;��H;��H;Y�H;��H;[�H;e�H;��H;u�H;��H;,�H;)�H;��H;��H;��H;��H;s�H;��H;C�H;R�H;ϳH;�H;��H;5�H;��H;�H;��H;��H;1zH;tH;�oH;^lH;!jH;      X�H;ǋH;H�H;��H;�H;��H;M�H;F�H;��H;
�H;��H;�H;a�H;k�H;6�H;z�H;~�H;(�H;l�H;E�H;��H;��H;��H;B�H;��H;��H;��H;S�H;��H;K�H;��H;��H;6�H;]�H;h�H;��H;��H;��H;h�H;]�H;6�H;��H;��H;K�H;��H;S�H;��H;��H;��H;B�H;��H;��H;��H;E�H;l�H;(�H;~�H;z�H;6�H;k�H;a�H;�H;��H;
�H;��H;F�H;M�H;��H;�H;��H;H�H;ǋH;      s�H;ѣH;ϤH;t�H;��H;��H;ĮH;g�H;:�H;9�H;N�H;J�H;#�H;��H;R�H;��H;��H;I�H;��H;��H;��H;H�H;��H;�H;��H;��H;j�H;�H;Y�H;��H;��H;)�H;a�H;o�H;��H;��H;��H;��H;��H;o�H;a�H;)�H;��H;��H;Y�H;�H;j�H;��H;��H;�H;��H;H�H;��H;��H;��H;I�H;��H;��H;R�H;��H;#�H;J�H;N�H;9�H;:�H;g�H;ĮH;��H;��H;t�H;ϤH;ѣH;      ��H;��H;��H;��H;��H;��H;�H;��H;q�H;`�H;M�H;5�H;�H;��H;t�H;��H;/�H;J�H;
�H;��H;��H;G�H;h�H;�H;��H;��H; �H;i�H;��H;��H;)�H;A�H;k�H;��H;��H;��H;��H;��H;��H;��H;k�H;A�H;)�H;��H;��H;i�H; �H;��H;��H;�H;h�H;G�H;��H;��H;
�H;J�H;/�H;��H;t�H;��H;�H;5�H;M�H;`�H;q�H;��H;�H;��H;��H;��H;��H;��H;      E�H;��H;�H;��H;3�H;��H;e�H;7�H;J�H;n�H;��H;��H;��H;�H;�H;��H;��H;��H;[�H;��H;��H;��H;c�H;�H;��H;,�H;}�H;��H;��H;6�H;a�H;k�H;{�H;��H;��H;��H;��H;��H;��H;��H;{�H;k�H;a�H;6�H;��H;��H;}�H;,�H;��H;�H;c�H;��H;��H;��H;[�H;��H;��H;��H;�H;�H;��H;��H;��H;n�H;J�H;7�H;e�H;��H;3�H;��H;�H;��H;      ��H;��H;b�H;��H;��H;�H;e�H;��H;��H;+�H;��H;��H;(�H;��H;.�H;��H;��H;(�H;<�H;6�H;��H;��H;O�H;��H;=�H;~�H;��H;�H;5�H;]�H;o�H;��H;��H;��H;��H;��H;��H;��H;��H;��H;��H;��H;o�H;]�H;5�H;�H;��H;~�H;=�H;��H;O�H;��H;��H;6�H;<�H;(�H;��H;��H;.�H;��H;(�H;��H;��H;+�H;��H;��H;e�H;�H;��H;��H;b�H;��H;      �H;��H;��H;��H;E�H;2�H;*�H;P�H;��H;��H;<�H;��H;��H;1�H;k�H;��H;��H;��H;W�H;�H;��H;p�H;��H;H�H;��H;��H;�H;E�H;e�H;h�H;��H;��H;��H;��H;��H;��H;��H;��H;��H;��H;��H;��H;��H;h�H;e�H;E�H;�H;��H;��H;H�H;��H;p�H;��H;�H;W�H;��H;��H;��H;k�H;1�H;��H;��H;<�H;��H;��H;P�H;*�H;2�H;E�H;��H;��H;��H;      ��H;��H;#�H;��H;7�H;�H;��H;��H;��H;�H;(�H;B�H;i�H;��H;��H;��H;��H;G�H;
�H;��H;^�H;��H;(�H;��H;��H;�H;;�H;[�H;o�H;��H;��H;��H;��H;��H;��H;��H;��H;��H;��H;��H;��H;��H;��H;��H;o�H;[�H;;�H;�H;��H;��H;(�H;��H;^�H;��H;
�H;G�H;��H;��H;��H;��H;i�H;B�H;(�H;�H;��H;��H;��H;�H;7�H;��H;#�H;��H;      ��H;��H; �H;�H;�H;��H;��H;��H;��H;��H;��H;�H;%�H;�H;��H;��H;��H;��H;��H;�H;b�H;��H;P�H;��H;��H;�H;Y�H;M�H;b�H;��H;��H;��H;��H;��H;��H;��H;��H;��H;��H;��H;��H;��H;��H;��H;b�H;M�H;Y�H;�H;��H;��H;P�H;��H;b�H;�H;��H;��H;��H;��H;��H;�H;%�H;�H;��H;��H;��H;��H;��H;��H;�H;�H; �H;��H;      ��H;��H;#�H;��H;7�H;�H;��H;��H;��H;�H;(�H;B�H;i�H;��H;��H;��H;��H;G�H;
�H;��H;^�H;��H;(�H;��H;��H;�H;;�H;[�H;o�H;��H;��H;��H;��H;��H;��H;��H;��H;��H;��H;��H;��H;��H;��H;��H;o�H;[�H;;�H;�H;��H;��H;(�H;��H;^�H;��H;
�H;G�H;��H;��H;��H;��H;i�H;B�H;(�H;�H;��H;��H;��H;�H;7�H;��H;#�H;��H;      �H;��H;��H;��H;E�H;2�H;*�H;P�H;��H;��H;<�H;��H;��H;1�H;k�H;��H;��H;��H;W�H;�H;��H;p�H;��H;H�H;��H;��H;�H;E�H;e�H;h�H;��H;��H;��H;��H;��H;��H;��H;��H;��H;��H;��H;��H;��H;h�H;e�H;E�H;�H;��H;��H;H�H;��H;p�H;��H;�H;W�H;��H;��H;��H;k�H;1�H;��H;��H;<�H;��H;��H;P�H;*�H;2�H;E�H;��H;��H;��H;      ��H;��H;b�H;��H;��H;�H;e�H;��H;��H;+�H;��H;��H;(�H;��H;.�H;��H;��H;(�H;<�H;6�H;��H;��H;O�H;��H;=�H;~�H;��H;�H;5�H;]�H;o�H;��H;��H;��H;��H;��H;��H;��H;��H;��H;��H;��H;o�H;]�H;5�H;�H;��H;~�H;=�H;��H;O�H;��H;��H;6�H;<�H;(�H;��H;��H;.�H;��H;(�H;��H;��H;+�H;��H;��H;e�H;�H;��H;��H;b�H;��H;      E�H;��H;�H;��H;3�H;��H;e�H;7�H;J�H;n�H;��H;��H;��H;�H;�H;��H;��H;��H;[�H;��H;��H;��H;c�H;�H;��H;,�H;}�H;��H;��H;6�H;a�H;k�H;{�H;��H;��H;��H;��H;��H;��H;��H;{�H;k�H;a�H;6�H;��H;��H;}�H;,�H;��H;�H;c�H;��H;��H;��H;[�H;��H;��H;��H;�H;�H;��H;��H;��H;n�H;J�H;7�H;e�H;��H;3�H;��H;�H;��H;      ��H;��H;��H;��H;��H;��H;�H;��H;q�H;`�H;M�H;5�H;�H;��H;t�H;��H;/�H;J�H;
�H;��H;��H;G�H;h�H;�H;��H;��H; �H;i�H;��H;��H;)�H;A�H;k�H;��H;��H;��H;��H;��H;��H;��H;k�H;A�H;)�H;��H;��H;i�H; �H;��H;��H;�H;h�H;G�H;��H;��H;
�H;J�H;/�H;��H;t�H;��H;�H;5�H;M�H;`�H;q�H;��H;�H;��H;��H;��H;��H;��H;      s�H;ѣH;ϤH;t�H;��H;��H;ĮH;g�H;:�H;9�H;N�H;J�H;#�H;��H;R�H;��H;��H;I�H;��H;��H;��H;H�H;��H;�H;��H;��H;j�H;�H;Y�H;��H;��H;)�H;a�H;o�H;��H;��H;��H;��H;��H;o�H;a�H;)�H;��H;��H;Y�H;�H;j�H;��H;��H;�H;��H;H�H;��H;��H;��H;I�H;��H;��H;R�H;��H;#�H;J�H;N�H;9�H;:�H;g�H;ĮH;��H;��H;t�H;ϤH;ѣH;      X�H;ǋH;H�H;��H;�H;��H;M�H;F�H;��H;
�H;��H;�H;a�H;k�H;6�H;z�H;~�H;(�H;l�H;E�H;��H;��H;��H;B�H;��H;��H;��H;S�H;��H;K�H;��H;��H;6�H;]�H;h�H;��H;��H;��H;h�H;]�H;6�H;��H;��H;K�H;��H;S�H;��H;��H;��H;B�H;��H;��H;��H;E�H;l�H;(�H;~�H;z�H;6�H;k�H;a�H;�H;��H;
�H;��H;F�H;M�H;��H;�H;��H;H�H;ǋH;      tiH;!jH;^lH;�oH;tH;1zH;��H;��H;�H;��H;5�H;��H;�H;ϳH;R�H;C�H;��H;s�H;��H;��H;��H;��H;)�H;,�H;��H;u�H;��H;e�H;[�H;��H;Y�H;��H;��H;5�H;e�H;o�H;b�H;o�H;e�H;5�H;��H;��H;Y�H;��H;[�H;e�H;��H;u�H;��H;,�H;)�H;��H;��H;��H;��H;s�H;��H;C�H;R�H;ϳH;�H;��H;5�H;��H;�H;��H;��H;1zH;tH;�oH;^lH;!jH;      5/H;�0H;Q5H;J<H;5EH;hOH;ZH;eH;�oH;�zH;��H;�H;�H;h�H;�H;�H;k�H;��H;��H;��H;��H;��H;�H;��H;��H;��H;J�H;��H;e�H;S�H;�H;i�H;��H;�H;E�H;[�H;M�H;[�H;E�H;�H;��H;i�H;�H;S�H;e�H;��H;J�H;��H;��H;��H;�H;��H;��H;��H;��H;��H;k�H;�H;�H;h�H;�H;�H;��H;�zH;�oH;eH;ZH;hOH;5EH;J<H;Q5H;�0H;      �G;�G;��G;��G;/�G;,�G;�H;)H;)?H;�RH;�cH;�rH;��H;��H;��H;[�H;
�H;��H;{�H;!�H;��H;��H;��H;W�H;O�H;��H;��H;J�H;��H;��H;j�H; �H;}�H;��H;�H;;�H;Y�H;;�H;�H;��H;}�H; �H;j�H;��H;��H;J�H;��H;��H;O�H;W�H;��H;��H;��H;!�H;{�H;��H;
�H;[�H;��H;��H;��H;�rH;�cH;�RH;)?H;)H;�H;,�G;/�G;��G;��G;�G;      ?ZF;�cF;5�F;��F;�F;�!G;EaG;�G;��G;iH; )H;�FH;�]H;�pH;5�H;�H; �H;��H;��H;��H;	�H;e�H;��H;E�H;�H;5�H;��H;��H;u�H;��H;��H;��H;,�H;~�H;��H;�H;�H;�H;��H;~�H;,�H;��H;��H;��H;u�H;��H;��H;5�H;�H;E�H;��H;e�H;	�H;��H;��H;��H; �H;�H;5�H;�pH;�]H;�FH; )H;iH;��G;�G;EaG;�!G;�F;��F;5�F;�cF;      �VC; nC; �C;�D;|�D;V4E;)�E;�ZF;��F;�KG;,�G;��G;c H;^EH;D`H;=uH;#�H;��H;��H;b�H;<�H;��H;�H;I�H;�H;�H;O�H;��H;��H;��H;��H;��H;��H;=�H;��H;��H;��H;��H;��H;=�H;��H;��H;��H;��H;��H;��H;O�H;�H;�H;I�H;�H;��H;<�H;b�H;��H;��H;#�H;=uH;D`H;^EH;c H;��G;,�G;�KG;��F;�ZF;)�E;V4E;|�D;�D; �C; nC;      ��<;M�<;P\=;�N>;�?;��@;�6B;u�C;-�D;ͱE;��F;�!G;�G;1�G;
)H;iOH;FjH;gH;W�H;Y�H;�H;߷H;��H;H�H;I�H;E�H;W�H;��H;,�H;B�H;�H;�H;�H;��H;H�H;��H;��H;��H;H�H;��H;�H;�H;�H;B�H;,�H;��H;W�H;E�H;I�H;H�H;��H;߷H;�H;Y�H;W�H;gH;FjH;iOH;
)H;1�G;�G;�!G;��F;ͱE;-�D;u�C;�6B;��@;�?;�N>;P\=;M�<;      Y.;�.;�0;2;��4;�7;�{:;v\=;��?;�6B;�D;rnE;fwF;e4G;ߵG;
H;?H;aH;�yH;��H;.�H;ܫH;`�H;��H;�H;��H;��H;�H;)�H;��H;��H;h�H;c�H;O�H;��H;(�H;P�H;(�H;��H;O�H;c�H;h�H;��H;��H;)�H;�H;��H;��H;�H;��H;`�H;ܫH;.�H;��H;�yH;aH;?H;
H;ߵG;e4G;fwF;rnE;�D;�6B;��?;v\=;�{:;�7;��4;2;�0;�.;      ^;��;Ml;VZ;�_;%;+;8�0;G6;��:;��>;��A;�D;�E;`�F;PzG;t�G;1H;ZH;�uH;��H;g�H;ܫH;߷H;��H;e�H;��H;��H;��H;��H;H�H;G�H;��H;��H;p�H;��H;��H;��H;p�H;��H;��H;G�H;H�H;��H;��H;��H;��H;e�H;��H;߷H;ܫH;g�H;��H;�uH;ZH;1H;t�G;PzG;`�F;�E;�D;��A;��>;��:;G6;8�0;+;%;�_;VZ;Ml;��;      ��:B,�:#f�:���:~�:^;��;��;��#;y�,;��4;Q�:;�W?;.�B;��D;�ZF;FG;�G;}'H;VH;�tH;��H;.�H;�H;<�H;	�H;��H;��H;��H;��H;��H;��H;��H;��H;��H;^�H;b�H;^�H;��H;��H;��H;��H;��H;��H;��H;��H;��H;	�H;<�H;�H;.�H;��H;�tH;VH;}'H;�G;FG;�ZF;��D;.�B;�W?;Q�:;��4;y�,;��#;��;��;^;~�:���:#f�:B,�:      %�e9��9��9�:��Y:�x�:v:�:��:0^;8�;�";r-;(G6;��<;2>A;0D;�F;f"G;�G;$H;VH;�uH;��H;Y�H;b�H;��H;!�H;��H;��H;E�H;��H;��H;��H;6�H;�H;��H;�H;��H;�H;6�H;��H;��H;��H;E�H;��H;��H;!�H;��H;b�H;Y�H;��H;�uH;VH;$H;�G;f"G;�F;0D;2>A;��<;(G6;r-;�";8�;0^;��:v:�:�x�:��Y:�:��9��9      �����뺸кh����Y����k89w5:O.�:�c�:�A;�l;@?&;~2;�{:;` @;��C;�E;�G;�G;}'H;ZH;�yH;W�H;��H;��H;{�H;��H;��H;l�H;��H;
�H;[�H;<�H;W�H;
�H;��H;
�H;W�H;<�H;[�H;
�H;��H;l�H;��H;��H;{�H;��H;��H;W�H;�yH;ZH;}'H;�G;�G;�E;��C;` @;�{:;~2;@?&;�l;�A;�c�:O.�:w5:�k89���Y�h����к���      暩�\���4J��Y��T�b�)�-�3��YJx�-��#:��:?��:9�;� ;��.;/�8;��?;2�C;�E;f"G;�G;1H;aH;gH;��H;��H;��H;��H;s�H;(�H;I�H;J�H;��H;(�H;��H;G�H;��H;G�H;��H;(�H;��H;J�H;I�H;(�H;s�H;��H;��H;��H;��H;gH;aH;1H;�G;f"G;�E;2�C;��?;/�8;��.;� ;9�;?��:��:#:-��YJx�3��)�-�T�b�Y��4J��\���      �B(��%�����_�}����˻	��.�b�x&�c ��@���Y:�:T^;B�;��,;Z_8;��?;��C;�F;FG;t�G;?H;FjH;#�H; �H;
�H;k�H;��H;~�H;��H;/�H;��H;��H;��H;��H;��H;��H;��H;��H;��H;/�H;��H;~�H;��H;k�H;
�H; �H;#�H;FjH;?H;t�G;FG;�F;��C;��?;Z_8;��,;B�;T^;�:��Y:@�c ��x&�.�b�	���˻}����_�����%�      �����x���#��(F{���]��E<����J�뻲���bd\���]�-2:��:���:�Z;��,;/�8;` @;0D;�ZF;PzG;
H;iOH;=uH;�H;[�H;�H;C�H;z�H;��H;��H;��H;��H;��H;��H;��H;��H;��H;��H;��H;��H;��H;z�H;C�H;�H;[�H;�H;=uH;iOH;
H;PzG;�ZF;0D;` @;/�8;��,;�Z;���:��:-2:]���bd\�����J�뻛���E<���]�(F{��#���x��      >�Ｘ���o�Wrμ����bv��="���]N�����?ݻf^��z��.�Y�a�9��:���:B�;��.;�{:;2>A;��D;`�F;ߵG;
)H;D`H;5�H;��H;�H;R�H;6�H;R�H;t�H;�H;.�H;k�H;��H;��H;��H;k�H;.�H;�H;t�H;R�H;6�H;R�H;�H;��H;5�H;D`H;
)H;ߵG;`�F;��D;2>A;�{:;��.;B�;���:��:a�9.�Y�z��f^���?ݻ����]N�="��bv������Wrμ�o༸��      Gn;�`\8��s/�(�!�h��>���Prμ��������E<�������N3��Ix�a�9��:T^;� ;~2;��<;.�B;�E;e4G;1�G;^EH;�pH;��H;h�H;ϳH;k�H;��H;��H;�H;��H;1�H;��H;�H;��H;1�H;��H;�H;��H;��H;k�H;ϳH;h�H;��H;�pH;^EH;1�G;e4G;�E;.�B;��<;~2;� ;T^;��:a�9�Ix��N3�������E<��������Prμ>���h��(�!��s/�`\8�      ���������Ȅ�KSt���Y�Dn;�O�P#���Oļ�����&R��_������N3�.�Y�-2:�:9�;@?&;(G6;�W?;�D;fwF;�G;c H;�]H;��H;�H;�H;a�H;#�H;�H;��H;(�H;��H;i�H;%�H;i�H;��H;(�H;��H;�H;#�H;a�H;�H;�H;��H;�]H;c H;�G;fwF;�D;�W?;(G6;@?&;9�;�:-2:.�Y��N3������_��&R������OļP#��O�Dn;���Y�KSt��Ȅ�����      ��ѽ�[νa�ý�㳽&����L��r�d�Z\8�c���ټWv����Y��_����z��]���Y:?��:�l;r-;Q�:;��A;rnE;�!G;��G;�FH;�rH;�H;��H;�H;J�H;5�H;��H;��H;��H;B�H;�H;B�H;��H;��H;��H;5�H;J�H;�H;��H;�H;�rH;�FH;��G;�!G;rnE;��A;Q�:;r-;�l;?��:��Y:]�z������_���Y�Wv���ټc��Z\8�r�d��L��&����㳽a�ý�[ν      ��]�È�a}�q�_�ý�u�������K����o�Wv���&R���f^����@���:�A;�";��4;��>;�D;��F;,�G; )H;�cH;��H;5�H;��H;N�H;M�H;��H;��H;<�H;(�H;��H;(�H;<�H;��H;��H;M�H;N�H;��H;5�H;��H;�cH; )H;,�G;��F;�D;��>;��4;�";�A;��:@���f^�����&R�Wv���o����K������u��_�ýq�a}�È�]�      j+X��T��nH�ؕ6�� �Y��(��㳽����mR����ټ�����E<��?ݻbd\�c ��#:�c�:8�;y�,;��:;�6B;ͱE;�KG;iH;�RH;�zH;��H;
�H;9�H;`�H;n�H;+�H;��H;�H;��H;�H;��H;+�H;n�H;`�H;9�H;
�H;��H;�zH;�RH;iH;�KG;ͱE;�6B;��:;y�,;8�;�c�:#:c ��bd\��?ݻ�E<������ټ���mR�����㳽(�Y��� �ؕ6��nH��T�      Ѱ������n���*|�4S\�� :����Z�U$������K�c���Oļ����������x&�-��O.�:0^;��#;G6;��?;-�D;��F;��G;)?H;�oH;�H;��H;:�H;q�H;J�H;��H;��H;��H;��H;��H;��H;��H;J�H;q�H;:�H;��H;�H;�oH;)?H;��G;��F;-�D;��?;G6;��#;0^;O.�:-��x&������������Oļc���K����U$���Z���� :�4S\��*|�n������      -�; 9ɾi㼾�A�������Mw��nH�����Z��㳽����Z\8�P#�������]N�J��.�b�YJx�w5:��:��;8�0;v\=;u�C;�ZF;�G;)H;eH;��H;F�H;g�H;��H;7�H;��H;P�H;��H;��H;��H;P�H;��H;7�H;��H;g�H;F�H;��H;eH;)H;�G;�ZF;u�C;v\=;8�0;��;��:w5:YJx�.�b�J���]N�����P#��Z\8������㳽�Z񽞯��nH��Mw������A��i㼾 9ɾ      #y��v�R���-�߾����0��1����nH���(Ὁu��r�d�O�Prμ="�����	��3���k89v:�:��;+;�{:;�6B;)�E;EaG;�H;ZH;��H;M�H;ĮH;�H;e�H;e�H;*�H;��H;��H;��H;*�H;e�H;e�H;�H;ĮH;M�H;��H;ZH;�H;EaG;)�E;�6B;�{:;+;��;v:�:�k893��	�����="��PrμO�r�d��u��(����nH�1���0������-�߾R����v�      �O/�aM+�I�����1W�� 9ɾ0���Mw�� :�Y��_�ý�L��Dn;�>���bv���E<��˻)�-����x�:^;%;�7;��@;V4E;�!G;,�G;hOH;1zH;��H;��H;��H;��H;�H;2�H;�H;��H;�H;2�H;�H;��H;��H;��H;��H;1zH;hOH;,�G;�!G;V4E;��@;�7;%;^;�x�:��)�-��˻�E<�bv��>���Dn;��L��_�ýY��� :��Mw�0�� 9ɾ1W�����I��aM+�      $�X�EvS�%E��O/��S�1W����������4S\�� �q�&�����Y�h��������]�}���T�b��Y���Y:~�:�_;��4;�?;|�D;�F;/�G;5EH;tH;�H;��H;��H;3�H;��H;E�H;7�H;�H;7�H;E�H;��H;3�H;��H;��H;�H;tH;5EH;/�G;�F;|�D;�?;��4;�_;~�:��Y:�Y�T�b�}�����]�����h����Y�&���q�� �4S\���������1W���S��O/�%E�EvS�      � ����y�M�h�ބN��O/����-�߾�A���*|�ؕ6�a}��㳽KSt�(�!�Wrμ(F{��_�Y��h����:���:VZ;2;�N>;�D;��F;��G;J<H;�oH;��H;t�H;��H;��H;��H;��H;��H;�H;��H;��H;��H;��H;��H;t�H;��H;�oH;J<H;��G;��F;�D;�N>;2;VZ;���:�:h���Y���_�(F{�Wrμ(�!�KSt��㳽a}�ؕ6��*|��A��-�߾����O/�ބN�M�h���y�      1v��V���L ��M�h�%E�I��R���i㼾n���nH�È�a�ý�Ȅ��s/��o༼#�����4J���к��9#f�:Ml;�0;P\=; �C;5�F;��G;Q5H;^lH;H�H;ϤH;��H;�H;b�H;��H;#�H; �H;#�H;��H;b�H;�H;��H;ϤH;H�H;^lH;Q5H;��G;5�F; �C;P\=;�0;Ml;#f�:��9�к4J������#���o��s/��Ȅ�a�ýÈ��nH�n��i㼾R���I��%E�M�h�L ��V���      ph��"���V�����y�EvS�aM+��v� 9ɾ�����T�]��[ν����`\8�����x���%�\��������9B,�:��;�.;M�<; nC;�cF;�G;�0H;!jH;ǋH;ѣH;��H;��H;��H;��H;��H;��H;��H;��H;��H;��H;��H;ѣH;ǋH;!jH;�0H;�G;�cF; nC;M�<;�.;��;B,�:��9���\����%��x�����`\8������[ν]��T����� 9ɾ�v�aM+�EvS���y�V���"���      Vܿ%�ֿ�aǿ2^��&���Io���7����iþ�(���-=��` ��@����_�&]�&p����I�r�ѻ��)��R�[�:��
;*;C�:;�B;UHF;=�G;�kH;3�H;��H;h�H;��H;��H;o�H;��H;(�H;��H;(�H;��H;o�H;��H;��H;h�H;��H;3�H;�kH;=�G;UHF;�B;C�:;*;��
;[�:�R���)�r�ѻ��I�&p��&]���_��@���` ��-=��(���iþ����7�Io�&���2^���aǿ%�ֿ      %�ֿ5pѿ֊¿������PXi�Õ3��
�GD��;l��1�9�j.���R��\� �\x��1�E��ͻ��$�� ����:��;��*;[�:;.�B;3TF;��G;ZmH;ϠH;ܶH;��H;��H;��H;�H;��H;<�H;��H;<�H;��H;�H;��H;��H;��H;ܶH;ϠH;ZmH;��G;3TF;.�B;[�:;��*;��;���:� ���$��ͻ1�E�\x�� �\��R��j.��1�9�;l��GD���
�Õ3�PXi�������֊¿5pѿ      �aǿ֊¿���������s"Y��f'�����)o���.}��k/�m��ڟ�<Q�%#�ע��(;�P������/�7���:I�;�,;��;;�C;RvF;/�G;�qH;[�H;��H;=�H;�H;�H;��H;��H;j�H;��H;j�H;��H;��H;�H;�H;=�H;��H;[�H;�qH;/�G;RvF;�C;��;;�,;I�;��:/�7����P����(;�ע�%#�<Q�ڟ�m���k/��.}�)o�������f'�s"Y����������֊¿      2^������b���Io���@���޾����&ce�"����ڽ绒��f@������R���O*�mG�����u<^9Ѳ�:[;�c.;'�<;ՏC;F�F;��G;�xH;äH;8�H;I�H;��H;��H;��H;�H;��H;6�H;��H;�H;��H;��H;��H;I�H;8�H;äH;�xH;��G;F�F;ՏC;'�<;�c.;[;Ѳ�:u<^9���mG���O*��R�������f@�绒���ڽ"��&ce������޾���@�Io�b�������      &����������Io��!J�@�#��\��HD������jPH�����b��C��t +�u�ټ%��������������:���:��;�X1;3>;�/D;��F;�H;r�H;��H;)�H;��H;��H;)�H;��H;p�H;��H;~�H;��H;p�H;��H;)�H;��H;��H;)�H;��H;r�H;�H;��F;�/D;3>;�X1;��;���:��:����������%��u�ټt +�C���b�����jPH�����HD���\��@�#��!J�Io��������      Io�PXi�s"Y���@�@�#��
��о�A�� �i���(�i��gr����_��5��ɺ�o�`��<����d�@�\�M�X:OO�:6`;#�4;�?;��D;�7G;�/H;ȊH;��H;��H;.�H;��H;��H;�H;��H;-�H;��H;-�H;��H;�H;��H;��H;.�H;��H;��H;ȊH;�/H;�7G;��D;�?;#�4;6`;OO�:M�X:@�\���d��<��o�`��ɺ��5���_�gr��i����(� �i��A���о�
�@�#���@�s"Y�PXi�      ��7�Õ3��f'���\���о�����.}��-=�o
�y�ĽO��:����������7�@GĻ+�$�S�����:�z;�C&;E+8;EIA;0�E;��G;�KH;�H;��H;R�H;�H;(�H;��H;��H;@�H;��H;5�H;��H;@�H;��H;��H;(�H;�H;R�H;��H;�H;�KH;��G;0�E;EIA;E+8;�C&;�z;���:S��+�$�@GĻ�7���������:�O��y�Ľo
��-=��.}������о�\����f'�Õ3�      ���
������޾HD���A���.}��D�[t���ڽ�!��\����P�ļ�
v�F�����Jɺ�N�9���:h';�-;ӊ;;��B;�HF;��G;?eH;ʜH;�H;N�H;��H;��H;��H;{�H;��H;�H;��H;�H;��H;{�H;��H;��H;��H;N�H;�H;ʜH;?eH;��G;�HF;��B;ӊ;;�-;h';���:�N�9�Jɺ��F���
v�P�ļ���\��!����ڽ[t��D��.}��A��HD���޾�����
�      �iþGD��)o���������� �i��-=�[t����R��Tys�m +����s񗼗(;�H�ѻt@�χ!��1j:�O�:3�;�C3;}�>;CED;��F;�H;_{H;��H;��H;V�H;�H;�H;��H;9�H;R�H;��H;�H;��H;R�H;9�H;��H;�H;�H;V�H;��H;��H;_{H;�H;��F;CED;}�>;�C3;3�;�O�:�1j:χ!�t@�H�ѻ�(;�s����m +�Tys��R����[t��-=� �i���������)o��GD��      �(��;l���.}�&ce�jPH���(�o
���ڽ�R����{�4�6�� �$p��\�`�ר�-��JҺ�C^9`��:=�;�}(;t�8;IA;5{E;FiG;�<H;i�H; �H;H�H;�H;N�H;��H;��H;��H;��H;�H;i�H;�H;��H;��H;��H;��H;N�H;�H;H�H; �H;i�H;�<H;FiG;5{E;IA;t�8;�}(;=�;`��:�C^9JҺ-��ר�\�`�$p��� �4�6���{��R����ڽo
���(�jPH�&ce��.}�;l��      �-=�1�9��k/�"�����i��y�Ľ�!��Tys�4�6�#��ɺ��vz����c^��̃$������r:���:7�;�X1;>H=;jwC;WvF;R�G;/eH;m�H;��H;��H;��H;u�H;�H;��H;��H;��H;��H;��H;��H;��H;��H;��H;�H;u�H;��H;��H;��H;m�H;/eH;R�G;WvF;jwC;>H=;�X1;7�;���:��r:���̃$�c^������vz��ɺ�#�4�6�Tys��!��y�Ľi���"���k/�1�9�      �` �j.��m��ڽ�b��gr��O��\�m +�� ��ɺ�=��O*�bͻQ6R��ǅ���:���:ڃ;�);6t8;��@;�)E;�7G;t#H;p�H;c�H;�H;I�H;��H;��H;��H;�H;m�H;�H; �H;>�H; �H;�H;m�H;�H;��H;��H;��H;I�H;�H;c�H;p�H;t#H;�7G;�)E;��@;6t8;�);ڃ;���:��:�ǅ�Q6R�bͻ�O*�=��ɺ�� �m +�\�O��gr���b����ڽm��j.��      �@���R��ڟ�绒�C����_�:�������$p���vz��O*�5ֻfk������09�:_0;�� ;�C3;��=;�C;kF;��G;�[H;H;o�H;%�H;b�H;��H;��H;��H;�H;'�H;��H;n�H;��H;n�H;��H;'�H;�H;��H;��H;��H;b�H;%�H;o�H;H;�[H;��G;kF;�C;��=;�C3;�� ;_0;�:��09���fk�5ֻ�O*��vz�$p����輙��:���_�C��绒�ڟ��R��      ��_�\�<Q��f@�t +��5�����P�ļs�\�`����bͻfk��IɺB
7��:�O�:x�;%d.;��:;Z�A;c{E;�MG;q&H;/�H;�H;��H;��H;I�H;n�H;|�H;R�H;�H;��H;*�H;��H;�H;��H;*�H;��H;�H;R�H;|�H;n�H;I�H;��H;��H;�H;/�H;q&H;�MG;c{E;Z�A;��:;%d.;x�;�O�:�:B
7��Iɺfk�bͻ���\�`�s�P�ļ�����5�t +��f@�<Q�\�      &]� �%#�����u�ټ�ɺ������
v��(;�ר�c^��Q6R����B
7����:���:N�;k�*;+8;� @;��D;��F;'�G; eH;��H;��H;ľH;��H;�H;��H;B�H;��H;��H;��H;��H;B�H;u�H;B�H;��H;��H;��H;��H;B�H;��H;�H;��H;ľH;��H;��H; eH;'�G;��F;��D;� @;+8;k�*;N�;���:���:B
7����Q6R�c^��ר��(;��
v������ɺ�u�ټ����%#� �      &p��\x��ע��R��%��o�`��7�F��H�ѻ-��̃$��ǅ���09�:���:�; ~(;�Y6;��>;�C;&HF;�G;DH;s�H;�H;θH;2�H;K�H;2�H;�H;��H;��H;��H;,�H;�H;��H;��H;��H;�H;,�H;��H;��H;��H;�H;2�H;K�H;2�H;θH;�H;s�H;DH;�G;&HF;�C;��>;�Y6; ~(;�;���:�:��09�ǅ�̃$�-��H�ѻF���7�o�`�%���R��ע�\x��      ��I�1�E��(;��O*�����<��@GĻ��t@�JҺ���:�:�O�:N�; ~(;R�5;>;pC;k�E;�bG;k#H;"{H;^�H;I�H;��H;��H;Y�H;��H;:�H;w�H;��H;h�H;��H;Y�H;��H;�H;��H;Y�H;��H;h�H;��H;w�H;:�H;��H;Y�H;��H;��H;I�H;^�H;"{H;k#H;�bG;k�E;pC;>;R�5; ~(;N�;�O�:�:��:���JҺt@���@GĻ�<������O*��(;�1�E�      r�ѻ�ͻP���mG�������d�+�$��Jɺχ!��C^9��r:���:_0;x�;k�*;�Y6;>;n�B;��E;8G;�H;,mH;A�H;m�H;μH;��H;��H;��H;g�H;�H;��H;��H;�H;�H;��H;�H;<�H;�H;��H;�H;�H;��H;��H;�H;g�H;��H;��H;��H;μH;m�H;A�H;,mH;�H;8G;��E;n�B;>;�Y6;k�*;x�;_0;���:��r:�C^9χ!��Jɺ+�$���d����mG��P����ͻ      ��)���$�����������@�\�S���N�9�1j:`��:���:ڃ;�� ;%d.;+8;��>;pC;��E;�(G;��G;>cH;��H;��H;��H;��H;T�H;��H;��H;��H;��H;��H;a�H;��H;w�H;�H;I�H;b�H;I�H;�H;w�H;��H;a�H;��H;��H;��H;��H;��H;T�H;��H;��H;��H;��H;>cH;��G;�(G;��E;pC;��>;+8;%d.;�� ;ڃ;���:`��:�1j:�N�9S��@�\�������������$�      �R�� �/�7�u<^9��:M�X:���:���:�O�:=�;7�;�);�C3;��:;� @;�C;k�E;8G;��G;�_H;��H;?�H;?�H;��H;d�H;Q�H;i�H;w�H;��H;��H;��H;$�H;��H;��H;@�H;{�H;{�H;{�H;@�H;��H;��H;$�H;��H;��H;��H;w�H;i�H;Q�H;d�H;��H;?�H;?�H;��H;�_H;��G;8G;k�E;�C;� @;��:;�C3;�);7�;=�;�O�:���:���:M�X:��:u<^9/�7�� �      [�:���:��:Ѳ�:���:OO�:�z;h';3�;�}(;�X1;6t8;��=;Z�A;��D;&HF;�bG;�H;>cH;��H;m�H;��H;R�H;�H;��H;Y�H;d�H;��H;<�H;��H;��H;��H;l�H;��H;X�H;��H;��H;��H;X�H;��H;l�H;��H;��H;��H;<�H;��H;d�H;Y�H;��H;�H;R�H;��H;m�H;��H;>cH;�H;�bG;&HF;��D;Z�A;��=;6t8;�X1;�}(;3�;h';�z;OO�:���:Ѳ�:��:���:      ��
;��;I�;[;��;6`;�C&;�-;�C3;t�8;>H=;��@;�C;c{E;��F;�G;k#H;,mH;��H;?�H;��H;��H;Y�H;:�H;��H;��H;��H;��H;~�H;�H;4�H;�H;��H;1�H;r�H;��H;��H;��H;r�H;1�H;��H;�H;4�H;�H;~�H;��H;��H;��H;��H;:�H;Y�H;��H;��H;?�H;��H;,mH;k#H;�G;��F;c{E;�C;��@;>H=;t�8;�C3;�-;�C&;6`;��;[;I�;��;      *;��*;�,;�c.;�X1;#�4;E+8;ӊ;;}�>;IA;jwC;�)E;kF;�MG;'�G;DH;"{H;A�H;��H;?�H;R�H;Y�H;��H;�H;�H;w�H;#�H;�H;��H;��H;��H;��H;��H;L�H;��H;��H;��H;��H;��H;L�H;��H;��H;��H;��H;��H;�H;#�H;w�H;�H;�H;��H;Y�H;R�H;?�H;��H;A�H;"{H;DH;'�G;�MG;kF;�)E;jwC;IA;}�>;ӊ;;E+8;#�4;�X1;�c.;�,;��*;      C�:;[�:;��;;'�<;3>;�?;EIA;��B;CED;5{E;WvF;�7G;��G;q&H; eH;s�H;^�H;m�H;��H;��H;�H;:�H;�H;��H;5�H;��H;��H;G�H;��H;~�H;(�H;��H;,�H;l�H;��H;��H;��H;��H;��H;l�H;,�H;��H;(�H;~�H;��H;G�H;��H;��H;5�H;��H;�H;:�H;�H;��H;��H;m�H;^�H;s�H; eH;q&H;��G;�7G;WvF;5{E;CED;��B;EIA;�?;3>;'�<;��;;[�:;      �B;.�B;�C;ՏC;�/D;��D;0�E;�HF;��F;FiG;R�G;t#H;�[H;/�H;��H;�H;I�H;μH;��H;d�H;��H;��H;�H;5�H;��H;��H;�H;T�H;8�H;�H;��H;��H;=�H;��H;��H;��H;��H;��H;��H;��H;=�H;��H;��H;�H;8�H;T�H;�H;��H;��H;5�H;�H;��H;��H;d�H;��H;μH;I�H;�H;��H;/�H;�[H;t#H;R�G;FiG;��F;�HF;0�E;��D;�/D;ՏC;�C;.�B;      UHF;3TF;RvF;F�F;��F;�7G;��G;��G;�H;�<H;/eH;p�H;H;�H;��H;θH;��H;��H;T�H;Q�H;Y�H;��H;w�H;��H;��H;	�H;9�H;�H;��H;R�H;��H;.�H;C�H;}�H;��H;��H;��H;��H;��H;}�H;C�H;.�H;��H;R�H;��H;�H;9�H;	�H;��H;��H;w�H;��H;Y�H;Q�H;T�H;��H;��H;θH;��H;�H;H;p�H;/eH;�<H;�H;��G;��G;�7G;��F;F�F;RvF;3TF;      =�G;��G;/�G;��G;�H;�/H;�KH;?eH;_{H;i�H;m�H;c�H;o�H;��H;ľH;2�H;��H;��H;��H;i�H;d�H;��H;#�H;��H;�H;9�H;�H;��H;[�H;��H;��H;<�H;\�H;�H;��H;��H;��H;��H;��H;�H;\�H;<�H;��H;��H;[�H;��H;�H;9�H;�H;��H;#�H;��H;d�H;i�H;��H;��H;��H;2�H;ľH;��H;o�H;c�H;m�H;i�H;_{H;?eH;�KH;�/H;�H;��G;/�G;��G;      �kH;ZmH;�qH;�xH;r�H;ȊH;�H;ʜH;��H; �H;��H;�H;%�H;��H;��H;K�H;Y�H;��H;��H;w�H;��H;��H;�H;G�H;T�H;�H;��H;B�H;��H;��H;�H;B�H;k�H;l�H;��H;��H;��H;��H;��H;l�H;k�H;B�H;�H;��H;��H;B�H;��H;�H;T�H;G�H;�H;��H;��H;w�H;��H;��H;Y�H;K�H;��H;��H;%�H;�H;��H; �H;��H;ʜH;�H;ȊH;r�H;�xH;�qH;ZmH;      3�H;ϠH;[�H;äH;��H;��H;��H;�H;��H;H�H;��H;I�H;b�H;I�H;�H;2�H;��H;g�H;��H;��H;<�H;~�H;��H;��H;8�H;��H;[�H;��H;��H;�H;6�H;S�H;j�H;k�H;j�H;u�H;u�H;u�H;j�H;k�H;j�H;S�H;6�H;�H;��H;��H;[�H;��H;8�H;��H;��H;~�H;<�H;��H;��H;g�H;��H;2�H;�H;I�H;b�H;I�H;��H;H�H;��H;�H;��H;��H;��H;äH;[�H;ϠH;      ��H;ܶH;��H;8�H;)�H;��H;R�H;N�H;V�H;�H;��H;��H;��H;n�H;��H;�H;:�H;�H;��H;��H;��H;�H;��H;~�H;�H;R�H;��H;��H;�H;+�H;J�H;I�H;X�H;h�H;P�H;b�H;{�H;b�H;P�H;h�H;X�H;I�H;J�H;+�H;�H;��H;��H;R�H;�H;~�H;��H;�H;��H;��H;��H;�H;:�H;�H;��H;n�H;��H;��H;��H;�H;V�H;N�H;R�H;��H;)�H;8�H;��H;ܶH;      h�H;��H;=�H;I�H;��H;.�H;�H;��H;�H;N�H;u�H;��H;��H;|�H;B�H;��H;w�H;��H;��H;��H;��H;4�H;��H;(�H;��H;��H;��H;�H;6�H;J�H;a�H;T�H;E�H;E�H;c�H;U�H;6�H;U�H;c�H;E�H;E�H;T�H;a�H;J�H;6�H;�H;��H;��H;��H;(�H;��H;4�H;��H;��H;��H;��H;w�H;��H;B�H;|�H;��H;��H;u�H;N�H;�H;��H;�H;.�H;��H;I�H;=�H;��H;      ��H;��H;�H;��H;��H;��H;(�H;��H;�H;��H;�H;��H;��H;R�H;��H;��H;��H;��H;a�H;$�H;��H;�H;��H;��H;��H;.�H;<�H;B�H;S�H;I�H;T�H;Z�H;C�H;=�H;O�H;4�H;+�H;4�H;O�H;=�H;C�H;Z�H;T�H;I�H;S�H;B�H;<�H;.�H;��H;��H;��H;�H;��H;$�H;a�H;��H;��H;��H;��H;R�H;��H;��H;�H;��H;�H;��H;(�H;��H;��H;��H;�H;��H;      ��H;��H;�H;��H;)�H;��H;��H;��H;��H;��H;��H;�H;�H;�H;��H;��H;h�H;�H;��H;��H;l�H;��H;��H;,�H;=�H;C�H;\�H;k�H;j�H;X�H;E�H;C�H;G�H;C�H;"�H;#�H;S�H;#�H;"�H;C�H;G�H;C�H;E�H;X�H;j�H;k�H;\�H;C�H;=�H;,�H;��H;��H;l�H;��H;��H;�H;h�H;��H;��H;�H;�H;�H;��H;��H;��H;��H;��H;��H;)�H;��H;�H;��H;      o�H;�H;��H;��H;��H;�H;��H;{�H;9�H;��H;��H;m�H;'�H;��H;��H;,�H;��H;�H;w�H;��H;��H;1�H;L�H;l�H;��H;}�H;�H;l�H;k�H;h�H;E�H;=�H;C�H;-�H;�H;$�H;)�H;$�H;�H;-�H;C�H;=�H;E�H;h�H;k�H;l�H;�H;}�H;��H;l�H;L�H;1�H;��H;��H;w�H;�H;��H;,�H;��H;��H;'�H;m�H;��H;��H;9�H;{�H;��H;�H;��H;��H;��H;�H;      ��H;��H;��H;�H;p�H;��H;@�H;��H;R�H;��H;��H;�H;��H;*�H;��H;�H;Y�H;��H;�H;@�H;X�H;r�H;��H;��H;��H;��H;��H;��H;j�H;P�H;c�H;O�H;"�H;�H;'�H;�H;�H;�H;'�H;�H;"�H;O�H;c�H;P�H;j�H;��H;��H;��H;��H;��H;��H;r�H;X�H;@�H;�H;��H;Y�H;�H;��H;*�H;��H;�H;��H;��H;R�H;��H;@�H;��H;p�H;�H;��H;��H;      (�H;<�H;j�H;��H;��H;-�H;��H;�H;��H;�H;��H; �H;n�H;��H;B�H;��H;��H;�H;I�H;{�H;��H;��H;��H;��H;��H;��H;��H;��H;u�H;b�H;U�H;4�H;#�H;$�H;�H;�H;�H;�H;�H;$�H;#�H;4�H;U�H;b�H;u�H;��H;��H;��H;��H;��H;��H;��H;��H;{�H;I�H;�H;��H;��H;B�H;��H;n�H; �H;��H;�H;��H;�H;��H;-�H;��H;��H;j�H;<�H;      ��H;��H;��H;6�H;~�H;��H;5�H;��H;�H;i�H;��H;>�H;��H;�H;u�H;��H;�H;<�H;b�H;{�H;��H;��H;��H;��H;��H;��H;��H;��H;u�H;{�H;6�H;+�H;S�H;)�H;�H;�H;�H;�H;�H;)�H;S�H;+�H;6�H;{�H;u�H;��H;��H;��H;��H;��H;��H;��H;��H;{�H;b�H;<�H;�H;��H;u�H;�H;��H;>�H;��H;i�H;�H;��H;5�H;��H;~�H;6�H;��H;��H;      (�H;<�H;j�H;��H;��H;-�H;��H;�H;��H;�H;��H; �H;n�H;��H;B�H;��H;��H;�H;I�H;{�H;��H;��H;��H;��H;��H;��H;��H;��H;u�H;b�H;U�H;4�H;#�H;$�H;�H;�H;�H;�H;�H;$�H;#�H;4�H;U�H;b�H;u�H;��H;��H;��H;��H;��H;��H;��H;��H;{�H;I�H;�H;��H;��H;B�H;��H;n�H; �H;��H;�H;��H;�H;��H;-�H;��H;��H;j�H;<�H;      ��H;��H;��H;�H;p�H;��H;@�H;��H;R�H;��H;��H;�H;��H;*�H;��H;�H;Y�H;��H;�H;@�H;X�H;r�H;��H;��H;��H;��H;��H;��H;j�H;P�H;c�H;O�H;"�H;�H;'�H;�H;�H;�H;'�H;�H;"�H;O�H;c�H;P�H;j�H;��H;��H;��H;��H;��H;��H;r�H;X�H;@�H;�H;��H;Y�H;�H;��H;*�H;��H;�H;��H;��H;R�H;��H;@�H;��H;p�H;�H;��H;��H;      o�H;�H;��H;��H;��H;�H;��H;{�H;9�H;��H;��H;m�H;'�H;��H;��H;,�H;��H;�H;w�H;��H;��H;1�H;L�H;l�H;��H;}�H;�H;l�H;k�H;h�H;E�H;=�H;C�H;-�H;�H;$�H;)�H;$�H;�H;-�H;C�H;=�H;E�H;h�H;k�H;l�H;�H;}�H;��H;l�H;L�H;1�H;��H;��H;w�H;�H;��H;,�H;��H;��H;'�H;m�H;��H;��H;9�H;{�H;��H;�H;��H;��H;��H;�H;      ��H;��H;�H;��H;)�H;��H;��H;��H;��H;��H;��H;�H;�H;�H;��H;��H;h�H;�H;��H;��H;l�H;��H;��H;,�H;=�H;C�H;\�H;k�H;j�H;X�H;E�H;C�H;G�H;C�H;"�H;#�H;S�H;#�H;"�H;C�H;G�H;C�H;E�H;X�H;j�H;k�H;\�H;C�H;=�H;,�H;��H;��H;l�H;��H;��H;�H;h�H;��H;��H;�H;�H;�H;��H;��H;��H;��H;��H;��H;)�H;��H;�H;��H;      ��H;��H;�H;��H;��H;��H;(�H;��H;�H;��H;�H;��H;��H;R�H;��H;��H;��H;��H;a�H;$�H;��H;�H;��H;��H;��H;.�H;<�H;B�H;S�H;I�H;T�H;Z�H;C�H;=�H;O�H;4�H;+�H;4�H;O�H;=�H;C�H;Z�H;T�H;I�H;S�H;B�H;<�H;.�H;��H;��H;��H;�H;��H;$�H;a�H;��H;��H;��H;��H;R�H;��H;��H;�H;��H;�H;��H;(�H;��H;��H;��H;�H;��H;      h�H;��H;=�H;I�H;��H;.�H;�H;��H;�H;N�H;u�H;��H;��H;|�H;B�H;��H;w�H;��H;��H;��H;��H;4�H;��H;(�H;��H;��H;��H;�H;6�H;J�H;a�H;T�H;E�H;E�H;c�H;U�H;6�H;U�H;c�H;E�H;E�H;T�H;a�H;J�H;6�H;�H;��H;��H;��H;(�H;��H;4�H;��H;��H;��H;��H;w�H;��H;B�H;|�H;��H;��H;u�H;N�H;�H;��H;�H;.�H;��H;I�H;=�H;��H;      ��H;ܶH;��H;8�H;)�H;��H;R�H;N�H;V�H;�H;��H;��H;��H;n�H;��H;�H;:�H;�H;��H;��H;��H;�H;��H;~�H;�H;R�H;��H;��H;�H;+�H;J�H;I�H;X�H;h�H;P�H;b�H;{�H;b�H;P�H;h�H;X�H;I�H;J�H;+�H;�H;��H;��H;R�H;�H;~�H;��H;�H;��H;��H;��H;�H;:�H;�H;��H;n�H;��H;��H;��H;�H;V�H;N�H;R�H;��H;)�H;8�H;��H;ܶH;      3�H;ϠH;[�H;äH;��H;��H;��H;�H;��H;H�H;��H;I�H;b�H;I�H;�H;2�H;��H;g�H;��H;��H;<�H;~�H;��H;��H;8�H;��H;[�H;��H;��H;�H;6�H;S�H;j�H;k�H;j�H;u�H;u�H;u�H;j�H;k�H;j�H;S�H;6�H;�H;��H;��H;[�H;��H;8�H;��H;��H;~�H;<�H;��H;��H;g�H;��H;2�H;�H;I�H;b�H;I�H;��H;H�H;��H;�H;��H;��H;��H;äH;[�H;ϠH;      �kH;ZmH;�qH;�xH;r�H;ȊH;�H;ʜH;��H; �H;��H;�H;%�H;��H;��H;K�H;Y�H;��H;��H;w�H;��H;��H;�H;G�H;T�H;�H;��H;B�H;��H;��H;�H;B�H;k�H;l�H;��H;��H;��H;��H;��H;l�H;k�H;B�H;�H;��H;��H;B�H;��H;�H;T�H;G�H;�H;��H;��H;w�H;��H;��H;Y�H;K�H;��H;��H;%�H;�H;��H; �H;��H;ʜH;�H;ȊH;r�H;�xH;�qH;ZmH;      =�G;��G;/�G;��G;�H;�/H;�KH;?eH;_{H;i�H;m�H;c�H;o�H;��H;ľH;2�H;��H;��H;��H;i�H;d�H;��H;#�H;��H;�H;9�H;�H;��H;[�H;��H;��H;<�H;\�H;�H;��H;��H;��H;��H;��H;�H;\�H;<�H;��H;��H;[�H;��H;�H;9�H;�H;��H;#�H;��H;d�H;i�H;��H;��H;��H;2�H;ľH;��H;o�H;c�H;m�H;i�H;_{H;?eH;�KH;�/H;�H;��G;/�G;��G;      UHF;3TF;RvF;F�F;��F;�7G;��G;��G;�H;�<H;/eH;p�H;H;�H;��H;θH;��H;��H;T�H;Q�H;Y�H;��H;w�H;��H;��H;	�H;9�H;�H;��H;R�H;��H;.�H;C�H;}�H;��H;��H;��H;��H;��H;}�H;C�H;.�H;��H;R�H;��H;�H;9�H;	�H;��H;��H;w�H;��H;Y�H;Q�H;T�H;��H;��H;θH;��H;�H;H;p�H;/eH;�<H;�H;��G;��G;�7G;��F;F�F;RvF;3TF;      �B;.�B;�C;ՏC;�/D;��D;0�E;�HF;��F;FiG;R�G;t#H;�[H;/�H;��H;�H;I�H;μH;��H;d�H;��H;��H;�H;5�H;��H;��H;�H;T�H;8�H;�H;��H;��H;=�H;��H;��H;��H;��H;��H;��H;��H;=�H;��H;��H;�H;8�H;T�H;�H;��H;��H;5�H;�H;��H;��H;d�H;��H;μH;I�H;�H;��H;/�H;�[H;t#H;R�G;FiG;��F;�HF;0�E;��D;�/D;ՏC;�C;.�B;      C�:;[�:;��;;'�<;3>;�?;EIA;��B;CED;5{E;WvF;�7G;��G;q&H; eH;s�H;^�H;m�H;��H;��H;�H;:�H;�H;��H;5�H;��H;��H;G�H;��H;~�H;(�H;��H;,�H;l�H;��H;��H;��H;��H;��H;l�H;,�H;��H;(�H;~�H;��H;G�H;��H;��H;5�H;��H;�H;:�H;�H;��H;��H;m�H;^�H;s�H; eH;q&H;��G;�7G;WvF;5{E;CED;��B;EIA;�?;3>;'�<;��;;[�:;      *;��*;�,;�c.;�X1;#�4;E+8;ӊ;;}�>;IA;jwC;�)E;kF;�MG;'�G;DH;"{H;A�H;��H;?�H;R�H;Y�H;��H;�H;�H;w�H;#�H;�H;��H;��H;��H;��H;��H;L�H;��H;��H;��H;��H;��H;L�H;��H;��H;��H;��H;��H;�H;#�H;w�H;�H;�H;��H;Y�H;R�H;?�H;��H;A�H;"{H;DH;'�G;�MG;kF;�)E;jwC;IA;}�>;ӊ;;E+8;#�4;�X1;�c.;�,;��*;      ��
;��;I�;[;��;6`;�C&;�-;�C3;t�8;>H=;��@;�C;c{E;��F;�G;k#H;,mH;��H;?�H;��H;��H;Y�H;:�H;��H;��H;��H;��H;~�H;�H;4�H;�H;��H;1�H;r�H;��H;��H;��H;r�H;1�H;��H;�H;4�H;�H;~�H;��H;��H;��H;��H;:�H;Y�H;��H;��H;?�H;��H;,mH;k#H;�G;��F;c{E;�C;��@;>H=;t�8;�C3;�-;�C&;6`;��;[;I�;��;      [�:���:��:Ѳ�:���:OO�:�z;h';3�;�}(;�X1;6t8;��=;Z�A;��D;&HF;�bG;�H;>cH;��H;m�H;��H;R�H;�H;��H;Y�H;d�H;��H;<�H;��H;��H;��H;l�H;��H;X�H;��H;��H;��H;X�H;��H;l�H;��H;��H;��H;<�H;��H;d�H;Y�H;��H;�H;R�H;��H;m�H;��H;>cH;�H;�bG;&HF;��D;Z�A;��=;6t8;�X1;�}(;3�;h';�z;OO�:���:Ѳ�:��:���:      �R�� �/�7�u<^9��:M�X:���:���:�O�:=�;7�;�);�C3;��:;� @;�C;k�E;8G;��G;�_H;��H;?�H;?�H;��H;d�H;Q�H;i�H;w�H;��H;��H;��H;$�H;��H;��H;@�H;{�H;{�H;{�H;@�H;��H;��H;$�H;��H;��H;��H;w�H;i�H;Q�H;d�H;��H;?�H;?�H;��H;�_H;��G;8G;k�E;�C;� @;��:;�C3;�);7�;=�;�O�:���:���:M�X:��:u<^9/�7�� �      ��)���$�����������@�\�S���N�9�1j:`��:���:ڃ;�� ;%d.;+8;��>;pC;��E;�(G;��G;>cH;��H;��H;��H;��H;T�H;��H;��H;��H;��H;��H;a�H;��H;w�H;�H;I�H;b�H;I�H;�H;w�H;��H;a�H;��H;��H;��H;��H;��H;T�H;��H;��H;��H;��H;>cH;��G;�(G;��E;pC;��>;+8;%d.;�� ;ڃ;���:`��:�1j:�N�9S��@�\�������������$�      r�ѻ�ͻP���mG�������d�+�$��Jɺχ!��C^9��r:���:_0;x�;k�*;�Y6;>;n�B;��E;8G;�H;,mH;A�H;m�H;μH;��H;��H;��H;g�H;�H;��H;��H;�H;�H;��H;�H;<�H;�H;��H;�H;�H;��H;��H;�H;g�H;��H;��H;��H;μH;m�H;A�H;,mH;�H;8G;��E;n�B;>;�Y6;k�*;x�;_0;���:��r:�C^9χ!��Jɺ+�$���d����mG��P����ͻ      ��I�1�E��(;��O*�����<��@GĻ��t@�JҺ���:�:�O�:N�; ~(;R�5;>;pC;k�E;�bG;k#H;"{H;^�H;I�H;��H;��H;Y�H;��H;:�H;w�H;��H;h�H;��H;Y�H;��H;�H;��H;Y�H;��H;h�H;��H;w�H;:�H;��H;Y�H;��H;��H;I�H;^�H;"{H;k#H;�bG;k�E;pC;>;R�5; ~(;N�;�O�:�:��:���JҺt@���@GĻ�<������O*��(;�1�E�      &p��\x��ע��R��%��o�`��7�F��H�ѻ-��̃$��ǅ���09�:���:�; ~(;�Y6;��>;�C;&HF;�G;DH;s�H;�H;θH;2�H;K�H;2�H;�H;��H;��H;��H;,�H;�H;��H;��H;��H;�H;,�H;��H;��H;��H;�H;2�H;K�H;2�H;θH;�H;s�H;DH;�G;&HF;�C;��>;�Y6; ~(;�;���:�:��09�ǅ�̃$�-��H�ѻF���7�o�`�%���R��ע�\x��      &]� �%#�����u�ټ�ɺ������
v��(;�ר�c^��Q6R����B
7����:���:N�;k�*;+8;� @;��D;��F;'�G; eH;��H;��H;ľH;��H;�H;��H;B�H;��H;��H;��H;��H;B�H;u�H;B�H;��H;��H;��H;��H;B�H;��H;�H;��H;ľH;��H;��H; eH;'�G;��F;��D;� @;+8;k�*;N�;���:���:B
7����Q6R�c^��ר��(;��
v������ɺ�u�ټ����%#� �      ��_�\�<Q��f@�t +��5�����P�ļs�\�`����bͻfk��IɺB
7��:�O�:x�;%d.;��:;Z�A;c{E;�MG;q&H;/�H;�H;��H;��H;I�H;n�H;|�H;R�H;�H;��H;*�H;��H;�H;��H;*�H;��H;�H;R�H;|�H;n�H;I�H;��H;��H;�H;/�H;q&H;�MG;c{E;Z�A;��:;%d.;x�;�O�:�:B
7��Iɺfk�bͻ���\�`�s�P�ļ�����5�t +��f@�<Q�\�      �@���R��ڟ�绒�C����_�:�������$p���vz��O*�5ֻfk������09�:_0;�� ;�C3;��=;�C;kF;��G;�[H;H;o�H;%�H;b�H;��H;��H;��H;�H;'�H;��H;n�H;��H;n�H;��H;'�H;�H;��H;��H;��H;b�H;%�H;o�H;H;�[H;��G;kF;�C;��=;�C3;�� ;_0;�:��09���fk�5ֻ�O*��vz�$p����輙��:���_�C��绒�ڟ��R��      �` �j.��m��ڽ�b��gr��O��\�m +�� ��ɺ�=��O*�bͻQ6R��ǅ���:���:ڃ;�);6t8;��@;�)E;�7G;t#H;p�H;c�H;�H;I�H;��H;��H;��H;�H;m�H;�H; �H;>�H; �H;�H;m�H;�H;��H;��H;��H;I�H;�H;c�H;p�H;t#H;�7G;�)E;��@;6t8;�);ڃ;���:��:�ǅ�Q6R�bͻ�O*�=��ɺ�� �m +�\�O��gr���b����ڽm��j.��      �-=�1�9��k/�"�����i��y�Ľ�!��Tys�4�6�#��ɺ��vz����c^��̃$������r:���:7�;�X1;>H=;jwC;WvF;R�G;/eH;m�H;��H;��H;��H;u�H;�H;��H;��H;��H;��H;��H;��H;��H;��H;��H;�H;u�H;��H;��H;��H;m�H;/eH;R�G;WvF;jwC;>H=;�X1;7�;���:��r:���̃$�c^������vz��ɺ�#�4�6�Tys��!��y�Ľi���"���k/�1�9�      �(��;l���.}�&ce�jPH���(�o
���ڽ�R����{�4�6�� �$p��\�`�ר�-��JҺ�C^9`��:=�;�}(;t�8;IA;5{E;FiG;�<H;i�H; �H;H�H;�H;N�H;��H;��H;��H;��H;�H;i�H;�H;��H;��H;��H;��H;N�H;�H;H�H; �H;i�H;�<H;FiG;5{E;IA;t�8;�}(;=�;`��:�C^9JҺ-��ר�\�`�$p��� �4�6���{��R����ڽo
���(�jPH�&ce��.}�;l��      �iþGD��)o���������� �i��-=�[t����R��Tys�m +����s񗼗(;�H�ѻt@�χ!��1j:�O�:3�;�C3;}�>;CED;��F;�H;_{H;��H;��H;V�H;�H;�H;��H;9�H;R�H;��H;�H;��H;R�H;9�H;��H;�H;�H;V�H;��H;��H;_{H;�H;��F;CED;}�>;�C3;3�;�O�:�1j:χ!�t@�H�ѻ�(;�s����m +�Tys��R����[t��-=� �i���������)o��GD��      ���
������޾HD���A���.}��D�[t���ڽ�!��\����P�ļ�
v�F�����Jɺ�N�9���:h';�-;ӊ;;��B;�HF;��G;?eH;ʜH;�H;N�H;��H;��H;��H;{�H;��H;�H;��H;�H;��H;{�H;��H;��H;��H;N�H;�H;ʜH;?eH;��G;�HF;��B;ӊ;;�-;h';���:�N�9�Jɺ��F���
v�P�ļ���\��!����ڽ[t��D��.}��A��HD���޾�����
�      ��7�Õ3��f'���\���о�����.}��-=�o
�y�ĽO��:����������7�@GĻ+�$�S�����:�z;�C&;E+8;EIA;0�E;��G;�KH;�H;��H;R�H;�H;(�H;��H;��H;@�H;��H;5�H;��H;@�H;��H;��H;(�H;�H;R�H;��H;�H;�KH;��G;0�E;EIA;E+8;�C&;�z;���:S��+�$�@GĻ�7���������:�O��y�Ľo
��-=��.}������о�\����f'�Õ3�      Io�PXi�s"Y���@�@�#��
��о�A�� �i���(�i��gr����_��5��ɺ�o�`��<����d�@�\�M�X:OO�:6`;#�4;�?;��D;�7G;�/H;ȊH;��H;��H;.�H;��H;��H;�H;��H;-�H;��H;-�H;��H;�H;��H;��H;.�H;��H;��H;ȊH;�/H;�7G;��D;�?;#�4;6`;OO�:M�X:@�\���d��<��o�`��ɺ��5���_�gr��i����(� �i��A���о�
�@�#���@�s"Y�PXi�      &����������Io��!J�@�#��\��HD������jPH�����b��C��t +�u�ټ%��������������:���:��;�X1;3>;�/D;��F;�H;r�H;��H;)�H;��H;��H;)�H;��H;p�H;��H;~�H;��H;p�H;��H;)�H;��H;��H;)�H;��H;r�H;�H;��F;�/D;3>;�X1;��;���:��:����������%��u�ټt +�C���b�����jPH�����HD���\��@�#��!J�Io��������      2^������b���Io���@���޾����&ce�"����ڽ绒��f@������R���O*�mG�����u<^9Ѳ�:[;�c.;'�<;ՏC;F�F;��G;�xH;äH;8�H;I�H;��H;��H;��H;�H;��H;6�H;��H;�H;��H;��H;��H;I�H;8�H;äH;�xH;��G;F�F;ՏC;'�<;�c.;[;Ѳ�:u<^9���mG���O*��R�������f@�绒���ڽ"��&ce������޾���@�Io�b�������      �aǿ֊¿���������s"Y��f'�����)o���.}��k/�m��ڟ�<Q�%#�ע��(;�P������/�7���:I�;�,;��;;�C;RvF;/�G;�qH;[�H;��H;=�H;�H;�H;��H;��H;j�H;��H;j�H;��H;��H;�H;�H;=�H;��H;[�H;�qH;/�G;RvF;�C;��;;�,;I�;��:/�7����P����(;�ע�%#�<Q�ڟ�m���k/��.}�)o�������f'�s"Y����������֊¿      %�ֿ5pѿ֊¿������PXi�Õ3��
�GD��;l��1�9�j.���R��\� �\x��1�E��ͻ��$�� ����:��;��*;[�:;.�B;3TF;��G;ZmH;ϠH;ܶH;��H;��H;��H;�H;��H;<�H;��H;<�H;��H;�H;��H;��H;��H;ܶH;ϠH;ZmH;��G;3TF;.�B;[�:;��*;��;���:� ���$��ͻ1�E�\x�� �\��R��j.��1�9�;l��GD���
�Õ3�PXi�������֊¿5pѿ      ���$������꿥�ſ�ޞ�3s��2�/����� j���nHͽ������'�B<ͼ��n������Q^�0.��:�V;�R%;~n8;��A;mCF;�H;��H;��H;��H;L�H;>�H;C�H;��H;��H;��H;+�H;��H;��H;��H;C�H;>�H;L�H;��H;��H;��H;�H;mCF;��A;~n8;�R%;�V;�:0.��Q^�������n�B<ͼ��'�����nHͽ�� j���/����2�3s��ޞ���ſ������$�      $��������~�����cm�L�-�����Fh��Ide�-�̪ɽ�v��#�$���ɼ�mj�o����X�8��mĆ:�w;i�%;M�8;B;{QF;H;5�H;U�H;�H;p�H;B�H;5�H;��H;��H;��H;$�H;��H;��H;��H;5�H;B�H;p�H;�H;U�H;5�H;H;{QF;B;M�8;i�%;�w;mĆ:8���X�o����mj���ɼ#�$��v��̪ɽ-�Ide�Fh������L�-�cm����~���忖����      ������{���ԿBw�����/�\��"����b��M0X�}���;����w����������]�X��VF�2��nȒ:0�;^�';׎9;1oB;�yF;� H;��H;7�H;�H;��H;F�H;:�H;��H;��H;��H;�H;��H;��H;��H;:�H;F�H;��H;�H;7�H;��H;� H;�yF;1oB;׎9;^�';0�;nȒ:2��VF�X�黼�]����������w��;��}��M0X�b������"�/�\����Bw���Կ{�𿖏�      ������Կp���ޞ�RF�]�C�$E��;�I��sD�|�"��]�c�y��֯���J�P�ѻ]�)���K����:P�
;M*;��:;�C;�F;�7H;Z�H;��H;w�H;��H;>�H;9�H;��H;��H;��H;��H;��H;��H;��H;9�H;>�H;��H;w�H;��H;Z�H;�7H;�F;�C;��:;M*;P�
;���:��K�]�)�P�ѻ��J��֯�y�]�c�"��|�sD��I���;$E�]�C�RF��ޞ�p���Կ��      ��ſ~��Bw���ޞ�|���3�W�,�%�����^ɰ��|x�\{+�ű����J��  �Ҷ��n�1�f����+�
9q�:�;4�-;��<;��C;�G;�SH;Q�H;��H;��H;��H;V�H;2�H;��H;��H;��H;��H;��H;��H;��H;2�H;V�H;��H;��H;��H;Q�H;�SH;�G;��C;��<;4�-;�;q�:
9�+�f���n�1�Ҷ���  ��J���ű�\{+��|x�^ɰ�����,�%�3�W�|����ޞ�Bw��~��      �ޞ�������RF�3�W�M�-���4Kɾ�G����O�z��ƽ����Ȅ-���ۼㄼL4�[ǐ�-ж��Z:n��:�;ʕ1;
c>;{�D;�[G;KrH;��H;i�H;e�H;'�H;u�H;)�H;h�H;��H;|�H;��H;|�H;��H;h�H;)�H;u�H;'�H;e�H;i�H;��H;KrH;�[G;{�D;
c>;ʕ1;�;n��:�Z:-ж�[ǐ�L4�ㄼ��ۼȄ-�����ƽz����O��G��4Kɾ��M�-�3�W�RF�������      3s�cm�/�\�]�C�,�%����TҾa����i��C(����UP����[�x������Y�l���X���<���k:���:)� ;�5;ZQ@;otE;�G;9�H;L�H;��H;�H;I�H;l�H;$�H;c�H;s�H;W�H;��H;W�H;s�H;c�H;$�H;l�H;I�H;�H;��H;L�H;9�H;�G;otE;ZQ@;�5;)� ;���:��k:��<��X�l����Y����x���[�UP����콡C(���i�a���TҾ��,�%�]�C�/�\�cm�      �2�L�-��"�$E�����4Kɾa��w�s�.�5�y�k㻽�v��z0��;��+��-�*�S����6�LjS� L�:��	;��(;5�9;�.B;�CF;YH;ԪH;��H;��H;��H;w�H;��H;�H;0�H;C�H;<�H;Y�H;<�H;C�H;0�H;�H;��H;w�H;��H;��H;��H;ԪH;YH;�CF;�.B;5�9;��(;��	; L�:LjS��6�S���-�*��+���;�z0��v��k㻽y�.�5�w�s�a��4Kɾ����$E��"�L�-�      /�����������;^ɰ��G����i�.�5��	�ĪɽR����J�p���沼��]�J���V
x��
��~k:4��:v;��/;�,=;��C;M�F;#HH;��H;(�H;��H;#�H;��H;��H;��H;�H;�H;�H;$�H;�H;�H;�H;��H;��H;��H;#�H;��H;(�H;��H;#HH;M�F;��C;�,=;��/;v;4��:~k:�
��V
x�J�����]��沼p���J�R���Īɽ�	�.�5���i��G��^ɰ��;��徨���      ��Fh��b���I���|x���O��C(�y�Īɽ����JDX�D��'<ͼㄼ�X!�t��hX��K����:�x;7�#;$H6;IQ@;�OE;��G;��H;��H;1�H;��H;��H;��H;v�H;��H;��H;��H;��H;��H;��H;��H;��H;��H;v�H;��H;��H;��H;1�H;��H;��H;��G;�OE;IQ@;$H6;7�#;�x;���:�K�hX�t���X!�ㄼ'<ͼD��JDX�����Īɽy��C(���O��|x��I��b��Fh��       j�Ide�M0X�sD�\{+�z�����k㻽R���JDX������ۼо����;�>ۻ�X���y�;<":I��:��;��-;��;;�B;�yF;�H;��H;|�H;&�H;��H;��H;��H;m�H;��H;��H;��H;��H;z�H;��H;��H;��H;��H;m�H;��H;��H;��H;&�H;|�H;��H;�H;�yF;�B;��;;��-;��;I��:;<":��y��X�>ۻ��;�о����ۼ���JDX�R���k㻽���z��\{+�sD�M0X�Ide�      ��-�}��|�ű�ƽUP���v���J�D����ۼ��v�J������+���sѺ$
9eL�:�;�$;#�5;�?;��D;j[G;eH;��H;��H;��H;��H;!�H;��H;T�H;n�H;Y�H;T�H;a�H;7�H;a�H;T�H;Y�H;n�H;T�H;��H;!�H;��H;��H;��H;��H;eH;j[G;��D;�?;#�5;�$;�;eL�:$
9�sѺ�+������v�J�����ۼD���J��v��UP��ƽű�|�}��-�      nHͽ̪ɽ�;��"����������[�z0�p��'<ͼо��v�J���k��+��(����:�`�:|�;�/;�K<; C;9lF;��G;�H;
�H;�H;�H;A�H;T�H;��H;%�H;/�H;�H;�H;�H;��H;�H;�H;�H;/�H;%�H;��H;T�H;A�H;�H;�H;
�H;�H;��G;9lF; C;�K<;�/;|�;�`�:���:�(�+�k����v�J�о��'<ͼp��z0���[�������"���;��̪ɽ      �����v����w�]�c��J�Ȅ-�x��;缈沼ㄼ��;�����k��66�i��K<Q:գ�:�h;M*;��8;��@;�OE;�tG;DhH;��H;��H;�H;#�H;��H;y�H;��H;��H;��H;��H;��H;��H;��H;��H;��H;��H;��H;��H;��H;y�H;��H;#�H;�H;��H;��H;DhH;�tG;�OE;��@;��8;M*;�h;գ�:K<Q:i��66�k��������;�ㄼ�沼�;�x�Ȅ-��J�]�c���w��v��      ��'�#�$����y��  ���ۼ����+����]��X!�>ۻ�+��+�i���>:\��:@�;Z�%;	�5;��>;�'D;�F;� H;8�H;[�H;��H;��H;��H;��H;k�H;��H;��H;��H;��H;g�H;K�H;m�H;K�H;g�H;��H;��H;��H;��H;k�H;��H;��H;��H;��H;[�H;8�H;� H;�F;�'D;��>;	�5;Z�%;@�;\��:�>:i��+��+��>ۻ�X!���]��+�������ۼ�  �y����#�$�      B<ͼ��ɼ�����֯�Ҷ��ㄼ��Y�-�*�J���t���X��sѺ�(�K<Q:\��:��
;u�#;��3;�b=;#C;3CF;�G;�H;��H;�H;8�H;��H;W�H;!�H;d�H;��H;b�H;5�H;O�H;	�H;��H;�H;��H;	�H;O�H;5�H;b�H;��H;d�H;!�H;W�H;��H;8�H;�H;��H;�H;�G;3CF;#C;�b=;��3;u�#;��
;\��:K<Q:�(��sѺ�X�t��J���-�*���Y�ㄼҶ���֯�������ɼ      ��n��mj���]���J�n�1�L4�l��S���V
x�hX���y�$
9���:գ�:@�;u�#;v�2;�<;�oB;7�E;��G;�dH;��H;8�H;��H;��H;��H;��H;9�H;F�H;7�H;�H;��H;��H;��H;��H;��H;��H;��H;��H;��H;�H;7�H;F�H;9�H;��H;��H;��H;��H;8�H;��H;�dH;��G;7�E;�oB;�<;v�2;u�#;@�;գ�:���:$
9��y�hX�V
x�S���l��L4�n�1���J���]��mj�      ����o���X��P�ѻf���[ǐ��X��6��
���K�;<":eL�:�`�:�h;Z�%;��3;�<;X/B;��E;�[G;�GH;M�H;��H;a�H;�H;7�H;=�H;��H;�H;�H;��H;��H;��H;]�H;O�H;K�H;'�H;K�H;O�H;]�H;��H;��H;��H;�H;�H;��H;=�H;7�H;�H;a�H;��H;M�H;�GH;�[G;��E;X/B;�<;��3;Z�%;�h;�`�:eL�:;<":�K��
���6��X�[ǐ�f���P�ѻX��o���      �Q^��X�VF�]�)��+�-ж���<�LjS�~k:���:I��:�;|�;M*;	�5;�b=;�oB;��E;�IG;\7H;s�H;��H;�H;,�H;��H;��H;��H;��H;��H;��H;��H;t�H;P�H;��H;��H;��H;��H;��H;��H;��H;P�H;t�H;��H;��H;��H;��H;��H;��H;��H;,�H;�H;��H;s�H;\7H;�IG;��E;�oB;�b=;	�5;M*;|�;�;I��:���:~k:LjS���<�-ж��+�]�)�VF��X�      0.�8��2�깦�K�
9�Z:��k: L�:4��:�x;��;�$;�/;��8;��>;#C;7�E;�[G;\7H;̤H;�H;&�H;��H;5�H;��H;P�H;��H;��H;��H;z�H;5�H;�H;��H;��H;��H;��H;u�H;��H;��H;��H;��H;�H;5�H;z�H;��H;��H;��H;P�H;��H;5�H;��H;&�H;�H;̤H;\7H;�[G;7�E;#C;��>;��8;�/;�$;��;�x;4��: L�:��k:�Z:
9��K�2��8��      �:mĆ:nȒ:���:q�:n��:���:��	;v;7�#;��-;#�5;�K<;��@;�'D;3CF;��G;�GH;s�H;�H;��H;O�H;��H;\�H;"�H;��H;��H;��H;[�H;�H;��H;��H;m�H;[�H;)�H;�H;�H;�H;)�H;[�H;m�H;��H;��H;�H;[�H;��H;��H;��H;"�H;\�H;��H;O�H;��H;�H;s�H;�GH;��G;3CF;�'D;��@;�K<;#�5;��-;7�#;v;��	;���:n��:q�:���:nȒ:mĆ:      �V;�w;0�;P�
;�;�;)� ;��(;��/;$H6;��;;�?; C;�OE;�F;�G;�dH;M�H;��H;&�H;O�H;��H;0�H;��H;e�H;�H;��H;a�H;��H;��H;��H;A�H;�H;�H;��H;��H;��H;��H;��H;�H;�H;A�H;��H;��H;��H;a�H;��H;�H;e�H;��H;0�H;��H;O�H;&�H;��H;M�H;�dH;�G;�F;�OE; C;�?;��;;$H6;��/;��(;)� ;�;�;P�
;0�;�w;      �R%;i�%;^�';M*;4�-;ʕ1;�5;5�9;�,=;IQ@;�B;��D;9lF;�tG;� H;�H;��H;��H;�H;��H;��H;0�H;�H;a�H;��H;r�H;5�H;��H;��H;��H;�H;��H;��H;��H;|�H;e�H;L�H;e�H;|�H;��H;��H;��H;�H;��H;��H;��H;5�H;r�H;��H;a�H;�H;0�H;��H;��H;�H;��H;��H;�H;� H;�tG;9lF;��D;�B;IQ@;�,=;5�9;�5;ʕ1;4�-;M*;^�';i�%;      ~n8;M�8;׎9;��:;��<;
c>;ZQ@;�.B;��C;�OE;�yF;j[G;��G;DhH;8�H;��H;8�H;a�H;,�H;5�H;\�H;��H;a�H;k�H;i�H;D�H;��H;��H;e�H;	�H;��H;��H;Y�H;(�H;"�H;�H;��H;�H;"�H;(�H;Y�H;��H;��H;	�H;e�H;��H;��H;D�H;i�H;k�H;a�H;��H;\�H;5�H;,�H;a�H;8�H;��H;8�H;DhH;��G;j[G;�yF;�OE;��C;�.B;ZQ@;
c>;��<;��:;׎9;M�8;      ��A;B;1oB;�C;��C;{�D;otE;�CF;M�F;��G;�H;eH;�H;��H;[�H;�H;��H;�H;��H;��H;"�H;e�H;��H;i�H;-�H;��H;��H;i�H; �H;��H;r�H;@�H;
�H;��H;��H;��H;��H;��H;��H;��H;
�H;@�H;r�H;��H; �H;i�H;��H;��H;-�H;i�H;��H;e�H;"�H;��H;��H;�H;��H;�H;[�H;��H;�H;eH;�H;��G;M�F;�CF;otE;{�D;��C;�C;1oB;B;      mCF;{QF;�yF;�F;�G;�[G;�G;YH;#HH;��H;��H;��H;
�H;��H;��H;8�H;��H;7�H;��H;P�H;��H;�H;r�H;D�H;��H;��H;_�H;��H;��H;`�H;�H;��H;��H;��H;o�H;\�H;n�H;\�H;o�H;��H;��H;��H;�H;`�H;��H;��H;_�H;��H;��H;D�H;r�H;�H;��H;P�H;��H;7�H;��H;8�H;��H;��H;
�H;��H;��H;��H;#HH;YH;�G;�[G;�G;�F;�yF;{QF;      �H;H;� H;�7H;�SH;KrH;9�H;ԪH;��H;��H;|�H;��H;�H;�H;��H;��H;��H;=�H;��H;��H;��H;��H;5�H;��H;��H;_�H;��H;��H;H�H;�H;��H;��H;b�H;C�H;(�H;�H;�H;�H;(�H;C�H;b�H;��H;��H;�H;H�H;��H;��H;_�H;��H;��H;5�H;��H;��H;��H;��H;=�H;��H;��H;��H;�H;�H;��H;|�H;��H;��H;ԪH;9�H;KrH;�SH;�7H;� H;H;      ��H;5�H;��H;Z�H;Q�H;��H;L�H;��H;(�H;1�H;&�H;��H;�H;#�H;��H;W�H;��H;��H;��H;��H;��H;a�H;��H;��H;i�H;��H;��H;W�H;�H;��H;u�H;F�H; �H;��H;��H;��H;��H;��H;��H;��H; �H;F�H;u�H;��H;�H;W�H;��H;��H;i�H;��H;��H;a�H;��H;��H;��H;��H;��H;W�H;��H;#�H;�H;��H;&�H;1�H;(�H;��H;L�H;��H;Q�H;Z�H;��H;5�H;      ��H;U�H;7�H;��H;��H;i�H;��H;��H;��H;��H;��H;��H;A�H;��H;��H;!�H;9�H;�H;��H;��H;[�H;��H;��H;e�H; �H;��H;H�H;�H;��H;k�H;7�H;��H;��H;��H;��H;��H;�H;��H;��H;��H;��H;��H;7�H;k�H;��H;�H;H�H;��H; �H;e�H;��H;��H;[�H;��H;��H;�H;9�H;!�H;��H;��H;A�H;��H;��H;��H;��H;��H;��H;i�H;��H;��H;7�H;U�H;      ��H;�H;�H;w�H;��H;e�H;�H;��H;#�H;��H;��H;!�H;T�H;y�H;k�H;d�H;F�H;�H;��H;z�H;�H;��H;��H;	�H;��H;`�H;�H;��H;k�H;-�H;��H;��H;��H;��H;c�H;K�H;A�H;K�H;c�H;��H;��H;��H;��H;-�H;k�H;��H;�H;`�H;��H;	�H;��H;��H;�H;z�H;��H;�H;F�H;d�H;k�H;y�H;T�H;!�H;��H;��H;#�H;��H;�H;e�H;��H;w�H;�H;�H;      L�H;p�H;��H;��H;��H;'�H;I�H;w�H;��H;��H;��H;��H;��H;��H;��H;��H;7�H;��H;��H;5�H;��H;��H;�H;��H;r�H;�H;��H;u�H;7�H;��H;��H;��H;w�H;?�H;�H;'�H;(�H;'�H;�H;?�H;w�H;��H;��H;��H;7�H;u�H;��H;�H;r�H;��H;�H;��H;��H;5�H;��H;��H;7�H;��H;��H;��H;��H;��H;��H;��H;��H;w�H;I�H;'�H;��H;��H;��H;p�H;      >�H;B�H;F�H;>�H;V�H;u�H;l�H;��H;��H;v�H;m�H;T�H;%�H;��H;��H;b�H;�H;��H;t�H;�H;��H;A�H;��H;��H;@�H;��H;��H;F�H;��H;��H;��H;_�H;A�H;�H;��H;��H;��H;��H;��H;�H;A�H;_�H;��H;��H;��H;F�H;��H;��H;@�H;��H;��H;A�H;��H;�H;t�H;��H;�H;b�H;��H;��H;%�H;T�H;m�H;v�H;��H;��H;l�H;u�H;V�H;>�H;F�H;B�H;      C�H;5�H;:�H;9�H;2�H;)�H;$�H;�H;��H;��H;��H;n�H;/�H;��H;��H;5�H;��H;��H;P�H;��H;m�H;�H;��H;Y�H;
�H;��H;b�H; �H;��H;��H;w�H;A�H;��H;��H;��H;��H;��H;��H;��H;��H;��H;A�H;w�H;��H;��H; �H;b�H;��H;
�H;Y�H;��H;�H;m�H;��H;P�H;��H;��H;5�H;��H;��H;/�H;n�H;��H;��H;��H;�H;$�H;)�H;2�H;9�H;:�H;5�H;      ��H;��H;��H;��H;��H;h�H;c�H;0�H;�H;��H;��H;Y�H;�H;��H;��H;O�H;��H;]�H;��H;��H;[�H;�H;��H;(�H;��H;��H;C�H;��H;��H;��H;?�H;�H;��H;��H;��H;��H;��H;��H;��H;��H;��H;�H;?�H;��H;��H;��H;C�H;��H;��H;(�H;��H;�H;[�H;��H;��H;]�H;��H;O�H;��H;��H;�H;Y�H;��H;��H;�H;0�H;c�H;h�H;��H;��H;��H;��H;      ��H;��H;��H;��H;��H;��H;s�H;C�H;�H;��H;��H;T�H;�H;��H;g�H;	�H;��H;O�H;��H;��H;)�H;��H;|�H;"�H;��H;o�H;(�H;��H;��H;c�H;�H;��H;��H;��H;��H;��H;��H;��H;��H;��H;��H;��H;�H;c�H;��H;��H;(�H;o�H;��H;"�H;|�H;��H;)�H;��H;��H;O�H;��H;	�H;g�H;��H;�H;T�H;��H;��H;�H;C�H;s�H;��H;��H;��H;��H;��H;      ��H;��H;��H;��H;��H;|�H;W�H;<�H;�H;��H;��H;a�H;�H;��H;K�H;��H;��H;K�H;��H;��H;�H;��H;e�H;�H;��H;\�H;�H;��H;��H;K�H;'�H;��H;��H;��H;��H;��H;��H;��H;��H;��H;��H;��H;'�H;K�H;��H;��H;�H;\�H;��H;�H;e�H;��H;�H;��H;��H;K�H;��H;��H;K�H;��H;�H;a�H;��H;��H;�H;<�H;W�H;|�H;��H;��H;��H;��H;      +�H;$�H;�H;��H;��H;��H;��H;Y�H;$�H;��H;z�H;7�H;��H;��H;m�H;�H;��H;'�H;��H;u�H;�H;��H;L�H;��H;��H;n�H;�H;��H;�H;A�H;(�H;��H;��H;��H;��H;��H;~�H;��H;��H;��H;��H;��H;(�H;A�H;�H;��H;�H;n�H;��H;��H;L�H;��H;�H;u�H;��H;'�H;��H;�H;m�H;��H;��H;7�H;z�H;��H;$�H;Y�H;��H;��H;��H;��H;�H;$�H;      ��H;��H;��H;��H;��H;|�H;W�H;<�H;�H;��H;��H;a�H;�H;��H;K�H;��H;��H;K�H;��H;��H;�H;��H;e�H;�H;��H;\�H;�H;��H;��H;K�H;'�H;��H;��H;��H;��H;��H;��H;��H;��H;��H;��H;��H;'�H;K�H;��H;��H;�H;\�H;��H;�H;e�H;��H;�H;��H;��H;K�H;��H;��H;K�H;��H;�H;a�H;��H;��H;�H;<�H;W�H;|�H;��H;��H;��H;��H;      ��H;��H;��H;��H;��H;��H;s�H;C�H;�H;��H;��H;T�H;�H;��H;g�H;	�H;��H;O�H;��H;��H;)�H;��H;|�H;"�H;��H;o�H;(�H;��H;��H;c�H;�H;��H;��H;��H;��H;��H;��H;��H;��H;��H;��H;��H;�H;c�H;��H;��H;(�H;o�H;��H;"�H;|�H;��H;)�H;��H;��H;O�H;��H;	�H;g�H;��H;�H;T�H;��H;��H;�H;C�H;s�H;��H;��H;��H;��H;��H;      ��H;��H;��H;��H;��H;h�H;c�H;0�H;�H;��H;��H;Y�H;�H;��H;��H;O�H;��H;]�H;��H;��H;[�H;�H;��H;(�H;��H;��H;C�H;��H;��H;��H;?�H;�H;��H;��H;��H;��H;��H;��H;��H;��H;��H;�H;?�H;��H;��H;��H;C�H;��H;��H;(�H;��H;�H;[�H;��H;��H;]�H;��H;O�H;��H;��H;�H;Y�H;��H;��H;�H;0�H;c�H;h�H;��H;��H;��H;��H;      C�H;5�H;:�H;9�H;2�H;)�H;$�H;�H;��H;��H;��H;n�H;/�H;��H;��H;5�H;��H;��H;P�H;��H;m�H;�H;��H;Y�H;
�H;��H;b�H; �H;��H;��H;w�H;A�H;��H;��H;��H;��H;��H;��H;��H;��H;��H;A�H;w�H;��H;��H; �H;b�H;��H;
�H;Y�H;��H;�H;m�H;��H;P�H;��H;��H;5�H;��H;��H;/�H;n�H;��H;��H;��H;�H;$�H;)�H;2�H;9�H;:�H;5�H;      >�H;B�H;F�H;>�H;V�H;u�H;l�H;��H;��H;v�H;m�H;T�H;%�H;��H;��H;b�H;�H;��H;t�H;�H;��H;A�H;��H;��H;@�H;��H;��H;F�H;��H;��H;��H;_�H;A�H;�H;��H;��H;��H;��H;��H;�H;A�H;_�H;��H;��H;��H;F�H;��H;��H;@�H;��H;��H;A�H;��H;�H;t�H;��H;�H;b�H;��H;��H;%�H;T�H;m�H;v�H;��H;��H;l�H;u�H;V�H;>�H;F�H;B�H;      L�H;p�H;��H;��H;��H;'�H;I�H;w�H;��H;��H;��H;��H;��H;��H;��H;��H;7�H;��H;��H;5�H;��H;��H;�H;��H;r�H;�H;��H;u�H;7�H;��H;��H;��H;w�H;?�H;�H;'�H;(�H;'�H;�H;?�H;w�H;��H;��H;��H;7�H;u�H;��H;�H;r�H;��H;�H;��H;��H;5�H;��H;��H;7�H;��H;��H;��H;��H;��H;��H;��H;��H;w�H;I�H;'�H;��H;��H;��H;p�H;      ��H;�H;�H;w�H;��H;e�H;�H;��H;#�H;��H;��H;!�H;T�H;y�H;k�H;d�H;F�H;�H;��H;z�H;�H;��H;��H;	�H;��H;`�H;�H;��H;k�H;-�H;��H;��H;��H;��H;c�H;K�H;A�H;K�H;c�H;��H;��H;��H;��H;-�H;k�H;��H;�H;`�H;��H;	�H;��H;��H;�H;z�H;��H;�H;F�H;d�H;k�H;y�H;T�H;!�H;��H;��H;#�H;��H;�H;e�H;��H;w�H;�H;�H;      ��H;U�H;7�H;��H;��H;i�H;��H;��H;��H;��H;��H;��H;A�H;��H;��H;!�H;9�H;�H;��H;��H;[�H;��H;��H;e�H; �H;��H;H�H;�H;��H;k�H;7�H;��H;��H;��H;��H;��H;�H;��H;��H;��H;��H;��H;7�H;k�H;��H;�H;H�H;��H; �H;e�H;��H;��H;[�H;��H;��H;�H;9�H;!�H;��H;��H;A�H;��H;��H;��H;��H;��H;��H;i�H;��H;��H;7�H;U�H;      ��H;5�H;��H;Z�H;Q�H;��H;L�H;��H;(�H;1�H;&�H;��H;�H;#�H;��H;W�H;��H;��H;��H;��H;��H;a�H;��H;��H;i�H;��H;��H;W�H;�H;��H;u�H;F�H; �H;��H;��H;��H;��H;��H;��H;��H; �H;F�H;u�H;��H;�H;W�H;��H;��H;i�H;��H;��H;a�H;��H;��H;��H;��H;��H;W�H;��H;#�H;�H;��H;&�H;1�H;(�H;��H;L�H;��H;Q�H;Z�H;��H;5�H;      �H;H;� H;�7H;�SH;KrH;9�H;ԪH;��H;��H;|�H;��H;�H;�H;��H;��H;��H;=�H;��H;��H;��H;��H;5�H;��H;��H;_�H;��H;��H;H�H;�H;��H;��H;b�H;C�H;(�H;�H;�H;�H;(�H;C�H;b�H;��H;��H;�H;H�H;��H;��H;_�H;��H;��H;5�H;��H;��H;��H;��H;=�H;��H;��H;��H;�H;�H;��H;|�H;��H;��H;ԪH;9�H;KrH;�SH;�7H;� H;H;      mCF;{QF;�yF;�F;�G;�[G;�G;YH;#HH;��H;��H;��H;
�H;��H;��H;8�H;��H;7�H;��H;P�H;��H;�H;r�H;D�H;��H;��H;_�H;��H;��H;`�H;�H;��H;��H;��H;o�H;\�H;n�H;\�H;o�H;��H;��H;��H;�H;`�H;��H;��H;_�H;��H;��H;D�H;r�H;�H;��H;P�H;��H;7�H;��H;8�H;��H;��H;
�H;��H;��H;��H;#HH;YH;�G;�[G;�G;�F;�yF;{QF;      ��A;B;1oB;�C;��C;{�D;otE;�CF;M�F;��G;�H;eH;�H;��H;[�H;�H;��H;�H;��H;��H;"�H;e�H;��H;i�H;-�H;��H;��H;i�H; �H;��H;r�H;@�H;
�H;��H;��H;��H;��H;��H;��H;��H;
�H;@�H;r�H;��H; �H;i�H;��H;��H;-�H;i�H;��H;e�H;"�H;��H;��H;�H;��H;�H;[�H;��H;�H;eH;�H;��G;M�F;�CF;otE;{�D;��C;�C;1oB;B;      ~n8;M�8;׎9;��:;��<;
c>;ZQ@;�.B;��C;�OE;�yF;j[G;��G;DhH;8�H;��H;8�H;a�H;,�H;5�H;\�H;��H;a�H;k�H;i�H;D�H;��H;��H;e�H;	�H;��H;��H;Y�H;(�H;"�H;�H;��H;�H;"�H;(�H;Y�H;��H;��H;	�H;e�H;��H;��H;D�H;i�H;k�H;a�H;��H;\�H;5�H;,�H;a�H;8�H;��H;8�H;DhH;��G;j[G;�yF;�OE;��C;�.B;ZQ@;
c>;��<;��:;׎9;M�8;      �R%;i�%;^�';M*;4�-;ʕ1;�5;5�9;�,=;IQ@;�B;��D;9lF;�tG;� H;�H;��H;��H;�H;��H;��H;0�H;�H;a�H;��H;r�H;5�H;��H;��H;��H;�H;��H;��H;��H;|�H;e�H;L�H;e�H;|�H;��H;��H;��H;�H;��H;��H;��H;5�H;r�H;��H;a�H;�H;0�H;��H;��H;�H;��H;��H;�H;� H;�tG;9lF;��D;�B;IQ@;�,=;5�9;�5;ʕ1;4�-;M*;^�';i�%;      �V;�w;0�;P�
;�;�;)� ;��(;��/;$H6;��;;�?; C;�OE;�F;�G;�dH;M�H;��H;&�H;O�H;��H;0�H;��H;e�H;�H;��H;a�H;��H;��H;��H;A�H;�H;�H;��H;��H;��H;��H;��H;�H;�H;A�H;��H;��H;��H;a�H;��H;�H;e�H;��H;0�H;��H;O�H;&�H;��H;M�H;�dH;�G;�F;�OE; C;�?;��;;$H6;��/;��(;)� ;�;�;P�
;0�;�w;      �:mĆ:nȒ:���:q�:n��:���:��	;v;7�#;��-;#�5;�K<;��@;�'D;3CF;��G;�GH;s�H;�H;��H;O�H;��H;\�H;"�H;��H;��H;��H;[�H;�H;��H;��H;m�H;[�H;)�H;�H;�H;�H;)�H;[�H;m�H;��H;��H;�H;[�H;��H;��H;��H;"�H;\�H;��H;O�H;��H;�H;s�H;�GH;��G;3CF;�'D;��@;�K<;#�5;��-;7�#;v;��	;���:n��:q�:���:nȒ:mĆ:      0.�8��2�깦�K�
9�Z:��k: L�:4��:�x;��;�$;�/;��8;��>;#C;7�E;�[G;\7H;̤H;�H;&�H;��H;5�H;��H;P�H;��H;��H;��H;z�H;5�H;�H;��H;��H;��H;��H;u�H;��H;��H;��H;��H;�H;5�H;z�H;��H;��H;��H;P�H;��H;5�H;��H;&�H;�H;̤H;\7H;�[G;7�E;#C;��>;��8;�/;�$;��;�x;4��: L�:��k:�Z:
9��K�2��8��      �Q^��X�VF�]�)��+�-ж���<�LjS�~k:���:I��:�;|�;M*;	�5;�b=;�oB;��E;�IG;\7H;s�H;��H;�H;,�H;��H;��H;��H;��H;��H;��H;��H;t�H;P�H;��H;��H;��H;��H;��H;��H;��H;P�H;t�H;��H;��H;��H;��H;��H;��H;��H;,�H;�H;��H;s�H;\7H;�IG;��E;�oB;�b=;	�5;M*;|�;�;I��:���:~k:LjS���<�-ж��+�]�)�VF��X�      ����o���X��P�ѻf���[ǐ��X��6��
���K�;<":eL�:�`�:�h;Z�%;��3;�<;X/B;��E;�[G;�GH;M�H;��H;a�H;�H;7�H;=�H;��H;�H;�H;��H;��H;��H;]�H;O�H;K�H;'�H;K�H;O�H;]�H;��H;��H;��H;�H;�H;��H;=�H;7�H;�H;a�H;��H;M�H;�GH;�[G;��E;X/B;�<;��3;Z�%;�h;�`�:eL�:;<":�K��
���6��X�[ǐ�f���P�ѻX��o���      ��n��mj���]���J�n�1�L4�l��S���V
x�hX���y�$
9���:գ�:@�;u�#;v�2;�<;�oB;7�E;��G;�dH;��H;8�H;��H;��H;��H;��H;9�H;F�H;7�H;�H;��H;��H;��H;��H;��H;��H;��H;��H;��H;�H;7�H;F�H;9�H;��H;��H;��H;��H;8�H;��H;�dH;��G;7�E;�oB;�<;v�2;u�#;@�;գ�:���:$
9��y�hX�V
x�S���l��L4�n�1���J���]��mj�      B<ͼ��ɼ�����֯�Ҷ��ㄼ��Y�-�*�J���t���X��sѺ�(�K<Q:\��:��
;u�#;��3;�b=;#C;3CF;�G;�H;��H;�H;8�H;��H;W�H;!�H;d�H;��H;b�H;5�H;O�H;	�H;��H;�H;��H;	�H;O�H;5�H;b�H;��H;d�H;!�H;W�H;��H;8�H;�H;��H;�H;�G;3CF;#C;�b=;��3;u�#;��
;\��:K<Q:�(��sѺ�X�t��J���-�*���Y�ㄼҶ���֯�������ɼ      ��'�#�$����y��  ���ۼ����+����]��X!�>ۻ�+��+�i���>:\��:@�;Z�%;	�5;��>;�'D;�F;� H;8�H;[�H;��H;��H;��H;��H;k�H;��H;��H;��H;��H;g�H;K�H;m�H;K�H;g�H;��H;��H;��H;��H;k�H;��H;��H;��H;��H;[�H;8�H;� H;�F;�'D;��>;	�5;Z�%;@�;\��:�>:i��+��+��>ۻ�X!���]��+�������ۼ�  �y����#�$�      �����v����w�]�c��J�Ȅ-�x��;缈沼ㄼ��;�����k��66�i��K<Q:գ�:�h;M*;��8;��@;�OE;�tG;DhH;��H;��H;�H;#�H;��H;y�H;��H;��H;��H;��H;��H;��H;��H;��H;��H;��H;��H;��H;��H;y�H;��H;#�H;�H;��H;��H;DhH;�tG;�OE;��@;��8;M*;�h;գ�:K<Q:i��66�k��������;�ㄼ�沼�;�x�Ȅ-��J�]�c���w��v��      nHͽ̪ɽ�;��"����������[�z0�p��'<ͼо��v�J���k��+��(����:�`�:|�;�/;�K<; C;9lF;��G;�H;
�H;�H;�H;A�H;T�H;��H;%�H;/�H;�H;�H;�H;��H;�H;�H;�H;/�H;%�H;��H;T�H;A�H;�H;�H;
�H;�H;��G;9lF; C;�K<;�/;|�;�`�:���:�(�+�k����v�J�о��'<ͼp��z0���[�������"���;��̪ɽ      ��-�}��|�ű�ƽUP���v���J�D����ۼ��v�J������+���sѺ$
9eL�:�;�$;#�5;�?;��D;j[G;eH;��H;��H;��H;��H;!�H;��H;T�H;n�H;Y�H;T�H;a�H;7�H;a�H;T�H;Y�H;n�H;T�H;��H;!�H;��H;��H;��H;��H;eH;j[G;��D;�?;#�5;�$;�;eL�:$
9�sѺ�+������v�J�����ۼD���J��v��UP��ƽű�|�}��-�       j�Ide�M0X�sD�\{+�z�����k㻽R���JDX������ۼо����;�>ۻ�X���y�;<":I��:��;��-;��;;�B;�yF;�H;��H;|�H;&�H;��H;��H;��H;m�H;��H;��H;��H;��H;z�H;��H;��H;��H;��H;m�H;��H;��H;��H;&�H;|�H;��H;�H;�yF;�B;��;;��-;��;I��:;<":��y��X�>ۻ��;�о����ۼ���JDX�R���k㻽���z��\{+�sD�M0X�Ide�      ��Fh��b���I���|x���O��C(�y�Īɽ����JDX�D��'<ͼㄼ�X!�t��hX��K����:�x;7�#;$H6;IQ@;�OE;��G;��H;��H;1�H;��H;��H;��H;v�H;��H;��H;��H;��H;��H;��H;��H;��H;��H;v�H;��H;��H;��H;1�H;��H;��H;��G;�OE;IQ@;$H6;7�#;�x;���:�K�hX�t���X!�ㄼ'<ͼD��JDX�����Īɽy��C(���O��|x��I��b��Fh��      /�����������;^ɰ��G����i�.�5��	�ĪɽR����J�p���沼��]�J���V
x��
��~k:4��:v;��/;�,=;��C;M�F;#HH;��H;(�H;��H;#�H;��H;��H;��H;�H;�H;�H;$�H;�H;�H;�H;��H;��H;��H;#�H;��H;(�H;��H;#HH;M�F;��C;�,=;��/;v;4��:~k:�
��V
x�J�����]��沼p���J�R���Īɽ�	�.�5���i��G��^ɰ��;��徨���      �2�L�-��"�$E�����4Kɾa��w�s�.�5�y�k㻽�v��z0��;��+��-�*�S����6�LjS� L�:��	;��(;5�9;�.B;�CF;YH;ԪH;��H;��H;��H;w�H;��H;�H;0�H;C�H;<�H;Y�H;<�H;C�H;0�H;�H;��H;w�H;��H;��H;��H;ԪH;YH;�CF;�.B;5�9;��(;��	; L�:LjS��6�S���-�*��+���;�z0��v��k㻽y�.�5�w�s�a��4Kɾ����$E��"�L�-�      3s�cm�/�\�]�C�,�%����TҾa����i��C(����UP����[�x������Y�l���X���<���k:���:)� ;�5;ZQ@;otE;�G;9�H;L�H;��H;�H;I�H;l�H;$�H;c�H;s�H;W�H;��H;W�H;s�H;c�H;$�H;l�H;I�H;�H;��H;L�H;9�H;�G;otE;ZQ@;�5;)� ;���:��k:��<��X�l����Y����x���[�UP����콡C(���i�a���TҾ��,�%�]�C�/�\�cm�      �ޞ�������RF�3�W�M�-���4Kɾ�G����O�z��ƽ����Ȅ-���ۼㄼL4�[ǐ�-ж��Z:n��:�;ʕ1;
c>;{�D;�[G;KrH;��H;i�H;e�H;'�H;u�H;)�H;h�H;��H;|�H;��H;|�H;��H;h�H;)�H;u�H;'�H;e�H;i�H;��H;KrH;�[G;{�D;
c>;ʕ1;�;n��:�Z:-ж�[ǐ�L4�ㄼ��ۼȄ-�����ƽz����O��G��4Kɾ��M�-�3�W�RF�������      ��ſ~��Bw���ޞ�|���3�W�,�%�����^ɰ��|x�\{+�ű����J��  �Ҷ��n�1�f����+�
9q�:�;4�-;��<;��C;�G;�SH;Q�H;��H;��H;��H;V�H;2�H;��H;��H;��H;��H;��H;��H;��H;2�H;V�H;��H;��H;��H;Q�H;�SH;�G;��C;��<;4�-;�;q�:
9�+�f���n�1�Ҷ���  ��J���ű�\{+��|x�^ɰ�����,�%�3�W�|����ޞ�Bw��~��      ������Կp���ޞ�RF�]�C�$E��;�I��sD�|�"��]�c�y��֯���J�P�ѻ]�)���K����:P�
;M*;��:;�C;�F;�7H;Z�H;��H;w�H;��H;>�H;9�H;��H;��H;��H;��H;��H;��H;��H;9�H;>�H;��H;w�H;��H;Z�H;�7H;�F;�C;��:;M*;P�
;���:��K�]�)�P�ѻ��J��֯�y�]�c�"��|�sD��I���;$E�]�C�RF��ޞ�p���Կ��      ������{���ԿBw�����/�\��"����b��M0X�}���;����w����������]�X��VF�2��nȒ:0�;^�';׎9;1oB;�yF;� H;��H;7�H;�H;��H;F�H;:�H;��H;��H;��H;�H;��H;��H;��H;:�H;F�H;��H;�H;7�H;��H;� H;�yF;1oB;׎9;^�';0�;nȒ:2��VF�X�黼�]����������w��;��}��M0X�b������"�/�\����Bw���Կ{�𿖏�      $��������~�����cm�L�-�����Fh��Ide�-�̪ɽ�v��#�$���ɼ�mj�o����X�8��mĆ:�w;i�%;M�8;B;{QF;H;5�H;U�H;�H;p�H;B�H;5�H;��H;��H;��H;$�H;��H;��H;��H;5�H;B�H;p�H;�H;U�H;5�H;H;{QF;B;M�8;i�%;�w;mĆ:8���X�o����mj���ɼ#�$��v��̪ɽ-�Ide�Fh������L�-�cm����~���忖����      �>���8���*�O������˿�o��<�b�=\�+m־^��K�:��J�&��F�B�F���������/��������>:�r�:do ;�I6;DA;�HF;�MH;�H;!I;�I;I;�I;mI;I;q�H;��H;*�H;��H;q�H;I;mI;�I;I;�I;!I;�H;�MH;�HF;DA;�I6;do ;�r�:��>:�����/���������F��F�B�&���J�K�:�^��+m־=\�<�b��o���˿����O���*���8�      ��8��4��g&�0��2����<ƿ벗��>]����G�Ѿ�p���*7����"W��MR?�	}鼀8����s������7�G:���: !;&�6;'kA;�XF;�SH;s�H;!I;�I;�I;�I;FI;�I;e�H;��H;�H;��H;e�H;�I;FI;�I;�I;�I;!I;s�H;�SH;�XF;'kA;&�6; !;���:7�G:���s������8��	}�MR?�"W�����*7��p��G�Ѿ����>]�벗��<ƿ2���0���g&��4�      ��*��g&��#�o�K[�jL�������M�l5��>ľ
����,��D�撐��5�<�ݼ���q
���x��wk�~�b:�j�:#;ږ7;��A;�F;�cH;�I;\!I;I;oI;AI;�I;�I; �H;x�H;��H;x�H; �H;�I;�I;AI;oI;I;\!I;�I;�cH;�F;��A;ږ7;#;�j�:~�b:�wk���x��q
���<�ݼ�5�撐��Dὤ�,�
���>ľl5���M����jL��K[�o��#��g&�      O�0��o����˿:1��-�y���6��z �����)�l�+��ͽ!�����&���˼_�k�q���l�X��� �ϳ�:o�;)&;�9;��B;�F;�|H;�I;e!I;5I;�I;�
I;qI;FI;��H;"�H;��H;"�H;��H;FI;qI;�
I;�I;5I;e!I;�I;�|H;�F;��B;�9;)&;o�;ϳ�:�� �l�X�q���_�k���˼��&�!����ͽ+�)�l������z ���6�-�y�:1���˿���o�0��      ����2���K[忭˿�T��蟉�s�R�����E۾̗����M�~�	������j��3�"d��ɆO���׻c�/��
�����:��	;%*;k;;�iC;�&G;�H;�I;
!I;�I;�I;�	I;�I;� I;I�H;��H;��H;��H;I�H;� I;�I;�	I;�I;�I;
!I;�I;�H;�&G;�iC;k;;%*;��	;���:�
��c�/���׻ɆO�"d���3���j����~�	���M�̗���E۾���s�R�蟉��T���˿K[�2���      �˿�<ƿjL��:1��蟉��>]���)��$���ճ���{���,�j��$��Q`I��J��-��4/�T,��˻ ��!69	3�:�;o.;0-=;o`D;�G;o�H;�I;? I;`I;SI;�I;�I;��H;��H;�H;d�H;�H;��H;��H;�I;�I;SI;`I;? I;�I;o�H;�G;o`D;0-=;o.;�;	3�:�!69˻ �T,��4/�-���J��Q`I�$��j�齞�,���{��ճ��$����)��>]�蟉�:1��jL���<ƿ      �o��벗����-�y�s�R���)�iv��>ľ�]����I�Tl�~��������&�߮Ҽ
�}�VB�"���������!:>)�:Vy;�3;li?;�[E;��G;��H;tI;�I;�I;�I;|I;�I;�H;��H;c�H;��H;c�H;��H;�H;�I;|I;�I;�I;�I;tI;��H;��G;�[E;li?;�3;Vy;>)�:��!:����"���VB�
�}�߮Ҽ��&����~���Tl���I��]���>ľiv���)�s�R�-�y����벗�      <�b��>]���M���6�����$���>ľq��q�Z�+�K9ݽW����L����0F��&�G�\�׻�;�u�Ǌ:�h;5O$;�7;y�A;IF;9BH;��H;�I;mI;wI;I;-I;�I;�H;��H;��H;�H;��H;��H;�H;�I;-I;I;wI;mI;�I;��H;9BH;IF;y�A;�7;5O$;�h;Ǌ:u칹;�\�׻&�G�0F�������L�W��K9ݽ+�q�Z�q���>ľ�$�������6���M��>]�      =\����l5��z ��E۾�ճ��]��q�Z�F?#����A����j�(��Pϼ��������Tnۺj3�9�2�:o�;y�,;��;;C�C;�G;Q�H;�
I;� I;�I;FI;.
I;�I;> I;�H;�H;��H;!�H;��H;�H;�H;> I;�I;.
I;FI;�I;� I;�
I;Q�H;�G;C�C;��;;y�,;o�;�2�:j3�9Tnۺ��������Pϼ(����j��A�����F?#�q�Z��]���ճ��E۾�z �l5����      +m־G�Ѿ�>ľ����̗����{���I�+����V���{�?�/�.���,��c=���һ�@�=� ���k:B�:#a;��3;@i?;v1E;��G;p�H;7I;wI;�I;�I;%I;�I;��H;��H;��H;��H;V�H;��H;��H;��H;��H;�I;%I;�I;�I;wI;7I;p�H;��G;v1E;@i?;��3;#a;B�:��k:=� ��@���һc=��,��.��?�/��{��V�����+���I���{�̗�������>ľG�Ѿ      ^���p��
��)�l���M���,�Tl�K9ݽ�A���{���5��J��;���T[�J?������Q���I�9�:��;9*;4�9;ijB;چF;�MH;��H;I;�I;�I;!I;I;@I;^�H;��H;��H;��H;i�H;��H;��H;��H;^�H;@I;I;!I;�I;�I;I;��H;�MH;چF;ijB;4�9;9*;��;�:�I�9�Q������J?��T[�;���J����5��{��A��K9ݽTl���,���M�)�l�
���p��      K�:��*7���,�+�~�	�j��~���W����j�?�/��J���I��&�k���c.������:Ǌ:�m�:';mq3;1�>;8�D;t�G;R�H;I;. I;�I;�I;�	I;�I;`�H;��H;��H;��H;��H;^�H;��H;��H;��H;��H;`�H;�I;�	I;�I;�I;. I;I;R�H;t�G;8�D;1�>;mq3;';�m�::Ǌ:����c.����&�k��I���J��?�/���j�W��~���j��~�	�+���,��*7�      �J���D��ͽ���$�������L�(��.��;��&�k����I����/��"/�(�>:���:�A;v�,;��:;=�B;�wF;�;H;��H;	I;�I;�I;AI;�I;�I;��H;s�H;4�H;n�H;��H;l�H;��H;n�H;4�H;s�H;��H;�I;�I;AI;�I;�I;	I;��H;�;H;�wF;=�B;��:;v�,;�A;���:(�>:�"/���/��I����&�k�;��.��(����L����$������ͽ�Dὼ��      &��"W��撐�!�����j�Q`I���&����Pϼ�,���T[����I��;��qk�j:h3�:� ; &;�6;� @;C1E;�G;��H;�I;�I;OI;I;�	I;:I;t�H;��H;�H;��H;^�H;��H;D�H;��H;^�H;��H;�H;��H;t�H;:I;�	I;I;OI;�I;�I;��H;�G;C1E;� @;�6; &;� ;h3�:j:�qk�;��I�����T[��,��Pϼ�����&�Q`I���j�!���撐�"W��      F�B�MR?��5���&��3��J��߮Ҽ0F����c=�J?�c.����/��qk����9�ճ:�;J!;l3;��=;��C;*�F;cH;��H;�I;I;�I;$I;�I;�I;C�H;��H;��H;|�H;?�H;|�H;3�H;|�H;?�H;|�H;��H;��H;C�H;�I;�I;$I;�I;I;�I;��H;cH;*�F;��C;��=;l3;J!;�;�ճ:���9�qk���/�c.��J?�c=���0F��߮Ҽ�J���3���&��5�MR?�      F��	}�<�ݼ��˼"d��-��
�}�&�G������һ�������"/�j:�ճ:"�;�a;â0;�<;��B;�HF;uH;,�H;�I;yI;I;8I;Y	I;�I;�H;/�H;T�H;�H;#�H;�H;r�H;5�H;r�H;�H;#�H;�H;T�H;/�H;�H;�I;Y	I;8I;I;yI;�I;,�H;uH;�HF;��B;�<;â0;�a;"�;�ճ:j:�"/���������һ���&�G�
�}�-��"d����˼<�ݼ	}�      �����8����_�k�ɆO�4/�VB�\�׻����@��Q����(�>:h3�:�;�a;��/;=;;J�A;��E;ɾG;��H;�	I;gI;I;�I;�I;�I;� I;��H;;�H;��H;��H;��H;�H;c�H;)�H;c�H;�H;��H;��H;��H;;�H;��H;� I;�I;�I;�I;I;gI;�	I;��H;ɾG;��E;J�A;=;;��/;�a;�;h3�:(�>:���Q���@����\�׻VB�4/�ɆO�_�k����8��      ������q
�q�����׻T,��"����;�Tnۺ=� ��I�9:Ǌ:���:� ;J!;â0;=;;̒A;�oE;|�G;ӍH;��H;�I;9I;ZI; I;�I;oI;��H;=�H;x�H;�H;�H;��H;��H;[�H;1�H;[�H;��H;��H;�H;�H;x�H;=�H;��H;oI;�I; I;ZI;9I;�I;��H;ӍH;|�G;�oE;̒A;=;;â0;J!;� ;���::Ǌ:�I�9=� �Tnۺ�;�"���T,����׻q����q
���      �/��s�����x�l�X�c�/�˻ �����u�j3�9��k:�:�m�:�A; &;l3;�<;J�A;�oE;hsG;�{H;-�H;,I;rI;CI;�I;i	I;�I;L�H;I�H;�H;��H;x�H;��H;��H;��H;l�H;\�H;l�H;��H;��H;��H;x�H;��H;�H;I�H;L�H;�I;i	I;�I;CI;rI;,I;-�H;�{H;hsG;�oE;J�A;�<;l3; &;�A;�m�:�:��k:j3�9u칋���˻ �c�/�l�X���x�s���      ��������wk��� ��
���!69��!:Ǌ:�2�:B�:��;';v�,;�6;��=;��B;��E;|�G;�{H;��H;zI;I;�I;WI;�
I;"I;� I;A�H;��H;4�H;��H;�H;��H;��H;��H;}�H;k�H;}�H;��H;��H;��H;�H;��H;4�H;��H;A�H;� I;"I;�
I;WI;�I;I;zI;��H;�{H;|�G;��E;��B;��=;�6;v�,;';��;B�:�2�:Ǌ:��!:�!69�
���� ��wk����      ��>:7�G:~�b:ϳ�:���:	3�:>)�:�h;o�;#a;9*;mq3;��:;� @;��C;�HF;ɾG;ӍH;-�H;zI;I;BI;9I;�I;I;VI;�H;��H;��H;o�H;B�H;��H;��H;��H;	�H;��H;y�H;��H;	�H;��H;��H;��H;B�H;o�H;��H;��H;�H;VI;I;�I;9I;BI;I;zI;-�H;ӍH;ɾG;�HF;��C;� @;��:;mq3;9*;#a;o�;�h;>)�:	3�:���:ϳ�:~�b:7�G:      �r�:���:�j�:o�;��	;�;Vy;5O$;y�,;��3;4�9;1�>;=�B;C1E;*�F;uH;��H;��H;,I;I;BI;�I;6I;�I;�I;��H;�H;F�H;��H;��H;��H;��H;��H;��H;)�H;��H;��H;��H;)�H;��H;��H;��H;��H;��H;��H;F�H;�H;��H;�I;�I;6I;�I;BI;I;,I;��H;��H;uH;*�F;C1E;=�B;1�>;4�9;��3;y�,;5O$;Vy;�;��	;o�;�j�:���:      do ; !;#;)&;%*;o.;�3;�7;��;;@i?;ijB;8�D;�wF;�G;cH;,�H;�	I;�I;rI;�I;9I;6I;�I;QI;4�H;��H;��H; �H;��H;�H;��H;x�H;��H;��H;E�H;�H;��H;�H;E�H;��H;��H;x�H;��H;�H;��H; �H;��H;��H;4�H;QI;�I;6I;9I;�I;rI;�I;�	I;,�H;cH;�G;�wF;8�D;ijB;@i?;��;;�7;�3;o.;%*;)&;#; !;      �I6;&�6;ږ7;�9;k;;0-=;li?;y�A;C�C;v1E;چF;t�G;�;H;��H;��H;�I;gI;9I;CI;WI;�I;�I;QI;E�H;��H;��H;Y�H;$�H;0�H;��H;~�H;e�H;��H;�H;��H;]�H;:�H;]�H;��H;�H;��H;e�H;~�H;��H;0�H;$�H;Y�H;��H;��H;E�H;QI;�I;�I;WI;CI;9I;gI;�I;��H;��H;�;H;t�G;چF;v1E;C�C;y�A;li?;0-=;k;;�9;ږ7;&�6;      DA;'kA;��A;��B;�iC;o`D;�[E;IF;�G;��G;�MH;R�H;��H;�I;�I;yI;I;ZI;�I;�
I;I;�I;4�H;��H;��H;w�H;-�H;@�H;��H;��H;`�H;u�H;��H;O�H;��H;��H;��H;��H;��H;O�H;��H;u�H;`�H;��H;��H;@�H;-�H;w�H;��H;��H;4�H;�I;I;�
I;�I;ZI;I;yI;�I;�I;��H;R�H;�MH;��G;�G;IF;�[E;o`D;�iC;��B;��A;'kA;      �HF;�XF;�F;�F;�&G;�G;��G;9BH;Q�H;p�H;��H;I;	I;�I;I;I;�I; I;i	I;"I;VI;��H;��H;��H;w�H;S�H;Z�H;��H;��H;i�H;X�H;��H;&�H;��H;@�H;"�H;�H;"�H;@�H;��H;&�H;��H;X�H;i�H;��H;��H;Z�H;S�H;w�H;��H;��H;��H;VI;"I;i	I; I;�I;I;I;�I;	I;I;��H;p�H;Q�H;9BH;��G;�G;�&G;�F;�F;�XF;      �MH;�SH;�cH;�|H;�H;o�H;��H;��H;�
I;7I;I;. I;�I;OI;�I;8I;�I;�I;�I;� I;�H;�H;��H;Y�H;-�H;Z�H;��H;��H;X�H;Z�H;��H;��H;d�H;��H;��H;��H;��H;��H;��H;��H;d�H;��H;��H;Z�H;X�H;��H;��H;Z�H;-�H;Y�H;��H;�H;�H;� I;�I;�I;�I;8I;�I;OI;�I;. I;I;7I;�
I;��H;��H;o�H;�H;�|H;�cH;�SH;      �H;s�H;�I;�I;�I;�I;tI;�I;� I;wI;�I;�I;�I;I;$I;Y	I;�I;oI;L�H;A�H;��H;F�H; �H;$�H;@�H;��H;��H;k�H;O�H;��H;��H;;�H;��H;{�H;9�H;
�H;�H;
�H;9�H;{�H;��H;;�H;��H;��H;O�H;k�H;��H;��H;@�H;$�H; �H;F�H;��H;A�H;L�H;oI;�I;Y	I;$I;I;�I;�I;�I;wI;� I;�I;tI;�I;�I;�I;�I;s�H;      !I;!I;\!I;e!I;
!I;? I;�I;mI;�I;�I;�I;�I;AI;�	I;�I;�I;� I;��H;I�H;��H;��H;��H;��H;0�H;��H;��H;X�H;O�H;��H;��H;/�H;��H;M�H;��H;��H;��H;��H;��H;��H;��H;M�H;��H;/�H;��H;��H;O�H;X�H;��H;��H;0�H;��H;��H;��H;��H;I�H;��H;� I;�I;�I;�	I;AI;�I;�I;�I;�I;mI;�I;? I;
!I;e!I;\!I;!I;      �I;�I;I;5I;�I;`I;�I;wI;FI;�I;!I;�	I;�I;:I;�I;�H;��H;=�H;�H;4�H;o�H;��H;�H;��H;��H;i�H;Z�H;��H;��H;�H;��H;C�H;��H;��H;f�H;J�H;9�H;J�H;f�H;��H;��H;C�H;��H;�H;��H;��H;Z�H;i�H;��H;��H;�H;��H;o�H;4�H;�H;=�H;��H;�H;�I;:I;�I;�	I;!I;�I;FI;wI;�I;`I;�I;5I;I;�I;      I;�I;oI;�I;�I;SI;�I;I;.
I;%I;I;�I;�I;t�H;C�H;/�H;;�H;x�H;��H;��H;B�H;��H;��H;~�H;`�H;X�H;��H;��H;/�H;��H;'�H;��H;v�H;<�H;	�H;��H;��H;��H;	�H;<�H;v�H;��H;'�H;��H;/�H;��H;��H;X�H;`�H;~�H;��H;��H;B�H;��H;��H;x�H;;�H;/�H;C�H;t�H;�I;�I;I;%I;.
I;I;�I;SI;�I;�I;oI;�I;      �I;�I;AI;�
I;�	I;�I;|I;-I;�I;�I;@I;`�H;��H;��H;��H;T�H;��H;�H;x�H;�H;��H;��H;x�H;e�H;u�H;��H;��H;;�H;��H;C�H;��H;R�H;!�H;��H;��H;��H;��H;��H;��H;��H;!�H;R�H;��H;C�H;��H;;�H;��H;��H;u�H;e�H;x�H;��H;��H;�H;x�H;�H;��H;T�H;��H;��H;��H;`�H;@I;�I;�I;-I;|I;�I;�	I;�
I;AI;�I;      mI;FI;�I;qI;�I;�I;�I;�I;> I;��H;^�H;��H;s�H;�H;��H;�H;��H;�H;��H;��H;��H;��H;��H;��H;��H;&�H;d�H;��H;M�H;��H;v�H;!�H;��H;��H;��H;m�H;f�H;m�H;��H;��H;��H;!�H;v�H;��H;M�H;��H;d�H;&�H;��H;��H;��H;��H;��H;��H;��H;�H;��H;�H;��H;�H;s�H;��H;^�H;��H;> I;�I;�I;�I;�I;qI;�I;FI;      I;�I;�I;FI;� I;��H;�H;�H;�H;��H;��H;��H;4�H;��H;|�H;#�H;��H;��H;��H;��H;��H;��H;��H;�H;O�H;��H;��H;{�H;��H;��H;<�H;��H;��H;n�H;V�H;J�H;9�H;J�H;V�H;n�H;��H;��H;<�H;��H;��H;{�H;��H;��H;O�H;�H;��H;��H;��H;��H;��H;��H;��H;#�H;|�H;��H;4�H;��H;��H;��H;�H;�H;�H;��H;� I;FI;�I;�I;      q�H;e�H; �H;��H;I�H;��H;��H;��H;�H;��H;��H;��H;n�H;^�H;?�H;�H;�H;��H;��H;��H;	�H;)�H;E�H;��H;��H;@�H;��H;9�H;��H;f�H;	�H;��H;��H;V�H;1�H;&�H;(�H;&�H;1�H;V�H;��H;��H;	�H;f�H;��H;9�H;��H;@�H;��H;��H;E�H;)�H;	�H;��H;��H;��H;�H;�H;?�H;^�H;n�H;��H;��H;��H;�H;��H;��H;��H;I�H;��H; �H;e�H;      ��H;��H;x�H;"�H;��H;�H;c�H;��H;��H;��H;��H;��H;��H;��H;|�H;r�H;c�H;[�H;l�H;}�H;��H;��H;�H;]�H;��H;"�H;��H;
�H;��H;J�H;��H;��H;m�H;J�H;&�H;
�H;�H;
�H;&�H;J�H;m�H;��H;��H;J�H;��H;
�H;��H;"�H;��H;]�H;�H;��H;��H;}�H;l�H;[�H;c�H;r�H;|�H;��H;��H;��H;��H;��H;��H;��H;c�H;�H;��H;"�H;x�H;��H;      *�H;�H;��H;��H;��H;d�H;��H;�H;!�H;V�H;i�H;^�H;l�H;D�H;3�H;5�H;)�H;1�H;\�H;k�H;y�H;��H;��H;:�H;��H;�H;��H;�H;��H;9�H;��H;��H;f�H;9�H;(�H;�H;�H;�H;(�H;9�H;f�H;��H;��H;9�H;��H;�H;��H;�H;��H;:�H;��H;��H;y�H;k�H;\�H;1�H;)�H;5�H;3�H;D�H;l�H;^�H;i�H;V�H;!�H;�H;��H;d�H;��H;��H;��H;�H;      ��H;��H;x�H;"�H;��H;�H;c�H;��H;��H;��H;��H;��H;��H;��H;|�H;r�H;c�H;[�H;l�H;}�H;��H;��H;�H;]�H;��H;"�H;��H;
�H;��H;J�H;��H;��H;m�H;J�H;&�H;
�H;�H;
�H;&�H;J�H;m�H;��H;��H;J�H;��H;
�H;��H;"�H;��H;]�H;�H;��H;��H;}�H;l�H;[�H;c�H;r�H;|�H;��H;��H;��H;��H;��H;��H;��H;c�H;�H;��H;"�H;x�H;��H;      q�H;e�H; �H;��H;I�H;��H;��H;��H;�H;��H;��H;��H;n�H;^�H;?�H;�H;�H;��H;��H;��H;	�H;)�H;E�H;��H;��H;@�H;��H;9�H;��H;f�H;	�H;��H;��H;V�H;1�H;&�H;(�H;&�H;1�H;V�H;��H;��H;	�H;f�H;��H;9�H;��H;@�H;��H;��H;E�H;)�H;	�H;��H;��H;��H;�H;�H;?�H;^�H;n�H;��H;��H;��H;�H;��H;��H;��H;I�H;��H; �H;e�H;      I;�I;�I;FI;� I;��H;�H;�H;�H;��H;��H;��H;4�H;��H;|�H;#�H;��H;��H;��H;��H;��H;��H;��H;�H;O�H;��H;��H;{�H;��H;��H;<�H;��H;��H;n�H;V�H;J�H;9�H;J�H;V�H;n�H;��H;��H;<�H;��H;��H;{�H;��H;��H;O�H;�H;��H;��H;��H;��H;��H;��H;��H;#�H;|�H;��H;4�H;��H;��H;��H;�H;�H;�H;��H;� I;FI;�I;�I;      mI;FI;�I;qI;�I;�I;�I;�I;> I;��H;^�H;��H;s�H;�H;��H;�H;��H;�H;��H;��H;��H;��H;��H;��H;��H;&�H;d�H;��H;M�H;��H;v�H;!�H;��H;��H;��H;m�H;f�H;m�H;��H;��H;��H;!�H;v�H;��H;M�H;��H;d�H;&�H;��H;��H;��H;��H;��H;��H;��H;�H;��H;�H;��H;�H;s�H;��H;^�H;��H;> I;�I;�I;�I;�I;qI;�I;FI;      �I;�I;AI;�
I;�	I;�I;|I;-I;�I;�I;@I;`�H;��H;��H;��H;T�H;��H;�H;x�H;�H;��H;��H;x�H;e�H;u�H;��H;��H;;�H;��H;C�H;��H;R�H;!�H;��H;��H;��H;��H;��H;��H;��H;!�H;R�H;��H;C�H;��H;;�H;��H;��H;u�H;e�H;x�H;��H;��H;�H;x�H;�H;��H;T�H;��H;��H;��H;`�H;@I;�I;�I;-I;|I;�I;�	I;�
I;AI;�I;      I;�I;oI;�I;�I;SI;�I;I;.
I;%I;I;�I;�I;t�H;C�H;/�H;;�H;x�H;��H;��H;B�H;��H;��H;~�H;`�H;X�H;��H;��H;/�H;��H;'�H;��H;v�H;<�H;	�H;��H;��H;��H;	�H;<�H;v�H;��H;'�H;��H;/�H;��H;��H;X�H;`�H;~�H;��H;��H;B�H;��H;��H;x�H;;�H;/�H;C�H;t�H;�I;�I;I;%I;.
I;I;�I;SI;�I;�I;oI;�I;      �I;�I;I;5I;�I;`I;�I;wI;FI;�I;!I;�	I;�I;:I;�I;�H;��H;=�H;�H;4�H;o�H;��H;�H;��H;��H;i�H;Z�H;��H;��H;�H;��H;C�H;��H;��H;f�H;J�H;9�H;J�H;f�H;��H;��H;C�H;��H;�H;��H;��H;Z�H;i�H;��H;��H;�H;��H;o�H;4�H;�H;=�H;��H;�H;�I;:I;�I;�	I;!I;�I;FI;wI;�I;`I;�I;5I;I;�I;      !I;!I;\!I;e!I;
!I;? I;�I;mI;�I;�I;�I;�I;AI;�	I;�I;�I;� I;��H;I�H;��H;��H;��H;��H;0�H;��H;��H;X�H;O�H;��H;��H;/�H;��H;M�H;��H;��H;��H;��H;��H;��H;��H;M�H;��H;/�H;��H;��H;O�H;X�H;��H;��H;0�H;��H;��H;��H;��H;I�H;��H;� I;�I;�I;�	I;AI;�I;�I;�I;�I;mI;�I;? I;
!I;e!I;\!I;!I;      �H;s�H;�I;�I;�I;�I;tI;�I;� I;wI;�I;�I;�I;I;$I;Y	I;�I;oI;L�H;A�H;��H;F�H; �H;$�H;@�H;��H;��H;k�H;O�H;��H;��H;;�H;��H;{�H;9�H;
�H;�H;
�H;9�H;{�H;��H;;�H;��H;��H;O�H;k�H;��H;��H;@�H;$�H; �H;F�H;��H;A�H;L�H;oI;�I;Y	I;$I;I;�I;�I;�I;wI;� I;�I;tI;�I;�I;�I;�I;s�H;      �MH;�SH;�cH;�|H;�H;o�H;��H;��H;�
I;7I;I;. I;�I;OI;�I;8I;�I;�I;�I;� I;�H;�H;��H;Y�H;-�H;Z�H;��H;��H;X�H;Z�H;��H;��H;d�H;��H;��H;��H;��H;��H;��H;��H;d�H;��H;��H;Z�H;X�H;��H;��H;Z�H;-�H;Y�H;��H;�H;�H;� I;�I;�I;�I;8I;�I;OI;�I;. I;I;7I;�
I;��H;��H;o�H;�H;�|H;�cH;�SH;      �HF;�XF;�F;�F;�&G;�G;��G;9BH;Q�H;p�H;��H;I;	I;�I;I;I;�I; I;i	I;"I;VI;��H;��H;��H;w�H;S�H;Z�H;��H;��H;i�H;X�H;��H;&�H;��H;@�H;"�H;�H;"�H;@�H;��H;&�H;��H;X�H;i�H;��H;��H;Z�H;S�H;w�H;��H;��H;��H;VI;"I;i	I; I;�I;I;I;�I;	I;I;��H;p�H;Q�H;9BH;��G;�G;�&G;�F;�F;�XF;      DA;'kA;��A;��B;�iC;o`D;�[E;IF;�G;��G;�MH;R�H;��H;�I;�I;yI;I;ZI;�I;�
I;I;�I;4�H;��H;��H;w�H;-�H;@�H;��H;��H;`�H;u�H;��H;O�H;��H;��H;��H;��H;��H;O�H;��H;u�H;`�H;��H;��H;@�H;-�H;w�H;��H;��H;4�H;�I;I;�
I;�I;ZI;I;yI;�I;�I;��H;R�H;�MH;��G;�G;IF;�[E;o`D;�iC;��B;��A;'kA;      �I6;&�6;ږ7;�9;k;;0-=;li?;y�A;C�C;v1E;چF;t�G;�;H;��H;��H;�I;gI;9I;CI;WI;�I;�I;QI;E�H;��H;��H;Y�H;$�H;0�H;��H;~�H;e�H;��H;�H;��H;]�H;:�H;]�H;��H;�H;��H;e�H;~�H;��H;0�H;$�H;Y�H;��H;��H;E�H;QI;�I;�I;WI;CI;9I;gI;�I;��H;��H;�;H;t�G;چF;v1E;C�C;y�A;li?;0-=;k;;�9;ږ7;&�6;      do ; !;#;)&;%*;o.;�3;�7;��;;@i?;ijB;8�D;�wF;�G;cH;,�H;�	I;�I;rI;�I;9I;6I;�I;QI;4�H;��H;��H; �H;��H;�H;��H;x�H;��H;��H;E�H;�H;��H;�H;E�H;��H;��H;x�H;��H;�H;��H; �H;��H;��H;4�H;QI;�I;6I;9I;�I;rI;�I;�	I;,�H;cH;�G;�wF;8�D;ijB;@i?;��;;�7;�3;o.;%*;)&;#; !;      �r�:���:�j�:o�;��	;�;Vy;5O$;y�,;��3;4�9;1�>;=�B;C1E;*�F;uH;��H;��H;,I;I;BI;�I;6I;�I;�I;��H;�H;F�H;��H;��H;��H;��H;��H;��H;)�H;��H;��H;��H;)�H;��H;��H;��H;��H;��H;��H;F�H;�H;��H;�I;�I;6I;�I;BI;I;,I;��H;��H;uH;*�F;C1E;=�B;1�>;4�9;��3;y�,;5O$;Vy;�;��	;o�;�j�:���:      ��>:7�G:~�b:ϳ�:���:	3�:>)�:�h;o�;#a;9*;mq3;��:;� @;��C;�HF;ɾG;ӍH;-�H;zI;I;BI;9I;�I;I;VI;�H;��H;��H;o�H;B�H;��H;��H;��H;	�H;��H;y�H;��H;	�H;��H;��H;��H;B�H;o�H;��H;��H;�H;VI;I;�I;9I;BI;I;zI;-�H;ӍH;ɾG;�HF;��C;� @;��:;mq3;9*;#a;o�;�h;>)�:	3�:���:ϳ�:~�b:7�G:      ��������wk��� ��
���!69��!:Ǌ:�2�:B�:��;';v�,;�6;��=;��B;��E;|�G;�{H;��H;zI;I;�I;WI;�
I;"I;� I;A�H;��H;4�H;��H;�H;��H;��H;��H;}�H;k�H;}�H;��H;��H;��H;�H;��H;4�H;��H;A�H;� I;"I;�
I;WI;�I;I;zI;��H;�{H;|�G;��E;��B;��=;�6;v�,;';��;B�:�2�:Ǌ:��!:�!69�
���� ��wk����      �/��s�����x�l�X�c�/�˻ �����u�j3�9��k:�:�m�:�A; &;l3;�<;J�A;�oE;hsG;�{H;-�H;,I;rI;CI;�I;i	I;�I;L�H;I�H;�H;��H;x�H;��H;��H;��H;l�H;\�H;l�H;��H;��H;��H;x�H;��H;�H;I�H;L�H;�I;i	I;�I;CI;rI;,I;-�H;�{H;hsG;�oE;J�A;�<;l3; &;�A;�m�:�:��k:j3�9u칋���˻ �c�/�l�X���x�s���      ������q
�q�����׻T,��"����;�Tnۺ=� ��I�9:Ǌ:���:� ;J!;â0;=;;̒A;�oE;|�G;ӍH;��H;�I;9I;ZI; I;�I;oI;��H;=�H;x�H;�H;�H;��H;��H;[�H;1�H;[�H;��H;��H;�H;�H;x�H;=�H;��H;oI;�I; I;ZI;9I;�I;��H;ӍH;|�G;�oE;̒A;=;;â0;J!;� ;���::Ǌ:�I�9=� �Tnۺ�;�"���T,����׻q����q
���      �����8����_�k�ɆO�4/�VB�\�׻����@��Q����(�>:h3�:�;�a;��/;=;;J�A;��E;ɾG;��H;�	I;gI;I;�I;�I;�I;� I;��H;;�H;��H;��H;��H;�H;c�H;)�H;c�H;�H;��H;��H;��H;;�H;��H;� I;�I;�I;�I;I;gI;�	I;��H;ɾG;��E;J�A;=;;��/;�a;�;h3�:(�>:���Q���@����\�׻VB�4/�ɆO�_�k����8��      F��	}�<�ݼ��˼"d��-��
�}�&�G������һ�������"/�j:�ճ:"�;�a;â0;�<;��B;�HF;uH;,�H;�I;yI;I;8I;Y	I;�I;�H;/�H;T�H;�H;#�H;�H;r�H;5�H;r�H;�H;#�H;�H;T�H;/�H;�H;�I;Y	I;8I;I;yI;�I;,�H;uH;�HF;��B;�<;â0;�a;"�;�ճ:j:�"/���������һ���&�G�
�}�-��"d����˼<�ݼ	}�      F�B�MR?��5���&��3��J��߮Ҽ0F����c=�J?�c.����/��qk����9�ճ:�;J!;l3;��=;��C;*�F;cH;��H;�I;I;�I;$I;�I;�I;C�H;��H;��H;|�H;?�H;|�H;3�H;|�H;?�H;|�H;��H;��H;C�H;�I;�I;$I;�I;I;�I;��H;cH;*�F;��C;��=;l3;J!;�;�ճ:���9�qk���/�c.��J?�c=���0F��߮Ҽ�J���3���&��5�MR?�      &��"W��撐�!�����j�Q`I���&����Pϼ�,���T[����I��;��qk�j:h3�:� ; &;�6;� @;C1E;�G;��H;�I;�I;OI;I;�	I;:I;t�H;��H;�H;��H;^�H;��H;D�H;��H;^�H;��H;�H;��H;t�H;:I;�	I;I;OI;�I;�I;��H;�G;C1E;� @;�6; &;� ;h3�:j:�qk�;��I�����T[��,��Pϼ�����&�Q`I���j�!���撐�"W��      �J���D��ͽ���$�������L�(��.��;��&�k����I����/��"/�(�>:���:�A;v�,;��:;=�B;�wF;�;H;��H;	I;�I;�I;AI;�I;�I;��H;s�H;4�H;n�H;��H;l�H;��H;n�H;4�H;s�H;��H;�I;�I;AI;�I;�I;	I;��H;�;H;�wF;=�B;��:;v�,;�A;���:(�>:�"/���/��I����&�k�;��.��(����L����$������ͽ�Dὼ��      K�:��*7���,�+�~�	�j��~���W����j�?�/��J���I��&�k���c.������:Ǌ:�m�:';mq3;1�>;8�D;t�G;R�H;I;. I;�I;�I;�	I;�I;`�H;��H;��H;��H;��H;^�H;��H;��H;��H;��H;`�H;�I;�	I;�I;�I;. I;I;R�H;t�G;8�D;1�>;mq3;';�m�::Ǌ:����c.����&�k��I���J��?�/���j�W��~���j��~�	�+���,��*7�      ^���p��
��)�l���M���,�Tl�K9ݽ�A���{���5��J��;���T[�J?������Q���I�9�:��;9*;4�9;ijB;چF;�MH;��H;I;�I;�I;!I;I;@I;^�H;��H;��H;��H;i�H;��H;��H;��H;^�H;@I;I;!I;�I;�I;I;��H;�MH;چF;ijB;4�9;9*;��;�:�I�9�Q������J?��T[�;���J����5��{��A��K9ݽTl���,���M�)�l�
���p��      +m־G�Ѿ�>ľ����̗����{���I�+����V���{�?�/�.���,��c=���һ�@�=� ���k:B�:#a;��3;@i?;v1E;��G;p�H;7I;wI;�I;�I;%I;�I;��H;��H;��H;��H;V�H;��H;��H;��H;��H;�I;%I;�I;�I;wI;7I;p�H;��G;v1E;@i?;��3;#a;B�:��k:=� ��@���һc=��,��.��?�/��{��V�����+���I���{�̗�������>ľG�Ѿ      =\����l5��z ��E۾�ճ��]��q�Z�F?#����A����j�(��Pϼ��������Tnۺj3�9�2�:o�;y�,;��;;C�C;�G;Q�H;�
I;� I;�I;FI;.
I;�I;> I;�H;�H;��H;!�H;��H;�H;�H;> I;�I;.
I;FI;�I;� I;�
I;Q�H;�G;C�C;��;;y�,;o�;�2�:j3�9Tnۺ��������Pϼ(����j��A�����F?#�q�Z��]���ճ��E۾�z �l5����      <�b��>]���M���6�����$���>ľq��q�Z�+�K9ݽW����L����0F��&�G�\�׻�;�u�Ǌ:�h;5O$;�7;y�A;IF;9BH;��H;�I;mI;wI;I;-I;�I;�H;��H;��H;�H;��H;��H;�H;�I;-I;I;wI;mI;�I;��H;9BH;IF;y�A;�7;5O$;�h;Ǌ:u칹;�\�׻&�G�0F�������L�W��K9ݽ+�q�Z�q���>ľ�$�������6���M��>]�      �o��벗����-�y�s�R���)�iv��>ľ�]����I�Tl�~��������&�߮Ҽ
�}�VB�"���������!:>)�:Vy;�3;li?;�[E;��G;��H;tI;�I;�I;�I;|I;�I;�H;��H;c�H;��H;c�H;��H;�H;�I;|I;�I;�I;�I;tI;��H;��G;�[E;li?;�3;Vy;>)�:��!:����"���VB�
�}�߮Ҽ��&����~���Tl���I��]���>ľiv���)�s�R�-�y����벗�      �˿�<ƿjL��:1��蟉��>]���)��$���ճ���{���,�j��$��Q`I��J��-��4/�T,��˻ ��!69	3�:�;o.;0-=;o`D;�G;o�H;�I;? I;`I;SI;�I;�I;��H;��H;�H;d�H;�H;��H;��H;�I;�I;SI;`I;? I;�I;o�H;�G;o`D;0-=;o.;�;	3�:�!69˻ �T,��4/�-���J��Q`I�$��j�齞�,���{��ճ��$����)��>]�蟉�:1��jL���<ƿ      ����2���K[忭˿�T��蟉�s�R�����E۾̗����M�~�	������j��3�"d��ɆO���׻c�/��
�����:��	;%*;k;;�iC;�&G;�H;�I;
!I;�I;�I;�	I;�I;� I;I�H;��H;��H;��H;I�H;� I;�I;�	I;�I;�I;
!I;�I;�H;�&G;�iC;k;;%*;��	;���:�
��c�/���׻ɆO�"d���3���j����~�	���M�̗���E۾���s�R�蟉��T���˿K[�2���      O�0��o����˿:1��-�y���6��z �����)�l�+��ͽ!�����&���˼_�k�q���l�X��� �ϳ�:o�;)&;�9;��B;�F;�|H;�I;e!I;5I;�I;�
I;qI;FI;��H;"�H;��H;"�H;��H;FI;qI;�
I;�I;5I;e!I;�I;�|H;�F;��B;�9;)&;o�;ϳ�:�� �l�X�q���_�k���˼��&�!����ͽ+�)�l������z ���6�-�y�:1���˿���o�0��      ��*��g&��#�o�K[�jL�������M�l5��>ľ
����,��D�撐��5�<�ݼ���q
���x��wk�~�b:�j�:#;ږ7;��A;�F;�cH;�I;\!I;I;oI;AI;�I;�I; �H;x�H;��H;x�H; �H;�I;�I;AI;oI;I;\!I;�I;�cH;�F;��A;ږ7;#;�j�:~�b:�wk���x��q
���<�ݼ�5�撐��Dὤ�,�
���>ľl5���M����jL��K[�o��#��g&�      ��8��4��g&�0��2����<ƿ벗��>]����G�Ѿ�p���*7����"W��MR?�	}鼀8����s������7�G:���: !;&�6;'kA;�XF;�SH;s�H;!I;�I;�I;�I;FI;�I;e�H;��H;�H;��H;e�H;�I;FI;�I;�I;�I;!I;s�H;�SH;�XF;'kA;&�6; !;���:7�G:���s������8��	}�MR?�"W�����*7��p��G�Ѿ����>]�벗��<ƿ2���0���g&��4�      �Aq���i���U�A:�@�����6���q���uA�a5�� ��y^Z�����A���]�����d��|",�6��:�Ѻ���9'��:d�;dX4;p�@;�UF;��H;�FI;�aI;2NI;A9I;�(I;<I;�I;�I;�I;�
I;�I;�I;�I;<I;�(I;A9I;2NI;�aI;�FI;��H;�UF;p�@;dX4;d�;'��:���9:�Ѻ6��|",��d������]��A�����y^Z�� ��a5�uA�q���6�������@�A:���U���i�      ��i���b�T�O�.5�-i������������q<�����e��[
V�FE	�!���IY�s9�Z����(� S����Ⱥ��:���:'�;K�4;h�@;kgF;��H;4HI;�aI;�MI;�8I;�(I;I;~I;�I;{I;x
I;{I;�I;~I;I;�(I;�8I;�MI;�aI;4HI;��H;kgF;h�@;K�4;'�;���:��:��Ⱥ S���(�Z���s9��IY�!��FE	�[
V��e������q<������������-i�.5�T�O���b�      ��U�T�O�B-?�(�'���F�`欿Y�{�aa/���뾙���I����e���ZN�o5��Ǩ��nH�� ������ܧ":��:��;��5;�_A;ٚF;Z�H;;LI;aI;�LI;�7I;(I;aI;I;_I;&I;&
I;&I;_I;I;aI;(I;�7I;�LI;aI;;LI;Z�H;ٚF;�_A;��5;��;��:ܧ":����� ��nH�Ǩ��o5���ZN�e������I�������aa/�Y�{��欿F����(�'�B-?�T�O�      A:�.5�(�'��������dȿ���e$_���Q�Ҿؕ��
�6�����*���`=�P���)��{G��6��B����Q:�:/";�7;�%B;�F;��H;RI;�_I;�JI;C6I;�&I;ZI;7I;�I;�
I;�	I;�
I;�I;7I;ZI;�&I;C6I;�JI;�_I;RI;��H;�F;�%B;�7;/";�:��Q:B���6��{G��)��P���`=��*�����
�6�ؕ��Q�Ҿ��e$_����dȿ�������(�'�.5�      @�-i�������B�ѿf�������q<��:��a����q����Wн齅���'�ib̼�zl�/���X�{���:��;
�&;٪9;KC;vLG;�H;]XI;�]I;�GI;4I;�$I;I;'I;�I;�	I;�I;�	I;�I;'I;I;�$I;4I;�GI;�]I;]XI;�H;vLG;KC;٪9;
�&;��;�:{���X�/���zl�ib̼��'�齅��Wн����q��a���:��q<����f���B�ѿ������-i�      �������F��dȿf���������O���u]׾w���	�I�����A��C�d�v��֮�<RH�Kkλ �$�x5����:mM;˅+;�<;"3D;�G;�I;�]I;�ZI;	DI;H1I;�"I;`I;�I;�I;�I;�I;�I;�I;�I;`I;�"I;H1I;	DI;�ZI;�]I;�I;�G;"3D;�<;˅+;mM;���:x5� �$�Kkλ<RH��֮�v�C�d��A�����	�I�w���u]׾����O�����f���dȿF�ῢ��      6��������欿��������O�}x����� ���l���"��ܽ���`=�Ý��l"��R���ۺM��9�=�:�K;��0;͞>;�LE;|"H;�$I;�`I;(VI;�?I;.I;` I;[I;"I;/
I;lI;�I;lI;/
I;"I;[I;` I;.I;�?I;(VI;�`I;�$I;|"H;�LE;͞>;��0;�K;�=�:M��9�ۺ�R��l"����Ý��`=����ܽ��"��l�� �����}x���O��������欿����      q�������Y�{�e$_��q<�������}��w���6�����!��!�h��������� d��.��g_e�UL[���Z:���:�+ ;��5;�A;�UF;˃H;@I;�aI;�PI;;I;e*I;�I;+I;WI;�I;I;LI;I;�I;WI;+I;�I;e*I;;I;�PI;�aI;@I;˃H;�UF;�A;��5;�+ ;���:��Z:UL[�g_e��.��� d��������!�h�!�������6�w���}��������q<�e$_�Y�{�����      uA��q<�aa/����:�u]׾� ��w��>�BE	�����ܽ����3�r�꼰���>",�X��4��`AQ�خ�:�L
;�e);ބ:;D?C;?G;|�H;fSI;�^I;KJI;6I;t&I;�I;�I;ZI;�I;�I;�I;�I;�I;ZI;�I;�I;t&I;6I;KJI;�^I;fSI;|�H;?G;D?C;ބ:;�e);�L
;خ�:`AQ�4��X��>",�����r�꼠�3�ܽ������BE	�>�w��� ��u]׾�:���aa/��q<�      a5�������Q�Ҿ�a��w����l��6�BE	���Ƚk���aG����z֮�C�W����:�k����T`,:���:�;��1;m�>;^E;L�G;BI;G^I;hYI;ZCI;�0I;V"I;cI;I;#	I;,I;�I;=I;�I;,I;#	I;I;cI;V"I;�0I;ZCI;hYI;G^I;BI;L�G;^E;m�>;��1;�;���:T`,:���:�k����C�W�z֮�����aG�k����ȽBE	��6��l�w����a��Q�Ҿ������      � ���e�����ؕ����q�	�I���"���������k���ZN�c�6¼~�y��$�PR��]� ���[��:G/;J�&;
w8;��A;��F;��H;?I;aI;�QI;:<I;7+I;�I;I;uI;�I;WI;9I;� I;9I;WI;�I;uI;I;�I;7+I;:<I;�QI;aI;?I;��H;��F;��A;
w8;J�&;G/;�:��[�]� �PR���$�~�y�6¼c��ZN�k������������"�	�I���q�ؕ������e��      y^Z�[
V��I�
�6�������ܽ!��ܽ���aG�c��ȼ�)����(����H5���-�Z:j�:7R;/&1;��=;ПD;P�G;�H;�WI;9]I;�HI;5I;�%I;�I;�I;�	I;�I;mI;|�H;��H;|�H;mI;�I;�	I;�I;�I;�%I;5I;�HI;9]I;�WI;�H;P�G;ПD;��=;/&1;7R;j�:-�Z:��H5������(��)���ȼc��aG�ܽ��!���ܽ�����
�6��I�[
V�      ���FE	��������Wн�A����!�h���3����6¼�)��ax/�v�һD�X� %����9���:�=;[e);�_9;�%B;ډF;�|H;�5I;u`I;�TI;�?I;�-I; I;jI;DI;�I;jI;q�H;��H;�H;��H;q�H;jI;�I;DI;jI; I;�-I;�?I;�TI;u`I;�5I;�|H;ډF;�%B;�_9;[e);�=;���:��9 %��D�X�v�һax/��)��6¼�����3�!�h��󑽢A���Wн��콹��FE	�      �A��!��e���*��齅�C�d��`=����r��z֮�~�y���(�v�һk^e�������f9���:X�;m0";A�4;�l?; E;��G;��H;�VI;�]I;(JI;�6I;'I;�I;FI;�	I;=I;7 I;��H;��H;V�H;��H;��H;7 I;=I;�	I;FI;�I;'I;�6I;(JI;�]I;�VI;��H;��G; E;�l?;A�4;m0";X�;���:��f9����k^e�v�һ��(�~�y�z֮�r�꼠���`=�C�d�齅��*��e��!��      �]��IY��ZN��`=���'�v�Ý���������C�W��$����D�X������9�ޚ:���:��;ʷ0;�<;v�C;GG;�H;�>I;P`I;�SI;^?I;1.I;z I;�I;.I;�I;�I;��H;��H;&�H;��H;&�H;��H;��H;�I;�I;.I;�I;z I;1.I;^?I;�SI;P`I;�>I;�H;GG;v�C;�<;ʷ0;��;���:�ޚ:�9����D�X�����$�C�W���������Ý�v���'��`=��ZN��IY�      ���s9�o5��P��ib̼�֮����� d�>",����PR��H5� %����f9�ޚ:��:6�;��-;��:;KB;_UF;:JH; I;�[I;G[I;�GI;%5I;<&I;6I;�I;9	I;^I;�H;��H;��H;n�H;�H;n�H;��H;��H;�H;^I;9	I;�I;6I;<&I;%5I;�GI;G[I;�[I; I;:JH;_UF;KB;��:;��-;6�;��:�ޚ:��f9 %��H5�PR�����>",�� d�����֮�ib̼P��o5��s9�      �d��Z���Ǩ���)���zl�<RH�l"��.��X��:�k�]� �����9���:���:6�;�-;�9;j`A;۹E;J�G;��H;#RI;4_I;OI;�;I;�+I;�I;MI;)I;�I;p I;��H;��H;��H;��H;{�H;��H;��H;��H;��H;p I;�I;)I;MI;�I;�+I;�;I;OI;4_I;#RI;��H;J�G;۹E;j`A;�9;�-;6�;���:���:��9��]� �:�k�X���.��l"�<RH��zl��)��Ǩ��Z���      |",��(�nH�{G�/��Kkλ�R��g_e�4�������[�-�Z:���:X�;��;��-;�9;�A;�bE;D�G;��H;tFI;`I;�TI;bAI;�0I;#I;�I;I;�I;I;��H;a�H;��H;!�H;,�H;��H;,�H;!�H;��H;a�H;��H;I;�I;I;�I;#I;�0I;bAI;�TI;`I;tFI;��H;D�G;�bE;�A;�9;��-;��;X�;���:-�Z:��[����4��g_e��R��Kkλ/��{G�nH��(�      6�� S��� ���6���X� �$��ۺUL[�`AQ�T`,:�:j�:�=;m0";ʷ0;��:;j`A;�bE;�G;��H;�<I;N_I;�XI;FI;5I;�&I;I;�I;
I;�I;��H;�H;6�H;�H;��H;��H;S�H;��H;��H;�H;6�H;�H;��H;�I;
I;�I;I;�&I;5I;FI;�XI;N_I;�<I;��H;�G;�bE;j`A;��:;ʷ0;m0";�=;j�:�:T`,:`AQ�UL[��ۺ �$��X��6��� �� S��      :�Ѻ��Ⱥ����B��{��x5�M��9��Z:خ�:���:G/;7R;[e);A�4;�<;KB;۹E;D�G;��H;�9I;q^I;�ZI;?II;8I;�)I;�I;I;I;vI;$ I;��H;��H;%�H;C�H;�H;F�H;��H;F�H;�H;C�H;%�H;��H;��H;$ I;vI;I;I;�I;�)I;8I;?II;�ZI;q^I;�9I;��H;D�G;۹E;KB;�<;A�4;[e);7R;G/;���:خ�:��Z:M��9x5�{��B��������Ⱥ      ���9��:ܧ":��Q:�:���:�=�:���:�L
;�;J�&;/&1;�_9;�l?;v�C;_UF;J�G;��H;�<I;q^I;1[I;�JI;1:I;�+I;�I;I;�I;�I;`I;��H;K�H;��H;J�H;��H;��H;��H;��H;��H;��H;��H;J�H;��H;K�H;��H;`I;�I;�I;I;�I;�+I;1:I;�JI;1[I;q^I;�<I;��H;J�G;_UF;v�C;�l?;�_9;/&1;J�&;�;�L
;���:�=�:���:�:��Q:ܧ":��:      '��:���:��:�:��;mM;�K;�+ ;�e);��1;
w8;��=;�%B; E;GG;:JH;��H;tFI;N_I;�ZI;�JI;�:I;-I;H!I;QI;*I;0I;xI;��H;��H;��H;}�H;��H;-�H;R�H;��H;y�H;��H;R�H;-�H;��H;}�H;��H;��H;��H;xI;0I;*I;QI;H!I;-I;�:I;�JI;�ZI;N_I;tFI;��H;:JH;GG; E;�%B;��=;
w8;��1;�e);�+ ;�K;mM;��;�:��:���:      d�;'�;��;/";
�&;˅+;��0;��5;ބ:;m�>;��A;ПD;ډF;��G;�H; I;#RI;`I;�XI;?II;1:I;-I;�!I;I;�I;	I;BI;]�H;��H;j�H;��H;��H;�H;��H; �H;��H;p�H;��H; �H;��H;�H;��H;��H;j�H;��H;]�H;BI;	I;�I;I;�!I;-I;1:I;?II;�XI;`I;#RI; I;�H;��G;ډF;ПD;��A;m�>;ބ:;��5;��0;˅+;
�&;/";��;'�;      dX4;K�4;��5;�7;٪9;�<;͞>;�A;D?C;^E;��F;P�G;�|H;��H;�>I;�[I;4_I;�TI;FI;8I;�+I;H!I;I;8I;v	I;�I; �H;��H;��H;��H;��H;�H;��H;��H;��H;��H;u�H;��H;��H;��H;��H;�H;��H;��H;��H;��H; �H;�I;v	I;8I;I;H!I;�+I;8I;FI;�TI;4_I;�[I;�>I;��H;�|H;P�G;��F;^E;D?C;�A;͞>;�<;٪9;�7;��5;K�4;      p�@;h�@;�_A;�%B;KC;"3D;�LE;�UF;?G;L�G;��H;�H;�5I;�VI;P`I;G[I;OI;bAI;5I;�)I;�I;QI;�I;v	I;I;.�H;D�H;��H;0�H;��H;�H;��H;[�H;��H;��H;��H;r�H;��H;��H;��H;[�H;��H;�H;��H;0�H;��H;D�H;.�H;I;v	I;�I;QI;�I;�)I;5I;bAI;OI;G[I;P`I;�VI;�5I;�H;��H;L�G;?G;�UF;�LE;"3D;KC;�%B;�_A;h�@;      �UF;kgF;ٚF;�F;vLG;�G;|"H;˃H;|�H;BI;?I;�WI;u`I;�]I;�SI;�GI;�;I;�0I;�&I;�I;I;*I;	I;�I;.�H;V�H;'�H;i�H;��H;�H;��H;V�H;L�H;��H;�H;��H;��H;��H;�H;��H;L�H;V�H;��H;�H;��H;i�H;'�H;V�H;.�H;�I;	I;*I;I;�I;�&I;�0I;�;I;�GI;�SI;�]I;u`I;�WI;?I;BI;|�H;˃H;|"H;�G;vLG;�F;ٚF;kgF;      ��H;��H;Z�H;��H;�H;�I;�$I;@I;fSI;G^I;aI;9]I;�TI;(JI;^?I;%5I;�+I;#I;I;I;�I;0I;BI; �H;D�H;'�H;\�H;�H;7�H;|�H;6�H;�H;E�H;��H;@�H;��H;��H;��H;@�H;��H;E�H;�H;6�H;|�H;7�H;�H;\�H;'�H;D�H; �H;BI;0I;�I;I;I;#I;�+I;%5I;^?I;(JI;�TI;9]I;aI;G^I;fSI;@I;�$I;�I;�H;��H;Z�H;��H;      �FI;4HI;;LI;RI;]XI;�]I;�`I;�aI;�^I;hYI;�QI;�HI;�?I;�6I;1.I;<&I;�I;�I;�I;I;�I;xI;]�H;��H;��H;i�H;�H;�H;��H;2�H;�H;�H;p�H;��H;|�H;F�H;@�H;F�H;|�H;��H;p�H;�H;�H;2�H;��H;�H;�H;i�H;��H;��H;]�H;xI;�I;I;�I;�I;�I;<&I;1.I;�6I;�?I;�HI;�QI;hYI;�^I;�aI;�`I;�]I;]XI;RI;;LI;4HI;      �aI;�aI;aI;�_I;�]I;�ZI;(VI;�PI;KJI;ZCI;:<I;5I;�-I;'I;z I;6I;MI;I;
I;vI;`I;��H;��H;��H;0�H;��H;7�H;��H;)�H;�H; �H;B�H;��H;2�H;��H;��H;��H;��H;��H;2�H;��H;B�H; �H;�H;)�H;��H;7�H;��H;0�H;��H;��H;��H;`I;vI;
I;I;MI;6I;z I;'I;�-I;5I;:<I;ZCI;KJI;�PI;(VI;�ZI;�]I;�_I;aI;�aI;      2NI;�MI;�LI;�JI;�GI;	DI;�?I;;I;6I;�0I;7+I;�%I; I;�I;�I;�I;)I;�I;�I;$ I;��H;��H;j�H;��H;��H;�H;|�H;2�H;�H;�H;1�H;��H;��H;��H;H�H;(�H;%�H;(�H;H�H;��H;��H;��H;1�H;�H;�H;2�H;|�H;�H;��H;��H;j�H;��H;��H;$ I;�I;�I;)I;�I;�I;�I; I;�%I;7+I;�0I;6I;;I;�?I;	DI;�GI;�JI;�LI;�MI;      A9I;�8I;�7I;C6I;4I;H1I;.I;e*I;t&I;V"I;�I;�I;jI;FI;.I;9	I;�I;I;��H;��H;K�H;��H;��H;��H;�H;��H;6�H;�H; �H;1�H;��H;��H;d�H;�H;��H;��H;��H;��H;��H;�H;d�H;��H;��H;1�H; �H;�H;6�H;��H;�H;��H;��H;��H;K�H;��H;��H;I;�I;9	I;.I;FI;jI;�I;�I;V"I;t&I;e*I;.I;H1I;4I;C6I;�7I;�8I;      �(I;�(I;(I;�&I;�$I;�"I;` I;�I;�I;cI;I;�I;DI;�	I;�I;^I;p I;��H;�H;��H;��H;}�H;��H;�H;��H;V�H;�H;�H;B�H;��H;��H;{�H;��H;��H;z�H;T�H;>�H;T�H;z�H;��H;��H;{�H;��H;��H;B�H;�H;�H;V�H;��H;�H;��H;}�H;��H;��H;�H;��H;p I;^I;�I;�	I;DI;�I;I;cI;�I;�I;` I;�"I;�$I;�&I;(I;�(I;      <I;I;aI;ZI;I;`I;[I;+I;�I;I;uI;�	I;�I;=I;�I;�H;��H;a�H;6�H;%�H;J�H;��H;�H;��H;[�H;L�H;E�H;p�H;��H;��H;d�H;��H;��H;[�H;�H;�H;�H;�H;�H;[�H;��H;��H;d�H;��H;��H;p�H;E�H;L�H;[�H;��H;�H;��H;J�H;%�H;6�H;a�H;��H;�H;�I;=I;�I;�	I;uI;I;�I;+I;[I;`I;I;ZI;aI;I;      �I;~I;I;7I;'I;�I;"I;WI;ZI;#	I;�I;�I;jI;7 I;��H;��H;��H;��H;�H;C�H;��H;-�H;��H;��H;��H;��H;��H;��H;2�H;��H;�H;��H;[�H; �H;��H;��H;��H;��H;��H; �H;[�H;��H;�H;��H;2�H;��H;��H;��H;��H;��H;��H;-�H;��H;C�H;�H;��H;��H;��H;��H;7 I;jI;�I;�I;#	I;ZI;WI;"I;�I;'I;7I;I;~I;      �I;�I;_I;�I;�I;�I;/
I;�I;�I;,I;WI;mI;q�H;��H;��H;��H;��H;!�H;��H;�H;��H;R�H; �H;��H;��H;�H;@�H;|�H;��H;H�H;��H;z�H;�H;��H;��H;��H;��H;��H;��H;��H;�H;z�H;��H;H�H;��H;|�H;@�H;�H;��H;��H; �H;R�H;��H;�H;��H;!�H;��H;��H;��H;��H;q�H;mI;WI;,I;�I;�I;/
I;�I;�I;�I;_I;�I;      �I;{I;&I;�
I;�	I;�I;lI;I;�I;�I;9I;|�H;��H;��H;&�H;n�H;��H;,�H;��H;F�H;��H;��H;��H;��H;��H;��H;��H;F�H;��H;(�H;��H;T�H;�H;��H;��H;��H;}�H;��H;��H;��H;�H;T�H;��H;(�H;��H;F�H;��H;��H;��H;��H;��H;��H;��H;F�H;��H;,�H;��H;n�H;&�H;��H;��H;|�H;9I;�I;�I;I;lI;�I;�	I;�
I;&I;{I;      �
I;x
I;&
I;�	I;�I;�I;�I;LI;�I;=I;� I;��H;�H;V�H;��H;�H;{�H;��H;S�H;��H;��H;y�H;p�H;u�H;r�H;��H;��H;@�H;��H;%�H;��H;>�H;�H;��H;��H;}�H;��H;}�H;��H;��H;�H;>�H;��H;%�H;��H;@�H;��H;��H;r�H;u�H;p�H;y�H;��H;��H;S�H;��H;{�H;�H;��H;V�H;�H;��H;� I;=I;�I;LI;�I;�I;�I;�	I;&
I;x
I;      �I;{I;&I;�
I;�	I;�I;lI;I;�I;�I;9I;|�H;��H;��H;&�H;n�H;��H;,�H;��H;F�H;��H;��H;��H;��H;��H;��H;��H;F�H;��H;(�H;��H;T�H;�H;��H;��H;��H;}�H;��H;��H;��H;�H;T�H;��H;(�H;��H;F�H;��H;��H;��H;��H;��H;��H;��H;F�H;��H;,�H;��H;n�H;&�H;��H;��H;|�H;9I;�I;�I;I;lI;�I;�	I;�
I;&I;{I;      �I;�I;_I;�I;�I;�I;/
I;�I;�I;,I;WI;mI;q�H;��H;��H;��H;��H;!�H;��H;�H;��H;R�H; �H;��H;��H;�H;@�H;|�H;��H;H�H;��H;z�H;�H;��H;��H;��H;��H;��H;��H;��H;�H;z�H;��H;H�H;��H;|�H;@�H;�H;��H;��H; �H;R�H;��H;�H;��H;!�H;��H;��H;��H;��H;q�H;mI;WI;,I;�I;�I;/
I;�I;�I;�I;_I;�I;      �I;~I;I;7I;'I;�I;"I;WI;ZI;#	I;�I;�I;jI;7 I;��H;��H;��H;��H;�H;C�H;��H;-�H;��H;��H;��H;��H;��H;��H;2�H;��H;�H;��H;[�H; �H;��H;��H;��H;��H;��H; �H;[�H;��H;�H;��H;2�H;��H;��H;��H;��H;��H;��H;-�H;��H;C�H;�H;��H;��H;��H;��H;7 I;jI;�I;�I;#	I;ZI;WI;"I;�I;'I;7I;I;~I;      <I;I;aI;ZI;I;`I;[I;+I;�I;I;uI;�	I;�I;=I;�I;�H;��H;a�H;6�H;%�H;J�H;��H;�H;��H;[�H;L�H;E�H;p�H;��H;��H;d�H;��H;��H;[�H;�H;�H;�H;�H;�H;[�H;��H;��H;d�H;��H;��H;p�H;E�H;L�H;[�H;��H;�H;��H;J�H;%�H;6�H;a�H;��H;�H;�I;=I;�I;�	I;uI;I;�I;+I;[I;`I;I;ZI;aI;I;      �(I;�(I;(I;�&I;�$I;�"I;` I;�I;�I;cI;I;�I;DI;�	I;�I;^I;p I;��H;�H;��H;��H;}�H;��H;�H;��H;V�H;�H;�H;B�H;��H;��H;{�H;��H;��H;z�H;T�H;>�H;T�H;z�H;��H;��H;{�H;��H;��H;B�H;�H;�H;V�H;��H;�H;��H;}�H;��H;��H;�H;��H;p I;^I;�I;�	I;DI;�I;I;cI;�I;�I;` I;�"I;�$I;�&I;(I;�(I;      A9I;�8I;�7I;C6I;4I;H1I;.I;e*I;t&I;V"I;�I;�I;jI;FI;.I;9	I;�I;I;��H;��H;K�H;��H;��H;��H;�H;��H;6�H;�H; �H;1�H;��H;��H;d�H;�H;��H;��H;��H;��H;��H;�H;d�H;��H;��H;1�H; �H;�H;6�H;��H;�H;��H;��H;��H;K�H;��H;��H;I;�I;9	I;.I;FI;jI;�I;�I;V"I;t&I;e*I;.I;H1I;4I;C6I;�7I;�8I;      2NI;�MI;�LI;�JI;�GI;	DI;�?I;;I;6I;�0I;7+I;�%I; I;�I;�I;�I;)I;�I;�I;$ I;��H;��H;j�H;��H;��H;�H;|�H;2�H;�H;�H;1�H;��H;��H;��H;H�H;(�H;%�H;(�H;H�H;��H;��H;��H;1�H;�H;�H;2�H;|�H;�H;��H;��H;j�H;��H;��H;$ I;�I;�I;)I;�I;�I;�I; I;�%I;7+I;�0I;6I;;I;�?I;	DI;�GI;�JI;�LI;�MI;      �aI;�aI;aI;�_I;�]I;�ZI;(VI;�PI;KJI;ZCI;:<I;5I;�-I;'I;z I;6I;MI;I;
I;vI;`I;��H;��H;��H;0�H;��H;7�H;��H;)�H;�H; �H;B�H;��H;2�H;��H;��H;��H;��H;��H;2�H;��H;B�H; �H;�H;)�H;��H;7�H;��H;0�H;��H;��H;��H;`I;vI;
I;I;MI;6I;z I;'I;�-I;5I;:<I;ZCI;KJI;�PI;(VI;�ZI;�]I;�_I;aI;�aI;      �FI;4HI;;LI;RI;]XI;�]I;�`I;�aI;�^I;hYI;�QI;�HI;�?I;�6I;1.I;<&I;�I;�I;�I;I;�I;xI;]�H;��H;��H;i�H;�H;�H;��H;2�H;�H;�H;p�H;��H;|�H;F�H;@�H;F�H;|�H;��H;p�H;�H;�H;2�H;��H;�H;�H;i�H;��H;��H;]�H;xI;�I;I;�I;�I;�I;<&I;1.I;�6I;�?I;�HI;�QI;hYI;�^I;�aI;�`I;�]I;]XI;RI;;LI;4HI;      ��H;��H;Z�H;��H;�H;�I;�$I;@I;fSI;G^I;aI;9]I;�TI;(JI;^?I;%5I;�+I;#I;I;I;�I;0I;BI; �H;D�H;'�H;\�H;�H;7�H;|�H;6�H;�H;E�H;��H;@�H;��H;��H;��H;@�H;��H;E�H;�H;6�H;|�H;7�H;�H;\�H;'�H;D�H; �H;BI;0I;�I;I;I;#I;�+I;%5I;^?I;(JI;�TI;9]I;aI;G^I;fSI;@I;�$I;�I;�H;��H;Z�H;��H;      �UF;kgF;ٚF;�F;vLG;�G;|"H;˃H;|�H;BI;?I;�WI;u`I;�]I;�SI;�GI;�;I;�0I;�&I;�I;I;*I;	I;�I;.�H;V�H;'�H;i�H;��H;�H;��H;V�H;L�H;��H;�H;��H;��H;��H;�H;��H;L�H;V�H;��H;�H;��H;i�H;'�H;V�H;.�H;�I;	I;*I;I;�I;�&I;�0I;�;I;�GI;�SI;�]I;u`I;�WI;?I;BI;|�H;˃H;|"H;�G;vLG;�F;ٚF;kgF;      p�@;h�@;�_A;�%B;KC;"3D;�LE;�UF;?G;L�G;��H;�H;�5I;�VI;P`I;G[I;OI;bAI;5I;�)I;�I;QI;�I;v	I;I;.�H;D�H;��H;0�H;��H;�H;��H;[�H;��H;��H;��H;r�H;��H;��H;��H;[�H;��H;�H;��H;0�H;��H;D�H;.�H;I;v	I;�I;QI;�I;�)I;5I;bAI;OI;G[I;P`I;�VI;�5I;�H;��H;L�G;?G;�UF;�LE;"3D;KC;�%B;�_A;h�@;      dX4;K�4;��5;�7;٪9;�<;͞>;�A;D?C;^E;��F;P�G;�|H;��H;�>I;�[I;4_I;�TI;FI;8I;�+I;H!I;I;8I;v	I;�I; �H;��H;��H;��H;��H;�H;��H;��H;��H;��H;u�H;��H;��H;��H;��H;�H;��H;��H;��H;��H; �H;�I;v	I;8I;I;H!I;�+I;8I;FI;�TI;4_I;�[I;�>I;��H;�|H;P�G;��F;^E;D?C;�A;͞>;�<;٪9;�7;��5;K�4;      d�;'�;��;/";
�&;˅+;��0;��5;ބ:;m�>;��A;ПD;ډF;��G;�H; I;#RI;`I;�XI;?II;1:I;-I;�!I;I;�I;	I;BI;]�H;��H;j�H;��H;��H;�H;��H; �H;��H;p�H;��H; �H;��H;�H;��H;��H;j�H;��H;]�H;BI;	I;�I;I;�!I;-I;1:I;?II;�XI;`I;#RI; I;�H;��G;ډF;ПD;��A;m�>;ބ:;��5;��0;˅+;
�&;/";��;'�;      '��:���:��:�:��;mM;�K;�+ ;�e);��1;
w8;��=;�%B; E;GG;:JH;��H;tFI;N_I;�ZI;�JI;�:I;-I;H!I;QI;*I;0I;xI;��H;��H;��H;}�H;��H;-�H;R�H;��H;y�H;��H;R�H;-�H;��H;}�H;��H;��H;��H;xI;0I;*I;QI;H!I;-I;�:I;�JI;�ZI;N_I;tFI;��H;:JH;GG; E;�%B;��=;
w8;��1;�e);�+ ;�K;mM;��;�:��:���:      ���9��:ܧ":��Q:�:���:�=�:���:�L
;�;J�&;/&1;�_9;�l?;v�C;_UF;J�G;��H;�<I;q^I;1[I;�JI;1:I;�+I;�I;I;�I;�I;`I;��H;K�H;��H;J�H;��H;��H;��H;��H;��H;��H;��H;J�H;��H;K�H;��H;`I;�I;�I;I;�I;�+I;1:I;�JI;1[I;q^I;�<I;��H;J�G;_UF;v�C;�l?;�_9;/&1;J�&;�;�L
;���:�=�:���:�:��Q:ܧ":��:      :�Ѻ��Ⱥ����B��{��x5�M��9��Z:خ�:���:G/;7R;[e);A�4;�<;KB;۹E;D�G;��H;�9I;q^I;�ZI;?II;8I;�)I;�I;I;I;vI;$ I;��H;��H;%�H;C�H;�H;F�H;��H;F�H;�H;C�H;%�H;��H;��H;$ I;vI;I;I;�I;�)I;8I;?II;�ZI;q^I;�9I;��H;D�G;۹E;KB;�<;A�4;[e);7R;G/;���:خ�:��Z:M��9x5�{��B��������Ⱥ      6�� S��� ���6���X� �$��ۺUL[�`AQ�T`,:�:j�:�=;m0";ʷ0;��:;j`A;�bE;�G;��H;�<I;N_I;�XI;FI;5I;�&I;I;�I;
I;�I;��H;�H;6�H;�H;��H;��H;S�H;��H;��H;�H;6�H;�H;��H;�I;
I;�I;I;�&I;5I;FI;�XI;N_I;�<I;��H;�G;�bE;j`A;��:;ʷ0;m0";�=;j�:�:T`,:`AQ�UL[��ۺ �$��X��6��� �� S��      |",��(�nH�{G�/��Kkλ�R��g_e�4�������[�-�Z:���:X�;��;��-;�9;�A;�bE;D�G;��H;tFI;`I;�TI;bAI;�0I;#I;�I;I;�I;I;��H;a�H;��H;!�H;,�H;��H;,�H;!�H;��H;a�H;��H;I;�I;I;�I;#I;�0I;bAI;�TI;`I;tFI;��H;D�G;�bE;�A;�9;��-;��;X�;���:-�Z:��[����4��g_e��R��Kkλ/��{G�nH��(�      �d��Z���Ǩ���)���zl�<RH�l"��.��X��:�k�]� �����9���:���:6�;�-;�9;j`A;۹E;J�G;��H;#RI;4_I;OI;�;I;�+I;�I;MI;)I;�I;p I;��H;��H;��H;��H;{�H;��H;��H;��H;��H;p I;�I;)I;MI;�I;�+I;�;I;OI;4_I;#RI;��H;J�G;۹E;j`A;�9;�-;6�;���:���:��9��]� �:�k�X���.��l"�<RH��zl��)��Ǩ��Z���      ���s9�o5��P��ib̼�֮����� d�>",����PR��H5� %����f9�ޚ:��:6�;��-;��:;KB;_UF;:JH; I;�[I;G[I;�GI;%5I;<&I;6I;�I;9	I;^I;�H;��H;��H;n�H;�H;n�H;��H;��H;�H;^I;9	I;�I;6I;<&I;%5I;�GI;G[I;�[I; I;:JH;_UF;KB;��:;��-;6�;��:�ޚ:��f9 %��H5�PR�����>",�� d�����֮�ib̼P��o5��s9�      �]��IY��ZN��`=���'�v�Ý���������C�W��$����D�X������9�ޚ:���:��;ʷ0;�<;v�C;GG;�H;�>I;P`I;�SI;^?I;1.I;z I;�I;.I;�I;�I;��H;��H;&�H;��H;&�H;��H;��H;�I;�I;.I;�I;z I;1.I;^?I;�SI;P`I;�>I;�H;GG;v�C;�<;ʷ0;��;���:�ޚ:�9����D�X�����$�C�W���������Ý�v���'��`=��ZN��IY�      �A��!��e���*��齅�C�d��`=����r��z֮�~�y���(�v�һk^e�������f9���:X�;m0";A�4;�l?; E;��G;��H;�VI;�]I;(JI;�6I;'I;�I;FI;�	I;=I;7 I;��H;��H;V�H;��H;��H;7 I;=I;�	I;FI;�I;'I;�6I;(JI;�]I;�VI;��H;��G; E;�l?;A�4;m0";X�;���:��f9����k^e�v�һ��(�~�y�z֮�r�꼠���`=�C�d�齅��*��e��!��      ���FE	��������Wн�A����!�h���3����6¼�)��ax/�v�һD�X� %����9���:�=;[e);�_9;�%B;ډF;�|H;�5I;u`I;�TI;�?I;�-I; I;jI;DI;�I;jI;q�H;��H;�H;��H;q�H;jI;�I;DI;jI; I;�-I;�?I;�TI;u`I;�5I;�|H;ډF;�%B;�_9;[e);�=;���:��9 %��D�X�v�һax/��)��6¼�����3�!�h��󑽢A���Wн��콹��FE	�      y^Z�[
V��I�
�6�������ܽ!��ܽ���aG�c��ȼ�)����(����H5���-�Z:j�:7R;/&1;��=;ПD;P�G;�H;�WI;9]I;�HI;5I;�%I;�I;�I;�	I;�I;mI;|�H;��H;|�H;mI;�I;�	I;�I;�I;�%I;5I;�HI;9]I;�WI;�H;P�G;ПD;��=;/&1;7R;j�:-�Z:��H5������(��)���ȼc��aG�ܽ��!���ܽ�����
�6��I�[
V�      � ���e�����ؕ����q�	�I���"���������k���ZN�c�6¼~�y��$�PR��]� ���[��:G/;J�&;
w8;��A;��F;��H;?I;aI;�QI;:<I;7+I;�I;I;uI;�I;WI;9I;� I;9I;WI;�I;uI;I;�I;7+I;:<I;�QI;aI;?I;��H;��F;��A;
w8;J�&;G/;�:��[�]� �PR���$�~�y�6¼c��ZN�k������������"�	�I���q�ؕ������e��      a5�������Q�Ҿ�a��w����l��6�BE	���Ƚk���aG����z֮�C�W����:�k����T`,:���:�;��1;m�>;^E;L�G;BI;G^I;hYI;ZCI;�0I;V"I;cI;I;#	I;,I;�I;=I;�I;,I;#	I;I;cI;V"I;�0I;ZCI;hYI;G^I;BI;L�G;^E;m�>;��1;�;���:T`,:���:�k����C�W�z֮�����aG�k����ȽBE	��6��l�w����a��Q�Ҿ������      uA��q<�aa/����:�u]׾� ��w��>�BE	�����ܽ����3�r�꼰���>",�X��4��`AQ�خ�:�L
;�e);ބ:;D?C;?G;|�H;fSI;�^I;KJI;6I;t&I;�I;�I;ZI;�I;�I;�I;�I;�I;ZI;�I;�I;t&I;6I;KJI;�^I;fSI;|�H;?G;D?C;ބ:;�e);�L
;خ�:`AQ�4��X��>",�����r�꼠�3�ܽ������BE	�>�w��� ��u]׾�:���aa/��q<�      q�������Y�{�e$_��q<�������}��w���6�����!��!�h��������� d��.��g_e�UL[���Z:���:�+ ;��5;�A;�UF;˃H;@I;�aI;�PI;;I;e*I;�I;+I;WI;�I;I;LI;I;�I;WI;+I;�I;e*I;;I;�PI;�aI;@I;˃H;�UF;�A;��5;�+ ;���:��Z:UL[�g_e��.��� d��������!�h�!�������6�w���}��������q<�e$_�Y�{�����      6��������欿��������O�}x����� ���l���"��ܽ���`=�Ý��l"��R���ۺM��9�=�:�K;��0;͞>;�LE;|"H;�$I;�`I;(VI;�?I;.I;` I;[I;"I;/
I;lI;�I;lI;/
I;"I;[I;` I;.I;�?I;(VI;�`I;�$I;|"H;�LE;͞>;��0;�K;�=�:M��9�ۺ�R��l"����Ý��`=����ܽ��"��l�� �����}x���O��������欿����      �������F��dȿf���������O���u]׾w���	�I�����A��C�d�v��֮�<RH�Kkλ �$�x5����:mM;˅+;�<;"3D;�G;�I;�]I;�ZI;	DI;H1I;�"I;`I;�I;�I;�I;�I;�I;�I;�I;`I;�"I;H1I;	DI;�ZI;�]I;�I;�G;"3D;�<;˅+;mM;���:x5� �$�Kkλ<RH��֮�v�C�d��A�����	�I�w���u]׾����O�����f���dȿF�ῢ��      @�-i�������B�ѿf�������q<��:��a����q����Wн齅���'�ib̼�zl�/���X�{���:��;
�&;٪9;KC;vLG;�H;]XI;�]I;�GI;4I;�$I;I;'I;�I;�	I;�I;�	I;�I;'I;I;�$I;4I;�GI;�]I;]XI;�H;vLG;KC;٪9;
�&;��;�:{���X�/���zl�ib̼��'�齅��Wн����q��a���:��q<����f���B�ѿ������-i�      A:�.5�(�'��������dȿ���e$_���Q�Ҿؕ��
�6�����*���`=�P���)��{G��6��B����Q:�:/";�7;�%B;�F;��H;RI;�_I;�JI;C6I;�&I;ZI;7I;�I;�
I;�	I;�
I;�I;7I;ZI;�&I;C6I;�JI;�_I;RI;��H;�F;�%B;�7;/";�:��Q:B���6��{G��)��P���`=��*�����
�6�ؕ��Q�Ҿ��e$_����dȿ�������(�'�.5�      ��U�T�O�B-?�(�'���F�`欿Y�{�aa/���뾙���I����e���ZN�o5��Ǩ��nH�� ������ܧ":��:��;��5;�_A;ٚF;Z�H;;LI;aI;�LI;�7I;(I;aI;I;_I;&I;&
I;&I;_I;I;aI;(I;�7I;�LI;aI;;LI;Z�H;ٚF;�_A;��5;��;��:ܧ":����� ��nH�Ǩ��o5���ZN�e������I�������aa/�Y�{��欿F����(�'�B-?�T�O�      ��i���b�T�O�.5�-i������������q<�����e��[
V�FE	�!���IY�s9�Z����(� S����Ⱥ��:���:'�;K�4;h�@;kgF;��H;4HI;�aI;�MI;�8I;�(I;I;~I;�I;{I;x
I;{I;�I;~I;I;�(I;�8I;�MI;�aI;4HI;��H;kgF;h�@;K�4;'�;���:��:��Ⱥ S���(�Z���s9��IY�!��FE	�[
V��e������q<������������-i�.5�T�O���b�      ݶ��O���ά��(�_���7�w�}߿���~,b��V�*l¾Fx�c.���Ž��t�6�����*�?��N�����sx9���:��;��2;T?@;�eF;C�H;��I;��I;8{I;�ZI;�BI;#1I;�$I;�I;�I;NI;�I;�I;�$I;#1I;�BI;�ZI;8{I;��I;��I;C�H;�eF;T?@;��2;��;���:�sx9���N��*�?����6����t���Žc.�Fx�*l¾�V�~,b����}߿w���7�(�_�ά��O���      O���A���}��+Y��3�����$ڿ"����\����(���s��3�9�����p�p�p���<<����f������9{��:�;V$3;ho@;yF;��H;�I;�I;�zI;rZI;yBI;�0I;s$I;EI;tI; I;tI;EI;s$I;�0I;yBI;rZI;�zI;�I;�I;��H;yF;ho@;V$3;�;{��:���9f�������<<�p��p���p�9����3��s�(�������\�"���$ڿ����3��+Y�}�A���      ά��}�8tf��lG�Ң%��p�*�ʿV����>M����S����d�ɤ�̷�9�d��
��I��@�1�������ޤ�9���:M;�T4;��@;�F;@�H; �I;ۙI;�xI;�XI;bAI;�/I;�#I;�I;�I;�I;�I;�I;�#I;�/I;bAI;�XI;�xI;ۙI; �I;@�H;�F;��@;�T4;M;���:ޤ�9������@�1��I���
�9�d�̷�ɤ��d�S�������>M�V���*�ʿ�p�Ң%��lG�8tf�}�      (�_��+Y��lG�f.�w���꿭���J䂿��5���󾋰��M�N�W��V��-�Q�*�������;i!��g��-󳺍:��:�;e06;��A;tG;I;Z�I;��I;�uI;qVI;�?I;�.I;�"I;�I;'I;�I;'I;�I;�"I;�.I;�?I;qVI;�uI;��I;Z�I;I;tG;��A;e06;�;��:�:-��g��;i!�����*���-�Q�V��W��M�N���������5�J䂿�������w�f.��lG��+Y�      ��7��3�Ң%�w��<����ſ�����\�9����Ͼ����`�3����z����9�z�ἷ���z��8}�ht�F�^:�)�:΢#;��8;��B;ArG;�$I;јI;�I;#qI;6SI;=I;�,I;0!I;nI;I;�I;I;nI;0!I;�,I;=I;6SI;#qI;�I;јI;�$I;ArG;��B;��8;΢#;�)�:F�^:ht��8}��z����z�Ἁ�9��z����`�3�������Ͼ9����\������ſ�<��w�Ң%��3�      w�����p������ſ!��{Ps���1�-r���d���d�}I�҈Ž��}�l*�fC��W�^�RC�g�D�+N๩��:��;�);-6;;JD;e�G;kGI;ΜI;ǎI;�kI;OI;�9I;3*I;8I;�I;�I;KI;�I;�I;8I;3*I;�9I;OI;�kI;ǎI;ΜI;kGI;e�G;JD;-6;;�);��;���:+N�g�D�RC�W�^�fC��l*���}�҈Ž}I��d��d��-r����1�{Ps�!����ſ��꿀p����      }߿�$ڿ*�ʿ�������{Ps�MX:����#l¾�ǆ���7����<5��$�Q�����t��85���������8�Ǽ:��;��.;��=;�DE;�XH;�gI;G�I;ڇI;FeI;@JI;E6I;a'I;�I;I;�I;�I;�I;I;�I;a'I;E6I;@JI;FeI;ڇI;G�I;�gI;�XH;�DE;��=;��.;��;�Ǽ:��8������85��t�����$�Q�<5�������7��ǆ�#l¾���MX:�{Ps��������*�ʿ�$ڿ      ���"��V���J䂿��\���1�����J˾睒�C�N�y��L������c�'���Ҽ �|��z�ko�� z��&�&:�N�:˧;�V4;�@;HfF;��H;.�I;A�I;UI;=^I;�DI;%2I;<$I;bI;�I;I;�I;I;�I;bI;<$I;%2I;�DI;=^I;UI;A�I;.�I;��H;HfF;�@;�V4;˧;�N�:&�&: z��ko���z� �|���Ҽc�'����L���y��C�N�睒��J˾�����1���\�J䂿V���"��      ~,b���\��>M���5�9��-r��#l¾睒�"&W��3�<Sؽ�z��fG�����I���?��̻{�-����J��:��;ο&;B{9;�C;�cG;sI;\�I;r�I;ruI;�VI;O?I;�-I;� I;�I;yI;�I;�I;�I;yI;�I;� I;�-I;O?I;�VI;ruI;r�I;\�I;sI;�cG;�C;B{9;ο&;��;J��:���{�-��̻�?��I�����fG��z��<Sؽ�3�"&W�睒�#l¾-r��9����5��>M���\�      �V������������Ͼ�d���ǆ�C�N��3��c�[����\�@��EC��O�o�Ъ	�t숻1�I��9I��:�g;o�/;\�=;aE;2H;�VI;؜I;�I;�jI;�NI;F9I;)I;=I;�I;I;�I;�
I;�I;I;�I;=I;)I;F9I;�NI;�jI;�I;؜I;�VI;2H;aE;\�=;o�/;�g;I��:I��91�t숻Ъ	�O�o�EC��@����\�[���cཱ3�C�N��ǆ��d����Ͼ���������      *l¾(��S������������d���7�y��<Sؽ[�� �d�P*�kּI\����'�����S������
�:�Y;�#;Y<7;M�A;2�F;{�H;��I;�I;րI;	`I;�FI;3I;B$I;�I;�I;vI;h	I;iI;h	I;vI;�I;�I;B$I;3I;�FI;	`I;րI;�I;��I;{�H;2�F;M�A;Y<7;�#;�Y;�
�:�����S������'�I\��kּP*� �d�[��<Sؽy����7��d���������S���(��      Fx��s��d�M�N�`�3�}I����L����z����\�P*�'�ݼe���j<<���ڻ��V��gt�q�&:���:[B;�;/;nC=;��D;��G;8I;�I;ÓI;3sI;IUI;}>I;�,I;�I;�I;xI;�	I;I;.I;I;�	I;xI;�I;�I;�,I;}>I;IUI;3sI;ÓI;�I;8I;��G;��D;nC=;�;/;[B;���:q�&:�gt���V���ڻj<<�e���'�ݼP*���\��z��L������}I�`�3�M�N��d��s�      c.��3�ɤ�W����҈Ž<5�����fG�@��kּe���:yC�?�X7}�񮼺E�x9���:%	;N�&;�:8;��A;��F;ϸH;WxI;��I;�I;PeI;�JI;m6I;�&I;�I;�I;uI;/I;�I;�I;�I;/I;uI;�I;�I;�&I;m6I;�JI;PeI;�I;��I;WxI;ϸH;��F;��A;�:8;N�&;%	;���:E�x9񮼺X7}�?�:yC�e���kּ@��fG����<5��҈Ž��W��ɤ��3�      ��Ž9���̷�V���z����}�$�Q�c�'����EC��I\��j<<�?��n�� ��rU�b��:Y��:,�;�&3;��>;�E;�H;};I;�I;ÔI;�uI;�WI;�@I;�.I;� I;�I;I;oI;I;<I;�I;<I;I;oI;I;�I;� I;�.I;�@I;�WI;�uI;ÔI;�I;};I;�H;�E;��>;�&3;,�;Y��:b��:rU� ���n��?�j<<�I\��EC�����c�'�$�Q���}��z��V��̷�9���      ��t���p�9�d�-�Q���9�l*������Ҽ�I��O�o���'���ڻX7}� ��vH��߄:�k�:��;�.;5<;�nC;^6G;��H;�I;��I;�I;;eI;^KI;7I;�&I;�I;�I;h
I;cI;�I;��H;l�H;��H;�I;cI;h
I;�I;�I;�&I;7I;^KI;;eI;�I;��I;�I;��H;^6G;�nC;5<;�.;��;�k�:�߄:vH� ��X7}���ڻ��'�O�o��I����Ҽ���l*���9�-�Q�9�d���p�      6��p��
�*���z��fC���t�� �|��?�Ъ	������V�񮼺rU��߄:��:�g;6�+;�9;��A;�eF;w�H;�^I;��I;��I; rI;�UI;�?I;�-I; I;uI;'I;�I;�I;i�H;��H;�H;��H;i�H;�I;�I;'I;uI; I;�-I;�?I;�UI; rI;��I;��I;�^I;w�H;�eF;��A;�9;6�+;�g;��:�߄:rU�񮼺��V����Ъ	��?� �|��t��fC��z��*����
�p�      ���p���I���������W�^�85��z��̻t숻�S��gt�E�x9b��:�k�:�g;y�*;�8;�@;��E;W'H;�7I;ߒI;2�I;o}I;�_I;�GI;�4I;y%I;�I;QI;	I;�I;��H;�H;i�H;��H;i�H;�H;��H;�I;	I;QI;�I;y%I;�4I;�GI;�_I;o}I;2�I;ߒI;�7I;W'H;��E;�@;�8;y�*;�g;�k�:b��:E�x9�gt��S�t숻�̻�z�85�W�^���������I��p��      *�?��<<�@�1�;i!��z�RC����ko��{�-�1򳺵���q�&:���:Y��:��;6�+;�8;W�@;]E;��G;eI;	�I;l�I;P�I;�hI;TOI;";I;�*I;�I;�I;nI;EI;� I;��H;��H;d�H;��H;d�H;��H;��H;� I;EI;nI;�I;�I;�*I;";I;TOI;�hI;P�I;l�I;	�I;eI;��G;]E;W�@;�8;6�+;��;Y��:���:q�&:����1�{�-�ko�����RC��z�;i!�@�1��<<�      �N����������g���8}�g�D���� z�����I��9�
�:���:%	;,�;�.;�9;�@;]E;��G;\I;�~I;#�I;g�I;�oI;�UI;�@I;�/I;�!I;�I;I;I;�I;��H;s�H;��H;r�H;��H;r�H;��H;s�H;��H;�I;I;I;�I;�!I;�/I;�@I;�UI;�oI;g�I;#�I;�~I;\I;��G;]E;�@;�9;�.;,�;%	;���:�
�:I��9��� z�����g�D��8}��g���������      ��f�����-�ht�+N���8&�&:J��:I��:�Y;[B;N�&;�&3;5<;��A;��E;��G;\I;v{I;ߛI;��I;�tI;�ZI;*EI;�3I;D%I;�I;bI;�I;I;O�H;��H;I�H;��H;��H;1�H;��H;��H;I�H;��H;O�H;I;�I;bI;�I;D%I;�3I;*EI;�ZI;�tI;��I;ߛI;v{I;\I;��G;��E;��A;5<;�&3;N�&;[B;�Y;I��:J��:&�&:��8+N�ht�-���f���      �sx9���9ޤ�9�:F�^:���:�Ǽ:�N�:��;�g;�#;�;/;�:8;��>;�nC;�eF;W'H;eI;�~I;ߛI;ːI;wI;�]I;QHI;�6I;(I;"I;�I;�
I;\I;b�H;]�H;h�H;L�H;��H;��H;��H;��H;��H;L�H;h�H;]�H;b�H;\I;�
I;�I;"I;(I;�6I;QHI;�]I;wI;ːI;ߛI;�~I;eI;W'H;�eF;�nC;��>;�:8;�;/;�#;�g;��;�N�:�Ǽ:���:F�^:�:ޤ�9���9      ���:{��:���:��:�)�:��;��;˧;ο&;o�/;Y<7;nC=;��A;�E;^6G;w�H;�7I;	�I;#�I;��I;wI;�^I;�II;�8I;*I;I;LI;QI;�I;L I;�H;��H;*�H;M�H;��H;�H;��H;�H;��H;M�H;*�H;��H;�H;L I;�I;QI;LI;I;*I;�8I;�II;�^I;wI;��I;#�I;	�I;�7I;w�H;^6G;�E;��A;nC=;Y<7;o�/;ο&;˧;��;��;�)�:��:���:{��:      ��;�;M;�;΢#;�);��.;�V4;B{9;\�=;M�A;��D;��F;�H;��H;�^I;ߒI;l�I;g�I;�tI;�]I;�II;=9I;6+I;VI;�I;gI;�I;4I;��H;�H;F�H;�H;z�H;o�H;��H;b�H;��H;o�H;z�H;�H;F�H;�H;��H;4I;�I;gI;�I;VI;6+I;=9I;�II;�]I;�tI;g�I;l�I;ߒI;�^I;��H;�H;��F;��D;M�A;\�=;B{9;�V4;��.;�);΢#;�;M;�;      ��2;V$3;�T4;e06;��8;-6;;��=;�@;�C;aE;2�F;��G;ϸH;};I;�I;��I;2�I;P�I;�oI;�ZI;QHI;�8I;6+I;�I;5I;2I;iI;�I;Y�H;s�H;q�H;:�H;L�H;��H;��H;i�H;�H;i�H;��H;��H;L�H;:�H;q�H;s�H;Y�H;�I;iI;2I;5I;�I;6+I;�8I;QHI;�ZI;�oI;P�I;2�I;��I;�I;};I;ϸH;��G;2�F;aE;�C;�@;��=;-6;;��8;e06;�T4;V$3;      T?@;ho@;��@;��A;��B;JD;�DE;HfF;�cG;2H;{�H;8I;WxI;�I;��I;��I;o}I;�hI;�UI;*EI;�6I;*I;VI;5I;tI;�I;QI;��H;��H;��H;.�H;0�H;��H;}�H;��H;,�H;	�H;,�H;��H;}�H;��H;0�H;.�H;��H;��H;��H;QI;�I;tI;5I;VI;*I;�6I;*EI;�UI;�hI;o}I;��I;��I;�I;WxI;8I;{�H;2H;�cG;HfF;�DE;JD;��B;��A;��@;ho@;      �eF;yF;�F;tG;ArG;e�G;�XH;��H;sI;�VI;��I;�I;��I;ÔI;�I; rI;�_I;TOI;�@I;�3I;(I;I;�I;2I;�I;jI;��H;�H;��H;a�H;?�H;q�H;#�H;9�H;|�H;�H;�H;�H;|�H;9�H;#�H;q�H;?�H;a�H;��H;�H;��H;jI;�I;2I;�I;I;(I;�3I;�@I;TOI;�_I; rI;�I;ÔI;��I;�I;��I;�VI;sI;��H;�XH;e�G;ArG;tG;�F;yF;      C�H;��H;@�H;I;�$I;kGI;�gI;.�I;\�I;؜I;�I;ÓI;�I;�uI;;eI;�UI;�GI;";I;�/I;D%I;"I;LI;gI;iI;QI;��H;�H;��H;s�H;@�H;{�H; �H;��H;�H;q�H;�H;�H;�H;q�H;�H;��H; �H;{�H;@�H;s�H;��H;�H;��H;QI;iI;gI;LI;"I;D%I;�/I;";I;�GI;�UI;;eI;�uI;�I;ÓI;�I;؜I;\�I;.�I;�gI;kGI;�$I;I;@�H;��H;      ��I;�I; �I;Z�I;јI;ΜI;G�I;A�I;r�I;�I;րI;3sI;PeI;�WI;^KI;�?I;�4I;�*I;�!I;�I;�I;QI;�I;�I;��H;�H;��H;k�H;Q�H;j�H;��H;��H;��H;�H;��H;H�H;1�H;H�H;��H;�H;��H;��H;��H;j�H;Q�H;k�H;��H;�H;��H;�I;�I;QI;�I;�I;�!I;�*I;�4I;�?I;^KI;�WI;PeI;3sI;րI;�I;r�I;A�I;G�I;ΜI;јI;Z�I; �I;�I;      ��I;�I;ۙI;��I;�I;ǎI;ڇI;UI;ruI;�jI;	`I;IUI;�JI;�@I;7I;�-I;y%I;�I;�I;bI;�
I;�I;4I;Y�H;��H;��H;s�H;Q�H;i�H;��H;��H;��H;��H;,�H;��H;��H;Y�H;��H;��H;,�H;��H;��H;��H;��H;i�H;Q�H;s�H;��H;��H;Y�H;4I;�I;�
I;bI;�I;�I;y%I;�-I;7I;�@I;�JI;IUI;	`I;�jI;ruI;UI;ڇI;ǎI;�I;��I;ۙI;�I;      8{I;�zI;�xI;�uI;#qI;�kI;FeI;=^I;�VI;�NI;�FI;}>I;m6I;�.I;�&I; I;�I;�I;I;�I;\I;L I;��H;s�H;��H;a�H;@�H;j�H;��H;��H;��H;��H;�H;��H;�H;��H;��H;��H;�H;��H;�H;��H;��H;��H;��H;j�H;@�H;a�H;��H;s�H;��H;L I;\I;�I;I;�I;�I; I;�&I;�.I;m6I;}>I;�FI;�NI;�VI;=^I;FeI;�kI;#qI;�uI;�xI;�zI;      �ZI;rZI;�XI;qVI;6SI;OI;@JI;�DI;O?I;F9I;3I;�,I;�&I;� I;�I;uI;QI;nI;I;I;b�H;�H;�H;q�H;.�H;?�H;{�H;��H;��H;��H;��H;��H;_�H;��H;|�H;c�H;Z�H;c�H;|�H;��H;_�H;��H;��H;��H;��H;��H;{�H;?�H;.�H;q�H;�H;�H;b�H;I;I;nI;QI;uI;�I;� I;�&I;�,I;3I;F9I;O?I;�DI;@JI;OI;6SI;qVI;�XI;rZI;      �BI;yBI;bAI;�?I;=I;�9I;E6I;%2I;�-I;)I;B$I;�I;�I;�I;�I;'I;	I;EI;�I;O�H;]�H;��H;F�H;:�H;0�H;q�H; �H;��H;��H;��H;��H;I�H;��H;U�H;�H;��H;��H;��H;�H;U�H;��H;I�H;��H;��H;��H;��H; �H;q�H;0�H;:�H;F�H;��H;]�H;O�H;�I;EI;	I;'I;�I;�I;�I;�I;B$I;)I;�-I;%2I;E6I;�9I;=I;�?I;bAI;yBI;      #1I;�0I;�/I;�.I;�,I;3*I;a'I;<$I;� I;=I;�I;�I;�I;I;h
I;�I;�I;� I;��H;��H;h�H;*�H;�H;L�H;��H;#�H;��H;��H;��H;�H;_�H;��H;8�H;��H;��H;��H;t�H;��H;��H;��H;8�H;��H;_�H;�H;��H;��H;��H;#�H;��H;L�H;�H;*�H;h�H;��H;��H;� I;�I;�I;h
I;I;�I;�I;�I;=I;� I;<$I;a'I;3*I;�,I;�.I;�/I;�0I;      �$I;s$I;�#I;�"I;0!I;8I;�I;bI;�I;�I;�I;xI;uI;oI;cI;�I;��H;��H;s�H;I�H;L�H;M�H;z�H;��H;}�H;9�H;�H;�H;,�H;��H;��H;U�H;��H;��H;b�H;@�H;(�H;@�H;b�H;��H;��H;U�H;��H;��H;,�H;�H;�H;9�H;}�H;��H;z�H;M�H;L�H;I�H;s�H;��H;��H;�I;cI;oI;uI;xI;�I;�I;�I;bI;�I;8I;0!I;�"I;�#I;s$I;      �I;EI;�I;�I;nI;�I;I;�I;yI;I;vI;�	I;/I;I;�I;i�H;�H;��H;��H;��H;��H;��H;o�H;��H;��H;|�H;q�H;��H;��H;�H;|�H;�H;��H;b�H;�H;�H;�H;�H;�H;b�H;��H;�H;|�H;�H;��H;��H;q�H;|�H;��H;��H;o�H;��H;��H;��H;��H;��H;�H;i�H;�I;I;/I;�	I;vI;I;yI;�I;I;�I;nI;�I;�I;EI;      �I;tI;�I;'I;I;�I;�I;I;�I;�I;h	I;I;�I;<I;��H;��H;i�H;d�H;r�H;��H;��H;�H;��H;i�H;,�H;�H;�H;H�H;��H;��H;c�H;��H;��H;@�H;�H;��H;��H;��H;�H;@�H;��H;��H;c�H;��H;��H;H�H;�H;�H;,�H;i�H;��H;�H;��H;��H;r�H;d�H;i�H;��H;��H;<I;�I;I;h	I;�I;�I;I;�I;�I;I;'I;�I;tI;      NI; I;�I;�I;�I;KI;�I;�I;�I;�
I;iI;.I;�I;�I;l�H;�H;��H;��H;��H;1�H;��H;��H;b�H;�H;	�H;�H;�H;1�H;Y�H;��H;Z�H;��H;t�H;(�H;�H;��H;��H;��H;�H;(�H;t�H;��H;Z�H;��H;Y�H;1�H;�H;�H;	�H;�H;b�H;��H;��H;1�H;��H;��H;��H;�H;l�H;�I;�I;.I;iI;�
I;�I;�I;�I;KI;�I;�I;�I; I;      �I;tI;�I;'I;I;�I;�I;I;�I;�I;h	I;I;�I;<I;��H;��H;i�H;d�H;r�H;��H;��H;�H;��H;i�H;,�H;�H;�H;H�H;��H;��H;c�H;��H;��H;@�H;�H;��H;��H;��H;�H;@�H;��H;��H;c�H;��H;��H;H�H;�H;�H;,�H;i�H;��H;�H;��H;��H;r�H;d�H;i�H;��H;��H;<I;�I;I;h	I;�I;�I;I;�I;�I;I;'I;�I;tI;      �I;EI;�I;�I;nI;�I;I;�I;yI;I;vI;�	I;/I;I;�I;i�H;�H;��H;��H;��H;��H;��H;o�H;��H;��H;|�H;q�H;��H;��H;�H;|�H;�H;��H;b�H;�H;�H;�H;�H;�H;b�H;��H;�H;|�H;�H;��H;��H;q�H;|�H;��H;��H;o�H;��H;��H;��H;��H;��H;�H;i�H;�I;I;/I;�	I;vI;I;yI;�I;I;�I;nI;�I;�I;EI;      �$I;s$I;�#I;�"I;0!I;8I;�I;bI;�I;�I;�I;xI;uI;oI;cI;�I;��H;��H;s�H;I�H;L�H;M�H;z�H;��H;}�H;9�H;�H;�H;,�H;��H;��H;U�H;��H;��H;b�H;@�H;(�H;@�H;b�H;��H;��H;U�H;��H;��H;,�H;�H;�H;9�H;}�H;��H;z�H;M�H;L�H;I�H;s�H;��H;��H;�I;cI;oI;uI;xI;�I;�I;�I;bI;�I;8I;0!I;�"I;�#I;s$I;      #1I;�0I;�/I;�.I;�,I;3*I;a'I;<$I;� I;=I;�I;�I;�I;I;h
I;�I;�I;� I;��H;��H;h�H;*�H;�H;L�H;��H;#�H;��H;��H;��H;�H;_�H;��H;8�H;��H;��H;��H;t�H;��H;��H;��H;8�H;��H;_�H;�H;��H;��H;��H;#�H;��H;L�H;�H;*�H;h�H;��H;��H;� I;�I;�I;h
I;I;�I;�I;�I;=I;� I;<$I;a'I;3*I;�,I;�.I;�/I;�0I;      �BI;yBI;bAI;�?I;=I;�9I;E6I;%2I;�-I;)I;B$I;�I;�I;�I;�I;'I;	I;EI;�I;O�H;]�H;��H;F�H;:�H;0�H;q�H; �H;��H;��H;��H;��H;I�H;��H;U�H;�H;��H;��H;��H;�H;U�H;��H;I�H;��H;��H;��H;��H; �H;q�H;0�H;:�H;F�H;��H;]�H;O�H;�I;EI;	I;'I;�I;�I;�I;�I;B$I;)I;�-I;%2I;E6I;�9I;=I;�?I;bAI;yBI;      �ZI;rZI;�XI;qVI;6SI;OI;@JI;�DI;O?I;F9I;3I;�,I;�&I;� I;�I;uI;QI;nI;I;I;b�H;�H;�H;q�H;.�H;?�H;{�H;��H;��H;��H;��H;��H;_�H;��H;|�H;c�H;Z�H;c�H;|�H;��H;_�H;��H;��H;��H;��H;��H;{�H;?�H;.�H;q�H;�H;�H;b�H;I;I;nI;QI;uI;�I;� I;�&I;�,I;3I;F9I;O?I;�DI;@JI;OI;6SI;qVI;�XI;rZI;      8{I;�zI;�xI;�uI;#qI;�kI;FeI;=^I;�VI;�NI;�FI;}>I;m6I;�.I;�&I; I;�I;�I;I;�I;\I;L I;��H;s�H;��H;a�H;@�H;j�H;��H;��H;��H;��H;�H;��H;�H;��H;��H;��H;�H;��H;�H;��H;��H;��H;��H;j�H;@�H;a�H;��H;s�H;��H;L I;\I;�I;I;�I;�I; I;�&I;�.I;m6I;}>I;�FI;�NI;�VI;=^I;FeI;�kI;#qI;�uI;�xI;�zI;      ��I;�I;ۙI;��I;�I;ǎI;ڇI;UI;ruI;�jI;	`I;IUI;�JI;�@I;7I;�-I;y%I;�I;�I;bI;�
I;�I;4I;Y�H;��H;��H;s�H;Q�H;i�H;��H;��H;��H;��H;,�H;��H;��H;Y�H;��H;��H;,�H;��H;��H;��H;��H;i�H;Q�H;s�H;��H;��H;Y�H;4I;�I;�
I;bI;�I;�I;y%I;�-I;7I;�@I;�JI;IUI;	`I;�jI;ruI;UI;ڇI;ǎI;�I;��I;ۙI;�I;      ��I;�I; �I;Z�I;јI;ΜI;G�I;A�I;r�I;�I;րI;3sI;PeI;�WI;^KI;�?I;�4I;�*I;�!I;�I;�I;QI;�I;�I;��H;�H;��H;k�H;Q�H;j�H;��H;��H;��H;�H;��H;H�H;1�H;H�H;��H;�H;��H;��H;��H;j�H;Q�H;k�H;��H;�H;��H;�I;�I;QI;�I;�I;�!I;�*I;�4I;�?I;^KI;�WI;PeI;3sI;րI;�I;r�I;A�I;G�I;ΜI;јI;Z�I; �I;�I;      C�H;��H;@�H;I;�$I;kGI;�gI;.�I;\�I;؜I;�I;ÓI;�I;�uI;;eI;�UI;�GI;";I;�/I;D%I;"I;LI;gI;iI;QI;��H;�H;��H;s�H;@�H;{�H; �H;��H;�H;q�H;�H;�H;�H;q�H;�H;��H; �H;{�H;@�H;s�H;��H;�H;��H;QI;iI;gI;LI;"I;D%I;�/I;";I;�GI;�UI;;eI;�uI;�I;ÓI;�I;؜I;\�I;.�I;�gI;kGI;�$I;I;@�H;��H;      �eF;yF;�F;tG;ArG;e�G;�XH;��H;sI;�VI;��I;�I;��I;ÔI;�I; rI;�_I;TOI;�@I;�3I;(I;I;�I;2I;�I;jI;��H;�H;��H;a�H;?�H;q�H;#�H;9�H;|�H;�H;�H;�H;|�H;9�H;#�H;q�H;?�H;a�H;��H;�H;��H;jI;�I;2I;�I;I;(I;�3I;�@I;TOI;�_I; rI;�I;ÔI;��I;�I;��I;�VI;sI;��H;�XH;e�G;ArG;tG;�F;yF;      T?@;ho@;��@;��A;��B;JD;�DE;HfF;�cG;2H;{�H;8I;WxI;�I;��I;��I;o}I;�hI;�UI;*EI;�6I;*I;VI;5I;tI;�I;QI;��H;��H;��H;.�H;0�H;��H;}�H;��H;,�H;	�H;,�H;��H;}�H;��H;0�H;.�H;��H;��H;��H;QI;�I;tI;5I;VI;*I;�6I;*EI;�UI;�hI;o}I;��I;��I;�I;WxI;8I;{�H;2H;�cG;HfF;�DE;JD;��B;��A;��@;ho@;      ��2;V$3;�T4;e06;��8;-6;;��=;�@;�C;aE;2�F;��G;ϸH;};I;�I;��I;2�I;P�I;�oI;�ZI;QHI;�8I;6+I;�I;5I;2I;iI;�I;Y�H;s�H;q�H;:�H;L�H;��H;��H;i�H;�H;i�H;��H;��H;L�H;:�H;q�H;s�H;Y�H;�I;iI;2I;5I;�I;6+I;�8I;QHI;�ZI;�oI;P�I;2�I;��I;�I;};I;ϸH;��G;2�F;aE;�C;�@;��=;-6;;��8;e06;�T4;V$3;      ��;�;M;�;΢#;�);��.;�V4;B{9;\�=;M�A;��D;��F;�H;��H;�^I;ߒI;l�I;g�I;�tI;�]I;�II;=9I;6+I;VI;�I;gI;�I;4I;��H;�H;F�H;�H;z�H;o�H;��H;b�H;��H;o�H;z�H;�H;F�H;�H;��H;4I;�I;gI;�I;VI;6+I;=9I;�II;�]I;�tI;g�I;l�I;ߒI;�^I;��H;�H;��F;��D;M�A;\�=;B{9;�V4;��.;�);΢#;�;M;�;      ���:{��:���:��:�)�:��;��;˧;ο&;o�/;Y<7;nC=;��A;�E;^6G;w�H;�7I;	�I;#�I;��I;wI;�^I;�II;�8I;*I;I;LI;QI;�I;L I;�H;��H;*�H;M�H;��H;�H;��H;�H;��H;M�H;*�H;��H;�H;L I;�I;QI;LI;I;*I;�8I;�II;�^I;wI;��I;#�I;	�I;�7I;w�H;^6G;�E;��A;nC=;Y<7;o�/;ο&;˧;��;��;�)�:��:���:{��:      �sx9���9ޤ�9�:F�^:���:�Ǽ:�N�:��;�g;�#;�;/;�:8;��>;�nC;�eF;W'H;eI;�~I;ߛI;ːI;wI;�]I;QHI;�6I;(I;"I;�I;�
I;\I;b�H;]�H;h�H;L�H;��H;��H;��H;��H;��H;L�H;h�H;]�H;b�H;\I;�
I;�I;"I;(I;�6I;QHI;�]I;wI;ːI;ߛI;�~I;eI;W'H;�eF;�nC;��>;�:8;�;/;�#;�g;��;�N�:�Ǽ:���:F�^:�:ޤ�9���9      ��f�����-�ht�+N���8&�&:J��:I��:�Y;[B;N�&;�&3;5<;��A;��E;��G;\I;v{I;ߛI;��I;�tI;�ZI;*EI;�3I;D%I;�I;bI;�I;I;O�H;��H;I�H;��H;��H;1�H;��H;��H;I�H;��H;O�H;I;�I;bI;�I;D%I;�3I;*EI;�ZI;�tI;��I;ߛI;v{I;\I;��G;��E;��A;5<;�&3;N�&;[B;�Y;I��:J��:&�&:��8+N�ht�-���f���      �N����������g���8}�g�D���� z�����I��9�
�:���:%	;,�;�.;�9;�@;]E;��G;\I;�~I;#�I;g�I;�oI;�UI;�@I;�/I;�!I;�I;I;I;�I;��H;s�H;��H;r�H;��H;r�H;��H;s�H;��H;�I;I;I;�I;�!I;�/I;�@I;�UI;�oI;g�I;#�I;�~I;\I;��G;]E;�@;�9;�.;,�;%	;���:�
�:I��9��� z�����g�D��8}��g���������      *�?��<<�@�1�;i!��z�RC����ko��{�-�1򳺵���q�&:���:Y��:��;6�+;�8;W�@;]E;��G;eI;	�I;l�I;P�I;�hI;TOI;";I;�*I;�I;�I;nI;EI;� I;��H;��H;d�H;��H;d�H;��H;��H;� I;EI;nI;�I;�I;�*I;";I;TOI;�hI;P�I;l�I;	�I;eI;��G;]E;W�@;�8;6�+;��;Y��:���:q�&:����1�{�-�ko�����RC��z�;i!�@�1��<<�      ���p���I���������W�^�85��z��̻t숻�S��gt�E�x9b��:�k�:�g;y�*;�8;�@;��E;W'H;�7I;ߒI;2�I;o}I;�_I;�GI;�4I;y%I;�I;QI;	I;�I;��H;�H;i�H;��H;i�H;�H;��H;�I;	I;QI;�I;y%I;�4I;�GI;�_I;o}I;2�I;ߒI;�7I;W'H;��E;�@;�8;y�*;�g;�k�:b��:E�x9�gt��S�t숻�̻�z�85�W�^���������I��p��      6��p��
�*���z��fC���t�� �|��?�Ъ	������V�񮼺rU��߄:��:�g;6�+;�9;��A;�eF;w�H;�^I;��I;��I; rI;�UI;�?I;�-I; I;uI;'I;�I;�I;i�H;��H;�H;��H;i�H;�I;�I;'I;uI; I;�-I;�?I;�UI; rI;��I;��I;�^I;w�H;�eF;��A;�9;6�+;�g;��:�߄:rU�񮼺��V����Ъ	��?� �|��t��fC��z��*����
�p�      ��t���p�9�d�-�Q���9�l*������Ҽ�I��O�o���'���ڻX7}� ��vH��߄:�k�:��;�.;5<;�nC;^6G;��H;�I;��I;�I;;eI;^KI;7I;�&I;�I;�I;h
I;cI;�I;��H;l�H;��H;�I;cI;h
I;�I;�I;�&I;7I;^KI;;eI;�I;��I;�I;��H;^6G;�nC;5<;�.;��;�k�:�߄:vH� ��X7}���ڻ��'�O�o��I����Ҽ���l*���9�-�Q�9�d���p�      ��Ž9���̷�V���z����}�$�Q�c�'����EC��I\��j<<�?��n�� ��rU�b��:Y��:,�;�&3;��>;�E;�H;};I;�I;ÔI;�uI;�WI;�@I;�.I;� I;�I;I;oI;I;<I;�I;<I;I;oI;I;�I;� I;�.I;�@I;�WI;�uI;ÔI;�I;};I;�H;�E;��>;�&3;,�;Y��:b��:rU� ���n��?�j<<�I\��EC�����c�'�$�Q���}��z��V��̷�9���      c.��3�ɤ�W����҈Ž<5�����fG�@��kּe���:yC�?�X7}�񮼺E�x9���:%	;N�&;�:8;��A;��F;ϸH;WxI;��I;�I;PeI;�JI;m6I;�&I;�I;�I;uI;/I;�I;�I;�I;/I;uI;�I;�I;�&I;m6I;�JI;PeI;�I;��I;WxI;ϸH;��F;��A;�:8;N�&;%	;���:E�x9񮼺X7}�?�:yC�e���kּ@��fG����<5��҈Ž��W��ɤ��3�      Fx��s��d�M�N�`�3�}I����L����z����\�P*�'�ݼe���j<<���ڻ��V��gt�q�&:���:[B;�;/;nC=;��D;��G;8I;�I;ÓI;3sI;IUI;}>I;�,I;�I;�I;xI;�	I;I;.I;I;�	I;xI;�I;�I;�,I;}>I;IUI;3sI;ÓI;�I;8I;��G;��D;nC=;�;/;[B;���:q�&:�gt���V���ڻj<<�e���'�ݼP*���\��z��L������}I�`�3�M�N��d��s�      *l¾(��S������������d���7�y��<Sؽ[�� �d�P*�kּI\����'�����S������
�:�Y;�#;Y<7;M�A;2�F;{�H;��I;�I;րI;	`I;�FI;3I;B$I;�I;�I;vI;h	I;iI;h	I;vI;�I;�I;B$I;3I;�FI;	`I;րI;�I;��I;{�H;2�F;M�A;Y<7;�#;�Y;�
�:�����S������'�I\��kּP*� �d�[��<Sؽy����7��d���������S���(��      �V������������Ͼ�d���ǆ�C�N��3��c�[����\�@��EC��O�o�Ъ	�t숻1�I��9I��:�g;o�/;\�=;aE;2H;�VI;؜I;�I;�jI;�NI;F9I;)I;=I;�I;I;�I;�
I;�I;I;�I;=I;)I;F9I;�NI;�jI;�I;؜I;�VI;2H;aE;\�=;o�/;�g;I��:I��91�t숻Ъ	�O�o�EC��@����\�[���cཱ3�C�N��ǆ��d����Ͼ���������      ~,b���\��>M���5�9��-r��#l¾睒�"&W��3�<Sؽ�z��fG�����I���?��̻{�-����J��:��;ο&;B{9;�C;�cG;sI;\�I;r�I;ruI;�VI;O?I;�-I;� I;�I;yI;�I;�I;�I;yI;�I;� I;�-I;O?I;�VI;ruI;r�I;\�I;sI;�cG;�C;B{9;ο&;��;J��:���{�-��̻�?��I�����fG��z��<Sؽ�3�"&W�睒�#l¾-r��9����5��>M���\�      ���"��V���J䂿��\���1�����J˾睒�C�N�y��L������c�'���Ҽ �|��z�ko�� z��&�&:�N�:˧;�V4;�@;HfF;��H;.�I;A�I;UI;=^I;�DI;%2I;<$I;bI;�I;I;�I;I;�I;bI;<$I;%2I;�DI;=^I;UI;A�I;.�I;��H;HfF;�@;�V4;˧;�N�:&�&: z��ko���z� �|���Ҽc�'����L���y��C�N�睒��J˾�����1���\�J䂿V���"��      }߿�$ڿ*�ʿ�������{Ps�MX:����#l¾�ǆ���7����<5��$�Q�����t��85���������8�Ǽ:��;��.;��=;�DE;�XH;�gI;G�I;ڇI;FeI;@JI;E6I;a'I;�I;I;�I;�I;�I;I;�I;a'I;E6I;@JI;FeI;ڇI;G�I;�gI;�XH;�DE;��=;��.;��;�Ǽ:��8������85��t�����$�Q�<5�������7��ǆ�#l¾���MX:�{Ps��������*�ʿ�$ڿ      w�����p������ſ!��{Ps���1�-r���d���d�}I�҈Ž��}�l*�fC��W�^�RC�g�D�+N๩��:��;�);-6;;JD;e�G;kGI;ΜI;ǎI;�kI;OI;�9I;3*I;8I;�I;�I;KI;�I;�I;8I;3*I;�9I;OI;�kI;ǎI;ΜI;kGI;e�G;JD;-6;;�);��;���:+N�g�D�RC�W�^�fC��l*���}�҈Ž}I��d��d��-r����1�{Ps�!����ſ��꿀p����      ��7��3�Ң%�w��<����ſ�����\�9����Ͼ����`�3����z����9�z�ἷ���z��8}�ht�F�^:�)�:΢#;��8;��B;ArG;�$I;јI;�I;#qI;6SI;=I;�,I;0!I;nI;I;�I;I;nI;0!I;�,I;=I;6SI;#qI;�I;јI;�$I;ArG;��B;��8;΢#;�)�:F�^:ht��8}��z����z�Ἁ�9��z����`�3�������Ͼ9����\������ſ�<��w�Ң%��3�      (�_��+Y��lG�f.�w���꿭���J䂿��5���󾋰��M�N�W��V��-�Q�*�������;i!��g��-󳺍:��:�;e06;��A;tG;I;Z�I;��I;�uI;qVI;�?I;�.I;�"I;�I;'I;�I;'I;�I;�"I;�.I;�?I;qVI;�uI;��I;Z�I;I;tG;��A;e06;�;��:�:-��g��;i!�����*���-�Q�V��W��M�N���������5�J䂿�������w�f.��lG��+Y�      ά��}�8tf��lG�Ң%��p�*�ʿV����>M����S����d�ɤ�̷�9�d��
��I��@�1�������ޤ�9���:M;�T4;��@;�F;@�H; �I;ۙI;�xI;�XI;bAI;�/I;�#I;�I;�I;�I;�I;�I;�#I;�/I;bAI;�XI;�xI;ۙI; �I;@�H;�F;��@;�T4;M;���:ޤ�9������@�1��I���
�9�d�̷�ɤ��d�S�������>M�V���*�ʿ�p�Ң%��lG�8tf�}�      O���A���}��+Y��3�����$ڿ"����\����(���s��3�9�����p�p�p���<<����f������9{��:�;V$3;ho@;yF;��H;�I;�I;�zI;rZI;yBI;�0I;s$I;EI;tI; I;tI;EI;s$I;�0I;yBI;rZI;�zI;�I;�I;��H;yF;ho@;V$3;�;{��:���9f�������<<�p��p���p�9����3��s�(�������\�"���$ڿ����3��+Y�}�A���      ����,������Q���F�Q�Ù$�.���~�7�}�E(�>�׾�T���L+���սr����@L��jO�9�ͻ�����l8�m�:��;T�1;��?;uF;r�H;��I;��I;��I;�uI;�VI;�@I;1I;�&I;� I;I;� I;�&I;1I;�@I;�VI;�uI;��I;��I;��I;r�H;uF;��?;T�1;��;�m�:��l8���9�ͻjO�@L����r����ս�L+��T��>�׾E(�7�}�~�.���Ù$�F�Q�Q��������,��      �,��^�� P���{��K��x �����n�����w��$���Ҿf��� (���ѽٷ��7����%�K��ɻ��݀�8���:��;��1;@;��F;.I;�I;3�I;ĝI;�tI;NVI;�@I;�0I;�&I;� I;�I;� I;�&I;�0I;�@I;NVI;�tI;ĝI;3�I;�I;.I;��F;@;��1;��;���:݀�8���ɻ%�K����7�ٷ����ѽ (�f�����Ҿ�$���w�n��������x ��K��{� P��^��      ���� P�������d���;� ����㿰���#f�b��ž��z���C�ƽ40v�e5�R����o@�	���pj��Pu9]I�:=\;�63;?�@;�F;WI;��I;{�I;o�I;�rI;�TI;^?I;0I;&I;, I;LI;, I;&I;0I;^?I;�TI;�rI;o�I;{�I;��I;WI;�F;?�@;�63;=\;]I�:�Pu9pj�	����o@�R���e5�40v�C�ƽ����z�žb��#f�������� ����;���d���� P��      Q����{���d��F�Ù$�7����ɿ,蒿��K�O���j�� Zb�H�8�����a����`���&�.�!e��X�غè�9�W�:VW;�15;?�A;� G;Z6I;��I;k�I;m�I;�oI;�RI;�=I;�.I;�$I;AI;NI;AI;�$I;�.I;�=I;�RI;�oI;m�I;k�I;��I;Z6I;� G;?�A;�15;VW;�W�:è�9X�غ!e��&�.�`��������a�8���H� Zb��j��O����K�,蒿��ɿ7��Ù$��F���d��{�      F�Q��K���;�Ù$��;
��޿�����w�o,���澝���(�D������I��3�G�����N��Ǩ�2��;�����9:���:�m!;��7;ڸB;}�G;	YI;K�I;��I;ؑI;�kI;�OI;4;I;�,I;3#I;�I;�I;�I;3#I;�,I;4;I;�OI;�kI;ؑI;��I;K�I;	YI;}�G;ڸB;��7;�m!;���:��9:;���2��Ǩ��N�����3�G��I������(�D��������o,���w�����޿�;
�Ù$���;��K�      Ù$��x � ��7���޿m���ǅ����F�{�
��~����z��$���ս$���P2+���ϼXPp����K�]��*�!��:,�;�7';��:;�C;+H;�|I;?�I;��I;��I;�fI;�KI;98I;V*I;D!I;I;GI;I;D!I;V*I;98I;�KI;�fI;��I;��I;?�I;�|I;+H;�C;��:;�7';,�;!��:�*�K�]����XPp���ϼP2+�$�����ս�$���z��~��{�
���F�ǅ��m����޿7�� ���x �      .���������㿆�ɿ���ǅ����P�b��:�׾�`��U�H����@��a�a�"���"D�Hɻ�!������U�:�~;�H-;G{=;ABE;ȄH;)�I;��I;��I;ւI;�`I;BGI;�4I;�'I;�I; I;oI; I;�I;�'I;�4I;BGI;�`I;ւI;��I;��I;)�I;ȄH;ABE;G{=;�H-;�~;�U�:�����!�Hɻ"D��"��a�a��@����U�H��`��:�׾b����P�ǅ�������ɿ��㿯���      ~�n�������,蒿��w���F�b��Ȱ�����Yb�+����ѽ�%��'D4����@X��ʨ��H���轺G��9ap�:�; 93;:P@;�uF;8�H;%�I;��I;��I;�yI;�YI;2BI;�0I;�$I;dI;�I;@I;�I;dI;�$I;�0I;2BI;�YI;�yI;��I;��I;%�I;8�H;�uF;:P@; 93;�;ap�:G��9�轺�H��ʨ�@X�����'D4��%����ѽ+���Yb����Ȱ�b����F���w�,蒿����n���      7�}���w�#f���K�o,�{�
�:�׾�����k���'�lz꽥I���;V�LM�*����iO��G�opE����a�:S� ;��$;˳8;q�B;�G;UJI;1�I;9�I;a�I;*pI;�RI;�<I;�,I;%!I;�I;9I;�I;9I;�I;%!I;�,I;�<I;�RI;*pI;a�I;9�I;1�I;UJI;�G;q�B;˳8;��$;S� ;a�:���opE��G��iO�*���LM��;V��I��lz���'���k����:�׾{�
�o,���K�#f���w�      E(��$�b��O������~���`���Yb���'��U�N$��S�m�5����ϼ0�����`�����غ�0�9b��: F;�F.;3{=;aE;�[H;A�I;��I;��I;�I;%fI;%KI;7I;%(I;�I;�I;�I;DI;�I;�I;�I;%(I;7I;%KI;%fI;�I;��I;��I;A�I;�[H;aE;3{=;�F.; F;b��:�0�9��غ`������0����ϼ5��S�m�N$���U���'��Yb��`���~�����O��b���$�      >�׾��Ҿž�j��������z�U�H�+��lz�N$��0v�!2+����9�� �5�-ɻ54�0�����:���:Mn!;*O6;(kA;��F;��H;��I;��I;�I;j|I;�[I;~CI;%1I;�#I;�I;jI;�I;�I;�I;jI;�I;�#I;%1I;~CI;�[I;j|I;�I;��I;��I;��H;��F;(kA;*O6;Mn!;���:���:0��54�-ɻ �5�9�����!2+�0v�N$��lz�+��U�H���z������j��ž��Ҿ      �T��f�����z� Zb�(�D��$�����ѽ�I��S�m�!2+��������K��ﻚ�p�<������9KR�:�.;��-;��<;iyD;uH;�lI;�I;��I;��I;�nI;�QI;�;I;!+I;�I;*I;NI;�I;�I;�I;NI;*I;�I;!+I;�;I;�QI;�nI;��I;��I;�I;�lI;uH;iyD;��<;��-;�.;KR�:���9<�����p��ﻍ�K������!2+�S�m��I����ѽ���$�(�D� Zb���z�f���      �L+� (���H�������ս�@���%���;V�5���������MS�������{F��n8o�:�;��$;^7;J�A;��F;�H;��I;��I;��I;��I;uaI;�GI;-4I;A%I;HI;ZI;
I;�	I;	I;�	I;
I;ZI;HI;A%I;-4I;�GI;uaI;��I;��I;��I;��I;�H;��F;J�A;^7;��$;�;o�:�n8{F⺧������MS�������5���;V��%���@����ս����H��� (�      ��ս��ѽC�ƽ8����I��$���a�a�'D4�LM���ϼ9����K�����G��^g�w�o���:�@�:�X;��1;jk>;�
E;
/H;;pI;"�I;�I;��I; rI;�TI;>I;�,I;~I;�I;�I;�	I;.I;MI;.I;�	I;�I;�I;~I;�,I;>I;�TI; rI;��I;�I;"�I;;pI;
/H;�
E;jk>;��1;�X;�@�:��:w�o�^g��G�������K�9����ϼLM�'D4�a�a�$����I��8���C�ƽ��ѽ      r��ٷ��40v���a�3�G�P2+�"�����*���0�� �5��ﻧ��^g��ହ�g:]�:�;0H-;3f;;NC;)RG;�I;�I;@�I;�I;$�I;+bI;�HI;�4I;�%I;�I;PI;�
I;�I;eI;sI;eI;�I;�
I;PI;�I;�%I;�4I;�HI;+bI;$�I;�I;@�I;�I;�I;)RG;NC;3f;;0H-;�;]�:�g:�ହ^g������ �5�0��*������"��P2+�3�G���a�40v�ٷ��      ��7�e5���������ϼ�@X���iO����-ɻ��p�{F�w�o��g:^�:YF;�*;�9;��A;�tF;;�H;�I;��I;ȺI;d�I;�oI;SSI;n=I;9,I;�I;�I;I;pI;�I;�I;� I;�I;�I;pI;I;�I;�I;9,I;n=I;SSI;�oI;d�I;ȺI;��I;�I;;�H;�tF;��A;�9;�*;YF;^�:�g:w�o�{F⺚�p�-ɻ����iO�@X�����ϼ������e5�7�      @L�����R���`����N��XPp�"D�ʨ��G�`���54�<����n8��:]�:YF;�(;��7;u�@;��E;mPH;5lI;��I;�I;��I;B|I;�]I;�EI;�2I;�#I;zI;�I;		I;(I;� I; �H;g�H; �H;� I;(I;		I;�I;zI;�#I;�2I;�EI;�]I;B|I;��I;�I;��I;5lI;mPH;��E;u�@;��7;�(;YF;]�:��:�n8<���54�`����G�ʨ�"D�XPp��N��`���R������      jO�%�K��o@�&�.�Ǩ����Hɻ�H��opE���غ0�����9o�:�@�:�;�*;��7;�O@;�[E;H;�HI;��I;��I;)�I;|�I;YgI;�MI;z9I;W)I;�I;�I;�
I;,I;'I;G�H;r�H;��H;r�H;G�H;'I;,I;�
I;�I;�I;W)I;z9I;�MI;YgI;|�I;)�I;��I;��I;�HI;H;�[E;�O@;��7;�*;�;�@�:o�:���90����غopE��H��Hɻ���Ǩ�&�.��o@�%�K�      9�ͻ�ɻ	���!e��2��K�]��!��轺����0�9���:KR�:�;�X;0H-;�9;u�@;�[E;��G;P4I;ճI;d�I;��I;l�I;�oI;�TI;q?I;M.I;� I;�I;YI;�I;�I;6�H;��H;,�H;��H;,�H;��H;6�H;�I;�I;YI;�I;� I;M.I;q?I;�TI;�oI;l�I;��I;d�I;ճI;P4I;��G;�[E;u�@;�9;0H-;�X;�;KR�:���:�0�9����轺�!�K�]�2��!e��	����ɻ      �����pj�X�غ;����*�����G��9a�:b��:���:�.;��$;��1;3f;;��A;��E;H;P4I;W�I;��I;m�I;��I;�uI;sZI;xDI;�2I;K$I;�I;�I;hI;�I;��H;s�H;7�H;��H;��H;��H;7�H;s�H;��H;�I;hI;�I;�I;K$I;�2I;xDI;sZI;�uI;��I;m�I;��I;W�I;P4I;H;��E;��A;3f;;��1;��$;�.;���:b��:a�:G��9�����*�;���X�غpj���      ��l8݀�8�Pu9è�9��9:!��:�U�:ap�:S� ; F;Mn!;��-;^7;jk>;NC;�tF;mPH;�HI;ճI;��I;ϺI;әI;�yI;�^I;aHI;d6I;|'I;uI;�I;0
I;�I;>�H;��H;��H;�H;��H;��H;��H;�H;��H;��H;>�H;�I;0
I;�I;uI;|'I;d6I;aHI;�^I;�yI;әI;ϺI;��I;ճI;�HI;mPH;�tF;NC;jk>;^7;��-;Mn!; F;S� ;ap�:�U�:!��:��9:è�9�Pu9݀�8      �m�:���:]I�:�W�:���:,�;�~;�;��$;�F.;*O6;��<;J�A;�
E;)RG;;�H;5lI;��I;d�I;m�I;әI;�zI;�`I;�JI;�8I;�)I;�I;�I;�I;9I; I;�H;��H;{�H; �H;�H;��H;�H; �H;{�H;��H;�H; I;9I;�I;�I;�I;�)I;�8I;�JI;�`I;�zI;әI;m�I;d�I;��I;5lI;;�H;)RG;�
E;J�A;��<;*O6;�F.;��$;�;�~;,�;���:�W�:]I�:���:      ��;��;=\;VW;�m!;�7';�H-; 93;˳8;3{=;(kA;iyD;��F;
/H;�I;�I;��I;��I;��I;��I;�yI;�`I;�KI;4:I;+I;EI;8I;I;MI;� I;��H;�H;w�H;~�H;�H;a�H;2�H;a�H;�H;~�H;w�H;�H;��H;� I;MI;I;8I;EI;+I;4:I;�KI;�`I;�yI;��I;��I;��I;��I;�I;�I;
/H;��F;iyD;(kA;3{=;˳8; 93;�H-;�7';�m!;VW;=\;��;      T�1;��1;�63;�15;��7;��:;G{=;:P@;q�B;aE;��F;uH;�H;;pI;�I;��I;�I;)�I;l�I;�uI;�^I;�JI;4:I;�+I; I;+I;�I;*I;�I;�H;��H;~�H;4�H;��H;z�H;��H;��H;��H;z�H;��H;4�H;~�H;��H;�H;�I;*I;�I;+I; I;�+I;4:I;�JI;�^I;�uI;l�I;)�I;�I;��I;�I;;pI;�H;uH;��F;aE;q�B;:P@;G{=;��:;��7;�15;�63;��1;      ��?;@;?�@;?�A;ڸB;�C;ABE;�uF;�G;�[H;��H;�lI;��I;"�I;@�I;ȺI;��I;|�I;�oI;sZI;aHI;�8I;+I; I;�I;sI;�I;I;s�H;��H;��H;;�H;d�H;��H;��H;f�H;=�H;f�H;��H;��H;d�H;;�H;��H;��H;s�H;I;�I;sI;�I; I;+I;�8I;aHI;sZI;�oI;|�I;��I;ȺI;@�I;"�I;��I;�lI;��H;�[H;�G;�uF;ABE;�C;ڸB;?�A;?�@;@;      uF;��F;�F;� G;}�G;+H;ȄH;8�H;UJI;A�I;��I;�I;��I;�I;�I;d�I;B|I;YgI;�TI;xDI;d6I;�)I;EI;+I;sI;�I;ZI;��H;��H;��H;6�H;I�H;��H;j�H;��H;$�H;��H;$�H;��H;j�H;��H;I�H;6�H;��H;��H;��H;ZI;�I;sI;+I;EI;�)I;d6I;xDI;�TI;YgI;B|I;d�I;�I;�I;��I;�I;��I;A�I;UJI;8�H;ȄH;+H;}�G;� G;�F;��F;      r�H;.I;WI;Z6I;	YI;�|I;)�I;%�I;1�I;��I;��I;��I;��I;��I;$�I;�oI;�]I;�MI;q?I;�2I;|'I;�I;8I;�I;�I;ZI;��H;2�H;��H;@�H;1�H;s�H;%�H;#�H;��H;�H;��H;�H;��H;#�H;%�H;s�H;1�H;@�H;��H;2�H;��H;ZI;�I;�I;8I;�I;|'I;�2I;q?I;�MI;�]I;�oI;$�I;��I;��I;��I;��I;��I;1�I;%�I;)�I;�|I;	YI;Z6I;WI;.I;      ��I;�I;��I;��I;K�I;?�I;��I;��I;9�I;��I;�I;��I;��I; rI;+bI;SSI;�EI;z9I;M.I;K$I;uI;�I;I;*I;I;��H;2�H;�H;L�H;-�H;d�H;��H;��H;
�H;b�H;�H;��H;�H;b�H;
�H;��H;��H;d�H;-�H;L�H;�H;2�H;��H;I;*I;I;�I;uI;K$I;M.I;z9I;�EI;SSI;+bI; rI;��I;��I;�I;��I;9�I;��I;��I;?�I;K�I;��I;��I;�I;      ��I;3�I;{�I;k�I;��I;��I;��I;��I;a�I;�I;j|I;�nI;uaI;�TI;�HI;n=I;�2I;W)I;� I;�I;�I;�I;MI;�I;s�H;��H;��H;L�H;8�H;a�H;��H;��H;��H;�H;��H;<�H;4�H;<�H;��H;�H;��H;��H;��H;a�H;8�H;L�H;��H;��H;s�H;�I;MI;�I;�I;�I;� I;W)I;�2I;n=I;�HI;�TI;uaI;�nI;j|I;�I;a�I;��I;��I;��I;��I;k�I;{�I;3�I;      ��I;ĝI;o�I;m�I;ؑI;��I;ւI;�yI;*pI;%fI;�[I;�QI;�GI;>I;�4I;9,I;�#I;�I;�I;�I;0
I;9I;� I;�H;��H;��H;@�H;-�H;a�H;��H;��H;��H;��H;!�H;��H;��H;c�H;��H;��H;!�H;��H;��H;��H;��H;a�H;-�H;@�H;��H;��H;�H;� I;9I;0
I;�I;�I;�I;�#I;9,I;�4I;>I;�GI;�QI;�[I;%fI;*pI;�yI;ւI;��I;ؑI;m�I;o�I;ĝI;      �uI;�tI;�rI;�oI;�kI;�fI;�`I;�YI;�RI;%KI;~CI;�;I;-4I;�,I;�%I;�I;zI;�I;YI;hI;�I; I;��H;��H;��H;6�H;1�H;d�H;��H;��H;��H;��H;��H;c�H;�H;��H;��H;��H;�H;c�H;��H;��H;��H;��H;��H;d�H;1�H;6�H;��H;��H;��H; I;�I;hI;YI;�I;zI;�I;�%I;�,I;-4I;�;I;~CI;%KI;�RI;�YI;�`I;�fI;�kI;�oI;�rI;�tI;      �VI;NVI;�TI;�RI;�OI;�KI;BGI;2BI;�<I;7I;%1I;!+I;A%I;~I;�I;�I;�I;�
I;�I;�I;>�H;�H;�H;~�H;;�H;I�H;s�H;��H;��H;��H;��H;��H;K�H;��H;��H;J�H;P�H;J�H;��H;��H;K�H;��H;��H;��H;��H;��H;s�H;I�H;;�H;~�H;�H;�H;>�H;�I;�I;�
I;�I;�I;�I;~I;A%I;!+I;%1I;7I;�<I;2BI;BGI;�KI;�OI;�RI;�TI;NVI;      �@I;�@I;^?I;�=I;4;I;98I;�4I;�0I;�,I;%(I;�#I;�I;HI;�I;PI;I;		I;,I;�I;��H;��H;��H;w�H;4�H;d�H;��H;%�H;��H;��H;��H;��H;K�H;��H;d�H;�H;��H;��H;��H;�H;d�H;��H;K�H;��H;��H;��H;��H;%�H;��H;d�H;4�H;w�H;��H;��H;��H;�I;,I;		I;I;PI;�I;HI;�I;�#I;%(I;�,I;�0I;�4I;98I;4;I;�=I;^?I;�@I;      1I;�0I;0I;�.I;�,I;V*I;�'I;�$I;%!I;�I;�I;*I;ZI;�I;�
I;pI;(I;'I;6�H;s�H;��H;{�H;~�H;��H;��H;j�H;#�H;
�H;�H;!�H;c�H;��H;d�H;��H;��H;��H;��H;��H;��H;��H;d�H;��H;c�H;!�H;�H;
�H;#�H;j�H;��H;��H;~�H;{�H;��H;s�H;6�H;'I;(I;pI;�
I;�I;ZI;*I;�I;�I;%!I;�$I;�'I;V*I;�,I;�.I;0I;�0I;      �&I;�&I;&I;�$I;3#I;D!I;�I;dI;�I;�I;jI;NI;
I;�	I;�I;�I;� I;G�H;��H;7�H;�H; �H;�H;z�H;��H;��H;��H;b�H;��H;��H;�H;��H;�H;��H;��H;d�H;[�H;d�H;��H;��H;�H;��H;�H;��H;��H;b�H;��H;��H;��H;z�H;�H; �H;�H;7�H;��H;G�H;� I;�I;�I;�	I;
I;NI;jI;�I;�I;dI;�I;D!I;3#I;�$I;&I;�&I;      � I;� I;, I;AI;�I;I; I;�I;9I;�I;�I;�I;�	I;.I;eI;�I; �H;r�H;,�H;��H;��H;�H;a�H;��H;f�H;$�H;�H;�H;<�H;��H;��H;J�H;��H;��H;d�H;2�H;/�H;2�H;d�H;��H;��H;J�H;��H;��H;<�H;�H;�H;$�H;f�H;��H;a�H;�H;��H;��H;,�H;r�H; �H;�I;eI;.I;�	I;�I;�I;�I;9I;�I; I;I;�I;AI;, I;� I;      I;�I;LI;NI;�I;GI;oI;@I;�I;DI;�I;�I;	I;MI;sI;� I;g�H;��H;��H;��H;��H;��H;2�H;��H;=�H;��H;��H;��H;4�H;c�H;��H;P�H;��H;��H;[�H;/�H;�H;/�H;[�H;��H;��H;P�H;��H;c�H;4�H;��H;��H;��H;=�H;��H;2�H;��H;��H;��H;��H;��H;g�H;� I;sI;MI;	I;�I;�I;DI;�I;@I;oI;GI;�I;NI;LI;�I;      � I;� I;, I;AI;�I;I; I;�I;9I;�I;�I;�I;�	I;.I;eI;�I; �H;r�H;,�H;��H;��H;�H;a�H;��H;f�H;$�H;�H;�H;<�H;��H;��H;J�H;��H;��H;d�H;2�H;/�H;2�H;d�H;��H;��H;J�H;��H;��H;<�H;�H;�H;$�H;f�H;��H;a�H;�H;��H;��H;,�H;r�H; �H;�I;eI;.I;�	I;�I;�I;�I;9I;�I; I;I;�I;AI;, I;� I;      �&I;�&I;&I;�$I;3#I;D!I;�I;dI;�I;�I;jI;NI;
I;�	I;�I;�I;� I;G�H;��H;7�H;�H; �H;�H;z�H;��H;��H;��H;b�H;��H;��H;�H;��H;�H;��H;��H;d�H;[�H;d�H;��H;��H;�H;��H;�H;��H;��H;b�H;��H;��H;��H;z�H;�H; �H;�H;7�H;��H;G�H;� I;�I;�I;�	I;
I;NI;jI;�I;�I;dI;�I;D!I;3#I;�$I;&I;�&I;      1I;�0I;0I;�.I;�,I;V*I;�'I;�$I;%!I;�I;�I;*I;ZI;�I;�
I;pI;(I;'I;6�H;s�H;��H;{�H;~�H;��H;��H;j�H;#�H;
�H;�H;!�H;c�H;��H;d�H;��H;��H;��H;��H;��H;��H;��H;d�H;��H;c�H;!�H;�H;
�H;#�H;j�H;��H;��H;~�H;{�H;��H;s�H;6�H;'I;(I;pI;�
I;�I;ZI;*I;�I;�I;%!I;�$I;�'I;V*I;�,I;�.I;0I;�0I;      �@I;�@I;^?I;�=I;4;I;98I;�4I;�0I;�,I;%(I;�#I;�I;HI;�I;PI;I;		I;,I;�I;��H;��H;��H;w�H;4�H;d�H;��H;%�H;��H;��H;��H;��H;K�H;��H;d�H;�H;��H;��H;��H;�H;d�H;��H;K�H;��H;��H;��H;��H;%�H;��H;d�H;4�H;w�H;��H;��H;��H;�I;,I;		I;I;PI;�I;HI;�I;�#I;%(I;�,I;�0I;�4I;98I;4;I;�=I;^?I;�@I;      �VI;NVI;�TI;�RI;�OI;�KI;BGI;2BI;�<I;7I;%1I;!+I;A%I;~I;�I;�I;�I;�
I;�I;�I;>�H;�H;�H;~�H;;�H;I�H;s�H;��H;��H;��H;��H;��H;K�H;��H;��H;J�H;P�H;J�H;��H;��H;K�H;��H;��H;��H;��H;��H;s�H;I�H;;�H;~�H;�H;�H;>�H;�I;�I;�
I;�I;�I;�I;~I;A%I;!+I;%1I;7I;�<I;2BI;BGI;�KI;�OI;�RI;�TI;NVI;      �uI;�tI;�rI;�oI;�kI;�fI;�`I;�YI;�RI;%KI;~CI;�;I;-4I;�,I;�%I;�I;zI;�I;YI;hI;�I; I;��H;��H;��H;6�H;1�H;d�H;��H;��H;��H;��H;��H;c�H;�H;��H;��H;��H;�H;c�H;��H;��H;��H;��H;��H;d�H;1�H;6�H;��H;��H;��H; I;�I;hI;YI;�I;zI;�I;�%I;�,I;-4I;�;I;~CI;%KI;�RI;�YI;�`I;�fI;�kI;�oI;�rI;�tI;      ��I;ĝI;o�I;m�I;ؑI;��I;ւI;�yI;*pI;%fI;�[I;�QI;�GI;>I;�4I;9,I;�#I;�I;�I;�I;0
I;9I;� I;�H;��H;��H;@�H;-�H;a�H;��H;��H;��H;��H;!�H;��H;��H;c�H;��H;��H;!�H;��H;��H;��H;��H;a�H;-�H;@�H;��H;��H;�H;� I;9I;0
I;�I;�I;�I;�#I;9,I;�4I;>I;�GI;�QI;�[I;%fI;*pI;�yI;ւI;��I;ؑI;m�I;o�I;ĝI;      ��I;3�I;{�I;k�I;��I;��I;��I;��I;a�I;�I;j|I;�nI;uaI;�TI;�HI;n=I;�2I;W)I;� I;�I;�I;�I;MI;�I;s�H;��H;��H;L�H;8�H;a�H;��H;��H;��H;�H;��H;<�H;4�H;<�H;��H;�H;��H;��H;��H;a�H;8�H;L�H;��H;��H;s�H;�I;MI;�I;�I;�I;� I;W)I;�2I;n=I;�HI;�TI;uaI;�nI;j|I;�I;a�I;��I;��I;��I;��I;k�I;{�I;3�I;      ��I;�I;��I;��I;K�I;?�I;��I;��I;9�I;��I;�I;��I;��I; rI;+bI;SSI;�EI;z9I;M.I;K$I;uI;�I;I;*I;I;��H;2�H;�H;L�H;-�H;d�H;��H;��H;
�H;b�H;�H;��H;�H;b�H;
�H;��H;��H;d�H;-�H;L�H;�H;2�H;��H;I;*I;I;�I;uI;K$I;M.I;z9I;�EI;SSI;+bI; rI;��I;��I;�I;��I;9�I;��I;��I;?�I;K�I;��I;��I;�I;      r�H;.I;WI;Z6I;	YI;�|I;)�I;%�I;1�I;��I;��I;��I;��I;��I;$�I;�oI;�]I;�MI;q?I;�2I;|'I;�I;8I;�I;�I;ZI;��H;2�H;��H;@�H;1�H;s�H;%�H;#�H;��H;�H;��H;�H;��H;#�H;%�H;s�H;1�H;@�H;��H;2�H;��H;ZI;�I;�I;8I;�I;|'I;�2I;q?I;�MI;�]I;�oI;$�I;��I;��I;��I;��I;��I;1�I;%�I;)�I;�|I;	YI;Z6I;WI;.I;      uF;��F;�F;� G;}�G;+H;ȄH;8�H;UJI;A�I;��I;�I;��I;�I;�I;d�I;B|I;YgI;�TI;xDI;d6I;�)I;EI;+I;sI;�I;ZI;��H;��H;��H;6�H;I�H;��H;j�H;��H;$�H;��H;$�H;��H;j�H;��H;I�H;6�H;��H;��H;��H;ZI;�I;sI;+I;EI;�)I;d6I;xDI;�TI;YgI;B|I;d�I;�I;�I;��I;�I;��I;A�I;UJI;8�H;ȄH;+H;}�G;� G;�F;��F;      ��?;@;?�@;?�A;ڸB;�C;ABE;�uF;�G;�[H;��H;�lI;��I;"�I;@�I;ȺI;��I;|�I;�oI;sZI;aHI;�8I;+I; I;�I;sI;�I;I;s�H;��H;��H;;�H;d�H;��H;��H;f�H;=�H;f�H;��H;��H;d�H;;�H;��H;��H;s�H;I;�I;sI;�I; I;+I;�8I;aHI;sZI;�oI;|�I;��I;ȺI;@�I;"�I;��I;�lI;��H;�[H;�G;�uF;ABE;�C;ڸB;?�A;?�@;@;      T�1;��1;�63;�15;��7;��:;G{=;:P@;q�B;aE;��F;uH;�H;;pI;�I;��I;�I;)�I;l�I;�uI;�^I;�JI;4:I;�+I; I;+I;�I;*I;�I;�H;��H;~�H;4�H;��H;z�H;��H;��H;��H;z�H;��H;4�H;~�H;��H;�H;�I;*I;�I;+I; I;�+I;4:I;�JI;�^I;�uI;l�I;)�I;�I;��I;�I;;pI;�H;uH;��F;aE;q�B;:P@;G{=;��:;��7;�15;�63;��1;      ��;��;=\;VW;�m!;�7';�H-; 93;˳8;3{=;(kA;iyD;��F;
/H;�I;�I;��I;��I;��I;��I;�yI;�`I;�KI;4:I;+I;EI;8I;I;MI;� I;��H;�H;w�H;~�H;�H;a�H;2�H;a�H;�H;~�H;w�H;�H;��H;� I;MI;I;8I;EI;+I;4:I;�KI;�`I;�yI;��I;��I;��I;��I;�I;�I;
/H;��F;iyD;(kA;3{=;˳8; 93;�H-;�7';�m!;VW;=\;��;      �m�:���:]I�:�W�:���:,�;�~;�;��$;�F.;*O6;��<;J�A;�
E;)RG;;�H;5lI;��I;d�I;m�I;әI;�zI;�`I;�JI;�8I;�)I;�I;�I;�I;9I; I;�H;��H;{�H; �H;�H;��H;�H; �H;{�H;��H;�H; I;9I;�I;�I;�I;�)I;�8I;�JI;�`I;�zI;әI;m�I;d�I;��I;5lI;;�H;)RG;�
E;J�A;��<;*O6;�F.;��$;�;�~;,�;���:�W�:]I�:���:      ��l8݀�8�Pu9è�9��9:!��:�U�:ap�:S� ; F;Mn!;��-;^7;jk>;NC;�tF;mPH;�HI;ճI;��I;ϺI;әI;�yI;�^I;aHI;d6I;|'I;uI;�I;0
I;�I;>�H;��H;��H;�H;��H;��H;��H;�H;��H;��H;>�H;�I;0
I;�I;uI;|'I;d6I;aHI;�^I;�yI;әI;ϺI;��I;ճI;�HI;mPH;�tF;NC;jk>;^7;��-;Mn!; F;S� ;ap�:�U�:!��:��9:è�9�Pu9݀�8      �����pj�X�غ;����*�����G��9a�:b��:���:�.;��$;��1;3f;;��A;��E;H;P4I;W�I;��I;m�I;��I;�uI;sZI;xDI;�2I;K$I;�I;�I;hI;�I;��H;s�H;7�H;��H;��H;��H;7�H;s�H;��H;�I;hI;�I;�I;K$I;�2I;xDI;sZI;�uI;��I;m�I;��I;W�I;P4I;H;��E;��A;3f;;��1;��$;�.;���:b��:a�:G��9�����*�;���X�غpj���      9�ͻ�ɻ	���!e��2��K�]��!��轺����0�9���:KR�:�;�X;0H-;�9;u�@;�[E;��G;P4I;ճI;d�I;��I;l�I;�oI;�TI;q?I;M.I;� I;�I;YI;�I;�I;6�H;��H;,�H;��H;,�H;��H;6�H;�I;�I;YI;�I;� I;M.I;q?I;�TI;�oI;l�I;��I;d�I;ճI;P4I;��G;�[E;u�@;�9;0H-;�X;�;KR�:���:�0�9����轺�!�K�]�2��!e��	����ɻ      jO�%�K��o@�&�.�Ǩ����Hɻ�H��opE���غ0�����9o�:�@�:�;�*;��7;�O@;�[E;H;�HI;��I;��I;)�I;|�I;YgI;�MI;z9I;W)I;�I;�I;�
I;,I;'I;G�H;r�H;��H;r�H;G�H;'I;,I;�
I;�I;�I;W)I;z9I;�MI;YgI;|�I;)�I;��I;��I;�HI;H;�[E;�O@;��7;�*;�;�@�:o�:���90����غopE��H��Hɻ���Ǩ�&�.��o@�%�K�      @L�����R���`����N��XPp�"D�ʨ��G�`���54�<����n8��:]�:YF;�(;��7;u�@;��E;mPH;5lI;��I;�I;��I;B|I;�]I;�EI;�2I;�#I;zI;�I;		I;(I;� I; �H;g�H; �H;� I;(I;		I;�I;zI;�#I;�2I;�EI;�]I;B|I;��I;�I;��I;5lI;mPH;��E;u�@;��7;�(;YF;]�:��:�n8<���54�`����G�ʨ�"D�XPp��N��`���R������      ��7�e5���������ϼ�@X���iO����-ɻ��p�{F�w�o��g:^�:YF;�*;�9;��A;�tF;;�H;�I;��I;ȺI;d�I;�oI;SSI;n=I;9,I;�I;�I;I;pI;�I;�I;� I;�I;�I;pI;I;�I;�I;9,I;n=I;SSI;�oI;d�I;ȺI;��I;�I;;�H;�tF;��A;�9;�*;YF;^�:�g:w�o�{F⺚�p�-ɻ����iO�@X�����ϼ������e5�7�      r��ٷ��40v���a�3�G�P2+�"�����*���0�� �5��ﻧ��^g��ହ�g:]�:�;0H-;3f;;NC;)RG;�I;�I;@�I;�I;$�I;+bI;�HI;�4I;�%I;�I;PI;�
I;�I;eI;sI;eI;�I;�
I;PI;�I;�%I;�4I;�HI;+bI;$�I;�I;@�I;�I;�I;)RG;NC;3f;;0H-;�;]�:�g:�ହ^g������ �5�0��*������"��P2+�3�G���a�40v�ٷ��      ��ս��ѽC�ƽ8����I��$���a�a�'D4�LM���ϼ9����K�����G��^g�w�o���:�@�:�X;��1;jk>;�
E;
/H;;pI;"�I;�I;��I; rI;�TI;>I;�,I;~I;�I;�I;�	I;.I;MI;.I;�	I;�I;�I;~I;�,I;>I;�TI; rI;��I;�I;"�I;;pI;
/H;�
E;jk>;��1;�X;�@�:��:w�o�^g��G�������K�9����ϼLM�'D4�a�a�$����I��8���C�ƽ��ѽ      �L+� (���H�������ս�@���%���;V�5���������MS�������{F��n8o�:�;��$;^7;J�A;��F;�H;��I;��I;��I;��I;uaI;�GI;-4I;A%I;HI;ZI;
I;�	I;	I;�	I;
I;ZI;HI;A%I;-4I;�GI;uaI;��I;��I;��I;��I;�H;��F;J�A;^7;��$;�;o�:�n8{F⺧������MS�������5���;V��%���@����ս����H��� (�      �T��f�����z� Zb�(�D��$�����ѽ�I��S�m�!2+��������K��ﻚ�p�<������9KR�:�.;��-;��<;iyD;uH;�lI;�I;��I;��I;�nI;�QI;�;I;!+I;�I;*I;NI;�I;�I;�I;NI;*I;�I;!+I;�;I;�QI;�nI;��I;��I;�I;�lI;uH;iyD;��<;��-;�.;KR�:���9<�����p��ﻍ�K������!2+�S�m��I����ѽ���$�(�D� Zb���z�f���      >�׾��Ҿž�j��������z�U�H�+��lz�N$��0v�!2+����9�� �5�-ɻ54�0�����:���:Mn!;*O6;(kA;��F;��H;��I;��I;�I;j|I;�[I;~CI;%1I;�#I;�I;jI;�I;�I;�I;jI;�I;�#I;%1I;~CI;�[I;j|I;�I;��I;��I;��H;��F;(kA;*O6;Mn!;���:���:0��54�-ɻ �5�9�����!2+�0v�N$��lz�+��U�H���z������j��ž��Ҿ      E(��$�b��O������~���`���Yb���'��U�N$��S�m�5����ϼ0�����`�����غ�0�9b��: F;�F.;3{=;aE;�[H;A�I;��I;��I;�I;%fI;%KI;7I;%(I;�I;�I;�I;DI;�I;�I;�I;%(I;7I;%KI;%fI;�I;��I;��I;A�I;�[H;aE;3{=;�F.; F;b��:�0�9��غ`������0����ϼ5��S�m�N$���U���'��Yb��`���~�����O��b���$�      7�}���w�#f���K�o,�{�
�:�׾�����k���'�lz꽥I���;V�LM�*����iO��G�opE����a�:S� ;��$;˳8;q�B;�G;UJI;1�I;9�I;a�I;*pI;�RI;�<I;�,I;%!I;�I;9I;�I;9I;�I;%!I;�,I;�<I;�RI;*pI;a�I;9�I;1�I;UJI;�G;q�B;˳8;��$;S� ;a�:���opE��G��iO�*���LM��;V��I��lz���'���k����:�׾{�
�o,���K�#f���w�      ~�n�������,蒿��w���F�b��Ȱ�����Yb�+����ѽ�%��'D4����@X��ʨ��H���轺G��9ap�:�; 93;:P@;�uF;8�H;%�I;��I;��I;�yI;�YI;2BI;�0I;�$I;dI;�I;@I;�I;dI;�$I;�0I;2BI;�YI;�yI;��I;��I;%�I;8�H;�uF;:P@; 93;�;ap�:G��9�轺�H��ʨ�@X�����'D4��%����ѽ+���Yb����Ȱ�b����F���w�,蒿����n���      .���������㿆�ɿ���ǅ����P�b��:�׾�`��U�H����@��a�a�"���"D�Hɻ�!������U�:�~;�H-;G{=;ABE;ȄH;)�I;��I;��I;ւI;�`I;BGI;�4I;�'I;�I; I;oI; I;�I;�'I;�4I;BGI;�`I;ւI;��I;��I;)�I;ȄH;ABE;G{=;�H-;�~;�U�:�����!�Hɻ"D��"��a�a��@����U�H��`��:�׾b����P�ǅ�������ɿ��㿯���      Ù$��x � ��7���޿m���ǅ����F�{�
��~����z��$���ս$���P2+���ϼXPp����K�]��*�!��:,�;�7';��:;�C;+H;�|I;?�I;��I;��I;�fI;�KI;98I;V*I;D!I;I;GI;I;D!I;V*I;98I;�KI;�fI;��I;��I;?�I;�|I;+H;�C;��:;�7';,�;!��:�*�K�]����XPp���ϼP2+�$�����ս�$���z��~��{�
���F�ǅ��m����޿7�� ���x �      F�Q��K���;�Ù$��;
��޿�����w�o,���澝���(�D������I��3�G�����N��Ǩ�2��;�����9:���:�m!;��7;ڸB;}�G;	YI;K�I;��I;ؑI;�kI;�OI;4;I;�,I;3#I;�I;�I;�I;3#I;�,I;4;I;�OI;�kI;ؑI;��I;K�I;	YI;}�G;ڸB;��7;�m!;���:��9:;���2��Ǩ��N�����3�G��I������(�D��������o,���w�����޿�;
�Ù$���;��K�      Q����{���d��F�Ù$�7����ɿ,蒿��K�O���j�� Zb�H�8�����a����`���&�.�!e��X�غè�9�W�:VW;�15;?�A;� G;Z6I;��I;k�I;m�I;�oI;�RI;�=I;�.I;�$I;AI;NI;AI;�$I;�.I;�=I;�RI;�oI;m�I;k�I;��I;Z6I;� G;?�A;�15;VW;�W�:è�9X�غ!e��&�.�`��������a�8���H� Zb��j��O����K�,蒿��ɿ7��Ù$��F���d��{�      ���� P�������d���;� ����㿰���#f�b��ž��z���C�ƽ40v�e5�R����o@�	���pj��Pu9]I�:=\;�63;?�@;�F;WI;��I;{�I;o�I;�rI;�TI;^?I;0I;&I;, I;LI;, I;&I;0I;^?I;�TI;�rI;o�I;{�I;��I;WI;�F;?�@;�63;=\;]I�:�Pu9pj�	����o@�R���e5�40v�C�ƽ����z�žb��#f�������� ����;���d���� P��      �,��^�� P���{��K��x �����n�����w��$���Ҿf��� (���ѽٷ��7����%�K��ɻ��݀�8���:��;��1;@;��F;.I;�I;3�I;ĝI;�tI;NVI;�@I;�0I;�&I;� I;�I;� I;�&I;�0I;�@I;NVI;�tI;ĝI;3�I;�I;.I;��F;@;��1;��;���:݀�8���ɻ%�K����7�ٷ����ѽ (�f�����Ҿ�$���w�n��������x ��K��{� P��^��      A(��o'���o��L�d��X1�|x�Ŀ����3�v���x����4�s��b+���'�"�ü�yY�mlٻq&���p�W��:^;��0;��?;�F;tI;�I;��I;H�I;��I;ucI;�JI;�8I;�-I;�&I;�$I;�&I;�-I;�8I;�JI;ucI;��I;H�I;��I;�I;tI;�F;��?;��0;^;W��:��p�q&�mlٻ�yY�"�ü�'�b+��s����4��x��v���3����Ŀ|x��X1�d�L��o��o'��      o'���X��c^�������]]���,�N9�3g��S�����/����o��j1��hܽ���-$��l��,}U��Ի!���-���:;�41;��?;l�F;N&I;��I;6�I;Y�I;ąI;�bI;\JI;�8I;E-I;�&I;�$I;�&I;E-I;�8I;\JI;�bI;ąI;Y�I;6�I;��I;N&I;l�F;��?;�41;;��:��-�!��Ի,}U��l���-$����hܽj1��o���྘�/�S���3g��N9���,��]]�����c^���X��      �o��c^���ē��4z�1K�e��M��$ﱿQ�v��X#���Ѿń�	�&�x�нk̀�r��������I� ǻ�5��9�
�:W�; �2;��@;�F;:I;�I;�I;��I;��I;qaI;II;�7I;~,I;�%I;�#I;�%I;~,I;�7I;II;qaI;��I;��I;�I;�I;:I;�F;��@; �2;W�;�
�:�9�5� ǻ��I�����r��k̀�x�н	�&�ń���Ѿ�X#�Q�v�$ﱿM��e��1K��4z��ē�c^��      L������4z���V��X1��<�pؿ����RZ��	�(���KUo����fy��?l�l�S����7������𺞽�9��:��;\�4;�sA;�1G;�WI;��I;r�I;)�I;�I;�^I;GI;A6I;+I;�$I;�"I;�$I;+I;A6I;GI;�^I;�I;)�I;r�I;��I;�WI;�1G;�sA;\�4;��;��:���9�𺙼����7�S��l�?l�fy�����KUo�(����	��RZ����pؿ�<��X1���V��4z�����      d��]]�1K��X1�Xf���kQ��S���Z58��A���נ���O���h什�Q�,���cߓ��� �W��~谺�":��:# ;�/7;�B;`�G;{I;�I;��I;ԦI;\{I;Y[I;hDI;;4I;X)I;Q#I;G!I;Q#I;X)I;;4I;hDI;Y[I;\{I;ԦI;��I;�I;{I;`�G;�B;�/7;# ;��:�":~谺W���� �cߓ�,����Q�h什����O��נ��A��Z58�S���kQ����Xf��X1�1K��]]�      �X1���,�e���<���2g��c_���U�˂�ՌȾ	ń�-�-�q��Y ��8�2�/?ټ��{�G"��n��O���u:�O ;�&;5":;[�C;!%H;0�I;C�I;��I;�I;�uI;�VI;AI;�1I;3'I;c!I;|I;c!I;3'I;�1I;AI;�VI;�uI;�I;��I;C�I;0�I;!%H;[�C;5":;�&;�O ;��u:�O��n�G"���{�/?ټ8�2�Y ��q��-�-�	ń�ՌȾ˂��U�c_��2g���<�e����,�      |x�N9�M��pؿkQ��c_��4�_��X#�p���f��<�S�{�����-l�T�-w��f�M�#�Ի�+��LT���:�d;�[,;/=;�AE;|�H;��I;��I;��I;֕I;�nI;�QI;/=I;{.I;�$I;I;bI;I;�$I;{.I;/=I;�QI;�nI;֕I;��I;��I;��I;|�H;�AE;/=;�[,;�d;��:�LT��+�#�Իf�M�-w��T�-l�����{�<�S��f��p���X#�4�_�c_��kQ��pؿM��N9�      Ŀ3g��$ﱿ���S����U��X#�s��d���JUo�
�#��hܽ����n<����`���Ӊ �<❻K�Ժ�l�9q��:�U;�2;�@;s�F;�I;�I;b�I;J�I;��I;$gI;.LI;�8I;+I;�!I;�I;�I;�I;�!I;+I;�8I;.LI;$gI;��I;J�I;b�I;�I;�I;s�F;�@;�2;�U;q��:�l�9K�Ժ<❻Ӊ �`�������n<�����hܽ
�#�JUo�d���s���X#��U�S������$ﱿ3g��      ���S���Q�v��RZ�Z58�˂�p��d���hoy�`1�gO��d什�`�`��7����yY���컟�T��1���u:��:[~#;-88;�B;��G;lI;,�I;!�I;L�I;��I;�^I;!FI;4I;C'I;�I;�I;)I;�I;�I;C'I;4I;!FI;�^I;��I;L�I;!�I;,�I;lI;��G;�B;-88;[~#;��:��u:�1���T���컷yY�7���`���`�d什gO��`1�hoy�d���p��˂�Z58��RZ�Q�v�S���      �3���/��X#��	��A��ՌȾ�f��JUo�`1�Ӱ���n���x��'��>ټ�@��.l�T���'���39�!�::Q; d-;�.=;�E;~wH;��I;,�I;��I;�I;5uI;�VI;�?I;/I;B#I;_I;�I;SI;�I;_I;B#I;/I;�?I;�VI;5uI;�I;��I;,�I;��I;~wH;�E;�.=; d-;:Q;�!�:�39'��T���.l��@���>ټ�'��x��n��Ӱ��`1�JUo��f��ՌȾ�A���	��X#���/�      v���ྃ�Ѿ(����נ�	ń�<�S�
�#�gO���n��R̀��2�-������>���Ի��B��#�Wm:�E�:n ;��5;�EA;��F;�I;r�I;o�I;ĽI;��I;�iI;�MI;.9I;�)I;I;�I;�I;iI;�I;�I;I;�)I;.9I;�MI;�iI;��I;ĽI;o�I;r�I;�I;��F;�EA;��5;n ;�E�:Wm:�#���B���Ի��>���-���2�R̀��n��gO��
�#�<�S�	ń��נ�(�����Ѿ��      �x���o��ń�KUo���O�-�-�{��hܽd什�x��2��b��yR���|U��2�����%찺�m�9��:C;��,;�g<;�qD;g$H;�I;��I;��I;&�I;%I;�]I;(EI;r2I;�$I;�I;}I;�I;PI;�I;}I;�I;�$I;r2I;(EI;�]I;%I;&�I;��I;��I;�I;g$H;�qD;�g<;��,;C;��:�m�9%찺����2���|U�yR���b���2��x�d什�hܽ{�-�-���O�KUo�ń��o��      ��4�j1�	�&������q�ཌྷ�������`��'�-��yR����]�����V��
[����o����:z�;<~#;/�6;msA;r�F;�I;��I;��I;��I;6�I;�oI;�RI;�<I;�+I;�I;�I;�I;`I;VI;`I;�I;�I;�I;�+I;�<I;�RI;�oI;6�I;��I;��I;��I;�I;r�F;msA;/�6;<~#;z�;���:��o�
[���V�������]�yR��-��'��`��������q�������	�&�j1�      s�ཾhܽx�нfy��h什Y ��-l��n<�`���>ټ�𛼞|U����H᝻�2�������u:hj�:�;|61;j(>;rE;+IH;p�I;��I;��I;�I;��I;zaI;�GI;G4I;~%I;�I;�I;WI;<
I;6	I;<
I;WI;�I;�I;~%I;G4I;�GI;zaI;��I;�I;��I;��I;p�I;+IH;rE;j(>;|61;�;hj�:��u:�����2�H᝻����|U����>ټ`���n<�-l�Y ��h什fy��x�н�hܽ      b+����k̀�?l��Q�8�2�T����7����@����>��2���V���2���� R:���:�;�[,;P;;;C;�dG;w8I;��I;U�I;��I;^�I;�pI;�SI;=I;W,I;KI;�I;�I;�	I;+I;'I;+I;�	I;�I;�I;KI;W,I;=I;�SI;�pI;^�I;��I;U�I;��I;w8I;�dG;;C;P;;�[,;�;���: R:���2��V���2����>��@��7������T�8�2��Q�?l�k̀���      �'��-$�r��l�,���/?ټ-w��`����yY�.l���Ի���
[������ R:���:�Q;�);�8;��A;�F;R�H;I�I;��I;��I;ȨI;$�I;�_I;GI;�3I;�$I;cI;�I;�
I;�I;*I;]I;*I;�I;�
I;�I;cI;�$I;�3I;GI;�_I;$�I;ȨI;��I;��I;I�I;R�H;�F;��A;�8;�);�Q;���: R:����
[�������Ի.l��yY�`���-w��/?ټ,���l�r���-$�      "�ü�l������S��cߓ���{�f�M�Ӊ ����T�����B�%찺��o���u:���:�Q;D�';)07;Մ@;�E;�kH;M�I;��I;��I;+�I;��I;�kI;�PI;C;I;�*I;�I;�I;|I;�I;ZI;CI;� I;CI;ZI;�I;|I;�I;�I;�*I;C;I;�PI;�kI;��I;+�I;��I;��I;M�I;�kH;�E;Մ@;)07;D�';�Q;���:��u:��o�%찺��B�T������Ӊ �f�M���{�cߓ�S�������l��      �yY�,}U���I���7��� �G"�#�Ի<❻��T�'���#��m�9���:hj�:�;�);)07;C@;U\E;�#H;�jI;'�I;r�I;�I;L�I;�vI;�YI;�BI;�0I;g"I;CI;�I;EI;�I;N I;�H;�H;�H;N I;�I;EI;�I;CI;g"I;�0I;�BI;�YI;�vI;L�I;�I;r�I;'�I;�jI;�#H;U\E;C@;)07;�);�;hj�:���:�m�9�#�'���T�<❻#�ԻG"��� ���7���I�,}U�      mlٻ�Ի ǻ����W���n��+�K�Ժ�1��39Wm:��:z�;�;�[,;�8;Մ@;U\E;�	H;iUI;��I;	�I;�I;}�I;#�I;�aI;}II;>6I;�&I;�I;GI;�	I;NI;O I;{�H;��H;��H;��H;{�H;O I;NI;�	I;GI;�I;�&I;>6I;}II;�aI;#�I;}�I;�I;	�I;��I;iUI;�	H;U\E;Մ@;�8;�[,;�;z�;��:Wm:�39�1�K�Ժ�+��n�W������ ǻ�Ի      q&�!��5���~谺�O��LT��l�9��u:�!�:�E�:C;<~#;|61;P;;��A;�E;�#H;iUI;,�I;��I;0�I;��I;�I;-hI;BOI;6;I;+I;3I;�I;�I;�I;� I;F�H;��H;��H;�H;��H;��H;F�H;� I;�I;�I;�I;3I;+I;6;I;BOI;-hI;�I;��I;0�I;��I;,�I;iUI;�#H;�E;��A;P;;|61;<~#;C;�E�:�!�:��u:�l�9�LT��O�~谺���5�!�      ��p���-��9���9�":��u:��:q��:��::Q;n ;��,;/�6;j(>;;C;�F;�kH;�jI;��I;��I;��I;3�I;��I;�lI;�SI;>?I;�.I;8!I;nI;�I;�I;�I;��H;��H;��H;c�H;��H;c�H;��H;��H;��H;�I;�I;�I;nI;8!I;�.I;>?I;�SI;�lI;��I;3�I;��I;��I;��I;�jI;�kH;�F;;C;j(>;/�6;��,;n ;:Q;��:q��:��:��u:�":���9�9��-�      W��:��:�
�:��:��:�O ;�d;�U;[~#; d-;��5;�g<;msA;rE;�dG;R�H;M�I;'�I;	�I;0�I;3�I;�I;!oI;aVI;BI;X1I;�#I;�I;�I;VI;�I;�H;��H;�H;f�H;>�H;��H;>�H;f�H;�H;��H;�H;�I;VI;�I;�I;�#I;X1I;BI;aVI;!oI;�I;3�I;0�I;	�I;'�I;M�I;R�H;�dG;rE;msA;�g<;��5; d-;[~#;�U;�d;�O ;��:��:�
�:��:      ^;;W�;��;# ;�&;�[,;�2;-88;�.=;�EA;�qD;r�F;+IH;w8I;I�I;��I;r�I;�I;��I;��I;!oI;bWI;�CI;3I;r%I;7I;�I;�	I;�I;��H;��H;��H;��H;G�H;V�H;�H;V�H;G�H;��H;��H;��H;��H;�I;�	I;�I;7I;r%I;3I;�CI;bWI;!oI;��I;��I;�I;r�I;��I;I�I;w8I;+IH;r�F;�qD;�EA;�.=;-88;�2;�[,;�&;# ;��;W�;;      ��0;�41; �2;\�4;�/7;5":;/=;�@;�B;�E;��F;g$H;�I;p�I;��I;��I;��I;�I;}�I;�I;�lI;aVI;�CI;�3I;Y&I;DI;I;�
I;II;>�H;A�H;��H;��H;��H;o�H;��H;w�H;��H;o�H;��H;��H;��H;A�H;>�H;II;�
I;I;DI;Y&I;�3I;�CI;aVI;�lI;�I;}�I;�I;��I;��I;��I;p�I;�I;g$H;��F;�E;�B;�@;/=;5":;�/7;\�4; �2;�41;      ��?;��?;��@;�sA;�B;[�C;�AE;s�F;��G;~wH;�I;�I;��I;��I;U�I;��I;+�I;L�I;#�I;-hI;�SI;BI;3I;Y&I;�I;�I;(I;�I;��H;��H;%�H;z�H;p�H;��H;��H;5�H;�H;5�H;��H;��H;p�H;z�H;%�H;��H;��H;�I;(I;�I;�I;Y&I;3I;BI;�SI;-hI;#�I;L�I;+�I;��I;U�I;��I;��I;�I;�I;~wH;��G;s�F;�AE;[�C;�B;�sA;��@;��?;      �F;l�F;�F;�1G;`�G;!%H;|�H;�I;lI;��I;r�I;��I;��I;��I;��I;ȨI;��I;�vI;�aI;BOI;>?I;X1I;r%I;DI;�I;OI;1I; I;��H;T�H;��H;c�H;��H;4�H;e�H;��H;��H;��H;e�H;4�H;��H;c�H;��H;T�H;��H; I;1I;OI;�I;DI;r%I;X1I;>?I;BOI;�aI;�vI;��I;ȨI;��I;��I;��I;��I;r�I;��I;lI;�I;|�H;!%H;`�G;�1G;�F;l�F;      tI;N&I;:I;�WI;{I;0�I;��I;�I;,�I;,�I;o�I;��I;��I;�I;^�I;$�I;�kI;�YI;}II;6;I;�.I;�#I;7I;I;(I;1I; I;��H;}�H;��H;\�H;`�H;��H;��H;�H;��H;w�H;��H;�H;��H;��H;`�H;\�H;��H;}�H;��H; I;1I;(I;I;7I;�#I;�.I;6;I;}II;�YI;�kI;$�I;^�I;�I;��I;��I;o�I;,�I;,�I;�I;��I;0�I;{I;�WI;:I;N&I;      �I;��I;�I;��I;�I;C�I;��I;b�I;!�I;��I;ĽI;&�I;6�I;��I;�pI;�_I;�PI;�BI;>6I;+I;8!I;�I;�I;�
I;�I; I;��H;y�H;��H;c�H;a�H;��H;��H;��H;��H;��H;y�H;��H;��H;��H;��H;��H;a�H;c�H;��H;y�H;��H; I;�I;�
I;�I;�I;8!I;+I;>6I;�BI;�PI;�_I;�pI;��I;6�I;&�I;ĽI;��I;!�I;b�I;��I;C�I;�I;��I;�I;��I;      ��I;6�I;�I;r�I;��I;��I;��I;J�I;L�I;�I;��I;%I;�oI;zaI;�SI;GI;C;I;�0I;�&I;3I;nI;�I;�	I;II;��H;��H;}�H;��H;X�H;[�H;��H;Z�H;K�H;��H;��H;��H;��H;��H;��H;��H;K�H;Z�H;��H;[�H;X�H;��H;}�H;��H;��H;II;�	I;�I;nI;3I;�&I;�0I;C;I;GI;�SI;zaI;�oI;%I;��I;�I;L�I;J�I;��I;��I;��I;r�I;�I;6�I;      H�I;Y�I;��I;)�I;ԦI;�I;֕I;��I;��I;5uI;�iI;�]I;�RI;�GI;=I;�3I;�*I;g"I;�I;�I;�I;VI;�I;>�H;��H;T�H;��H;c�H;[�H;��H;5�H;�H;A�H;��H;�H;��H;��H;��H;�H;��H;A�H;�H;5�H;��H;[�H;c�H;��H;T�H;��H;>�H;�I;VI;�I;�I;�I;g"I;�*I;�3I;=I;�GI;�RI;�]I;�iI;5uI;��I;��I;֕I;�I;ԦI;)�I;��I;Y�I;      ��I;ąI;��I;�I;\{I;�uI;�nI;$gI;�^I;�VI;�MI;(EI;�<I;G4I;W,I;�$I;�I;CI;GI;�I;�I;�I;��H;A�H;%�H;��H;\�H;a�H;��H;5�H;�H;�H;\�H;��H;z�H;7�H;��H;7�H;z�H;��H;\�H;�H;�H;5�H;��H;a�H;\�H;��H;%�H;A�H;��H;�I;�I;�I;GI;CI;�I;�$I;W,I;G4I;�<I;(EI;�MI;�VI;�^I;$gI;�nI;�uI;\{I;�I;��I;ąI;      ucI;�bI;qaI;�^I;Y[I;�VI;�QI;.LI;!FI;�?I;.9I;r2I;�+I;~%I;KI;cI;�I;�I;�	I;�I;�I;�H;��H;��H;z�H;c�H;`�H;��H;Z�H;�H;�H;U�H;��H;,�H;��H;��H;��H;��H;��H;,�H;��H;U�H;�H;�H;Z�H;��H;`�H;c�H;z�H;��H;��H;�H;�I;�I;�	I;�I;�I;cI;KI;~%I;�+I;r2I;.9I;�?I;!FI;.LI;�QI;�VI;Y[I;�^I;qaI;�bI;      �JI;\JI;II;GI;hDI;AI;/=I;�8I;4I;/I;�)I;�$I;�I;�I;�I;�I;|I;EI;NI;� I;��H;��H;��H;��H;p�H;��H;��H;��H;K�H;A�H;\�H;��H;�H;��H;M�H;!�H;3�H;!�H;M�H;��H;�H;��H;\�H;A�H;K�H;��H;��H;��H;p�H;��H;��H;��H;��H;� I;NI;EI;|I;�I;�I;�I;�I;�$I;�)I;/I;4I;�8I;/=I;AI;hDI;GI;II;\JI;      �8I;�8I;�7I;A6I;;4I;�1I;{.I;+I;C'I;B#I;I;�I;�I;�I;�I;�
I;�I;�I;O I;F�H;��H;�H;��H;��H;��H;4�H;��H;��H;��H;��H;��H;,�H;��H;<�H;��H;��H;��H;��H;��H;<�H;��H;,�H;��H;��H;��H;��H;��H;4�H;��H;��H;��H;�H;��H;F�H;O I;�I;�I;�
I;�I;�I;�I;�I;I;B#I;C'I;+I;{.I;�1I;;4I;A6I;�7I;�8I;      �-I;E-I;~,I;+I;X)I;3'I;�$I;�!I;�I;_I;�I;}I;�I;WI;�	I;�I;ZI;N I;{�H;��H;��H;f�H;G�H;o�H;��H;e�H;�H;��H;��H;�H;z�H;��H;M�H;��H;��H;��H;�H;��H;��H;��H;M�H;��H;z�H;�H;��H;��H;�H;e�H;��H;o�H;G�H;f�H;��H;��H;{�H;N I;ZI;�I;�	I;WI;�I;}I;�I;_I;�I;�!I;�$I;3'I;X)I;+I;~,I;E-I;      �&I;�&I;�%I;�$I;Q#I;c!I;I;�I;�I;�I;�I;�I;`I;<
I;+I;*I;CI;�H;��H;��H;c�H;>�H;V�H;��H;5�H;��H;��H;��H;��H;��H;7�H;��H;!�H;��H;��H;k�H;q�H;k�H;��H;��H;!�H;��H;7�H;��H;��H;��H;��H;��H;5�H;��H;V�H;>�H;c�H;��H;��H;�H;CI;*I;+I;<
I;`I;�I;�I;�I;�I;�I;I;c!I;Q#I;�$I;�%I;�&I;      �$I;�$I;�#I;�"I;G!I;|I;bI;�I;)I;SI;iI;PI;VI;6	I;'I;]I;� I;�H;��H;�H;��H;��H;�H;w�H;�H;��H;w�H;y�H;��H;��H;��H;��H;3�H;��H;�H;q�H;w�H;q�H;�H;��H;3�H;��H;��H;��H;��H;y�H;w�H;��H;�H;w�H;�H;��H;��H;�H;��H;�H;� I;]I;'I;6	I;VI;PI;iI;SI;)I;�I;bI;|I;G!I;�"I;�#I;�$I;      �&I;�&I;�%I;�$I;Q#I;c!I;I;�I;�I;�I;�I;�I;`I;<
I;+I;*I;CI;�H;��H;��H;c�H;>�H;V�H;��H;5�H;��H;��H;��H;��H;��H;7�H;��H;!�H;��H;��H;k�H;q�H;k�H;��H;��H;!�H;��H;7�H;��H;��H;��H;��H;��H;5�H;��H;V�H;>�H;c�H;��H;��H;�H;CI;*I;+I;<
I;`I;�I;�I;�I;�I;�I;I;c!I;Q#I;�$I;�%I;�&I;      �-I;E-I;~,I;+I;X)I;3'I;�$I;�!I;�I;_I;�I;}I;�I;WI;�	I;�I;ZI;N I;{�H;��H;��H;f�H;G�H;o�H;��H;e�H;�H;��H;��H;�H;z�H;��H;M�H;��H;��H;��H;�H;��H;��H;��H;M�H;��H;z�H;�H;��H;��H;�H;e�H;��H;o�H;G�H;f�H;��H;��H;{�H;N I;ZI;�I;�	I;WI;�I;}I;�I;_I;�I;�!I;�$I;3'I;X)I;+I;~,I;E-I;      �8I;�8I;�7I;A6I;;4I;�1I;{.I;+I;C'I;B#I;I;�I;�I;�I;�I;�
I;�I;�I;O I;F�H;��H;�H;��H;��H;��H;4�H;��H;��H;��H;��H;��H;,�H;��H;<�H;��H;��H;��H;��H;��H;<�H;��H;,�H;��H;��H;��H;��H;��H;4�H;��H;��H;��H;�H;��H;F�H;O I;�I;�I;�
I;�I;�I;�I;�I;I;B#I;C'I;+I;{.I;�1I;;4I;A6I;�7I;�8I;      �JI;\JI;II;GI;hDI;AI;/=I;�8I;4I;/I;�)I;�$I;�I;�I;�I;�I;|I;EI;NI;� I;��H;��H;��H;��H;p�H;��H;��H;��H;K�H;A�H;\�H;��H;�H;��H;M�H;!�H;3�H;!�H;M�H;��H;�H;��H;\�H;A�H;K�H;��H;��H;��H;p�H;��H;��H;��H;��H;� I;NI;EI;|I;�I;�I;�I;�I;�$I;�)I;/I;4I;�8I;/=I;AI;hDI;GI;II;\JI;      ucI;�bI;qaI;�^I;Y[I;�VI;�QI;.LI;!FI;�?I;.9I;r2I;�+I;~%I;KI;cI;�I;�I;�	I;�I;�I;�H;��H;��H;z�H;c�H;`�H;��H;Z�H;�H;�H;U�H;��H;,�H;��H;��H;��H;��H;��H;,�H;��H;U�H;�H;�H;Z�H;��H;`�H;c�H;z�H;��H;��H;�H;�I;�I;�	I;�I;�I;cI;KI;~%I;�+I;r2I;.9I;�?I;!FI;.LI;�QI;�VI;Y[I;�^I;qaI;�bI;      ��I;ąI;��I;�I;\{I;�uI;�nI;$gI;�^I;�VI;�MI;(EI;�<I;G4I;W,I;�$I;�I;CI;GI;�I;�I;�I;��H;A�H;%�H;��H;\�H;a�H;��H;5�H;�H;�H;\�H;��H;z�H;7�H;��H;7�H;z�H;��H;\�H;�H;�H;5�H;��H;a�H;\�H;��H;%�H;A�H;��H;�I;�I;�I;GI;CI;�I;�$I;W,I;G4I;�<I;(EI;�MI;�VI;�^I;$gI;�nI;�uI;\{I;�I;��I;ąI;      H�I;Y�I;��I;)�I;ԦI;�I;֕I;��I;��I;5uI;�iI;�]I;�RI;�GI;=I;�3I;�*I;g"I;�I;�I;�I;VI;�I;>�H;��H;T�H;��H;c�H;[�H;��H;5�H;�H;A�H;��H;�H;��H;��H;��H;�H;��H;A�H;�H;5�H;��H;[�H;c�H;��H;T�H;��H;>�H;�I;VI;�I;�I;�I;g"I;�*I;�3I;=I;�GI;�RI;�]I;�iI;5uI;��I;��I;֕I;�I;ԦI;)�I;��I;Y�I;      ��I;6�I;�I;r�I;��I;��I;��I;J�I;L�I;�I;��I;%I;�oI;zaI;�SI;GI;C;I;�0I;�&I;3I;nI;�I;�	I;II;��H;��H;}�H;��H;X�H;[�H;��H;Z�H;K�H;��H;��H;��H;��H;��H;��H;��H;K�H;Z�H;��H;[�H;X�H;��H;}�H;��H;��H;II;�	I;�I;nI;3I;�&I;�0I;C;I;GI;�SI;zaI;�oI;%I;��I;�I;L�I;J�I;��I;��I;��I;r�I;�I;6�I;      �I;��I;�I;��I;�I;C�I;��I;b�I;!�I;��I;ĽI;&�I;6�I;��I;�pI;�_I;�PI;�BI;>6I;+I;8!I;�I;�I;�
I;�I; I;��H;y�H;��H;c�H;a�H;��H;��H;��H;��H;��H;y�H;��H;��H;��H;��H;��H;a�H;c�H;��H;y�H;��H; I;�I;�
I;�I;�I;8!I;+I;>6I;�BI;�PI;�_I;�pI;��I;6�I;&�I;ĽI;��I;!�I;b�I;��I;C�I;�I;��I;�I;��I;      tI;N&I;:I;�WI;{I;0�I;��I;�I;,�I;,�I;o�I;��I;��I;�I;^�I;$�I;�kI;�YI;}II;6;I;�.I;�#I;7I;I;(I;1I; I;��H;}�H;��H;\�H;`�H;��H;��H;�H;��H;w�H;��H;�H;��H;��H;`�H;\�H;��H;}�H;��H; I;1I;(I;I;7I;�#I;�.I;6;I;}II;�YI;�kI;$�I;^�I;�I;��I;��I;o�I;,�I;,�I;�I;��I;0�I;{I;�WI;:I;N&I;      �F;l�F;�F;�1G;`�G;!%H;|�H;�I;lI;��I;r�I;��I;��I;��I;��I;ȨI;��I;�vI;�aI;BOI;>?I;X1I;r%I;DI;�I;OI;1I; I;��H;T�H;��H;c�H;��H;4�H;e�H;��H;��H;��H;e�H;4�H;��H;c�H;��H;T�H;��H; I;1I;OI;�I;DI;r%I;X1I;>?I;BOI;�aI;�vI;��I;ȨI;��I;��I;��I;��I;r�I;��I;lI;�I;|�H;!%H;`�G;�1G;�F;l�F;      ��?;��?;��@;�sA;�B;[�C;�AE;s�F;��G;~wH;�I;�I;��I;��I;U�I;��I;+�I;L�I;#�I;-hI;�SI;BI;3I;Y&I;�I;�I;(I;�I;��H;��H;%�H;z�H;p�H;��H;��H;5�H;�H;5�H;��H;��H;p�H;z�H;%�H;��H;��H;�I;(I;�I;�I;Y&I;3I;BI;�SI;-hI;#�I;L�I;+�I;��I;U�I;��I;��I;�I;�I;~wH;��G;s�F;�AE;[�C;�B;�sA;��@;��?;      ��0;�41; �2;\�4;�/7;5":;/=;�@;�B;�E;��F;g$H;�I;p�I;��I;��I;��I;�I;}�I;�I;�lI;aVI;�CI;�3I;Y&I;DI;I;�
I;II;>�H;A�H;��H;��H;��H;o�H;��H;w�H;��H;o�H;��H;��H;��H;A�H;>�H;II;�
I;I;DI;Y&I;�3I;�CI;aVI;�lI;�I;}�I;�I;��I;��I;��I;p�I;�I;g$H;��F;�E;�B;�@;/=;5":;�/7;\�4; �2;�41;      ^;;W�;��;# ;�&;�[,;�2;-88;�.=;�EA;�qD;r�F;+IH;w8I;I�I;��I;r�I;�I;��I;��I;!oI;bWI;�CI;3I;r%I;7I;�I;�	I;�I;��H;��H;��H;��H;G�H;V�H;�H;V�H;G�H;��H;��H;��H;��H;�I;�	I;�I;7I;r%I;3I;�CI;bWI;!oI;��I;��I;�I;r�I;��I;I�I;w8I;+IH;r�F;�qD;�EA;�.=;-88;�2;�[,;�&;# ;��;W�;;      W��:��:�
�:��:��:�O ;�d;�U;[~#; d-;��5;�g<;msA;rE;�dG;R�H;M�I;'�I;	�I;0�I;3�I;�I;!oI;aVI;BI;X1I;�#I;�I;�I;VI;�I;�H;��H;�H;f�H;>�H;��H;>�H;f�H;�H;��H;�H;�I;VI;�I;�I;�#I;X1I;BI;aVI;!oI;�I;3�I;0�I;	�I;'�I;M�I;R�H;�dG;rE;msA;�g<;��5; d-;[~#;�U;�d;�O ;��:��:�
�:��:      ��p���-��9���9�":��u:��:q��:��::Q;n ;��,;/�6;j(>;;C;�F;�kH;�jI;��I;��I;��I;3�I;��I;�lI;�SI;>?I;�.I;8!I;nI;�I;�I;�I;��H;��H;��H;c�H;��H;c�H;��H;��H;��H;�I;�I;�I;nI;8!I;�.I;>?I;�SI;�lI;��I;3�I;��I;��I;��I;�jI;�kH;�F;;C;j(>;/�6;��,;n ;:Q;��:q��:��:��u:�":���9�9��-�      q&�!��5���~谺�O��LT��l�9��u:�!�:�E�:C;<~#;|61;P;;��A;�E;�#H;iUI;,�I;��I;0�I;��I;�I;-hI;BOI;6;I;+I;3I;�I;�I;�I;� I;F�H;��H;��H;�H;��H;��H;F�H;� I;�I;�I;�I;3I;+I;6;I;BOI;-hI;�I;��I;0�I;��I;,�I;iUI;�#H;�E;��A;P;;|61;<~#;C;�E�:�!�:��u:�l�9�LT��O�~谺���5�!�      mlٻ�Ի ǻ����W���n��+�K�Ժ�1��39Wm:��:z�;�;�[,;�8;Մ@;U\E;�	H;iUI;��I;	�I;�I;}�I;#�I;�aI;}II;>6I;�&I;�I;GI;�	I;NI;O I;{�H;��H;��H;��H;{�H;O I;NI;�	I;GI;�I;�&I;>6I;}II;�aI;#�I;}�I;�I;	�I;��I;iUI;�	H;U\E;Մ@;�8;�[,;�;z�;��:Wm:�39�1�K�Ժ�+��n�W������ ǻ�Ի      �yY�,}U���I���7��� �G"�#�Ի<❻��T�'���#��m�9���:hj�:�;�);)07;C@;U\E;�#H;�jI;'�I;r�I;�I;L�I;�vI;�YI;�BI;�0I;g"I;CI;�I;EI;�I;N I;�H;�H;�H;N I;�I;EI;�I;CI;g"I;�0I;�BI;�YI;�vI;L�I;�I;r�I;'�I;�jI;�#H;U\E;C@;)07;�);�;hj�:���:�m�9�#�'���T�<❻#�ԻG"��� ���7���I�,}U�      "�ü�l������S��cߓ���{�f�M�Ӊ ����T�����B�%찺��o���u:���:�Q;D�';)07;Մ@;�E;�kH;M�I;��I;��I;+�I;��I;�kI;�PI;C;I;�*I;�I;�I;|I;�I;ZI;CI;� I;CI;ZI;�I;|I;�I;�I;�*I;C;I;�PI;�kI;��I;+�I;��I;��I;M�I;�kH;�E;Մ@;)07;D�';�Q;���:��u:��o�%찺��B�T������Ӊ �f�M���{�cߓ�S�������l��      �'��-$�r��l�,���/?ټ-w��`����yY�.l���Ի���
[������ R:���:�Q;�);�8;��A;�F;R�H;I�I;��I;��I;ȨI;$�I;�_I;GI;�3I;�$I;cI;�I;�
I;�I;*I;]I;*I;�I;�
I;�I;cI;�$I;�3I;GI;�_I;$�I;ȨI;��I;��I;I�I;R�H;�F;��A;�8;�);�Q;���: R:����
[�������Ի.l��yY�`���-w��/?ټ,���l�r���-$�      b+����k̀�?l��Q�8�2�T����7����@����>��2���V���2���� R:���:�;�[,;P;;;C;�dG;w8I;��I;U�I;��I;^�I;�pI;�SI;=I;W,I;KI;�I;�I;�	I;+I;'I;+I;�	I;�I;�I;KI;W,I;=I;�SI;�pI;^�I;��I;U�I;��I;w8I;�dG;;C;P;;�[,;�;���: R:���2��V���2����>��@��7������T�8�2��Q�?l�k̀���      s�ཾhܽx�нfy��h什Y ��-l��n<�`���>ټ�𛼞|U����H᝻�2�������u:hj�:�;|61;j(>;rE;+IH;p�I;��I;��I;�I;��I;zaI;�GI;G4I;~%I;�I;�I;WI;<
I;6	I;<
I;WI;�I;�I;~%I;G4I;�GI;zaI;��I;�I;��I;��I;p�I;+IH;rE;j(>;|61;�;hj�:��u:�����2�H᝻����|U����>ټ`���n<�-l�Y ��h什fy��x�н�hܽ      ��4�j1�	�&������q�ཌྷ�������`��'�-��yR����]�����V��
[����o����:z�;<~#;/�6;msA;r�F;�I;��I;��I;��I;6�I;�oI;�RI;�<I;�+I;�I;�I;�I;`I;VI;`I;�I;�I;�I;�+I;�<I;�RI;�oI;6�I;��I;��I;��I;�I;r�F;msA;/�6;<~#;z�;���:��o�
[���V�������]�yR��-��'��`��������q�������	�&�j1�      �x���o��ń�KUo���O�-�-�{��hܽd什�x��2��b��yR���|U��2�����%찺�m�9��:C;��,;�g<;�qD;g$H;�I;��I;��I;&�I;%I;�]I;(EI;r2I;�$I;�I;}I;�I;PI;�I;}I;�I;�$I;r2I;(EI;�]I;%I;&�I;��I;��I;�I;g$H;�qD;�g<;��,;C;��:�m�9%찺����2���|U�yR���b���2��x�d什�hܽ{�-�-���O�KUo�ń��o��      v���ྃ�Ѿ(����נ�	ń�<�S�
�#�gO���n��R̀��2�-������>���Ի��B��#�Wm:�E�:n ;��5;�EA;��F;�I;r�I;o�I;ĽI;��I;�iI;�MI;.9I;�)I;I;�I;�I;iI;�I;�I;I;�)I;.9I;�MI;�iI;��I;ĽI;o�I;r�I;�I;��F;�EA;��5;n ;�E�:Wm:�#���B���Ի��>���-���2�R̀��n��gO��
�#�<�S�	ń��נ�(�����Ѿ��      �3���/��X#��	��A��ՌȾ�f��JUo�`1�Ӱ���n���x��'��>ټ�@��.l�T���'���39�!�::Q; d-;�.=;�E;~wH;��I;,�I;��I;�I;5uI;�VI;�?I;/I;B#I;_I;�I;SI;�I;_I;B#I;/I;�?I;�VI;5uI;�I;��I;,�I;��I;~wH;�E;�.=; d-;:Q;�!�:�39'��T���.l��@���>ټ�'��x��n��Ӱ��`1�JUo��f��ՌȾ�A���	��X#���/�      ���S���Q�v��RZ�Z58�˂�p��d���hoy�`1�gO��d什�`�`��7����yY���컟�T��1���u:��:[~#;-88;�B;��G;lI;,�I;!�I;L�I;��I;�^I;!FI;4I;C'I;�I;�I;)I;�I;�I;C'I;4I;!FI;�^I;��I;L�I;!�I;,�I;lI;��G;�B;-88;[~#;��:��u:�1���T���컷yY�7���`���`�d什gO��`1�hoy�d���p��˂�Z58��RZ�Q�v�S���      Ŀ3g��$ﱿ���S����U��X#�s��d���JUo�
�#��hܽ����n<����`���Ӊ �<❻K�Ժ�l�9q��:�U;�2;�@;s�F;�I;�I;b�I;J�I;��I;$gI;.LI;�8I;+I;�!I;�I;�I;�I;�!I;+I;�8I;.LI;$gI;��I;J�I;b�I;�I;�I;s�F;�@;�2;�U;q��:�l�9K�Ժ<❻Ӊ �`�������n<�����hܽ
�#�JUo�d���s���X#��U�S������$ﱿ3g��      |x�N9�M��pؿkQ��c_��4�_��X#�p���f��<�S�{�����-l�T�-w��f�M�#�Ի�+��LT���:�d;�[,;/=;�AE;|�H;��I;��I;��I;֕I;�nI;�QI;/=I;{.I;�$I;I;bI;I;�$I;{.I;/=I;�QI;�nI;֕I;��I;��I;��I;|�H;�AE;/=;�[,;�d;��:�LT��+�#�Իf�M�-w��T�-l�����{�<�S��f��p���X#�4�_�c_��kQ��pؿM��N9�      �X1���,�e���<���2g��c_���U�˂�ՌȾ	ń�-�-�q��Y ��8�2�/?ټ��{�G"��n��O���u:�O ;�&;5":;[�C;!%H;0�I;C�I;��I;�I;�uI;�VI;AI;�1I;3'I;c!I;|I;c!I;3'I;�1I;AI;�VI;�uI;�I;��I;C�I;0�I;!%H;[�C;5":;�&;�O ;��u:�O��n�G"���{�/?ټ8�2�Y ��q��-�-�	ń�ՌȾ˂��U�c_��2g���<�e����,�      d��]]�1K��X1�Xf���kQ��S���Z58��A���נ���O���h什�Q�,���cߓ��� �W��~谺�":��:# ;�/7;�B;`�G;{I;�I;��I;ԦI;\{I;Y[I;hDI;;4I;X)I;Q#I;G!I;Q#I;X)I;;4I;hDI;Y[I;\{I;ԦI;��I;�I;{I;`�G;�B;�/7;# ;��:�":~谺W���� �cߓ�,����Q�h什����O��נ��A��Z58�S���kQ����Xf��X1�1K��]]�      L������4z���V��X1��<�pؿ����RZ��	�(���KUo����fy��?l�l�S����7������𺞽�9��:��;\�4;�sA;�1G;�WI;��I;r�I;)�I;�I;�^I;GI;A6I;+I;�$I;�"I;�$I;+I;A6I;GI;�^I;�I;)�I;r�I;��I;�WI;�1G;�sA;\�4;��;��:���9�𺙼����7�S��l�?l�fy�����KUo�(����	��RZ����pؿ�<��X1���V��4z�����      �o��c^���ē��4z�1K�e��M��$ﱿQ�v��X#���Ѿń�	�&�x�нk̀�r��������I� ǻ�5��9�
�:W�; �2;��@;�F;:I;�I;�I;��I;��I;qaI;II;�7I;~,I;�%I;�#I;�%I;~,I;�7I;II;qaI;��I;��I;�I;�I;:I;�F;��@; �2;W�;�
�:�9�5� ǻ��I�����r��k̀�x�н	�&�ń���Ѿ�X#�Q�v�$ﱿM��e��1K��4z��ē�c^��      o'���X��c^�������]]���,�N9�3g��S�����/����o��j1��hܽ���-$��l��,}U��Ի!���-���:;�41;��?;l�F;N&I;��I;6�I;Y�I;ąI;�bI;\JI;�8I;E-I;�&I;�$I;�&I;E-I;�8I;\JI;�bI;ąI;Y�I;6�I;��I;N&I;l�F;��?;�41;;��:��-�!��Ի,}U��l���-$����hܽj1��o���྘�/�S���3g��N9���,��]]�����c^���X��   