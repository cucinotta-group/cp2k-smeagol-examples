H   �V�\V�/@                        �V�\V�/@                        �V�\V�/@H      H   H   H            l����������Т��/�j��5���	� �ȿ'8����7�C�꾂S���7�	3�}L���)���Ƽ��\���ݻ+��Tɸ��:"x;��0;��?;J�F;�+I;��I;��I;սI;#�I;�hI;�NI;�<I;�0I;�)I;�'I;�)I;�0I;�<I;�NI;�hI; �I;ٽI;��I;��I;�+I;X�F;��?;��0;x;��:`Uɸ+���ݻ��\���Ƽ�)�}L��	3��7��S��C�꾨�7�'8�� �ȿ��	��5�/�j�Т����������      ��������B��^�����c�621�%X��ÿiڇ�r�3��s��7��|74�_�=ى���&�Nü$�X���ػ��%���J�҃�:�b;~�0;x�?;�F;�2I;��I;:�I;�I;I�I;QhI;�NI;1<I;y0I;b)I;�'I;^)I;|0I;0<I;�NI;ShI;E�I;�I;<�I;��I;�2I;�F;x�?;|�0;�b;̃�:@�J���%���ػ$�X�Nü��&�=ى�_�|74��7���s�r�3�iڇ��ÿ%X�621���c�^����B�����      �����B����E��w�P���#�L�������x|��'�XD־�X��o�)�Խ�Ă�I<�8_��z-M���ʻS���'�8Г�:�;!K2;v@;Q�F;�FI;k�I;�I;+�I;�I;�fI;?MI;D;I;�/I;�(I;�&I;�(I;�/I;B;I;?MI;�fI;��I;.�I;�I;n�I;�FI;]�F;v@;K2;�;̓�:�&�8P����ʻz-M�8_��I<��Ă�Խo�)��X��XD־�'��x|����L�����#�w�P�E�����B��      Т��^���E���/]��5�M���,ݿ+8��qm_��K��t��W�s�#>����8�o��3��۩���:�hT�� ���X(�9�f�:�<;�_4;hA;8G;|dI;�I;+�I;]�I;`�I;'dI;KI;�9I;J.I;�'I;�%I;�'I;M.I;�9I;KI;)dI;\�I;^�I;-�I;�I;|dI;8G;hA;�_4;�<;�f�:((�9����jT����:��۩��3�8�o����#>�W�s��t���K�qm_�+8���,ݿM���5��/]�E��^���      /�j���c�w�P��5���r��H���hڇ�Gv<�'���p���_S��������+T��� �)$���G#�̒��`1��(�:���::�;47;s�B;~�G;ćI;�I;g�I;̮I;��I;�`I;JHI;�7I;b,I;&I; $I;&I;d,I;�7I;LHI;�`I;��I;ϮI;e�I;�I;ƇI;��G;u�B;17;7�;���:�:X1��̒���G#�($���� �+T���������_S�p��'���Gv<�hڇ�H���r�����5�w�P���c�      �5�621���#�M��r���ÿ�ҕ�Z������̾�X��~�0�3�/W����5�zܼ=��W��X�s��U\���n:���:ެ%;��9;��C;�.H; �I;�I;�I;��I;y{I;\I;�DI;�4I;(*I;$I;"I;$I;)*I;�4I;�DI;\I;u{I;��I;�I;�I;�I;�.H;��C;��9;߬%;���:l�n:xU\�X�s�V��=��zܼ��5�/W��3�~�0��X����̾���Z��ҕ��ÿr��M����#�621�      ��	�%X�L����,ݿH����ҕ��d��'�>��$���x�W����j���1�o��G��*���Q���ػ��0� �~���:��;5,;f=;;BE;��H;��I;��I;F�I;�I;btI;�VI;�@I;�1I;�'I;�!I;�I;�!I;�'I;�1I;�@I;�VI;`tI;�I;H�I;��I;��I;��H;>BE;g=;5,;��;��:��~���0���ػ�Q��*���G�0�o�j������x�W�$���>�꾌'��d��ҕ�H����,ݿL���%X�       �ȿ�ÿ���+8��hڇ�Z��'�����l8��W�s�,�&�V�/h??��V�琼SG#�^7��jTܺ��9#W�:��;L2;T@;�F;�I;��I;w�I;R�I;D�I;�lI;�PI;]<I;�-I;�$I;%I;FI;#I;�$I;�-I;[<I;�PI;�lI;H�I;S�I;y�I;��I;�I;�F;S@;$L2;��;W�:��9fTܺ^7��RG#�琼�V�h??�/V�,�&�W�s�l8�������'�Z�hڇ�+8������ÿ      '8��iڇ��x|�qm_�Gv<����>��l8��"6~�o74��l��z���6nc�3���^����\��9�@Z���=���n:T��:�#;�8;��B;w�G;�xI;r�I;��I;��I;݆I;7dI;zJI;�7I;*I;5!I;PI;�I;MI;6!I;*I;�7I;zJI;8dI;��I;��I;��I;r�I;�xI;{�G;��B;�8;�#;P��:�n:��=�BZ��9���\��^��3��6nc�z����l��o74�"6~�l8��>�꾎��Gv<�qm_��x|�iڇ�      ��7�r�3��'��K�'�����̾$���V�s�o74����!N��͇|�߁)�7zܼ�Y��< ����0���pT9���:(�;-;	=;�E;�H;L�I;3�I;��I;��I;{I;^[I;�CI;X2I;&I;�I;-I;�I;+I;�I;&I;X2I;�CI;a[I;!{I;��I;��I;1�I;K�I;�H;�E;=;-;'�;:�T90������< ��Y��6zܼ߁)�͇|�!N�����o74�V�s�$�����̾'����K��'�r�3�      C���s�XD־�t��p���X��x�W�,�&��l��!N���Ă�j�5�����{Q����A�>�ػ��G��!/�8f:b�:��;f�5;�9A;J�F;�*I;��I;��I;�I;[�I;/oI;gRI;�<I;-I;�!I;AI;I;�I;I;CI;�!I;-I;�<I;kRI;4oI;a�I;�I;��I;��I;�*I;J�F;�9A;j�5;��;b�:Hf:�!/���G�>�ػ��A�zQ������i�5��Ă�!N���l��,�&�x�W��X��p���t��XD־�s�      �S���7���X��W�s��_S�~�0����V�z���͇|�i�5�f���ک�2�X�c �t��3���9��:�;�,;�L<;XoD;.H;śI;��I;��I;T�I;N�I;7cI;[II;�5I;�'I;GI;�I;�I;�I;�I;�I;JI;�'I;�5I;^II;;cI;Z�I;Z�I;��I;��I;˛I;.H;]oD;�L<;�,;��; ��:�9�3��r�c �1�X��ک�e��i�5�͇|�z���Vར��~�0��_S�W�s��X���7��      �7�{74�o�)�#>����3�j���/6nc�߁)������ک�ua��Q�N���N���ȸ0��:��;�#;w�6;hA;��F;�I;6�I;`�I;�I;x�I;�uI;mWI;r@I;
/I;c"I;I;�I;gI;[I;gI;�I;I;d"I;/I;w@I;tWI;�uI;}�I;�I;]�I;?�I;�I;��F;hA;y�6;�#;��;*��:��ȸN�N����Q�ta��ک�����߁)�6nc�.j���3����#>�o�)�{74�      3�_�Խ�������/W��0�o�g??�3��6zܼzQ��1�X��Q��6�������Ϲ��n:�m�:>;��0;�>;2E;QSH;N�I;��I;a�I;@�I;U�I;�fI;"LI;�7I;e(I;I;�I;^I;I;>I;I;]I;�I;I;a(I;�7I;*LI;�fI;\�I;B�I;]�I;��I;N�I;USH;9E;�>;��0;>;�m�:��n:��Ϲ����6���Q�0�X�zQ��6zܼ3��g??�0�o�/W���������Խ^�      |L��=ى��Ă�7�o�+T���5��G��V��^���Y����A�c �P���������\�J:il�:�e;&,;��:;5C;lG;�DI;�I;��I;��I;��I;�vI;�XI;BAI;�/I;"I;�I;�I;�I;�I;HI;�I;�I;�I;�I;"I;�/I;IAI;�XI;�vI;��I;��I;��I;�I;�DI;lG;5C;��:;*,;�e;ul�:X�J:������N���c ���A��Y���^���V��G���5�	+T�7�o��Ă�=ى�      �)���&�H<��3��� �zܼ�*��琼��\�< �>�ػt�N���ϹX�J:�j�:n�;|�(;�e8;��A;�F;��H;!�I;m�I; �I;��I;_�I;\eI;�KI;7I;�'I;�I;I;�I;aI;�I;&I;�I;^I;�I;I;�I;�'I;7I;�KI;ceI;`�I;��I;�I;n�I;"�I;��H;�F;��A;�e8;x�(;s�;�j�:\�J:��ϹN�r�>�ػ< ���\�琼�*��~zܼ�� ��3�H<���&�      ��ƼNü8_���۩�($��=���Q�PG#��9�����G��3��`�ȸ��n:sl�:u�; �';�7;xv@;$�E;vH;��I;��I;��I;;�I;��I;�qI;sUI;*?I;�-I;y I;I;kI;�I;CI;�I;I;�I;@I;�I;kI;I;~ I;�-I;/?I;wUI;�qI;��I;B�I;��I;��I;��I;vH;+�E;zv@;�7;#�';u�;ul�:��n:@�ȸ�3����G�����9�PG#��Q�<��)$���۩�:_��Nü      ��\�"�X�z-M���:��G#�U����ػZ7��?Z�"����!/��9"��:�m�:�e;y�(;�7;�@;(]E;�-H;5wI;x�I;��I;��I;��I;�|I;�^I;�FI;�3I;J%I;�I;�I;D
I;?I;"I;- I;r�H;* I; I;=I;D
I;�I;�I;N%I;�3I;�FI;�^I;�|I;��I;��I;��I;{�I;8wI;�-H;+]E;�@;�7;x�(;�e;�m�:$��:�9�!/�"���8Z�Z7����ػT���G#���:�x-M�"�X�      �ݻ��ػ��ʻgT��͒��H�s��0�VTܺ��=��T9`f: ��:��;>;*,;�e8;xv@;/]E;4H;bI;�I;��I;A�I;��I;T�I;�fI;�MI;�9I;�)I;iI;mI;�I;2I;I;G�H;~�H;��H;{�H;D�H;I;2I;�I;qI;lI;�)I;�9I;�MI;�fI;\�I;��I;;�I;��I;�I;bI;6H;)]E;|v@;�e8;*,;>;��;&��:df:�T9��=�VTܺ�0�N�s�ʒ��lT����ʻ��ػ      �+���%�J������n1��pU\�p�~���9�n:쉹:b�:��;�#;��0;��:;��A;(�E;�-H;bI;��I;h�I;}�I;�I;��I;�mI;�SI;?I;3.I;� I;XI;�I;^I;uI;��H;p�H;�H;t�H;
�H;n�H;��H;xI;\I;�I;VI;� I;9.I;?I;�SI;�mI;��I;�I;~�I;l�I;��I;bI;�-H;(�E;��A;��:;��0;�#;��;b�:쉹:�n:��9��~�\U\�`1�����X����%�       Pɸ �J��$�8(�9��:x�n:��:#W�:P��:(�;��;�,;w�6;�>;5C;�F;vH;?wI;�I;h�I;7�I;øI;Y�I;�rI;�XI;4CI;�1I;)$I;�I;�I;�I;EI;=�H;0�H;��H;��H;s�H;��H;��H;-�H;=�H;@I;�I;�I;�I;,$I;�1I;3CI;�XI;�rI;T�I;ǸI;;�I;h�I;�I;;wI;vH;�F;5C;�>;w�6;�,;��;(�;H��:W�:��:h�n: �:((�9�%�8��J�      ��:ꃹ:��:�f�:���:���:��;��;#;
-;m�5;�L<;	hA;:E;lG;��H;��I;}�I;��I;��I;ǸI;�I;�tI;y[I;HFI;�4I;�&I;3I;�I;Q
I;iI;��H;�H;t�H;��H;��H;f�H;��H;��H;t�H;�H;��H;nI;Q
I;�I;6I;�&I;�4I;NFI;x[I;�tI;�I;ɸI;��I;��I;{�I;��I;��H;lG;5E;hA;�L<;n�5;-;#;��;��;���:ݱ�:�f�:ړ�:ԃ�:      4x;�b;�;�<;,�;�%;A,;0L2;�8;=;�9A;foD;��F;bSH;�DI;)�I;��I;��I;A�I;�I;X�I;�tI;a\I;�GI;6I;�(I;�I;@I;�I;NI;C I;s�H;L�H;�H;��H;��H;��H;��H;��H;�H;L�H;r�H;H I;MI;�I;DI;�I;�(I;�6I;�GI;[\I;�tI;Y�I;
�I;B�I;��I;��I;(�I;�DI;\SH;��F;coD;�9A;=;�8;,L2;?,;�%;=�;�<;�;�b;      ��0;��0;K2;�_4;&7;��9;_=;S@;��B;�E;E�F;.H;�I;Q�I;�I;n�I;��I;��I;��I;��I;�rI;q[I;�GI;#7I;p)I;�I;SI;�I;2I;� I;��H;��H;��H;��H;��H;	�H;��H;�H;��H;��H;��H;��H;��H;� I;/I;�I;PI;�I;v)I;!7I;�GI;t[I;�rI;��I;��I;��I;��I;m�I;�I;J�I;�I;.H;J�F;�E;��B;X@;_=;��9;07;�_4;K2;��0;      ˤ?;x�?;v@;hA;e�B;��C;@BE;�F;y�G;�H;�*I;ЛI;9�I;��I;��I;�I;F�I;ƢI;`�I;�mI;�XI;KFI;�6I;{)I;\I;�I;6I;�I;wI;4�H;��H;��H;��H;*�H;�H;o�H;2�H;i�H;�H;,�H;��H;��H;��H;5�H;qI;�I;2I;�I;_I;x)I;�6I;OFI;�XI;�mI;b�I;��I;H�I;�I;��I;��I;;�I;ЛI;�*I;�H;x�G;�F;BBE;��C;s�B;hA;v@;x�?;      J�F;�F;K�F;8G;t�G;�.H;��H;I;�xI;X�I;��I;��I;e�I;k�I;��I;��I;��I;�|I;�fI;�SI;7CI;�4I;�(I;�I;�I;tI;0I;�I;p�H;��H;��H;��H;��H;��H;��H;��H;��H;��H;��H;��H;��H;��H;��H;��H;m�H;�I;,I;xI;�I;�I;�(I;�4I;7CI;�SI; gI;�|I;��I; �I;��I;e�I;d�I;��I;��I;V�I;�xI;I;��H;�.H;��G;8G;K�F;�F;      ,I;�2I;�FI;dI;��I;�I;��I;��I;s�I;4�I;��I;��I;�I;D�I;��I;b�I;�qI;�^I;NI;
?I;�1I;�&I;�I;WI;4I;/I;�I;��H;�H;��H;��H;��H;8�H;�H;,�H;��H;��H;��H;*�H;�H;9�H;��H;��H;��H;�H;��H;�I;2I;9I;SI;�I;�&I;�1I;?I;NI;�^I;�qI;d�I;��I;@�I;�I;��I;��I;1�I;p�I;��I;��I;�I;·I;tdI;�FI;�2I;      ��I;��I;g�I;
�I;�I;�I;��I;w�I;��I;��I;�I;\�I;x�I;_�I;�vI;_eI;sUI;�FI;�9I;5.I;-$I;/I;@I;�I;�I;�I;��H;2�H;!�H;��H;�H; �H;��H;��H;"�H;��H;��H;��H;"�H;��H;��H;��H;��H;��H;�H;2�H;��H;�I;�I;�I;AI;0I;-$I;2.I;�9I;�FI;tUI;beI;�vI;_�I;z�I;^�I;�I;��I;��I;u�I;��I;�I;�I;�I;g�I;��I;      ��I;.�I;��I;;�I;Z�I;�I;K�I;Y�I;��I;��I;a�I;[�I;�uI;�fI;�XI;�KI;3?I;�3I;�)I;� I;�I;�I;�I;/I;pI;i�H;�H;�H;��H;~�H;��H;��H;O�H;��H;;�H;��H;��H;��H;9�H;��H;Q�H;��H;��H;{�H;��H;�H;�H;h�H;sI;+I;�I;�I;�I;� I;�)I;�3I;2?I;�KI;�XI;�fI;�uI;[�I;e�I;��I;��I;Y�I;M�I;��I;e�I;?�I;��I;+�I;      ؽI;�I;6�I;Z�I;ȮI;��I;�I;N�I;�I;#{I;7oI;GcI;tWI;-LI;IAI;7I;�-I;I%I;hI;XI;�I;M
I;LI;� I;6�H;��H;��H;��H;��H;��H;��H;G�H;^�H;��H;#�H;��H;��H;��H; �H;��H;\�H;F�H;��H;��H;�H;��H;��H;��H;9�H;� I;MI;N
I;�I;UI;hI;G%I;�-I;7I;IAI;*LI;rWI;BcI;7oI;%{I;��I;H�I;��I;��I;ȮI;d�I;5�I;�I;       �I;`�I;�I;i�I;��I;y{I;btI;�lI;>dI;j[I;qRI;jII;|@I;�7I;�/I;�'I;� I;�I;tI;I;�I;kI;B I;��H;��H;��H;��H;��H;��H;��H;9�H;6�H;��H;��H;m�H;E�H;2�H;D�H;k�H;��H;��H;6�H;:�H;��H;��H;��H;��H;��H;��H;��H;H I;lI;�I;�I;tI;�I;� I;�'I;�/I;�7I;|@I;hII;qRI;k[I;>dI;�lI;ltI;t{I;��I;k�I;�I;`�I;      �hI;]hI;�fI;dI;~`I;\I;�VI;�PI;�JI;�CI;�<I;�5I;/I;l(I;"I;�I;I;�I; I;dI;OI;��H;p�H;��H;��H;��H;��H;�H;��H;J�H;4�H;��H;��H;2�H;��H;��H;��H;��H;��H;4�H;��H;��H;2�H;G�H;��H;�H;��H;��H;��H;��H;u�H;��H;HI;`I; I;�I;I;�I;"I;k(I;/I;�5I;�<I;�CI;JI;�PI;�VI;\I;�`I;'dI;�fI;^hI;      �NI;�NI;?MI;KI;IHI;�DI;�@I;[<I;�7I;V2I;-I;�'I;g"I;I;�I;I;rI;G
I;:I;|I;H�H;�H;I�H;��H;��H;��H;8�H;��H;X�H;a�H;��H;��H;�H;��H;x�H;5�H;/�H;5�H;w�H;��H;�H;��H;��H;Z�H;T�H;��H;6�H;��H;��H;��H;M�H;�H;B�H;xI;:I;G
I;uI;I;�I;I;f"I;�'I;#-I;X2I;�7I;X<I;�@I;�DI;MHI;KI;MMI;�NI;      �<I;1<I;>;I;�9I;�7I;�4I;�1I;.I;*I; &I;�!I;UI;I;�I;�I;�I;�I;?I;I; �H;7�H;t�H;��H;��H;%�H;��H;�H;��H;��H;��H;��H;3�H;��H;Q�H;�H;��H;��H;��H;�H;R�H;��H;4�H;��H;��H;��H;��H;�H;��H;)�H;��H;�H;t�H;1�H;��H;I;BI;�I;�I;�I;�I;I;SI;�!I;"&I;*I;.I;�1I;�4I;�7I;�9I;I;I;?<I;      �0I;�0I;�/I;Q.I;o,I;'*I;�'I;�$I;=!I;�I;OI;�I;
I;jI;�I;gI;JI;"I;K�H;s�H;��H;��H;��H;��H;�H;~�H;&�H;"�H;@�H;&�H;g�H;��H;x�H;�H;��H;��H;��H;��H;��H;�H;z�H;��H;e�H;�H;9�H;�H;&�H;}�H;�H;��H;��H;��H;��H;o�H;I�H;%I;LI;iI;�I;kI;
I;�I;TI;�I;?!I;�$I;�'I;)*I;i,I;Y.I;�/I;�0I;      �)I;m)I;�(I;�'I;&I;$I;�!I;-I;PI;8I;I;�I;mI;&I;	I;�I;�I;* I;��H;�H;��H;��H;��H;��H;f�H;��H;��H;��H;��H;��H;D�H;��H;9�H;��H;��H;h�H;h�H;l�H;��H;��H;:�H;��H;B�H;��H;��H;��H;��H;��H;h�H;��H;��H;��H;��H;
�H;��H;. I;�I;�I;	I;)I;mI;�I;I;9I;SI;*I;�!I;$I;&I;�'I;�(I;z)I;      �'I;�'I;�&I;�%I;�#I;"I;�I;QI;�I;�I;�I;�I;cI;KI;TI;-I;(I;v�H;��H;|�H;~�H;g�H;��H;��H;.�H;��H;��H;��H;��H;��H;,�H;��H;/�H;��H;��H;e�H;J�H;f�H;��H;��H;2�H;��H;,�H;��H;��H;��H;��H;��H;/�H;��H;��H;g�H;w�H;x�H;��H;x�H;(I;1I;VI;LI;cI;�I;�I;�I;�I;PI;�I;"I;�#I;�%I;�&I;�'I;      �)I;o)I;�(I;�'I;&I;$I;�!I;-I;QI;9I;I;�I;nI;)I;	I;�I;�I;* I;��H;�H;��H;��H;��H;��H;h�H;��H;��H;��H;��H;��H;D�H;��H;:�H;��H;��H;h�H;h�H;l�H;��H;��H;:�H;��H;B�H;��H;��H;��H;��H;��H;h�H;��H;��H;��H;��H;�H;��H;. I;�I;�I;	I;'I;mI;�I;I;6I;SI;-I;�!I;$I;&I;�'I;�(I;v)I;      �0I;�0I;�/I;M.I;o,I;'*I;�'I;�$I;?!I;�I;QI;�I;
I;jI;�I;gI;JI;$I;K�H;u�H;��H;��H;��H;��H;�H;}�H;&�H;"�H;?�H;%�H;e�H;��H;z�H;�H;��H;��H;��H;��H;��H;�H;z�H;��H;e�H;�H;;�H;�H;&�H;~�H;�H;��H;��H;��H;��H;o�H;I�H;%I;MI;iI;�I;kI;
I;�I;TI;�I;?!I;�$I;�'I;'*I;n,I;V.I;�/I;�0I;      �<I;4<I;>;I;�9I;�7I;�4I;�1I;	.I;*I; &I;�!I;TI;I;�I;�I;�I;�I;CI;I; �H;8�H;v�H; �H;��H;)�H;��H;�H;��H;��H;��H;��H;3�H;��H;Q�H;�H;��H;��H;��H;�H;Q�H;��H;4�H;��H;��H;��H;��H;�H;��H;(�H;��H;�H;v�H;.�H;��H;I;BI;�I;�I;�I;�I;I;SI;�!I;!&I;*I;.I;�1I;�4I;�7I;�9I;G;I;7<I;      �NI;�NI;CMI;KI;HHI;�DI;�@I;b<I;�7I;X2I; -I;�'I;f"I;I;�I;I;tI;G
I;9I;|I;I�H;�H;I�H;��H;��H;��H;6�H;��H;Y�H;a�H;��H;��H;�H;��H;z�H;5�H;/�H;5�H;x�H;��H;�H;��H;��H;Z�H;Q�H;��H;6�H;��H;��H;��H;N�H;�H;@�H;{I;9I;F
I;rI;I;�I;I;i"I;�'I;!-I;V2I;�7I;^<I;�@I;�DI;LHI;(KI;TMI;�NI;      �hI;`hI;�fI; dI;�`I;\I;�VI;�PI;JI;�CI;�<I;�5I;/I;k(I;"I;�I;I;�I;�I;cI;PI;��H;r�H;��H;��H;��H;��H;�H;��H;H�H;2�H;��H;��H;0�H;��H;��H;��H;��H;��H;2�H;��H;��H;1�H;F�H;��H; �H;��H;��H;��H;��H;v�H;��H;GI;`I;�I;�I;I;�I;"I;l(I;/I;�5I;�<I;�CI;�JI;�PI;�VI;\I;�`I;,dI;�fI;[hI;      �I;b�I;�I;c�I;��I;{{I;etI;�lI;>dI;j[I;pRI;lII;|@I;�7I;�/I;�'I;� I;�I;tI;�I;�I;lI;C I;��H;��H;��H;��H;��H;��H;��H;9�H;8�H;��H;��H;o�H;D�H;2�H;G�H;j�H;��H;��H;8�H;7�H;��H;��H;��H;��H;��H;��H;��H;H I;lI;�I;�I;uI;�I;� I;�'I;�/I;�7I;|@I;hII;qRI;h[I;AdI;�lI;ltI;x{I;��I;n�I;	�I;d�I;      ޽I;��I;1�I;d�I;��I;��I;�I;Q�I;�I;&{I;4oI;EcI;tWI;-LI;MAI;7I;�-I;J%I;iI;XI;�I;O
I;JI;� I;9�H;��H;��H;��H;��H;��H;��H;H�H;[�H;��H;#�H;��H;��H;��H; �H;��H;^�H;H�H;��H;��H;~�H;��H;��H;��H;6�H;� I;PI;N
I;�I;UI;jI;G%I;�-I;7I;LAI;,LI;rWI;BcI;4oI;({I;��I;N�I;��I;��I;ƮI;l�I;9�I;�I;      ��I;0�I;�I;2�I;L�I;�I;I�I;Y�I;��I;��I;c�I;\�I;�uI;�fI;�XI;�KI;3?I;�3I;�)I;� I;�I;�I;�I;/I;sI;e�H;�H;�H;��H;{�H;��H;��H;O�H;��H;;�H;��H;��H;��H;9�H;��H;Q�H;��H;��H;{�H;��H;�H;�H;i�H;pI;(I;�I;�I;�I;� I;�)I;�3I;3?I;�KI;�XI;�fI;�uI;Z�I;e�I;��I;��I;Y�I;P�I;�I;\�I;5�I;�I;+�I;      ��I;��I;]�I;�I;�I; �I;��I;z�I;��I;��I;�I;_�I;z�I;_�I;�vI;beI;tUI;�FI;�9I;3.I;0$I;3I;@I;�I;�I;�I;��H;2�H;"�H;��H;�H;�H;��H;��H;"�H;��H;��H;��H;!�H;��H;��H;��H;��H;��H;�H;/�H;��H;�I;�I;�I;DI;0I;,$I;2.I;�9I;�FI;wUI;ceI;�vI;^�I;z�I;\�I;�I;��I;��I;u�I;��I;�I;�I;�I;g�I;��I;      �+I;�2I;�FI;�dI;ćI;"�I;��I;��I;s�I;4�I;��I;��I;�I;C�I;��I;c�I;�qI;�^I;NI;?I;�1I;�&I;�I;ZI;9I;,I;�I;��H;�H;��H;��H;��H;6�H;�H;-�H;��H;��H;��H;*�H;�H;8�H;��H;��H;��H;�H;��H;�I;2I;6I;TI;�I;�&I;�1I;
?I;NI;�^I;�qI;f�I;��I;C�I;�I;��I;��I;3�I;p�I;��I;��I;�I;̇I;�dI;�FI;�2I;      C�F;�F;X�F;8G;z�G;�.H;��H;I;�xI;U�I;��I;��I;e�I;h�I;��I; �I;��I;�|I; gI;�SI;;CI;�4I;�(I;�I;�I;sI;/I;�I;s�H;��H;��H;��H;��H;��H;��H;��H;��H;��H;��H;��H;��H;��H;��H;��H;l�H;�I;/I;xI;�I;�I;�(I;�4I;7CI;�SI;gI;�|I;��I;�I;��I;h�I;d�I;��I;��I;V�I;�xI; I;��H;�.H;��G;8G;=�F;�F;      ɤ?;v�?;v@;hA;g�B;��C;BBE;�F;|�G;�H;�*I;ӛI;;�I;��I;��I;�I;H�I;ǢI;b�I;�mI;�XI;NFI;�6I;})I;`I;�I;4I;�I;wI;2�H;��H;��H;��H;*�H;�H;l�H;2�H;l�H;�H;*�H;��H;��H;��H;4�H;pI;�I;5I;�I;]I;x)I;�6I;NFI;�XI;�mI;d�I;��I;I�I;�I;��I;��I;<�I;ϛI;�*I;	�H;w�G;�F;CBE;��C;r�B;hA;v@;v�?;      l�0;u�0;K2;�_4;"7;��9;_=;V@;��B;�E;H�F;.H;�I;M�I;�I;p�I;��I;��I;��I;��I;�rI;r[I;�GI;#7I;w)I;�I;QI;�I;2I;� I;��H;��H;��H;��H;��H;�H;��H;	�H;��H;��H;��H;��H;��H;� I;0I;�I;SI;�I;t)I;#7I;�GI;r[I;�rI;��I;��I;��I;��I;q�I;�I;M�I;�I;.H;J�F;�E;��B;P@;b=;��9;47;�_4;K2;`�0;      0x;�b;�;�<;,�;�%;;,;,L2;�8;=;�9A;doD;��F;_SH;�DI;+�I;��I;��I;B�I;�I;[�I;�tI;]\I;�GI;�6I;�(I;�I;BI;�I;JI;E I;v�H;L�H;�H;��H;��H;��H;��H;��H; �H;M�H;u�H;I I;PI;�I;@I;�I;�(I;�6I;�GI;^\I;�tI;Y�I;�I;E�I;��I;��I;+�I;�DI;\SH;��F;coD;�9A;=;�8;)L2;;,;�%;)�;�<;�;�b;      ��:胹:ܓ�:�f�:���:���:��;��;#;-;m�5;�L<;	hA;6E;lG;��H;��I;}�I;��I;��I;̸I;�I;�tI;x[I;OFI;�4I;�&I;4I;�I;O
I;kI;��H;�H;t�H;��H;��H;g�H;��H;��H;s�H;�H;��H;oI;R
I;�I;3I;�&I;�4I;KFI;{[I;�tI;�I;ǸI;��I;��I;z�I;��I;��H;lG;8E;hA;�L<;n�5;-;#;��;��;���:ױ�:�f�:֓�:҃�:      �Qɸ �J��&�8((�9�:��n:��:W�:T��:$�;��;�,;y�6;�>;5C;�F;vH;<wI;�I;k�I;:�I;ǸI;V�I;�rI;�XI;2CI;�1I;*$I;�I;�I;�I;GI;=�H;1�H;��H;��H;u�H;��H;��H;,�H;>�H;EI;�I;�I;�I;)$I;�1I;3CI;�XI;�rI;U�I;ŸI;:�I;l�I;�I;9wI;vH;�F;5C;�>;y�6;�,;��;(�;L��:#W�:��:��n:0�:@(�9 (�8@�J�      q+���%�N������p1��`U\���~���9 �n:쉹:b�:��;�#;��0;��:;��A;*�E;�-H;bI;��I;n�I;��I;�I;��I;�mI;�SI;?I;5.I;� I;TI;�I;^I;xI;��H;r�H;�H;u�H;�H;n�H;��H;wI;]I;�I;UI;� I;3.I;?I;�SI;�mI;��I;�I;~�I;k�I;��I;bI;�-H;+�E;��A;��:;��0;�#;��; b�:批:�n:��9p�~�|U\�b1������Q����%�      �ݻ��ػ��ʻgT��͒��G�s��0�VTܺ��=��T9`f:$��:��;>;.,;�e8;zv@;-]E;6H;bI;�I;��I;A�I;��I;\�I;�fI;�MI;�9I;�)I;iI;nI;�I;2I;I;H�H;}�H;��H;~�H;E�H;I;3I;�I;qI;jI;�)I;�9I;�MI;�fI;V�I;��I;?�I;��I;�I;bI;4H;+]E;|v@;�e8;,,;>;��;$��:`f:�T9��=�TTܺ�0�J�s�Β��fT����ʻ��ػ      ��\� �X�|-M���:��G#�R����ػV7��8Z�"����!/��9(��:�m�:�e;|�(;�7;�@;+]E;�-H;8wI;}�I;��I;��I;��I;�|I;�^I;�FI;�3I;I%I;�I;�I;D
I;@I;!I;, I;r�H;- I;I;=I;F
I;�I;�I;L%I;�3I;�FI;�^I;�|I;��I;��I;��I;x�I;5wI;�-H;+]E;�@;�7;y�(;�e;�m�:(��:�9�!/�$���;Z�X7����ػT���G#���:�~-M� �X�      ��ƼNü8_���۩�($��<���Q�PG#��9�����G��3��@�ȸ��n:{l�:z�;#�';�7;yv@;*�E;vH;��I;��I;��I;D�I;��I;�qI;qUI;2?I;�-I;| I;I;mI;�I;CI;�I; I;�I;?I;�I;jI;I;} I;�-I;/?I;qUI;�qI;��I;>�I;��I;��I;��I;vH;*�E;yv@;�7;!�';u�;wl�:��n:`�ȸ�3����G�����9�PG#��Q�<��)$���۩�:_��Nü      �)���&�H<��3��� �~zܼ�*��琼��\�= �>�ػr�N���Ϲd�J:�j�:p�;{�(;�e8;��A;�F;��H;(�I;n�I;�I;��I;]�I;^eI;�KI;7I;�'I;�I;I;�I;bI;�I;&I;�I;^I;�I;I;�I;�'I;7I;�KI;^eI;]�I;��I;�I;n�I;%�I;��H;�F;��A;�e8;x�(;q�;�j�:X�J:��ϹN�t�>�ػ= ���\�琼�*��~zܼ�� ��3�I<���&�      }L��=ى��Ă�7�o�+T���5��G��V��^���Y����A�c �N���������h�J:ul�:�e;),;��:;5C;lG;�DI;�I;��I;��I;��I;�vI;�XI;DAI;�/I;"I;�I;�I;�I;�I;HI;�I;�I;�I;�I;"I;�/I;BAI;�XI;�vI;��I;��I;��I;�I;�DI;lG;	5C;��:;&,;�e;ul�:X�J:������P���c ���A��Y���^���V��G���5�	+T�8�o��Ă�=ى�      3�^�Խ�������/W��0�o�g??�3��6zܼzQ��0�X��Q��6�����X�Ϲ��n:�m�:>;��0;�>;8E;WSH;P�I;��I;b�I;?�I;X�I;�fI;%LI;�7I;d(I;I;�I;^I;I;>I; I;\I;�I;I;a(I;�7I;%LI;�fI;X�I;=�I;^�I;��I;Q�I;[SH;6E;�>;��0;>;�m�:��n:��Ϲ����6���Q�1�X�zQ��6zܼ3��g??�0�o�/W���������Խ^�      �7�{74�o�)�#>����3�j���.6nc�߁)������ک�ta��Q�L���N�@�ȸ.��:��;�#;~�6;hA;��F;�I;?�I;`�I;�I;x�I;�uI;oWI;u@I;
/I;c"I;I;�I;gI;[I;gI;�I;I;d"I;/I;s@I;nWI;�uI;x�I;�I;]�I;8�I;�I;��F;	hA;r�6;�#;��;*��:@�ȸN�N����Q�va��ک�����߁)�6nc�/j���3����#>�o�)�{74�      �S���7���X��W�s��_S�~�0����V�z���͇|�i�5�e���ک�1�X�c �s��3����9��:��;�,;�L<;_oD;.H;̛I;��I;��I;T�I;U�I;7cI;_II;�5I;�'I;LI;�I;�I;�I;�I;�I;II;�'I;�5I;\II;7cI;W�I;T�I;��I;��I;śI;.H;boD;�L<; �,;��;��:��9�3��t�c �2�X��ک�e��i�5�͇|�z���Vར��~�0��_S�W�s��X���7��      C���s�XD־�t��p���X��x�W�,�&��l��!N���Ă�i�5�����zQ����A�>�ػ��G��!/�Df:b�:��;j�5;�9A;K�F;�*I;��I;��I;�I;a�I;0oI;jRI;�<I;-I;�!I;AI;I;�I;I;AI;�!I;-I;�<I;gRI;/oI;a�I;�I;��I;��I;�*I;L�F;�9A;g�5;��;b�:8f:�!/���G�>�ػ��A�zQ������i�5��Ă�!N���l��,�&�x�W��X��p���t��XD־�s�      ��7�r�3��'��K�'�����̾$���V�s�o74����!N��͇|�߁)�6zܼ�Y��< ����0����T9쉹:.�;-;=;�E;�H;N�I;1�I;��I;��I;{I;c[I;�CI;X2I;&I;�I;+I;�I;+I;�I;&I;X2I;�CI;a[I;{I;��I;��I;0�I;L�I;�H;�E;=;-;!�;쉹:pT92������< ��Y��6zܼ߁)�͇|�!N�����o74�W�s�$�����̾'����K��'�r�3�      '8��iڇ��x|�qm_�Gv<����>��l8��"6~�o74��l��z���6nc�3���^����\��9�CZ���=��n:^��:�#;�8;��B;|�G;�xI;r�I;��I;��I;݆I;;dI;wJI;�7I;*I;4!I;OI;�I;MI;5!I;*I;�7I;wJI;5dI;چI;��I;��I;p�I;�xI;y�G;��B;�8;�#;H��:�n:��=�BZ��9���\��^��3��6nc�z����l��o74�"6~�l8��>�꾎��Gv<�qm_��x|�iڇ�       �ȿ�ÿ���+8��hڇ�Z��'�����l8��W�s�,�&�V�/h??��V�琼RG#�`7��dTܺ��9)W�:��;$L2;W@;�F;�I;��I;u�I;S�I;D�I;�lI;�PI;[<I;�-I;�$I;"I;FI;"I;�$I;�-I;[<I;�PI;�lI;F�I;S�I;v�I;��I;�I;�F;V@;%L2;��;W�:��9jTܺ^7��RG#�琼�V�h??�/V�,�&�W�s�l8�������'�Z�hڇ�+8������ÿ      ��	�%X�L����,ݿH����ҕ��d��'�>��$���x�W����j���1�o��G��*���Q���ػ��0���~���:��;5,;i=;>BE;��H;��I;��I;I�I;�I;dtI;�VI;�@I;�1I;�'I;�!I;�I;�!I;�'I;�1I;�@I;�VI;atI;�I;H�I;��I;��I;��H;<BE;i=;:,;��;��:��~���0���ػ�Q��*���G�0�o�j������x�W�$���>�꾌'��d��ҕ�H����,ݿL���%X�      �5�621���#�M��r���ÿ�ҕ�Z������̾�X��~�0�3�/W����5�zܼ=��W��V�s�xU\���n:���:߬%;��9;��C;�.H;�I;�I;�I;��I;{{I;\I;�DI;�4I;(*I;$I;"I;$I;)*I;�4I;�DI;\I;v{I;��I;�I;�I;�I;�.H;��C;��9;�%;���:t�n:pU\�Y�s�W��=��zܼ��5�/W��3�~�0��X����̾���Z��ҕ��ÿr��M����#�621�      /�j���c�w�P��5���r��H���hڇ�Gv<�'���p���_S��������+T��� �($���G#�ʒ��Z1��,�:���:8�;37;v�B;z�G;ćI;�I;g�I;ʮI;��I;�`I;IHI;�7I;^,I;&I; $I;&I;b,I;�7I;LHI;�`I;��I;ͮI;g�I;�I;ƇI;��G;u�B;67;8�;���:�:X1��̒���G#�)$���� �+T���������_S�p��'���Gv<�hڇ�I���r�����5�w�P���c�      Т��^���E���/]��5�M���,ݿ+8��qm_��K��t��W�s�#>����8�o��3��۩���:�hT������h(�9�f�:�<;�_4;hA;8G;ydI;�I;-�I;Z�I;b�I;&dI;KI;�9I;H.I;�'I;�%I;�'I;K.I;�9I;KI;)dI;_�I;^�I;+�I;�I;{dI;8G;hA;�_4;�<;�f�: (�9����jT����:��۩��3�8�o����#>�W�s��t���K�qm_�+8���,ݿM���5��/]�E��^���      �����B����E��w�P���#�L�������x|��'�XD־�X��o�)�Խ�Ă�I<�8_��z-M���ʻQ���'�8Г�:�;!K2;v@;O�F;�FI;k�I;�I;*�I;�I;�fI;=MI;A;I;�/I;�(I;�&I;�(I;�/I;B;I;?MI;�fI;��I;-�I;�I;o�I;�FI;\�F;v@; K2;�;̓�:�&�8N����ʻz-M�7_��H<��Ă�Խo�)��X��XD־�'��x|����L�����#�w�P�E�����B��      ��������B��]�����c�621�%X��ÿiڇ�r�3��s��7��|74�_�=ى���&�Nü$�X���ػ��%� �J�҃�:�b;~�0;x�?;�F;�2I;��I;:�I;�I;I�I;QhI;�NI;1<I;z0I;_)I;�'I;\)I;z0I;1<I;�NI;ThI;E�I;�I;<�I;��I;�2I;�F;v�?;}�0;�b;̃�:@�J���%���ػ$�X�Nü��&�=ى�_�|74��7���s�r�3�iڇ��ÿ%X�621���c�]����B�����      E(��q'���o��N�d��X1�~x�	Ŀ����3�w���x����4�j��Y+���'���ü7yY��kٻp&� �p�V��:?;��0;��?;F;k I; �I;��I;/�I;n�I;OdI;�KI;�9I;n.I;�'I;�%I;�'I;n.I;�9I;�KI;PdI;j�I;3�I;��I;�I;k I;΀F;��?;��0;9;N��:��p�p&��kٻ7yY���ü�'�Y+��j�ཽ�4��x��w���3����	Ŀ~x��X1�d�N��o��q'��      q'���X��e^�������]]���,�P9�7g��U�����/����o��f1��hܽ���-$�]l���|U�b�Իx!� �,���:�;�51;��?;7�F;D'I;d�I;�I;@�I;��I;�cI;AKI;{9I; .I;}'I;�%I;y'I;".I;z9I;BKI;�cI;��I;C�I;�I;g�I;C'I;E�F;��?;�51;�;{�: �,�x!�b�Ի�|U�]l���-$����hܽf1��o���ྙ�/�U���7g��P9���,��]]�����e^���X��      �o��e^���ē��4z�5K�h��R��%ﱿT�v��X#���Ѿń��&�o�нc̀�^��t���H�I��ǻ�4��"9��::�;$�2;��@;��F;�:I;��I;��I;��I;z�I;NbI;�II;�8I;\-I;�&I;�$I;�&I;\-I;�8I;JI;NbI;u�I;��I;��I;��I;�:I;��F;��@; �2;6�;��:�"9�4��ǻH�I�t���^��c̀�o�н�&�ń���Ѿ�X#�T�v�%ﱿR��h��5K��4z��ē�e^��      N������4z���V��X1��<�sؿ����RZ��	�(���IUo����]y��,l�X��R��A�7������Ƴ9��:��;^�4;ntA;`2G;�XI;��I;O�I;�I;��I;�_I;�GI;%7I;�+I;�%I;�#I;�%I;�+I;"7I;�GI;�_I;�I;�I;O�I;��I;�XI;j2G;mtA;[�4;��;��:�ų9������@�7��R��X�,l�]y�����IUo�(����	��RZ����sؿ�<��X1���V��4z�����      d��]]�5K��X1�Zf��nQ��T���[58��A���נ���O���_什�Q����>ߓ��� ��V��x氺�":��:	 ;�07;�B;3�G;�{I;��I;��I;��I;<|I;:\I;MEI;5I;6*I;3$I;,"I;0$I;7*I;5I;NEI;8\I;7|I;��I;��I;��I;�{I;;�G;�B;�07; ;޸�:�":n氺�V���� �>ߓ�����Q�_什����O��נ��A��[58�T���nQ���Zf��X1�5K��]]�      �X1���,�h���<��6g��e_���U�͂�֌Ⱦń�*�-�h��O ��$�2�	?ټ_�{� "��n��O���u:�P ;�&;.#:;A�C;�%H;!�I;%�I;��I;�I;`vI;�WI;�AI;|2I;(I;F"I;a I;A"I;(I;x2I;�AI;�WI;]vI;�I;��I;(�I;�I;�%H;A�C;+#:;�&;�P ;��u:��O��n� "�_�{�	?ټ$�2�O ��h��*�-�ń�֌Ⱦ͂��U�e_��6g��<�h����,�      ~x�P9�R��sؿnQ��e_��6�_��X#�q���f��9�S�{�����l�A�w���M���Ի��+��<T���:�e;�\,;�/=;�BE;V�H;�I;��I;��I;��I;�oI;�RI;>I;^/I;�%I;�I;GI;�I;�%I;^/I;>I;�RI;�oI;��I;��I;��I;{�I;]�H;�BE;�/=;�\,;�e;��:`<T���+���Ի�M�w��A�l�����{�9�S��f��q���X#�6�_�e_��nQ��sؿR��P9�      	Ŀ7g��%ﱿ���T����U��X#�t��d���HUo��#��hܽ����n<����;����� ��᝻0�Ժ�t�9n��:�V;҇2;� @;X�F;�I;�I;E�I;+�I;l�I; hI;MI;�9I;�+I;�"I;lI;�I;iI;�"I;�+I;�9I;MI; hI;o�I;,�I;H�I;��I;�I;\�F;� @;ԇ2;�V;f��:�t�92�Ժ�᝻�� �;�������n<�����hܽ�#�HUo�d���t���X#��U�T������%ﱿ7g��      ���U���T�v��RZ�[58�͂�q��d���foy�]1�_O��[什�`�L�����myY��컌�T���1���u:
��:M#;98;�B;l�G;�lI;�I;�I;/�I;w�I;�_I;GI;�4I;%(I;�I;�I;I;�I;�I;&(I;�4I;GI;�_I;z�I;2�I;�I;�I;�lI;p�G;�B;98;O#;��:��u:�1���T���myY����L���`�[什_O��]1�foy�d���q��͂�[58��RZ�T�v�U���      �3���/��X#��	��A��֌Ⱦ�f��HUo�]1�ʰ��{n��Ҽx��'��>ټ�@���k�ʼ����P�39�#�:4R;e-;�/=;�	E;`xH;��I;�I;q�I;�I;vI;cWI;�@I;�/I;%$I;<I;�I;7I;�I;>I;%$I;�/I;�@I;eWI;vI;�I;v�I;�I;��I;dxH;�	E;�/=;e-;4R;�#�:��39��ȼ���k��@���>ټ�'�Ҽx�{n��ʰ��]1�HUo��f��ՌȾ�A���	��X#���/�      w���ྃ�Ѿ(����נ�ń�9�S��#�_O��{n��Ì���2���𛼀�>���Ի��B��#�Tm:�G�:c ;��5;�FA;��F;�I;R�I;U�I;��I;j�I;mjI;�NI;:I;�*I;�I;�I;�I;II;�I;�I;�I;�*I;:I;�NI;tjI;q�I;��I;W�I;P�I;�I;��F;�FA;��5;e ;�G�:dm:�#���B���Ի��>�������2�Ì�{n��_O���#�9�S�ń��נ�(�����Ѿ��      �x���o��ń�IUo���O�*�-�{��hܽ[什Ӽx���2�rb��TR��T|U�W2��4��갺�u�9��:D;��,;�h<;erD;S%H;ƏI;j�I;��I;�I;�I;�^I;FI;W3I;�%I;�I;_I;iI;4I;hI;^I;�I;�%I;S3I;FI;�^I;�I;�I;��I;g�I;ʏI;T%H;lrD;�h<;��,;D;��:�u�9갺4��W2��S|U�SR��rb����2�Ӽx�[什�hܽ{�*�-���O�IUo�ń��o��      ��4�f1��&���� ��h�ང�������`��'���SR��B�]�|��V���X���Fo����:p�;,#;�6;XtA;T�F;�	I;x�I;��I;q�I;�I;�pI;�SI;�=I;�,I;w I;�I;�I;GI;;I;GI;�I;�I;y I;�,I;�=I;�SI;�pI;�I;r�I;��I;}�I;�	I;X�F;]tA; �6;8#;v�;���:@Eo��X��V��{��B�]�SR����'��`��������h��������&�f1�      j�ཷhܽo�н]y��^什P ��l��n<�L���>ټ��T|U�}�������1�H�����u:el�:�;h71;Y)>;X	E;JH;Z�I;��I;��I;�I;׃I;YbI;�HI;$5I;c&I;gI;qI;<I;#I;
I;#I;:I;rI;gI;b&I;-5I;�HI;cbI;ރI;�I;��I;��I;Z�I;JH;^	E;\)>;s71;�;el�:�u:X����1�����|��S|U��𛼿>ټL���n<�l�O ��_什]y��o�н�hܽ      X+����b̀�,l��Q�$�2�A��������@����>�X2��V���1�`��$R:���:�;}\,;:;;�;C;�eG;[9I;��I;0�I;��I;D�I;�qI;�TI;`>I;5-I;1 I;zI;qI;�
I;I;
I;I;�
I;rI;{I;1 I;<-I;g>I;�TI;�qI;F�I;��I;7�I;��I;\9I;�eG;�;C;E;;�\,;�;���:$R:`��~1�V��V2���>��@��������A�$�2��Q�-l�c̀���      �'�-$�^��X����	?ټw��:���myY��k���Ի6���X��X���$R:���:�R;�);�8;��A;��F;7�H;,�I;��I;��I;��I;�I;�`I;�GI;�4I;�%I;JI;�I;�I;oI;I;CI;I;mI;�I;�I;HI;�%I;�4I;�GI;�`I;�I;��I;��I;��I;-�I;>�H;��F;��A;�8;�);�R;���: $R:X����X��3����Ի�k�lyY�:���w��?ټ���X�^��-$�      ��ü\l��v����R��=ߓ�_�{��M��� ���Ƽ����B�
갺@Fo��u:���:�R;7�'; 17;Å@;��E;�lH;2�I;l�I;��I;�I;x�I;�lI;�QI;&<I;�+I;�I;�I;eI;�I;EI;0I;�I;,I;AI;�I;cI;�I;�I;�+I;)<I;�QI;�lI;t�I;�I;��I;k�I;8�I;�lH;�E;ǅ@;17;9�';�R;���:�u:@Fo�갺{�B�ż���컈� ��M�^�{�>ߓ��R��v���[l��      0yY��|U�H�I�=�7��� ��!���Ի�᝻��T� ��#��u�9���:al�:�;�);17;6 @;A]E;�$H;kkI;�I;Y�I;��I;*�I;�wI;�ZI;�CI;w1I;N#I;%I;�I;-	I;rI;8I;m�H;��H;h�H;5I;rI;+	I;�I;,I;U#I;z1I;�CI;�ZI;�wI;2�I;��I;U�I;�I;mkI;�$H;E]E;5 @;17;�);�;el�:���:�u�9�#�����T��᝻��Ի�!��� �>�7�F�I��|U�      �kٻf�Ի�ǻ	����V���n���+�"�Ժ̷1���39xm:��:r�;�;�\,;�8;Å@;F]E;�
H;QVI;v�I;��I;��I;f�I;��I;�bI;cJI;&7I;�'I;�I;,I;�
I;8I;;I;i�H;��H;z�H;��H;f�H;8I;8I;�
I;2I;�I;�'I;*7I;cJI;�bI;�I;l�I;��I;��I;{�I;TVI;�
H;B]E;ȅ@;�8;�\,;�;v�;��:�m:��39ط1��Ժ��+��n��V������ǻf�Ի      p&�{!��4���氺��O� <T��t�9��u:�#�:�G�:D;1#;p71;D;;��A;�E;�$H;QVI;�I;��I;�I;��I;��I;	iI;,PI;<I;�+I;I;�I;�I;�I;�I;3�H;��H;��H;�H;��H;��H;2�H;�I;�I;�I;�I;I;�+I;<I;)PI;iI;�I;��I;�I;��I;�I;VVI;�$H;�E;��A;D;;n71;0#;D;�G�:�#�:��u:�t�90<T�ܬO�n氺���4��!�      @�p� �,�p!9�ų9��":��u:��:t��:��:6R;e ;��,;�6;Z)>;�;C;��F;�lH;rkI;y�I;��I;��I;�I;u�I;�mI;zTI;)@I;�/I;$"I;YI;�I;�I;�I;t�H;t�H;��H;W�H;��H;P�H;��H;t�H;t�H;�I;�I;�I;WI;("I;�/I;'@I;�TI;�mI;p�I;�I;��I;��I;{�I;lkI;�lH;��F;�;C;W)>;�6;��,;f ;4R; ��:h��:��:��u:�":�ų9�!9 �,�      H��:��:�:#��:и�:�P ;�e;�V;Q#;e-;��5;�h<;ZtA;`	E;�eG;>�H;8�I;�I;��I;�I;�I;��I;pI;OWI;�BI;C2I;�$I;tI;oI;B	I;tI;��H;��H;�H;Z�H;5�H;��H;/�H;W�H;�H;��H;��H;yI;D	I;oI;wI;�$I;G2I;�BI;OWI;pI;��I;�I;�I;��I;�I;9�I;=�H;�eG;[	E;YtA;�h<;��5;e-;Q#;�V;�e;�P ;��:��: �:��:      Q;�;6�;��;� ;�&;�\,;��2; 98;�/=;�FA;urD;[�F;JH;`9I;4�I;r�I;_�I;��I;��I;u�I;pI;LXI;�DI;�3I;_&I;!I;�I;�
I;oI;��H;��H;��H;��H;;�H;J�H;�H;E�H;8�H;��H;��H;��H;��H;oI;~
I;�I;I;b&I;�3I;�DI;HXI;pI;w�I;��I;��I;W�I;r�I;1�I;^9I;JH;X�F;rrD;�FA;�/=;98;݇2;�\,;�&; ;��;2�;�;      ��0;�51;�2;X�4;�07;3#:;�/=;� @;�B;�	E;��F;T%H;�	I;\�I;��I;��I;��I;��I;g�I;��I;�mI;GWI;�DI;�4I;>'I;0I; I;I;;I;. I;,�H;��H;{�H;��H;e�H;��H;j�H;��H;c�H;��H;|�H;��H;1�H;. I;8I;I;�I;4I;E'I;�4I;�DI;KWI;�mI;��I;f�I;��I;��I;��I;��I;U�I;�	I;T%H;��F;�	E;�B;� @;�/=;##:;�07;U�4;�2;�51;      ��?;��?;��@;ctA;��B;K�C;�BE;[�F;p�G;dxH;�I;яI;{�I;��I;:�I;��I;�I;5�I;	�I;iI;�TI;�BI;�3I;I'I;�I;�I;I;�I;� I;��H;�H;k�H;a�H;��H;��H;.�H;��H;(�H;��H;��H;a�H;g�H;�H;��H;� I;�I;I;�I;�I;G'I;�3I;�BI;�TI;iI;�I;1�I;�I;��I;8�I;��I;{�I;ҏI;�I;dxH;n�G;X�F;�BE;A�C;
�B;ftA;��@;��?;      ��F;E�F;��F;\2G;'�G;&H;[�H;�I;�lI;��I;X�I;u�I;��I;��I;��I;��I;}�I;�wI;�bI;*PI;,@I;=2I;]&I;4I;}I;;I;I;I;��H;F�H;x�H;V�H;|�H;(�H;]�H;��H;��H;��H;[�H;'�H;�H;S�H;z�H;F�H;��H;I;I;AI;�I;3I;]&I;C2I;,@I;)PI;�bI;�wI;�I;��I;��I;��I;��I;s�I;^�I;��I;�lI;�I;^�H;�%H;?�G;q2G;��F;F�F;      u I;N'I;�:I;�XI;�{I;�I;��I;�I;�I;�I;Z�I;��I;p�I;�I;F�I;	�I;�lI;�ZI;gJI;"<I;�/I;�$I;#I;I;I;I;I;��H;v�H;��H;L�H;U�H;��H;��H;�H;��H;q�H;��H;�H;��H;��H;R�H;M�H;��H;q�H;��H;I;!I;I;I;%I;�$I;�/I;<I;fJI;�ZI;�lI;�I;D�I;�I;p�I;��I;[�I;�I;�I;�I;{�I;�I;�{I;�XI;�:I;6'I;      ��I;i�I;��I;��I;��I;%�I;��I;E�I;�I;x�I;��I;�I;�I;�I;�qI;�`I;�QI;�CI;&7I;�+I;)"I;pI;�I;I;�I;� I;��H;m�H;��H;V�H;T�H;��H;��H;��H;��H;��H;p�H;��H;��H;��H;��H;��H;U�H;V�H;��H;l�H;��H;I;�I;I;�I;tI;)"I;�+I;(7I;�CI;�QI;�`I;�qI;��I;�I;�I;��I;x�I;�I;E�I;��I;�I;��I;��I;��I;_�I;      ��I;�I;��I;]�I;��I;��I;��I;0�I;*�I;�I;q�I;�I;�pI;cbI;�TI;�GI;.<I;~1I;�'I;!I;aI;iI;~
I;8I;� I;��H;o�H;��H;Q�H;O�H;��H;P�H;?�H;��H;��H;��H;��H;��H;��H;��H;C�H;N�H;��H;N�H;O�H;��H;m�H;��H;� I;6I;
I;lI;^I;I;�'I;{1I;.<I;�GI;�TI;bbI;�pI;�I;v�I;�I;.�I;0�I;��I;��I;��I;`�I;��I;��I;      0�I;?�I;��I;�I;��I;�I;��I;s�I;z�I;vI;ujI;�^I;�SI;�HI;d>I;�4I;�+I;N#I;�I;�I;�I;?	I;nI;- I;��H;?�H;��H;X�H;U�H;��H;)�H;�H;8�H;��H;�H;��H;��H;��H;�H;��H;8�H;�H;,�H;��H;T�H;Z�H;��H;C�H;��H;- I;pI;C	I;�I;�I;�I;N#I;�+I;�4I;g>I;�HI;�SI;�^I;xjI;vI;z�I;p�I;ÖI;�I;��I;�I;��I;?�I;      g�I;��I;z�I; �I;8|I;`vI;�oI;hI;�_I;mWI;�NI;FI;�=I;15I;?-I;�%I;�I;*I;2I;�I;�I;vI;��H;.�H;�H;w�H;O�H;[�H;��H;0�H;�H;�H;T�H;��H;v�H;/�H;��H;,�H;u�H;��H;W�H;�H;�H;,�H;��H;[�H;M�H;z�H;�H;.�H;��H;yI;�I;�I;5I;,I;�I;�%I;?-I;.5I;�=I;FI;�NI;oWI;�_I;hI;�oI;[vI;?|I;�I;y�I;��I;      PdI;�cI;FbI;�_I;,\I;�WI;�RI;MI;GI;�@I;:I;^3I;�,I;j&I;4 I;MI;�I;�I;�
I;�I;�I;��H;��H;��H;m�H;O�H;R�H;��H;U�H;�H;�H;O�H;��H;#�H;��H;��H;��H;��H;��H;&�H;��H;O�H;	�H;�H;N�H;��H;R�H;P�H;p�H;��H;��H;��H;�I;�I;�
I;�I;�I;RI;7 I;j&I;�,I;\3I;:I;�@I;	GI;MI;�RI;�WI;5\I;�_I;QbI;�cI;      �KI;PKI;JI;HI;LEI;�AI;>I;�9I;�4I;�/I;�*I;�%I;| I;mI;I;�I;lI;.	I;=I;�I;��H;��H;��H;x�H;b�H;u�H;��H;��H;J�H;<�H;S�H;��H;�H;��H;J�H;�H;.�H;�H;H�H;��H;�H;��H;P�H;5�H;F�H;��H;��H;w�H;e�H;w�H;��H;��H;{�H;�I;?I;/	I;mI;�I;�I;mI;z I;�%I;�*I;�/I;�4I;�9I;>I;�AI;PEI; HI;JI;OKI;      �9I;z9I;�8I;7I;5I;p2I;`/I;�+I;)(I;0$I; I;�I;�I;{I;{I;�I;�I;sI;=I;7�H;}�H;�H;��H;��H;��H;!�H;��H;��H;��H;��H;��H;(�H;��H;7�H;��H;��H;��H;��H;��H;9�H;��H;(�H;��H;��H;��H;��H;��H; �H;��H;��H;��H;�H;x�H;2�H;@I;wI;�I;�I;{I;yI;�I;�I;
 I;1$I;,(I;�+I;h/I;n2I;5I;!7I;�8I;�9I;      b.I;=.I;b-I;,I;A*I;(I;�%I;�"I;�I;LI;�I;oI;�I;GI;�
I;vI;LI;9I;m�H;��H;��H;V�H;5�H;W�H;��H;Q�H;�H;��H;��H;�H;q�H;��H;J�H;��H;��H;��H;}�H;��H;��H;��H;K�H;��H;o�H;�H;��H;��H;�H;S�H;��H;W�H;8�H;U�H;��H;��H;m�H;;I;MI;xI;�
I;HI;�I;oI;�I;OI;�I;�"I;�%I;(I;=*I;
,I;a-I;?.I;      �'I;�'I;�&I;�%I;'$I;C"I;�I;vI;�I;�I;�I;sI;MI;*I;I;I;3I;j�H;��H;��H;^�H;/�H;B�H;��H;(�H;��H;��H;��H;��H;��H;-�H;��H; �H;��H;��H;c�H;p�H;f�H;��H;��H; �H;��H;,�H;��H;��H;��H;��H;��H;'�H;��H;F�H;/�H;W�H;��H;��H;m�H;5I;I;I;/I;MI;sI;�I;�I;�I;qI; I;C"I;)$I;�%I;�&I;�'I;      �%I;�%I;�$I;�#I;$"I;[ I;MI;�I;I;:I;YI;BI;BI;'
I;I;JI;�I;��H;��H;�H;��H;��H;�H;\�H;��H;��H;k�H;t�H;��H;��H;��H;��H;0�H;��H;}�H;j�H;v�H;o�H;z�H;��H;3�H;��H;��H;��H;��H;p�H;m�H;��H;��H;\�H;�H;��H;��H;�H;��H;�H;�I;MI;I;)
I;CI;AI;]I;=I;I;�I;RI;[ I;!"I;�#I;�$I;�%I;      �'I;�'I;�&I;�%I;)$I;F"I;�I;tI;�I;�I;�I;sI;NI;,I;I;I;3I;j�H;��H;��H;`�H;0�H;A�H;��H;(�H;��H;��H;��H;��H;��H;-�H;��H;!�H;��H;��H;c�H;q�H;f�H;��H;��H; �H;��H;,�H;��H;��H;��H;��H;��H;'�H;��H;F�H;.�H;V�H;��H;��H;m�H;5I;I;I;-I;MI;sI;�I;�I;�I;sI; I;D"I;)$I;�%I;�&I;�'I;      Y.I;?.I;^-I;�+I;A*I;(I;�%I;�"I;�I;MI;�I;pI;�I;FI;�
I;vI;JI;;I;m�H;��H;��H;V�H;4�H;V�H;��H;P�H;�H;��H;��H;�H;o�H;��H;J�H;��H;��H;��H;}�H;��H;��H;��H;M�H;��H;o�H;�H;��H;��H;�H;T�H;��H;V�H;9�H;W�H;��H;��H;m�H;<I;OI;yI;�
I;HI;�I;qI;�I;MI;�I;�"I;�%I;(I;@*I;,I;b-I;@.I;      �9I;{9I;�8I;7I;5I;u2I;`/I;�+I;,(I;0$I; I;�I;�I;yI;}I;�I;�I;wI;?I;7�H;}�H;�H;��H;��H;��H; �H;��H;��H;��H;��H;��H;(�H;��H;7�H;��H;��H;��H;��H;��H;7�H;��H;(�H;��H;��H;��H;��H;��H;!�H;��H;��H;��H;�H;t�H;5�H;BI;vI;�I;�I;|I;{I;�I;�I;
 I;1$I;,(I;�+I;j/I;t2I; 5I;"7I;�8I;~9I;      �KI;VKI;JI;�GI;JEI;�AI;>I;�9I;�4I;�/I;�*I;�%I;| I;nI;�I;�I;mI;1	I;?I;�I;��H;��H;��H;w�H;e�H;t�H;��H;��H;M�H;<�H;Q�H;��H;�H;��H;K�H;�H;/�H;�H;H�H;��H;�H;��H;Q�H;6�H;C�H;��H;��H;w�H;b�H;t�H;��H;��H;w�H;�I;@I;/	I;mI;�I;�I;nI;~ I;�%I;�*I;�/I;�4I;�9I;>I;�AI;NEI;HI;JI;SKI;      EdI;�cI;<bI;�_I;-\I;�WI;�RI;MI;	GI;�@I;:I;`3I;�,I;j&I;8 I;OI;�I;�I;�
I;�I;�I;��H;��H;��H;q�H;O�H;R�H;��H;W�H;�H;�H;P�H;��H;%�H;��H;��H;��H;��H;��H;(�H;��H;O�H;	�H;�H;R�H;��H;Q�H;Q�H;m�H;��H;��H;��H;�I;�I;�
I;�I;�I;RI;8 I;j&I;�,I;^3I;:I;�@I;
GI;MI;�RI;�WI;-\I;�_I;AbI;�cI;      ]�I;��I;|�I;��I;<|I;`vI;�oI;hI;�_I;kWI;�NI;FI;�=I;15I;@-I;�%I;�I;-I;5I;�I;�I;{I;��H;.�H;�H;u�H;O�H;[�H;��H;0�H;�H;�H;W�H;��H;{�H;/�H;��H;2�H;v�H;��H;W�H;�H;	�H;,�H;��H;V�H;L�H;x�H;�H;*�H;��H;{I;�I;�I;6I;,I;�I;�%I;@-I;25I;�=I;FI;�NI;kWI;�_I;hI;�oI;]vI;E|I;�I;~�I;��I;      6�I;D�I;��I;�I;��I;�I;��I;v�I;}�I; vI;qjI;�^I;�SI;�HI;i>I;�4I;�+I;R#I;�I;�I;�I;C	I;nI;. I;��H;?�H;��H;[�H;X�H;��H;,�H;�H;8�H;��H;�H;��H;��H;��H;�H;��H;;�H;�H;,�H;��H;R�H;W�H;��H;B�H;��H;) I;uI;B	I;�I;�I;�I;N#I;�+I;�4I;i>I;�HI;�SI;�^I;wjI;!vI;z�I;u�I;��I;�I;��I;�I;��I;<�I;      ��I;�I; �I;U�I;��I;��I;��I;0�I;4�I;�I;o�I;�I;�pI;cbI;�TI;�GI;-<I;1I;�'I;I;dI;lI;|
I;9I;� I;��H;o�H;��H;Q�H;N�H;��H;U�H;A�H;��H;��H;��H;��H;��H;��H;��H;C�H;P�H;��H;O�H;M�H;��H;l�H;��H;� I;2I;�
I;lI;^I;I;�'I;{1I;-<I;�GI;�TI;bbI;�pI;�I;u�I;�I;.�I;3�I;��I;��I;��I;V�I;��I;��I;      �I;_�I;��I;��I;��I;0�I;��I;M�I;�I;x�I;��I;�I;�I;��I;�qI;�`I;�QI;�CI;&7I;�+I;,"I;vI;�I;�I;�I;� I;��H;l�H;��H;T�H;V�H;��H;��H;��H;��H;��H;q�H;��H;��H;��H;��H;��H;U�H;V�H;��H;i�H;��H;� I;�I;|I;�I;tI;'"I;�+I;)7I;�CI;�QI;�`I;�qI;��I;�I;�I;��I;{�I;�I;E�I;��I;!�I;��I;��I;��I;_�I;      g I;T'I;�:I;�XI;�{I;"�I;~�I;�I;�I;�I;W�I;��I;m�I;�I;G�I;�I;�lI;�ZI;fJI;<I;�/I;�$I;!I;I;I;I;I;��H;w�H;��H;L�H;X�H;��H;��H;�H;��H;r�H;��H;�H;��H;��H;U�H;M�H;��H;q�H;��H;I; I;I;I;&I;�$I;�/I;"<I;iJI;�ZI;�lI;�I;G�I;�I;n�I;��I;Z�I;�I;�I;�I;��I;�I;�{I;�XI;�:I;@'I;      ��F;C�F;��F;_2G;0�G;&H;[�H;�I;�lI;��I;X�I;w�I;��I;��I;��I;��I;{�I;�wI;�bI;'PI;.@I;A2I;\&I;5I;�I;8I;I;I;��H;D�H;z�H;X�H;|�H;(�H;^�H;��H;��H;��H;Z�H;'�H;|�H;V�H;{�H;D�H;��H;I;I;<I;�I;1I;_&I;A2I;,@I;*PI;�bI;�wI;�I;��I;��I;��I;��I;q�I;\�I;��I;�lI;�I;^�H;�%H;:�G;b2G;��F;8�F;      ��?;��?;��@;gtA;��B;Q�C;�BE;[�F;p�G;fxH;�I;ԏI;y�I;��I;=�I;��I;�I;5�I;�I;iI;�TI;�BI;�3I;I'I;�I;|I;I;�I;� I;}�H;�H;n�H;`�H;��H;��H;+�H;��H;+�H;��H;��H;a�H;k�H;�H;}�H;� I;�I;I;�I;�I;H'I;�3I;�BI;�TI;iI;�I;2�I;�I;��I;>�I;��I;}�I;яI;�I;fxH;l�G;X�F;�BE;A�C;�B;ftA;��@;��?;      ��0;{51;�2;_�4;�07;;#:;�/=;� @;�B;�	E;��F;U%H;�	I;X�I;��I;��I;��I;�I;g�I;��I;�mI;KWI;�DI;�4I;E'I;-I;�I;I;<I;- I;0�H;��H;|�H;��H;d�H;��H;k�H;��H;a�H;��H;�H;��H;1�H;. I;8I;|I;I;1I;A'I;�4I;�DI;IWI;�mI;��I;j�I;��I;��I;��I;��I;X�I;�	I;T%H;��F;�	E;	�B;� @;�/=;0#:;�07;u�4;�2;f51;      M;�;(�;��;� ;�&;�\,;݇2;#98;�/=;�FA;urD;Y�F;JH;e9I;7�I;s�I;`�I;��I;��I;w�I;
pI;IXI;�DI;�3I;[&I;I;�I;�
I;lI;��H;��H;��H;��H;;�H;I�H;�H;H�H;8�H;��H;��H;��H;��H;pI;~
I;�I;%I;_&I;�3I;�DI;IXI;pI;v�I;��I;��I;Y�I;u�I;5�I;c9I;JH;[�F;rrD;�FA;�/=; 98;ۇ2;�\,;�&;� ;��;(�;�;      N��:��:��:��:и�:�P ;�e;�V;Q#;e-;��5;�h<;ZtA;^	E;�eG;A�H;9�I;�I;��I;�I;!�I;��I;pI;OWI;�BI;A2I;�$I;wI;pI;B	I;xI;��H;��H;�H;W�H;0�H;��H;3�H;V�H;�H;��H;��H;{I;D	I;lI;vI;�$I;D2I;�BI;RWI;pI;��I;�I;�I;��I;�I;8�I;?�H;�eG;]	E;YtA;�h<;��5;e-;T#;�V;�e;�P ;���:���:��:��:      ��p� �,�`"9�ų9�":��u:��:p��:��:4R;g ;��,;�6;Y)>;�;C;��F;�lH;rkI;{�I;��I;��I;�I;u�I;�mI;�TI;%@I;�/I;%"I;ZI;�I;�I;�I;u�H;u�H;��H;T�H;��H;V�H;��H;o�H;u�H;�I;�I;�I;VI;%"I;�/I;'@I;}TI;�mI;s�I;�I;��I;��I;|�I;mkI;�lH;��F;�;C;Y)>;�6;��,;g ;6R;��:p��:��:��u:$�":�ų9 #9 �,�      �o&�u!��4���氺ܬO� <T�u�9��u:�#�:�G�:D;3#;o71;E;;��A;�E;�$H;SVI;�I;��I;�I;��I; �I;iI;'PI;<I;�+I;I;�I;�I;�I;�I;7�H;��H;��H;�H;��H;��H;/�H;�I;�I;�I;�I;I;�+I; <I;*PI;iI;�I;��I;�I;��I;�I;TVI;�$H;�E;��A;B;;o71;1#;D;�G�:�#�:��u:�t�9 <T� �O�t氺����4�{!�      �kٻf�Ի�ǻ	����V���n���+��Ժķ1���39xm:��:v�;�;�\,;�8;Ņ@;E]E;�
H;SVI;{�I;��I;��I;i�I;�I;�bI;`JI;&7I;�'I;�I;/I;�
I;9I;;I;j�H;��H;z�H;��H;f�H;8I;8I;�
I;0I;�I;�'I;%7I;fJI;�bI; �I;l�I;��I;��I;y�I;TVI;�
H;A]E;Ņ@;�8;�\,;�;t�;��:|m:��39Է1��Ժ��+��n��V������ǻc�Ի      4yY��|U�I�I�>�7��� ��!���Ի�᝻��T� ��#��u�9���:el�:�;�);17;6 @;B]E;�$H;lkI;�I;\�I;�I;2�I;�wI;�ZI;�CI;}1I;N#I;)I;�I;-	I;sI;6I;j�H;��H;k�H;4I;rI;-	I;�I;)I;P#I;x1I;�CI;�ZI;�wI;+�I;�I;Y�I;�I;kkI;�$H;A]E;3 @;17;�);�;al�:���:�u�9�#� ���T��᝻��Ի�!��� �>�7�K�I��|U�      ��ü\l��u����R��=ߓ�^�{��M��� ���ż��}�B�갺@Fo��u:���:�R;:�';17;ą@;�E;�lH;8�I;o�I;��I;�I;x�I;�lI;�QI;,<I;�+I;�I;�I;eI;�I;BI;.I;�I;.I;?I;�I;cI;�I;�I;�+I;'<I;�QI;�lI;x�I;	�I;��I;o�I;8�I;�lH;�E;ą@;17;9�';�R;���:�u:@Fo�갺{�B�Ƽ���컇� ��M�]�{�>ߓ��R��v���[l��      �'�-$�^��W����?ټw��:���lyY��k���Ի3���X��X���($R:���:�R;�);�8;��A;��F;>�H;3�I;��I;��I;��I;�I;�`I;�GI;�4I;�%I;KI;�I;�I;qI;I;CI;I;mI;�I;�I;GI;�%I;�4I;�GI;�`I;�I;��I;��I;��I;0�I;=�H;��F;��A;�8;�);�R;���:$R:X����X��4����Ի�k�myY�:���w��?ټ���X�^��-$�      Y+����c̀�,l��Q�$�2�A��������@����>�V2��V��~1�@��($R:���:�;�\,;?;;�;C;�eG;b9I;��I;7�I;��I;B�I;�qI;�TI;c>I;9-I;1 I;zI;uI;�
I;I;
I;I;�
I;rI;zI;. I;8-I;`>I;�TI;�qI;C�I;��I;3�I;��I;^9I;�eG;�;C;A;;}\,;�;���:$R:`��~1�V��W2����>��@��������A�$�2��Q�-l�c̀���      j�ྲྀhܽo�н]y��^什O ��l��n<�L���>ټ��S|U�|������{1�8��� �u:al�:�;n71;`)>;]	E;JH;[�I;��I;��I;�I;ڃI;]bI;�HI;(5I;c&I;dI;qI;:I;!I;
I;%I;9I;qI;gI;_&I;&5I;�HI;]bI;ڃI;�I;��I;��I;[�I;JH;[	E;S)>;o71;�;al�:�u:X����1�����|��T|U��𛼿>ټL���n<�l�O ��^什]y��o�н�hܽ      ��4�f1��&���� ��h�ང�������`��'���SR��B�]�{��V���X�� Fo����:r�;3#;#�6;\tA;[�F;�	I;�I;��I;n�I;�I;�pI;�SI;�=I;�,I;v I;�I;�I;FI;9I;FI;�I;�I;y I;�,I;�=I;�SI;�pI;�I;n�I;��I;y�I;�	I;Y�F;YtA;�6;4#;p�;���:�Eo��X��V��{��B�]�SR����'��`��������h��������&�f1�      �x���o��ń�IUo���O�*�-�{��hܽ[什Ҽx���2�rb��SR��T|U�V2��3��갺�u�9��:D;��,;�h<;nrD;U%H;ΏI;j�I;��I;�I;
�I;�^I;FI;U3I;�%I;�I;\I;eI;5I;fI;\I;�I;�%I;S3I;FI;�^I;�I;�I;��I;j�I;ƏI;T%H;orD;�h<;��,;D;��:�u�9갺5��W2��T|U�TR��rb����2�Ӽx�[什�hܽ{�*�-���O�IUo�ń��o��      w���ྃ�Ѿ(����נ�ń�9�S��#�_O��{n��Ì���2���𛼀�>���Ի��B��#�\m:�G�:j ;��5;�FA;��F;�I;R�I;S�I;��I;o�I;njI;�NI;:I;�*I;�I;�I;�I;II;�I;�I;�I;�*I;:I;�NI;pjI;o�I;��I;S�I;Q�I;�I;��F;�FA;��5;^ ;�G�:Tm:�#���B���Ի��>�������2�Ì�{n��_O���#�9�S�ń��נ�(�����Ѿ��      �3���/��X#��	��A��֌Ⱦ�f��HUo�]1�ʰ��{n��Ҽx��'��>ټ�@���k�ȼ�����39�#�::R;e-;�/=;�	E;fxH;��I;�I;q�I;�I;vI;eWI;�@I;�/I;%$I;;I;�I;5I;�I;;I;#$I;�/I;�@I;eWI;vI;�I;s�I;�I;��I;_xH;�	E;�/=;e-;,R;�#�:`�39��Ǽ���k��@���>ټ�'�Ӽx�{n��ʰ��]1�HUo��f��֌Ⱦ�A���	��X#���/�      ���U���T�v��RZ�[58�͂�q��d���foy�]1�_O��[什�`�L�����myY��컐�T��1���u:��:O#;98;�B;r�G;�lI;�I;�I;2�I;x�I;�_I;GI;�4I;'(I;�I;�I;I;�I;�I;%(I;�4I;GI;�_I;v�I;1�I;�I;�I;�lI;n�G;�B;98;J#; ��:��u:�1���T���myY����L���`�[什_O��]1�foy�d���q��͂�[58��RZ�T�v�U���      	Ŀ7g��%ﱿ���T����U��X#�s��d���HUo��#��hܽ����n<����;����� ��᝻0�Ժ�t�9z��:�V;ԇ2;� @;^�F;�I;��I;C�I;+�I;k�I;hI;MI;�9I;�+I;�"I;lI;�I;iI;�"I;�+I;�9I;MI;hI;l�I;+�I;D�I;��I;�I;X�F;� @;և2;�V;b��:�t�92�Ժ�᝻�� �;�������n<�����hܽ�#�HUo�d���s���X#��U�T������%ﱿ7g��      ~x�P9�R��sؿnQ��e_��6�_��X#�q���f��9�S�{�����l�A�w���M���Ի��+�P<T���:�e;�\,;�/=;�BE;W�H;z�I;��I;��I;��I;�oI;�RI;>I;^/I;~%I;�I;GI;�I;�%I;^/I;>I;�RI;�oI;��I;��I;��I;}�I;]�H;�BE;0=;�\,;�e;��:P<T���+���Ի�M�w��A�l�����{�9�S��f��q���X#�6�_�e_��nQ��sؿR��P9�      �X1���,�h���<��6g��e_���U�͂�֌Ⱦń�*�-�h��O ��$�2�?ټ^�{� "��n��O���u:�P ;�&;0#:;A�C;�%H;�I;$�I;��I;�I;bvI;�WI;�AI;{2I;(I;D"I;a I;D"I;(I;{2I;�AI;�WI;]vI;�I;��I;(�I;�I;�%H;A�C;1#:;�&;�P ;��u:��O��n� "�_�{�?ټ$�2�O ��h��*�-�ń�֌Ⱦ͂��U�e_��6g��<�h����,�      d��]]�5K��X1�Zf��nQ��T���[58��A���נ���O���_什�Q����>ߓ��� ��V��n氺 �":��: ;�07;�B;0�G;�{I;��I;��I;��I;;|I;8\I;LEI;5I;3*I;4$I;,"I;0$I;6*I;5I;MEI;8\I;8|I;��I;��I;��I;�{I;;�G;�B;�07; ;��:�":n氺�V���� �>ߓ�����Q�_什����O��נ��A��[58�T���nQ���Zf��X1�5K��]]�      N������4z���V��X1��<�sؿ����RZ��	�(���IUo����]y��-l�X��R��@�7�
������0Ƴ9��:��;\�4;ntA;\2G;�XI;��I;N�I;�I;��I;�_I;�GI;#7I;�+I;�%I;�#I;�%I;�+I;"7I;�GI;�_I;��I;�I;N�I;��I;�XI;i2G;mtA;^�4;��;��:�ų9������@�7��R��X�-l�]y�����IUo�(����	��RZ����sؿ�<��X1���V��4z�����      �o��e^���ē��4z�5K�h��R��%ﱿT�v��X#���Ѿń��&�o�нc̀�^��t���H�I��ǻ�4��"9��::�;%�2;��@;��F;�:I;��I;��I;��I;z�I;NbI;�II;�8I;Z-I;�&I;�$I;�&I;\-I;�8I;JI;NbI;v�I;��I;��I;��I;�:I;��F;��@;"�2;6�;��:�"9�4��ǻH�I�t���^��c̀�o�н�&�ń���Ѿ�X#�T�v�%ﱿR��h��5K��4z��ē�e^��      q'���X��e^�������]]���,�P9�7g��U�����/����o��f1��hܽ���-$�]l���|U�a�Իw!� �,���:�;�51;��?;5�F;D'I;c�I;�I;@�I;��I;�cI;AKI;{9I;!.I;|'I;�%I;y'I;".I;{9I;BKI;�cI;��I;C�I;�I;g�I;D'I;E�F;��?;�51;�;{�: �,�w!�b�Ի�|U�]l���-$����hܽf1��o���ྙ�/�U���7g��P9���,��]]�����e^���X��      ����,������T���J�Q�ƙ$�3�����;�}�H(�@�׾�T���L+���սj��
��L���iO���ͻ��� "m8po�:`�;X�1;��?;�uF;j I;i�I;��I;��I;\vI;�WI;�AI;�1I;�'I;�!I;�I;�!I;�'I;�1I;�AI;�WI;YvI;��I;��I;k�I;j I;�uF;��?;U�1;[�;jo�: !m8�����ͻ�iO�L��
��j����ս�L+��T��@�׾H(�;�}���3���ƙ$�J�Q�T��������,��      �,��a��#P���{���K��x �����p�����w��$���Ҿf���  (���ѽѷ��&����ޔK�Aɻ#��@��8���:~�;��1;�@;m�F;!I;߿I;�I;��I;�uI;(WI;iAI;�1I;�'I;�!I;�I;�!I;�'I;�1I;jAI;)WI;�uI;��I;
�I;�I;"I;y�F;�@;��1;z�;x��:���8"��AɻޔK����&�ѷ����ѽ  (�f�����Ҿ�$���w�p��������x ���K��{�#P��a��      ����#P�������d���;�#���㿲���#f�d��ž��z���<�ƽ$0v�S5�0����o@�����vi� au9KK�:];�73;"�@;��F;JI;��I;R�I;V�I;�sI;�UI;E@I;�0I;�&I;!I;4I;!I;�&I;�0I;C@I;�UI;�sI;Z�I;S�I;��I;II;��F;$�@;�73;];CK�:�`u9ri������o@�0���S5�$0v�<�ƽ����z�žd��#f�������#����;���d����#P��      T����{���d��F�ř$�;����ɿ.蒿��K�P���j���Yb�F�0���r�a����=�����.��d��b�غ ��9�Y�:2X;�25;$�A;\!G;M7I;v�I;D�I;T�I;�pI;�SI;�>I;|/I;�%I;' I;2I;" I;�%I;{/I;�>I;�SI;�pI;V�I;G�I;v�I;L7I;d!G;#�A;�25;.X;�Y�:ذ�9^�غ�d����.�=������r�a�0���F��Yb��j��P����K�.蒿��ɿ;��ř$��F���d��{�      J�Q���K���;�ř$��;
��޿�����w�q,���澝���'�D������I��"�G�����N��������H�����9:b��:�n!;��7;��B;P�G;�YI;,�I;Z�I;��I;�lI;wPI;<I;�-I;$I;�I;�I;�I;$I;�-I;<I;vPI;�lI;ÒI;Z�I;/�I;�YI;U�G;��B;��7;�n!;`��:��9:B����������N�����"�G��I������'�D��������q,���w�����޿�;
�ř$���;���K�      ƙ$��x �#��;���޿o���ʅ���F�}�
��~����z��$���ս���?2+���ϼPp�����G�]� �*�$��:�;�8';��:;��C; H;�}I;�I;v�I;ًI;mgI;�LI; 9I;:+I;""I;�I;-I;�I;$"I;7+I;!9I;�LI;jgI;݋I;t�I;"�I;�}I;H;��C;��:;�8';�;��:�*�G�]�����Pp���ϼ?2+������ս�$���z��~��}�
��F�ʅ��o����޿;��#���x �      3��������㿊�ɿ���ʅ����P�d��<�׾�`��S�H����@��Q�a���̡���D��ɻ� �@׭��W�:�;dI-;9|=;#CE;��H;�I;��I;v�I;��I;iaI;#HI;�5I;r(I;�I;�I;TI;�I;�I;r(I;�5I;#HI;haI;��I;w�I;��I;�I;��H;$CE;;|=;dI-;�;�W�: ׭�� ��ɻ�D�̡����Q�a��@����S�H��`��<�׾d����P�ʅ�������ɿ�㿳���      ��p�������.蒿��w� �F�d��ʰ� ����Yb�)����ѽ�%��D4�ן�X����� H���潺��9Rr�:��;�93;*Q@;�vF;�H;�I;��I;��I;�zI;�ZI;CI;�1I;c%I;BI;�I;#I;�I;DI;e%I;�1I;CI;�ZI;�zI;��I;��I;	�I;�H;�vF;'Q@;�93;��;Hr�:��9�潺 H�����X��ן�D4��%����ѽ)���Yb� ���ʰ�d�� �F���w�.蒿����p���      ;�}���w�#f���K�q,�}�
�<�׾ �����k���'�dz꽝I���;V�<M�����iO�fG�ioE����@��:I� ;��$;��8;_�B;��G;2KI;�I;�I;A�I;qI;�SI;�=I;�-I;"I;nI;I;�I;I;nI;"I;�-I;�=I;�SI;qI;D�I;�I;�I;2KI; �G;_�B;��8;��$;G� ;N��:���joE�eG໩iO����<M��;V��I��dz���'���k� ���<�׾}�
�q,���K�#f���w�      G(��$�d��P������~���`���Yb���'��U�H$��C�m�%����ϼ�/��<��������غ�8�9D��:�F;�G.;|=;LE;�\H; �I;y�I;z�I;��I;gI; LI;�7I;)I;nI;rI;rI;%I;qI;rI;pI;)I;�7I;LI;
gI;��I;}�I;v�I;�I;�\H;KE;|=;�G.;�F;R��:�8�9��غ����<���/����ϼ%��C�m�H$���U���'��Yb��`���~�����P��d���$�      @�׾��Ҿž�j��������z�S�H�)��ez�H$���/v�2+�ې�����5��ɻ24��'�����:f��:=o!;P6;
lA;��F;u�H;��I;��I;�I;I}I;�\I;]DI;2I;r$I;�I;HI;�I;�I;�I;II;�I;p$I;2I;^DI;�\I;N}I;�I;��I;��I;z�H;��F;lA;P6;?o!;|��:���: (��.4��ɻ��5���ې�2+��/v�H$��dz�)��S�H���z������j��ž��Ҿ      �T��f�����z��Yb�&�D��$�����ѽ�I��C�m�2+�������G�K��ﻎ�p�:�����97T�:�/;x�-;j�<;HzD;_H;�mI;��I;��I;��I;�oI;�RI;�<I;,I;�I;
I;/I;�I;�I;�I;/I;I;�I; ,I;�<I;�RI;�oI;��I;~�I;��I;�mI;`H;MzD;q�<;x�-;�/;;T�:��94�����p���F�K�������2+�C�m��I����ѽ���$�'�D��Yb���z�f���      �L+�  (���F�������ս�@���%���;V�%��ې�����|MS�K��"��jD�@�n8q�:�;i�$;_7;.�A;i�F;��H;b�I;d�I;��I;߃I;TbI;�HI;5I;'&I;/I;=I;�I;�
I;
I;�
I;�I;=I;-I;$&I;5I;�HI;[bI;�I;��I;b�I;h�I; �H;l�F;4�A;_7;u�$;�;q�:��n8bD�"��J��|MS�����ې�%���;V��%���@����ս����F���  (�      ��ս��ѽ<�ƽ0����I�����Q�a�D4�<M���ϼ��G�K�L��LG��Wf�@�o���:�B�:�Y;��1;Vl>;�E;�/H;"qI;��I;��I;ژI;�rI;�UI;�>I;�-I;b I;�I;I;�
I;I;/I;I;�
I;�I;�I;` I;�-I;�>I;�UI;sI;ݘI;��I;�I;"qI;�/H;�E;Vl>;��1;�Y;�B�:��:@�o�Vf�HG��L��F�K�����ϼ;M�D4�Q�a�����I��0���<�ƽ��ѽ      j��ѷ��$0v�r�a�"�G�?2+���֟�����/����5���$��Xf��ج��g:E�:�;I-;g;;OC;SG;�I;̶I;�I;��I;	�I;
cI;~II;�5I;n&I;�I;5I;�I;�I;NI;XI;MI;�I;�I;5I;�I;u&I;�5I;�II;cI;�I;��I; �I;϶I;�I;SG;OC;"g;;"I-;�;O�:�g:xج�Tf�"������5��/�����֟���>2+�#�G�r�a�$0v�ѷ��      	��&�S5���������ϼˡ��X���iO�<���ɻ��p�vD�P�o� �g:`�:JG;t*;v9;��A;�uF;!�H;ÔI;��I;��I;H�I;�pI;3TI;N>I;-I;�I;{I;�I;VI;�I;�I;�I;�I;�I;VI;�I;zI;�I;!-I;T>I;:TI;�pI;D�I;��I;��I;ǔI;%�H;�uF;��A;z9;r*;LG;`�:�g:P�o�tD⺎�p��ɻ<���iO�X��ˡ����ϼ������S5�%�      L�����1���=����N��Pp��D����cG�����+4�6�����n8��:M�:OG;
�(;��7;`�@;��E;RQH;mI;��I;��I;��I;&}I;�^I;�FI;�3I;�$I;[I;�I;�	I;I;�I;��H;N�H;��H;�I;I;�	I;�I;aI;�$I;�3I;�FI;�^I;!}I;��I;��I;��I;mI;UQH;��E;d�@;��7;�(;QG;S�:��: �n80���(4�����bGໄ���D�Pp��N��>���2������      �iO�ܔK��o@���.���������ɻ�G��eoE���غ�'��В�9q�:�B�:�;t*;��7;�P@;�\E;�H;�II;��I;j�I;�I;Y�I;?hI;�NI;b:I;9*I;xI;�I;�I;I;I;2�H;a�H;��H;^�H;/�H;I;I;�I;�I;~I;:*I;f:I;�NI;<hI;a�I;�I;h�I;��I;�II;�H;�\E;�P@;��7;r*;�;�B�:q�:��9�'����غ_oE��G���ɻ����~����.��o@�ܔK�      ��ͻFɻ�����d�����5�]�� ��潺����8�9���:7T�:�;�Y;"I-;z9;`�@;�\E;��G;65I;��I;G�I;ݵI;V�I;dpI;�UI;V@I;4/I;{!I;�I;?I;�I;�I;!�H;��H;�H;��H;�H;��H;�H;�I;�I;DI;�I;}!I;9/I;V@I;�UI;lpI;Z�I;ٵI;L�I;��I;:5I;��G;�\E;f�@;y9;"I-;�Y;�;?T�:���:�8�9����潺� �<�]�����d������Fɻ      ���&��ki�H�غT����*� ֭���9L��:P��:z��:�/;o�$;��1;"g;;��A;��E;�H;75I;=�I;��I;O�I;��I;�vI;O[I;aEI;�3I;5%I;�I;�I;P	I;�I;|�H;a�H;'�H;��H;n�H;��H;$�H;`�H;�H;�I;T	I;�I;�I;9%I;�3I;_EI;W[I;�vI;��I;S�I;��I;?�I;:5I;�H;��E;��A;#g;;��1;o�$;�/;~��:R��:R��:��9�֭�؇*�F���b�غyi�-��      �*m8���8�_u9���9t�9:��:�W�:Vr�:G� ;�F;@o!;v�-; _7;Vl>;OC;�uF;TQH;�II;��I;��I;��I;��I;zI;�_I;@II;L7I;d(I;aI;�I;I;�I;* I;r�H;��H;�H;��H;t�H;��H;�H;��H;s�H;' I;�I;!I;�I;dI;d(I;L7I;FII;�_I;{zI;��I;��I;��I;��I;�II;WQH;�uF;OC;Ul>;_7;x�-;Do!;�F;E� ;Nr�:�W�:��:��9:Ȱ�9@`u9���8      ho�:���:kK�:�Y�:T��:"�;�;��;��$;�G.;P6;n�<;1�A;�E;SG;%�H;mI;��I;N�I;T�I;��I;�{I;xaI;�KI;�9I;�*I;�I;�I;�I;%I;� I;��H;��H;k�H;��H;�H;��H;�H;��H;k�H;��H;��H;� I;(I;�I;�I;�I;�*I;�9I;�KI;saI;�{I;��I;S�I;L�I;��I;mI;$�H;SG;�E;2�A;r�<;P6;�G.;��$;��;�;�;���:�Y�:SK�:���:      s�;~�;];>X;�n!;�8';pI-;�93;��8;|=;lA;SzD;n�F;�/H;�I;͔I;��I;o�I;ߵI;��I;zI;taI;yLI;#;I;b,I;3 I; I;�I;=I;�I;v�H;��H;e�H;m�H;
�H;U�H;"�H;O�H;�H;p�H;g�H;��H;z�H;�I;9I;�I; I;4 I;h,I;!;I;uLI;xaI;�zI;��I;�I;k�I;��I;˔I;�I;�/H;l�F;SzD;lA;|=;��8;�93;nI-;�8';�n!;@X;];f�;      X�1;��1;�73;�25;��7;��:;4|=;(Q@;[�B;NE;��F;`H;��H;$qI;̶I;��I;��I;�I;U�I;�vI;�_I;�KI;;I;�,I;� I;I;�I;I;tI;��H;q�H;n�H;!�H;��H;n�H;��H;��H;��H;m�H;��H;#�H;m�H;x�H;��H;qI;I;�I;I;� I;�,I;;I;�KI;�_I;�vI;S�I;�I;��I;��I;ͶI;qI;��H;`H;��F;KE;]�B;.Q@;2|=;��:;��7;�25;�73;��1;      ��?;�@;�@;�A;��B;�C;*CE;�vF; �G;�\H;|�H;�mI;e�I;
�I;#�I;��I;��I;d�I;rpI;\[I;LII;�9I;h,I;� I;qI;aI;�I;�I;i�H;��H;��H;-�H;U�H;��H;��H;^�H;4�H;X�H;��H;��H;U�H;(�H;��H;��H;f�H;�I;�I;cI;uI;� I;h,I;�9I;LII;Y[I;rpI;a�I;��I;��I;$�I;�I;f�I;�mI;~�H;�\H;��G;�vF;(CE;��C;¹B; �A;�@;�@;      �uF;{�F;��F;[!G;C�G;H;��H;#�H;5KI;(�I;��I;��I;f�I;��I;�I;M�I;+}I;AhI;�UI;_EI;P7I;�*I;1 I;I;^I;�I;HI;��H;��H;��H;$�H;>�H;��H;]�H;��H;�H;��H;�H;��H;^�H;��H;;�H;'�H;��H;��H;��H;EI;�I;cI;I;0 I;�*I;P7I;_EI;�UI;>hI;-}I;O�I; �I;��I;f�I;��I;��I;'�I;5KI; �H;��H; H;Z�G;m!G;��F;|�F;      x I;-I;EI;M7I;�YI;�}I;�I;�I;�I;y�I;��I;��I;��I;��I;	�I;�pI;�^I;�NI;Z@I;�3I;n(I;�I;$I;�I;�I;EI;��H;%�H;��H;2�H;"�H;i�H;�H;�H;��H;�H;��H;�H;�H;�H;�H;f�H;#�H;2�H;��H;#�H;��H;KI;�I;�I;$I;�I;l(I;�3I;X@I;�NI;�^I;�pI;�I;ژI;��I;��I;��I;x�I;�I;�I;�I;�}I;�YI;F7I;CI;I;      h�I;�I;��I;{�I;�I;"�I;��I;��I;�I;��I;�I;��I;��I;sI;cI;8TI;�FI;b:I;7/I;6%I;gI;�I;�I;I;�I;��H;"�H;��H;D�H;�H;W�H;��H;��H;�H;[�H;�H;��H;��H;Z�H;�H;��H;��H;Z�H;!�H;B�H;��H;!�H;��H;�I;I;�I;�I;eI;6%I;7/I;_:I;�FI;:TI;cI;sI;�I;��I;�I;��I;�I;��I;��I;�I;(�I;��I;��I;ݿI;      ��I; �I;O�I;W�I;P�I;v�I;|�I;��I;=�I;��I;M}I;�oI;VbI;�UI;�II;T>I;�3I;?*I;�!I;�I;�I;�I;9I;rI;d�H;��H;��H;C�H;2�H;U�H;��H;��H;��H;��H;|�H;5�H;.�H;1�H;z�H;��H;��H;��H;��H;U�H;/�H;C�H;��H;��H;j�H;pI;;I;�I;�I;�I;�!I;=*I;�3I;V>I;�II;�UI;UbI;�oI;S}I;��I;A�I;��I;|�I;m�I;Z�I;[�I;M�I;��I;      ��I;��I;d�I;P�I;��I;ًI;��I;�zI;qI;gI;�\I;�RI;�HI;�>I;�5I;-I;�$I;xI;�I;�I;%I;"I;�I;��H;��H;��H;2�H;#�H;[�H;��H;��H;��H;��H;�H;��H;|�H;]�H;y�H;��H;�H;��H;��H;��H;��H;X�H;%�H;/�H;��H;��H;��H;�I;(I;"I;�I;�I;wI;�$I;!-I;�5I;�>I;�HI;�RI;�\I;gI;qI;�zI;��I;ۋI;��I;[�I;a�I;��I;      YvI;�uI;�sI;�pI;�lI;ngI;jaI;�ZI;�SI;LI;bDI;�<I;5I;�-I;x&I;�I;fI;�I;GI;[	I;�I;� I;v�H;u�H;��H;$�H;#�H;^�H;��H;��H;��H;��H;��H;Z�H;�H;��H;��H;��H;�H;^�H;��H;��H;��H;��H;��H;[�H;"�H;(�H;��H;u�H;}�H;� I;�I;U	I;HI;�I;iI;�I;x&I;�-I;5I;�<I;dDI;LI;�SI;�ZI;saI;egI;�lI;�pI;�sI;�uI;      �WI;2WI;�UI;�SI;iPI;�LI;#HI;CI;�=I;�7I;	2I;,I;+&I;i I;�I;~I;�I;�I;�I;�I;4 I;��H;��H;k�H;-�H;6�H;f�H;��H;��H;��H;��H;��H;B�H;��H;|�H;A�H;K�H;A�H;{�H;��H;H�H;��H;��H;��H;��H;��H;f�H;:�H;1�H;h�H;�H;��H;0 I;�I;�I;�I;�I;�I;�I;i I;)&I;,I;2I;�7I;�=I;CI;,HI;�LI;sPI;�SI;�UI;2WI;      �AI;wAI;H@I;�>I;<I;9I;�5I;�1I;�-I;	)I;u$I;�I;2I;�I;:I;�I;�	I;I;�I;��H;��H;��H;d�H; �H;W�H;��H;�H;��H;��H;��H;��H;E�H;��H;\�H;�H;��H;��H;��H;�H;_�H;��H;H�H;��H;��H;��H;��H;�H;��H;\�H; �H;j�H;��H;z�H;��H;�I;I;�	I;�I;<I;�I;2I;�I;y$I;)I;�-I;�1I;�5I;9I;<I;�>I;Q@I;wAI;      �1I;�1I;�0I;t/I;�-I;0+I;u(I;j%I;	"I;zI;�I;I;GI;�I;�I;]I;I;I;&�H;i�H;��H;m�H;l�H;��H;��H;W�H;�H;�H;�H; �H;W�H;��H;]�H;��H;��H;��H;�H;��H;��H;��H;`�H;��H;W�H;�H;��H;�H;�H;X�H;��H;��H;s�H;k�H;��H;a�H;&�H;I;I;^I;�I;�I;EI;I;�I;{I;"I;h%I;|(I;,+I;�-I;y/I;�0I;�1I;      �'I;�'I;�&I;�%I;$I;"I;�I;NI;tI;�I;TI;@I;�I;�
I;�I;�I;�I;2�H;��H;+�H;�H;��H;�H;d�H;��H;��H;|�H;^�H;��H;��H;�H;~�H;�H;��H;�H;\�H;W�H;\�H;}�H;��H;�H;�H;�H;��H;|�H;X�H;|�H;��H;��H;d�H;
�H;��H;�H;'�H;��H;6�H;�I;�I;�I;�
I;�I;@I;[I;�I;uI;MI;�I; "I;$I;�%I;�&I;�'I;      �!I;�!I;!I;% I;�I;�I;�I;�I;I;|I;�I;�I;�
I;I;TI;�I;��H;^�H;�H;��H;��H;�H;L�H;��H;Z�H;�H;�H;�H;;�H;��H;��H;D�H;��H;��H;a�H;*�H;-�H;-�H;\�H;��H;��H;H�H;��H;{�H;7�H; �H;�H;�H;W�H;��H;P�H;�H;��H;��H;�H;b�H;��H;�I;WI;I;�
I;�I;�I;I;I;�I;�I;�I;�I;& I;!I;�!I;      �I;�I;DI;0I;�I;&I;ZI;-I;�I;+I;�I;�I;
I;;I;dI;�I;Z�H;��H;��H;v�H;��H;��H;�H;��H;1�H;��H;��H;��H;4�H;a�H;��H;M�H;��H;}�H;X�H;(�H;�H;*�H;T�H;~�H;��H;O�H;��H;\�H;.�H;��H;��H;��H;.�H;��H;"�H;��H;z�H;r�H;��H;��H;Z�H;�I;eI;@I;
I;�I;�I;,I;�I;,I;_I;&I;�I;6I;AI;�I;      �!I;�!I;!I;" I;�I;�I;�I;�I;I;}I;�I;�I;�
I;I;UI;�I;��H;_�H;�H;��H;��H;�H;L�H;��H;Z�H;�H;�H;�H;<�H;�H;��H;G�H;��H;��H;c�H;+�H;-�H;.�H;^�H;��H;��H;H�H;��H;y�H;7�H;��H;�H;�H;W�H;��H;R�H;�H;��H;��H;�H;b�H;��H;�I;WI;I;�
I;�I;�I;|I; I;�I;�I;�I;�I;* I;!I;�!I;      �'I;�'I;�&I;�%I;$I;"I;�I;QI;uI;�I;VI;BI;�I;�
I;�I;�I;�I;4�H;��H;,�H;�H;��H;�H;c�H;��H;��H;|�H;\�H;��H;��H;�H;~�H;�H;��H;��H;_�H;X�H;_�H;�H;��H;�H;�H;�H;��H;|�H;W�H;|�H;��H;��H;c�H;�H;��H;�H;%�H;��H;6�H;�I;�I;�I;�
I;�I;BI;[I;�I;uI;SI;�I;"I;$I;�%I;�&I;�'I;      �1I;�1I;�0I;x/I;�-I;4+I;u(I;o%I;"I;zI;�I;I;EI;�I;�I;^I;I;I;(�H;g�H;��H;n�H;l�H;��H;��H;W�H;�H;�H;�H;�H;W�H;��H;`�H;��H;��H;��H;��H;��H;��H;��H;`�H;��H;W�H;�H;��H;�H;�H;Z�H;��H;��H;q�H;k�H;��H;b�H;(�H;I;I;`I;�I;�I;EI;I;�I;zI;"I;l%I;~(I;2+I;�-I;y/I;�0I;�1I;      �AI;~AI;J@I;�>I;<I;9I;�5I;�1I;�-I;	)I;u$I;�I;3I;�I;?I;�I;�	I;I;�I;��H;��H;��H;d�H; �H;\�H;��H;�H;��H;��H;��H;��H;G�H;��H;]�H;�H;��H;��H;��H;�H;\�H;��H;H�H;��H;��H;��H;��H;�H;��H;W�H;�H;j�H;��H;w�H;��H;�I;I;�	I;�I;<I;�I;4I;�I;z$I;)I;�-I;�1I;�5I;9I;<I;�>I;W@I;xAI;      �WI;6WI;�UI;�SI;iPI;�LI;)HI;CI;�=I;�7I;2I;,I;)&I;h I;�I;�I;�I;�I;�I;�I;7 I;��H;��H;j�H;1�H;7�H;f�H;��H;��H;��H;��H;��H;E�H;��H;��H;A�H;M�H;F�H;|�H;��H;E�H;��H;��H;��H;��H;��H;c�H;7�H;-�H;c�H;�H;��H;. I;�I;�I;�I;�I;�I;�I;i I;,&I;,I;2I;�7I;�=I;CI;*HI;�LI;kPI;�SI;�UI;0WI;      QvI;�uI;�sI;�pI;�lI;mgI;laI;�ZI;�SI;
LI;dDI;�<I;5I;�-I;z&I;�I;iI;�I;GI;W	I;�I;� I;w�H;u�H;��H;!�H;#�H;^�H;��H;��H;��H;��H;��H;^�H;�H;��H;��H;��H;�H;`�H;��H;��H;��H;��H;��H;Z�H;!�H;&�H;��H;r�H;~�H;� I;�I;W	I;JI;�I;jI;�I;{&I;�-I;5I;�<I;gDI;LI;�SI;�ZI;saI;jgI;�lI;�pI;�sI;�uI;      ��I;��I;\�I;[�I;��I;�I;��I;�zI;qI;gI;�\I;�RI;�HI;�>I;�5I;!-I;�$I;zI;�I;�I;(I;'I;�I;��H;��H;��H;4�H;&�H;^�H;��H;��H;��H;��H;�H;��H;|�H;^�H;}�H;��H;�H;��H;��H;��H;��H;W�H;#�H;1�H;��H;��H;��H;�I;%I;"I;�I;�I;wI;�$I;#-I;�5I;�>I;�HI;�RI;�\I;gI;qI;�zI;��I;֋I;��I;b�I;g�I;��I;      ��I; �I;^�I;N�I;B�I;{�I;y�I;��I;E�I;��I;M}I;�oI;VbI;�UI;�II;V>I;�3I;A*I;�!I;�I;�I;�I;7I;tI;i�H;��H;��H;D�H;2�H;T�H;��H;��H;��H;��H;|�H;5�H;0�H;5�H;z�H;��H;��H;��H;��H;T�H;,�H;B�H;��H;��H;f�H;mI;=I;�I;�I;�I;�!I;=*I;�3I;Y>I;�II;�UI;XbI;�oI;Q}I;��I;A�I;��I;��I;t�I;R�I;P�I;^�I;��I;      s�I;ۿI;��I;}�I;�I;-�I;��I;��I;�I;��I;�I;��I;�I;sI;cI;:TI;�FI;c:I;6/I;5%I;hI;�I;�I;I;�I;��H;"�H;��H;G�H;�H;X�H;��H;��H;�H;^�H; �H;��H; �H;[�H;�H;��H;��H;[�H;�H;C�H;��H;"�H;��H;�I;I;�I;�I;dI;6%I;9/I;_:I;�FI;:TI;cI;sI;�I;��I;�I;��I;�I;��I;��I;�I;'�I;��I;��I;ۿI;      f I;0I;BI;X7I;�YI;�}I;�I;�I;�I;y�I;��I;��I;��I;ݘI;
�I;�pI;�^I;�NI;X@I;�3I;o(I;�I; I;�I;�I;DI;��H;&�H;��H;1�H;"�H;j�H;�H;�H;��H;�H;��H;�H;�H;�H;�H;l�H;#�H;1�H;��H;#�H;��H;II;�I;�I;'I;�I;i(I;�3I;Z@I;�NI;�^I;�pI;
�I;ܘI;��I;~�I;��I;x�I;�I;�I;�I;�}I;�YI;[7I;BI;I;      �uF;x�F;��F;\!G;J�G;H;��H;'�H;6KI;%�I;��I;��I;g�I;��I;�I;O�I;*}I;ChI;�UI;^EI;S7I;�*I;- I;I;aI;�I;GI;��H;��H;��H;'�H;@�H;��H;^�H;��H;�H;��H;�H;��H;]�H;��H;@�H;(�H;��H;��H;��H;HI;�I;`I;I;1 I;�*I;P7I;aEI;�UI;?hI;-}I;P�I;�I;��I;f�I;��I;��I;(�I;/KI;�H;��H;H;S�G;_!G;��F;m�F;      ��?;�@;�@; �A;��B;
�C;(CE;�vF;�G;�\H;|�H;�mI;e�I;�I;'�I;��I;��I;f�I;spI;Z[I;MII;�9I;h,I;� I;vI;\I;�I;�I;k�H;��H;��H;1�H;U�H;��H;��H;[�H;3�H;[�H;��H;��H;V�H;.�H;��H;��H;f�H;�I;�I;`I;qI;� I;k,I;�9I;LII;\[I;upI;a�I;��I;��I;'�I;	�I;h�I;�mI;|�H;�\H;��G;�vF;-CE;��C;��B; �A;�@;�@;      9�1;��1;�73;�25;~�7;��:;4|=;+Q@;`�B;IE;��F;dH;��H;#qI;϶I;��I;��I;�I;U�I;�vI;�_I;�KI;;I;�,I;� I;I;�I;I;uI;��H;t�H;t�H;$�H;��H;p�H;��H;��H;��H;k�H;��H;&�H;o�H;w�H;��H;qI;I;�I;I;� I;�,I;;I;�KI;�_I;�vI;Y�I;�I;��I;��I;϶I;"qI;��H;`H;��F;LE;[�B;'Q@;7|=;��:;��7;�25;�73;��1;      l�;~�;];LX;�n!;�8';jI-;�93;��8;|=;lA;VzD;l�F;�/H;�I;ДI;��I;r�I;�I;��I;�zI;xaI;vLI;#;I;i,I;- I;I;�I;@I;�I;x�H;�H;g�H;m�H;�H;U�H;%�H;S�H;�H;l�H;e�H;�H;{�H;�I;9I;�I;$I;1 I;d,I;!;I;wLI;waI;�zI;��I;�I;j�I;��I;͔I;�I;�/H;o�F;RzD;lA;|=;��8;�93;jI-;�8';�n!;JX;];j�;      ho�:���:QK�:�Y�:V��:(�;�;��;��$;�G.;P6;u�<;2�A;�E;SG;)�H;mI;��I;L�I;V�I;��I;�{I;waI;�KI;�9I;�*I;�I;�I;�I;%I;� I;��H;��H;k�H;��H;�H;��H;�H;��H;j�H;��H;��H;� I;(I;�I;�I;�I;�*I;�9I;�KI;waI;�{I;��I;V�I;N�I;��I;mI;'�H;SG;�E;2�A;q�<;P6;�G.;��$;��;�;�;���:�Y�:OK�:���:       (m8���8�`u9ذ�9t�9:,��:�W�:Rr�:L� ;�F;Co!;y�-;_7;Vl>;
OC;�uF;WQH;�II;��I;��I;��I;��I;~zI;�_I;GII;I7I;a(I;bI;�I;I;�I;- I;u�H;��H;�H;��H;u�H;��H; �H;��H;s�H;* I;�I;I;�I;bI;g(I;L7I;BII;�_I;|zI;��I;��I;��I;��I;�II;WQH;�uF;OC;Vl>;_7;x�-;Do!;�F;H� ;\r�:�W�:$��:��9:��9pau9 ��8      t��"��ri�D�غV���؇*��֭�8��9\��:R��:~��:�/;p�$;��1;%g;;��A;��E;�H;75I;@�I;��I;T�I;��I;�vI;W[I;^EI;�3I;6%I;�I;�I;T	I;�I;�H;b�H;'�H;��H;p�H;��H;$�H;^�H;}�H;�I;T	I;�I;�I;5%I;�3I;_EI;R[I;�vI;��I;Q�I;��I;?�I;95I;�H;��E;��A;#g;;��1;p�$;�/;���:L��:R��:��9`֭��*�F���\�غsi�)��      ��ͻFɻ�����d�����5�]�� ��潺����8�9���:?T�:�;�Y;(I-;}9;c�@;�\E;��G;95I;��I;L�I;ߵI;V�I;npI;�UI;T@I;4/I;!I;�I;CI;�I;�I;"�H;��H;�H;��H;�H;��H;�H;�I;�I;DI;�I;{!I;4/I;W@I;�UI;gpI;Z�I;ݵI;J�I;��I;:5I;��G;�\E;a�@;w9;"I-;�Y;�;=T�:���:�8�9����潺� �9�]�����d������Cɻ      �iO�۔K��o@���.��������ɻ�G��aoE���غ�'����9q�:�B�:�;v*;��7;�P@;�\E;�H;�II;��I;n�I;�I;a�I;<hI;�NI;c:I;<*I;xI;�I;�I;I;I;0�H;^�H;��H;a�H;-�H;I;I;�I;�I;zI;9*I;c:I;�NI;>hI;Z�I;�I;k�I;��I;�II;�H;�\E;�P@;��7;t*;�;�B�:q�:��9�'����غboE��G���ɻ��������.��o@�۔K�      L�����1���=����N��Pp��D����cG�����)4�.�����n8��:U�:SG;�(;��7;`�@;��E;UQH;mI;��I;��I;��I;$}I;�^I;�FI;�3I;�$I;^I;�I;�	I;I;�I;��H;P�H;��H;�I;I;�	I;�I;_I;�$I;�3I;�FI;�^I;$}I;��I;��I;��I;mI;QQH;��E;`�@;��7;
�(;OG;S�:��:@�n84���(4�����bGໄ���D�Pp��N��>���2������      	��&�S5���������ϼˡ��X���iO�<���ɻ��p�pD�P�o��g:`�:KG;t*;w9;��A;�uF;'�H;ʔI;��I;��I;H�I;�pI;3TI;T>I;-I;�I;}I;�I;ZI;�I;�I;�I;�I;�I;TI;�I;zI;�I;-I;Q>I;5TI;�pI;F�I;��I;��I;ȔI;$�H;�uF;��A;u9;p*;KG;`�:�g:@�o�vD⺏�p��ɻ<���iO�X��̡����ϼ������T5�&�      j��ѷ��$0v�q�a�"�G�>2+���֟�����/����5���"��Vf�Xج��g:O�:�;I-; g;;OC;SG;�I;ͶI;!�I; �I;�I;cI;�II;�5I;q&I;�I;5I;�I;�I;LI;XI;MI;�I;�I;5I;�I;p&I;�5I;�II;cI;�I; �I;�I;϶I;�I;SG;�NC; g;;I-;�;O�:�g:xج�Vf�#������5��/�����֟���>2+�#�G�r�a�%0v�ѷ��      ��ս��ѽ<�ƽ0����I�����Q�a�D4�;M���ϼ��F�K�L��HG��Sf���o���:�B�:�Y;��1;Yl>;�E;�/H;#qI;�I;��I;ژI; sI;�UI;�>I;�-I;b I;�I;�I;�
I;I;/I;I;�
I;�I;�I;` I;�-I;�>I;�UI;sI;ژI;��I;��I;&qI;�/H;�E;Pl>;��1;�Y;�B�:��: �o�Wf�HG��L��G�K�����ϼ;M�D4�Q�a�����I��0���<�ƽ��ѽ      �L+�  (���F�������ս�@���%���;V�%��ڐ�����{MS�J����fD�@�n8q�:�;p�$;_7;2�A;o�F; �H;i�I;c�I;��I;��I;XbI;�HI;5I;'&I;/I;@I;�I;�
I;
I;�
I;�I;=I;-I;"&I;5I;�HI;XbI;��I;��I;c�I;c�I;��H;n�F;1�A;�^7;r�$;�;q�:@�n8hD�!��J��|MS�����ڐ�%���;V��%���@����ս����F���  (�      �T��f�����z��Yb�&�D��$�����ѽ�I��C�m�2+�������F�K��ﻋ�p�:���В�9;T�:�/;|�-;n�<;OzD;cH;�mI;��I;|�I;��I;�oI;�RI;�<I;,I;�I;I;/I;�I;�I;�I;-I;I;�I; ,I;�<I;�RI;�oI;��I;z�I;��I;�mI;`H;PzD;m�<;r�-;�/;7T�:���94�����p���G�K�������2+�C�m��I����ѽ���$�'�D��Yb���z�f���      @�׾��Ҿž�j��������z�S�H�)��ez�H$���/v�2+�ې�����5��ɻ24� (�����:t��:Do!;P6;lA;��F;z�H;��I;��I;�I;L}I;�\I;^DI;2I;r$I;�I;FI;�I;�I;�I;FI;�I;p$I;2I;]DI;�\I;L}I;�I;��I;��I;t�H;��F;lA;P6;9o!;t��:���:(��.4��ɻ��5���ې�2+��/v�H$��dz�)��S�H���z������j��ž��Ҿ      G(��$�d��P������~���`���Yb���'��U�H$��C�m�%����ϼ�/��<��������غ�8�9P��:�F;�G.;|=;OE;�\H; �I;v�I;y�I;��I;gI;LI;�7I;)I;qI;oI;qI;'I;qI;qI;nI;)I;�7I;LI;gI;��I;|�I;u�I;�I;�\H;NE;|=;�G.;�F;P��:�8�9��غ����<���/����ϼ%��C�m�H$���U���'��Yb��`���~�����P��d���$�      ;�}���w�#f���K�q,�}�
�<�׾ �����k���'�dz꽝I���;V�<M�����iO�eG�joE����L��:N� ;��$;��8;b�B;�G;/KI;�I;�I;D�I;	qI;�SI;�=I;�-I;"I;jI;I;�I;I;kI;"I;�-I;�=I;�SI;	qI;D�I;�I;�I;3KI;��G;c�B;��8;��$;D� ;R��:���hoE�eG໨iO����<M��;V��I��dz���'���k� ���<�׾}�
�q,���K�#f���w�      ��p�������.蒿��w� �F�d��ʰ� ����Yb�)����ѽ�%��D4�ן�X�����H���潺 ��9\r�:��;�93;.Q@;�vF;�H;	�I;��I;��I;�zI;�ZI;CI;�1I;c%I;@I;�I;"I;�I;BI;b%I;�1I;CI;�ZI;�zI;��I;��I;�I;�H;~vF;+Q@;�93;��;Dr�:��9�潺 H�����X��ן�D4��%����ѽ)���Yb� ���ʰ�d�� �F���w�.蒿����p���      3��������㿊�ɿ���ʅ����P�d��<�׾�`��S�H����@��Q�a���̡���D��ɻ� ��֭��W�:�;fI-;>|=;$CE;��H;�I;��I;w�I;��I;laI;#HI;�5I;r(I;�I;�I;SI;�I;�I;r(I;�5I;%HI;iaI;��I;v�I;��I;�I;��H;!CE;>|=;jI-;�;�W�:�֭�� ��ɻ�D�̡����Q�a��@����S�H��`��<�׾d����P�ʅ�������ɿ�㿳���      ƙ$��x �#��;���޿o���ʅ���F�}�
��~����z��$���ս���?2+���ϼPp�����F�]��*�&��:�;�8';��:;��C;�H;�}I;�I;t�I;ۋI;ogI;�LI;9I;:+I;!"I;�I;-I;�I;""I;9+I; 9I;�LI;kgI;ڋI;s�I;"�I;�}I;H;��C;��:;�8';�;��:�*�G�]�����Pp���ϼ?2+������ս�$���z��~��}�
��F�ʅ��o����޿;��#���x �      J�Q���K���;�ř$��;
��޿�����w�q,���澝���'�D������I��"�G�����N��������B�����9:h��:�n!;��7;��B;J�G;�YI;+�I;\�I;��I;�lI;vPI;<I;�-I;$I;�I;�I;�I;$I;�-I;<I;uPI;�lI;��I;\�I;.�I;�YI;U�G;��B;��7;�n!;b��:��9:@����������N�����"�G��I������'�D��������q,���w�����޿�;
�ř$���;���K�      T����{���d��F�ř$�;����ɿ.蒿��K�P���j���Yb�F�0���r�a����=�����.��d��\�غ��9�Y�:0X;�25;$�A;X!G;I7I;t�I;D�I;S�I;�pI;�SI;�>I;}/I;�%I;& I;3I;# I;�%I;y/I;�>I;�SI;�pI;W�I;F�I;w�I;L7I;d!G;#�A;�25;.X;�Y�:ذ�9\�غ�d����.�=������r�a�0���F��Yb��j��P����K�.蒿��ɿ;��ř$��F���d��{�      ����#P�������d���;�#���㿲���#f�d��ž��z���<�ƽ$0v�S5�0����o@�����ui� au9IK�:];�73;%�@;��F;II;��I;R�I;V�I;�sI;�UI;B@I;�0I;�&I;!I;4I;!I;�&I;�0I;C@I;�UI;�sI;Z�I;S�I;��I;JI;��F;$�@;�73;];CK�:�`u9qi������o@�0���S5�$0v�<�ƽ����z�žd��#f�������#����;���d����#P��      �,��a��#P���{���K��x �����p�����w��$���Ҿf���  (���ѽѷ��&����ߔK�@ɻ"��`��8���:~�;��1;�@;k�F;!I;߿I;�I;��I;�uI;(WI;iAI;�1I;�'I;�!I;�I;�!I;�'I;�1I;jAI;*WI;�uI;��I;�I;�I;#I;{�F;�@;��1;z�;z��:���8 ��BɻޔK����&�ѷ����ѽ  (�f�����Ҿ�$���w�p��������x ���K��{�#P��a��      ඕ�S���Ѭ��-�_���7�z�}߿����,b��V�,l¾Hx�c.���Ž��t�)��d����?�N��!����x9���:R�;��2;3@@;`fF;9�H;��I;S�I;!|I;�[I;�CI;2I;�%I;_I;�I;4I;�I;^I;�%I;	2I;�CI;�[I;&|I;R�I;��I;<�H;mfF;3@@;��2;J�;���:`�x9��N����?�d��)����t���Žc.�Hx�,l¾�V��,b����}߿z���7�-�_�Ѭ��S���      S���D���#}��+Y��3�����$ڿ%��ý\����(���s��3�5����p�b�S���<<�5���������9O��:һ;R%3;Ep@;�yF;��H;��I;�I;�{I;O[I;RCI;�1I;U%I;!I;[I;I;WI;#I;T%I;�1I;SCI;K[I;�{I;�I;��I;��H;�yF;Gp@;O%3;˻;I��:`��9����5���<<�S��b��p�5����3��s�(�����Ľ\�$���$ڿ����3��+Y�#}�D���      Ѭ��#}�>tf��lG�ע%��p�.�ʿZ����>M����T�����d�Ȥ�̷�-�d��
��I���1�c���X��Ь�9���:;�U4;��@;ӱF;4�H;܎I;��I;�yI;�YI;<BI;�0I;�$I;�I;�I;�I;�I;�I;�$I;�0I;<BI;�YI;�yI;��I;ގI;4�H;߱F;��@;�U4;;���:���9P��d����1��I���
�.�d�̷�Ȥ���d�T�������>M�Z���.�ʿ�p�ע%��lG�>tf�#}�      -�_��+Y��lG�f.�z���꿱���M䂿��5���󾍰��N�N�V��R�� �Q����|����h!��g��`�|	:_
�:��;`16;��A;;G;I;9�I;x�I;nvI;LWI;n@I;o/I;�#I;�I;I;�I;	I;�I;�#I;n/I;n@I;HWI;qvI;{�I;9�I; I;DG;��A;\16;��;[
�:d	:Z񳺉g���h!�|������ �Q�R��V��N�N���������5�M䂿�������z�f.��lG��+Y�      ��7��3�ע%�z��<����ſ	���½\�<����Ͼ����`�3��轻z��|�9�^�Ἒ���z��7}��dt�(�^:e+�:��#;��8;��B;sG;q%I;��I;�I;
rI;TI;�=I;t-I;"I;MI;�I;~I;�I;NI;"I;t-I;�=I;TI;rI;�I;��I;q%I;sG;��B;��8;��#;c+�:�^:xdt��7}��z����^��|�9��z����`�3�������Ͼ<��½\�	�����ſ�<��z�ע%��3�      z�����p������ſ$���Ps���1�1r���d���d�|I�ΈŽ��}�_*�IC���^��B�v�D��F๘ �:��;p);7;;*D;4�G;WHI;��I;��I;�lI;�OI;�:I;+I; I;�I;}I;/I;yI;�I; I;+I;�:I;�OI;�lI;��I;��I;THI;=�G;*D;7;;n);��;� �:�F�w�D��B��^�IC��_*���}�ΈŽ|I��d��d��1r����1��Ps�$����ſ��꿃p����      }߿�$ڿ.�ʿ����	����Ps�PX:����%l¾�ǆ���7����75���Q�����t���75�f�����@�8�ɼ:��;��.;��=;�EE;�YH;�hI;$�I;��I;(fI;KI;&7I;H(I;�I;�I;�I;xI;�I;�I;�I;H(I;%7I;KI;,fI;��I;$�I;�hI;�YH;�EE;��=;��.;��;�ɼ:��8���h���75��t������Q�75�������7��ǆ�%l¾���PX:��Ps�	�������.�ʿ�$ڿ      ���$��Z���M䂿½\���1�����J˾青�D�N�x��H������U�'�c�Ҽ��|��z��n��>x����&:�P�:��;�W4;Ҡ@;%gF;c�H;�I; �I;2�I;_I;�EI;3I;!%I;DI;�I;�I;�I;�I;�I;GI;#%I;3I;�EI;#_I;2�I;"�I;�I;e�H;(gF;͠@;�W4;��;�P�:��&:>x���n���z���|�c�ҼU�'����H���x��D�N�青��J˾�����1�½\�M䂿Z���$��      �,b�ý\��>M���5�<��1r��%l¾蝒�"&W��3�8Sؽ�z��YG����zI����?���̻��-�h
����:��;��&;|9;�C;�dG;KI;A�I;Q�I;RvI;}WI;*@I;�.I;�!I;�I;XI;�I;�I;�I;XI;�I;�!I;�.I;*@I;�WI;SvI;T�I;?�I;NI;�dG;�C;!|9;��&;��;"��:h
����-���̻��?�zI�����YG��z��8Sؽ�3�"&W�青�%l¾1r��<����5��>M�ý\�      �V������������Ͼ�d���ǆ�D�N��3��c�[����\�2��(C���o���	��눻H����9��:�h;R�/;7�=;IE;�2H;�WI;��I;��I;�kI;�OI;":I;�)I;$I;�I;�I;�I;yI;�I;�I;�I;$I;�)I;$:I;�OI;�kI;��I;��I;�WI;�2H;HE;=�=;T�/;�h;#��:���9L��눻��	��o�(C��2����\�[���c཰3�D�N��ǆ��d����Ͼ���������      ,l¾(��T������������d���7�x��8Sؽ[���d�C*�bkּ,\����'�'���R�~��|�:�Z;ԣ#;==7;*�A;�F;V�H;o�I;�I;��I;�`I;�GI;�3I;&%I;rI;�I;SI;K
I;J	I;M
I;UI;�I;tI;$%I;�3I;�GI;�`I;��I;�I;l�I;[�H;�F;.�A;@=7;ӣ#;�Z;��:~���R�&����'�+\��bkּC*��d�[��8Sؽx����7��d���������T���(��      Gx��s���d�N�N�`�3�|I����H����z����\�C*�
�ݼH���.<<��ڻ�V�0dt�@�&:���:=C;�</;QD=;ԈD;��G;�8I;ǘI;��I;tI;'VI;\?I;�-I;b I;�I;YI;�
I;�I;I;�I;�
I;\I;�I;a I;�-I;a?I;/VI;tI;��I;ŘI;�8I;��G;ڈD;VD=;�</;IC;���:8�&: dt��V��ڻ,<<�H���
�ݼB*���\��z��H������|I�`�3�N�N���d��s�      c.��3�Ȥ�V����ΈŽ75�����YG�2��bkּH����xC��>�c6}���� �x9p��:	;/�&;�;8;��A;��F;��H;0yI;��I;��I;1fI;�KI;K7I;|'I;�I;�I;WI;I;�I;�I;�I;I;WI;�I;�I;�'I;S7I;�KI;4fI;��I;��I;7yI;��H;��F;��A;�;8;:�&;	;j��:`�x9���b6}��>��xC�H���bkּ2��YG����75��ΈŽ��V��Ȥ��3�      ��Ž4���̷�R���z����}��Q�U�'����(C��+\��-<<��>n��8����6��:6��:�;�'3;��>;�E;fH;a<I;˗I;��I;�vI;�XI;�AI;u/I;�!I;�I;�I;Q	I;bI;"I;rI;"I;aI;S	I;�I;�I;�!I;/I;�AI;�XI;�vI;��I;җI;a<I;kH;�E;��>;�'3;�;6��:D��:@�6�຀n���>�,<<�+\��(C�����U�'��Q���}��z��R��̷�4���      ��t��p�-�d� �Q�|�9�^*����a�ҼzI���o���'��ڻe6}�:��@9���:^m�:��;��.;<;�oC;?7G;��H;ՁI;ӜI;҅I;"fI;<LI;�7I;�'I;�I;tI;LI;GI;�I;� I;O I;� I;�I;HI;NI;rI;�I;�'I;�7I;ELI;"fI;ЅI;ٜI;ցI;��H;C7G;�oC;<;��.;��;hm�:��: 9�2��b6}��ڻ��'��o�yI��b�Ҽ���^*�}�9� �Q�.�d��p�      '��b��
����^��IC���t����|���?���	�&���V���� ���:��:�h;$�+;��9;��A;|fF;X�H;t_I;��I;��I;sI;�VI;r@I;�.I;� I;TI;I;�I;hI;M I;|�H;�H;{�H;J I;hI;�I;I;[I;� I;�.I;y@I;�VI;�rI;��I;��I;w_I;]�H;fF;��A;��9;!�+;�h;��:��:������V�$����	���?���|��t��HC��^������
�a�      b��R���I��|�������^��75��z���̻�눻�R�(dt�P�x9>��:fm�:�h;_�*;ߍ8;��@;�E;:(H;g8I;��I;�I;H~I;�`I;�HI;�5I;[&I;tI;2I;�	I;�I;� I;��H;V�H;��H;Q�H;��H;� I;�I;�	I;8I;xI;]&I;�5I;�HI;�`I;Q~I;�I;��I;k8I;=(H;�E;��@;ۍ8;c�*;�h;nm�:F��:0�x9 dt��R��눻��̻�z��75��^����|����I��P��      ��?��<<��1��h!��z��B�a���n����-�>��}��0�&:`��:0��:��;�+;׍8;A�@;�]E;h�G;GI;�I;Q�I;8�I;jiI;:PI;<I;�+I;�I;nI;OI;)I;qI;��H;��H;O�H;��H;M�H;��H;��H;pI;)I;VI;uI;�I;�+I;<I;7PI;riI;8�I;O�I;�I;JI;n�G;�]E;@�@;܍8; �+;��;6��:f��:8�&:�}��>𳺁�-��n��b���B黳z��h!��1��<<�      
N��:��b����g���7}�e�D����.x��8
�����9��:���:	;�;��.;��9;��@;�]E;l�G;?I;�I;�I;M�I;�pI;�VI;�AI;}0I;�"I;�I;�I;�I;�I;��H;^�H;w�H;^�H;��H;^�H;t�H;]�H;��H;�I;�I;�I;�I;�"I;~0I;�AI;�VI;�pI;J�I;
�I;�I;DI;p�G;�]E;��@;��9;��.;�;	;���:��:���98
��0x�����k�D��7}��g��b���:��      !������:��@񳺔dt��F๠�8��&:"��:%��:�Z;FC;6�&;�'3;<;��A;�E;p�G;@I;[|I;ÜI;��I;~uI;r[I;FI;�4I;+&I;�I;II;�	I;�I;9�H;��H;6�H;t�H;~�H;�H;x�H;q�H;5�H;��H;7�H;�I;�	I;II;�I;,&I;�4I;FI;u[I;}uI;��I;ʜI;_|I;FI;n�G;�E;��A;<;�'3;5�&;KC;�Z;%��:&��:��&:@�8�F�xdt�Z�V�ິ���      ��x9��9��9`	:��^:� �:�ɼ:�P�:��;�h;ԣ#;�</;�;8;��>;�oC;�fF;<(H;NI;�I;��I;��I;�wI;p^I;;II;�7I;)I;	I;�I;�I;GI;J I;I�H;S�H;:�H;��H;��H;��H;��H;��H;9�H;S�H;E�H;P I;LI;�I;�I;	I;)I;�7I;;II;m^I;�wI;��I;ĜI;�I;LI;>(H;�fF;�oC;��>;�;8;�</;ڣ#;�h;��;�P�:�ɼ:� �:(�^:l	:x��98��9      ���:s��:���:y
�:Y+�:��;��;��;��&;V�/;C=7;SD=;��A;�E;C7G;_�H;l8I;��I;
�I;��I;�wI;�_I;�JI;�9I;�*I;�I;5I;<I;I;9I;��H;��H;�H;<�H;��H;�H;��H;�H;��H;=�H;�H;��H;�H;<I;I;?I;5I;�I;�*I;�9I;�JI;�_I; xI;��I;�I;�I;o8I;^�H;F7G;�E;��A;XD=;F=7;T�/;��&;��;��;��;�+�:i
�:���:_��:      h�;һ;;��;��#;z);��.;�W4;(|9;>�=;4�A;ވD;��F;tH;��H;|_I;œI;U�I;M�I;�uI;p^I;�JI;':I;#,I;8 I;�I;OI;�I;!I;��H;��H;4�H;�H;k�H;c�H;��H;U�H;��H;c�H;n�H;�H;3�H;�H;��H;I;�I;OI;�I;< I; ,I;$:I;�JI;t^I;�uI;Q�I;Q�I;œI;{_I;��H;nH;��F;ވD;9�A;<�=;'|9;�W4;��.;t);��#;��;;��;      ��2;]%3;�U4;Y16;��8;!7;;��=;Р@;�C;JE;�F;��G;��H;d<I;ӁI;��I;�I;9�I;�pI;o[I;9II;�9I;,I;� I;I;I;TI;�I;H�H;d�H;\�H;*�H;:�H;��H;��H;a�H;�H;[�H;��H;��H;;�H;(�H;a�H;d�H;G�H;�I;QI;I;I;� I;,I;�9I;9II;n[I;�pI;5�I;�I;��I;ՁI;_<I;��H;��G;�F;IE;�C;֠@;��=;7;;��8;Z16;�U4;V%3;      W@@;Hp@;��@;��A;��B;5D;�EE;(gF;�dG;�2H;_�H;�8I;5yI;ؗI;ݜI;��I;U~I;viI;�VI;FI;�7I;�*I;> I;&I;]I;�I;@I;��H;��H;��H;�H;"�H;��H;o�H;��H;%�H;��H;�H;��H;r�H;��H;�H; �H;��H;��H;��H;;I;�I;aI;#I;< I;�*I;�7I;FI;�VI;siI;X~I;��I;ݜI;֗I;6yI;�8I;a�H;�2H;�dG;&gF;�EE;,D;��B;��A;��@;Hp@;      _fF;�yF;ֱF;8G;sG;A�G;�YH;o�H;NI;�WI;t�I;јI;��I;��I;ՅI;sI;�`I;;PI;�AI;�4I;)I;�I;�I;#I;�I;SI;��H;�H;��H;T�H;-�H;h�H;�H;-�H;t�H;�H;�H;�H;q�H;-�H;�H;c�H;0�H;U�H;��H;�H;��H;YI;�I;I;I;�I;)I;�4I;�AI;7PI;�`I;
sI;ՅI;��I;��I;ϘI;|�I;�WI;QI;n�H;�YH;6�G;sG;JG;ֱF;�yF;      J�H;��H;/�H;I;g%I;WHI;�hI;�I;D�I;��I;�I;��I;�I;�vI; fI;�VI;�HI;<I;�0I;/&I;I;4I;QI;ZI;;I;��H;�H;��H;j�H;2�H;l�H;��H;��H;�H;j�H;�H;�H;�H;h�H;	�H;��H;��H;o�H;2�H;f�H;��H;�H;��H;AI;VI;RI;8I;I;,&I;�0I;<I;�HI;�VI; fI;�vI;�I;��I;�I;��I;A�I;�I;�hI;QHI;|%I;�I;.�H;��H;      ��I; �I;׎I;=�I;��I;��I;.�I;"�I;U�I;��I;��I;tI;0fI;�XI;?LI;y@I;�5I;�+I;�"I;�I;�I;9I;�I;�I;��H;��H;��H;a�H;H�H;\�H;��H;��H;��H;��H;��H;B�H;'�H;>�H;��H; �H;��H;��H;��H;^�H;E�H;a�H;��H; �H;��H;�I;�I;<I;�I;�I;�"I;�+I;�5I;z@I;ALI;�XI;2fI;tI;��I; �I;U�I;"�I;.�I;��I;��I;C�I;׎I;��I;      Q�I;ޛI;��I;��I;ڔI;��I;��I;7�I;LvI;�kI;�`I;/VI;�KI;�AI;�7I;�.I;d&I;�I;�I;NI;�I;|I; I;J�H;��H;��H;b�H;H�H;b�H;��H;��H;��H;��H;&�H;��H;��H;R�H;�H;��H;'�H;��H;��H;��H;��H;_�H;H�H;b�H;��H;��H;G�H;"I;~I;�I;LI;�I;�I;d&I;�.I;�7I;�AI;�KI;/VI;�`I;�kI;PvI;8�I;��I;��I;�I;��I;��I;ٛI;      !|I;�{I;�yI;hvI;rI;�lI;)fI;#_I;�WI;�OI;�GI;g?I;R7I;�/I;�'I;� I;{I;nI;�I;�	I;QI;6I;��H;d�H;��H;M�H;2�H;a�H;��H;��H;��H;��H;��H;��H;�H;��H;��H;��H;�H;��H;��H;��H;��H;��H;��H;a�H;0�H;T�H;��H;c�H;��H;<I;MI;�	I;�I;nI;~I;� I;�'I;}/I;R7I;d?I;�GI;�OI;�WI;"_I;/fI;�lI;rI;svI;�yI;�{I;      �[I;d[I;�YI;UWI;TI;�OI;KI;�EI;0@I;):I;�3I;�-I;�'I;�!I;�I;\I;=I;WI;�I;�I;X I;�H;�H;`�H;�H;,�H;o�H;��H;��H;��H;~�H;��H;V�H;��H;x�H;\�H;U�H;Y�H;u�H;��H;Z�H;��H;��H;��H;��H;��H;m�H;2�H;#�H;`�H;�H;�H;V I;�I;�I;WI;@I;`I;�I;�!I;�'I;�-I;�3I;,:I;3@I;�EI;(KI;�OI;TI;WWI;�YI;d[I;      �CI;YCI;:BI;e@I;�=I;�:I;%7I;
3I;�.I;�)I;'%I;k I;�I;�I;wI;I;
I;/I;�I;A�H;S�H;��H;3�H;(�H;"�H;^�H;��H;��H;��H;��H;��H;D�H;��H;N�H;�H;��H;��H;��H;�H;Q�H;��H;B�H;��H;��H;��H;��H;��H;c�H;&�H;$�H;9�H;��H;O�H;=�H;�I;2I;
I;I;zI;�I;�I;h I;.%I;�)I;�.I;
3I;/7I;�:I;�=I;n@I;ABI;YCI;      2I;�1I;�0I;q/I;s-I;+I;C(I; %I;�!I;!I;wI;�I;�I;�I;PI;�I;�I;wI;��H;��H;b�H;�H;�H;9�H;��H;�H;��H;��H;��H;�H;S�H;��H;3�H;��H;��H;~�H;o�H;�H;��H;��H;5�H;��H;S�H;��H;��H;��H;��H;�H;��H;:�H;�H;�H;[�H;��H;��H;wI;�I;�I;SI;�I;�I;�I;{I;$I;�!I;%I;H(I;	+I;x-I;o/I;�0I;�1I;      �%I;S%I;�$I;�#I;"I; I;�I;LI;�I;�I;�I;eI;aI;\	I;OI;oI;� I;��H;e�H;?�H;D�H;?�H;j�H;��H;n�H;&�H;�H;�H;*�H;��H;��H;Q�H;��H;��H;^�H;8�H;&�H;8�H;\�H;��H;��H;R�H;��H;��H;&�H; �H;�H;*�H;o�H;��H;o�H;?�H;@�H;8�H;d�H;��H;� I;rI;RI;[	I;`I;dI;�I;�I;�I;II;�I; I;"I;�#I;�$I;_%I;      TI;9I;�I;�I;YI;�I;�I;�I;]I;�I;aI;�
I;I;oI;�I;T I;��H;��H;{�H;{�H;��H;��H;`�H;��H;��H;i�H;e�H;��H;��H;�H;q�H;�H;��H;\�H;�H;�H;�H;�H;�H;^�H;��H;�H;p�H;�H;��H;��H;f�H;k�H;��H;��H;d�H;��H;��H;t�H;z�H;��H;��H;X I;�I;mI;I;�
I;cI;�I;`I;�I;�I;�I;VI;�I;�I;;I;      �I;`I;�I;I;�I;vI;�I;�I;�I;�I;T
I;I;�I;*I;� I;��H;[�H;Q�H;e�H;��H;��H;�H;��H;Q�H;�H;�H;�H;B�H;��H;��H;X�H;��H;��H;9�H;	�H;��H;��H;��H;�H;=�H;��H;��H;V�H;��H;��H;?�H;�H;�H;�H;S�H;��H;�H;��H;{�H;d�H;T�H;^�H;��H;� I;-I;�I; I;X
I;�I;�I;�I;�I;wI;�I;I;�I;nI;      ;I;I;�I;�I;wI;(I;~I;�I;�I;{I;W	I;I;�I;�I;[ I;�H;��H;��H;��H;$�H;��H;��H;Q�H;��H;��H;	�H;�H;-�H;Y�H;��H;N�H;��H;p�H;!�H;�H;��H;��H;��H;�H;#�H;s�H;��H;N�H;��H;R�H;)�H;�H;�H;��H;��H;T�H;��H;��H; �H;��H;��H;��H;�H;] I;�I;�I;I;\	I;}I;�I;�I;�I;(I;vI;�I;�I;I;      �I;bI;�I;	I;�I;yI;�I;�I;�I;�I;R
I;I;�I;-I;� I;��H;[�H;Q�H;e�H;��H;��H;�H;��H;Q�H;�H;�H;�H;B�H;��H;��H;Y�H;��H;��H;9�H;�H;��H;��H;��H;�H;<�H;��H;��H;X�H;��H;��H;>�H;�H;	�H;�H;Q�H;��H;�H;��H;{�H;d�H;T�H;]�H;��H;� I;*I;�I; I;Y
I;�I;�I;�I;�I;wI;�I;I;�I;iI;      LI;<I;�I;�I;YI;�I;�I;�I;_I;�I;_I;�
I;I;oI;�I;V I;��H;��H;{�H;{�H;��H;��H;`�H;��H;��H;g�H;f�H;��H;��H;�H;q�H;�H;��H;_�H;�H;�H;�H;�H;�H;_�H;��H;�H;p�H;
�H;��H;��H;f�H;k�H;��H;��H;c�H;��H;��H;t�H;z�H;��H;��H;X I;�I;pI;I;�
I;eI;�I;_I;�I;�I;�I;YI;�I;�I;=I;      �%I;T%I;�$I;�#I;"I; I;�I;OI;�I;�I;�I;dI;`I;[	I;RI;qI;� I;��H;e�H;=�H;E�H;@�H;j�H;��H;r�H;(�H;	�H;�H;-�H;��H;��H;R�H;��H;��H;b�H;9�H;&�H;9�H;^�H;��H;��H;R�H;��H;��H;%�H;��H;�H;)�H;o�H;��H;n�H;=�H;=�H;9�H;e�H;��H;� I;tI;TI;\	I;`I;dI;�I;�I;�I;NI;�I; I;"I;�#I;�$I;U%I;      2I;�1I;�0I;n/I;q-I;+I;B(I;'%I;�!I;!I;wI;�I;�I;�I;SI;�I;�I;wI;��H;��H;b�H;�H;�H;:�H;��H;�H;��H;��H;��H;�H;S�H;��H;3�H;��H;��H;��H;q�H;��H;��H;��H;2�H;��H;R�H;��H;��H;��H;��H;�H;��H;6�H;�H;�H;X�H;��H;��H;vI;�I;�I;SI;�I;�I;�I;{I;"I;�!I;#%I;J(I;+I;v-I;u/I;�0I;�1I;      �CI;]CI;+BI;e@I;�=I;�:I;,7I;	3I;�.I;�)I;+%I;k I;�I;�I;zI;I;
I;2I;�I;@�H;V�H;��H;4�H;'�H;&�H;a�H;��H;��H;��H;��H;��H;D�H;��H;N�H;�H;��H;��H;��H;�H;O�H;��H;D�H;��H;��H;��H;��H;��H;a�H;"�H; �H;:�H;��H;M�H;=�H;�I;/I;
I;I;{I;�I;�I;k I;.%I;�)I;�.I;3I;,7I;�:I;�=I;p@I;2BI;WCI;      �[I;d[I;�YI;PWI;TI;�OI;!KI;�EI;0@I;):I;�3I;�-I;�'I;�!I;�I;_I;@I;XI;�I;�I;Z I;�H;�H;`�H;#�H;,�H;m�H;��H;��H;��H;��H;��H;Y�H;��H;|�H;\�H;V�H;_�H;u�H;��H;Z�H;��H;��H;��H;��H;��H;m�H;/�H;�H;]�H;�H;�H;S I;�I;�I;VI;BI;_I;�I;�!I;�'I;�-I;�3I;+:I;3@I;�EI;&KI;�OI;TI;ZWI;�YI;e[I;      ,|I;�{I;�yI;uvI;�qI;�lI;+fI;)_I;�WI;�OI;�GI;g?I;R7I;}/I;�'I;� I;|I;pI;�I;�	I;SI;;I;��H;c�H;��H;M�H;2�H;b�H;��H;��H;��H;��H;��H;��H;�H;��H;��H;��H;�H;��H;��H;��H;��H;��H;��H;a�H;0�H;Q�H;��H;`�H;��H;;I;MI;�	I;�I;lI;|I;� I;�'I;/I;S7I;d?I;�GI;�OI;�WI;&_I;/fI;�lI;rI;|vI;�yI;�{I;      ]�I;ߛI;��I;��I;ϔI;��I;��I;8�I;TvI;�kI;�`I;0VI;�KI;�AI;�7I;�.I;c&I;�I;�I;LI;�I;~I;I;J�H;��H;��H;b�H;I�H;c�H;��H;��H;��H;��H;'�H;��H;��H;S�H;��H;��H;&�H;��H;��H;��H;��H;_�H;G�H;c�H;��H;��H;D�H;$I;I;�I;LI;�I;�I;c&I;�.I;�7I;�AI;�KI;.VI;�`I;�kI;RvI;9�I;��I;��I;ޔI;��I;��I;כI;      ��I;��I;ˎI;@�I;��I;��I;/�I;)�I;T�I;��I;��I;tI;2fI;�XI;BLI;z@I;�5I;�+I;�"I;�I;�I;<I;�I;�I;��H;��H;��H;a�H;K�H;\�H;��H;��H;��H;��H;��H;?�H;,�H;B�H;��H; �H;��H;��H;��H;^�H;G�H;_�H;��H;��H;��H;�I;�I;;I;�I;�I;�"I;�+I;�5I;z@I;BLI;�XI;2fI;tI;��I; �I;S�I;"�I;/�I;��I;��I;C�I;֎I;��I;      <�H;��H;,�H;I;t%I;ZHI;�hI;�I;D�I;��I;�I;��I;�I;�vI;"fI;�VI;�HI;
<I;�0I;+&I;I;8I;OI;]I;>I;��H;�H;��H;j�H;2�H;m�H;��H;��H;�H;l�H;�H;�H;�H;h�H;	�H;��H;��H;p�H;3�H;f�H;��H;�H;��H;>I;VI;UI;6I;I;.&I;�0I;<I;�HI;�VI;"fI;�vI;�I;��I;�I;��I;A�I;�I;�hI;THI;{%I;I;.�H;��H;      VfF;�yF;ݱF;9G;	sG;K�G;�YH;s�H;RI;�WI;x�I;ҘI;��I;��I;ׅI;
sI;�`I;<PI;�AI;�4I;)I;�I;I;#I;�I;SI;��H;�H;��H;T�H;0�H;i�H;�H;-�H;u�H;�H;�H;�H;p�H;,�H;�H;h�H;3�H;U�H;��H;�H;��H;UI;�I;I;�I;�I;)I;�4I;�AI;8PI;�`I;sI;؅I;��I;��I;ϘI;{�I;�WI;KI;k�H;�YH;6�G;sG;<G;ñF;�yF;      T@@;Ep@;��@;��A;��B;;D;�EE;(gF;�dG;�2H;_�H;�8I;6yI;֗I;��I;��I;V~I;yiI;�VI;FI;�7I;�*I;< I;&I;cI;�I;;I;��H;��H;��H;�H;%�H;��H;p�H;��H;"�H;��H;"�H;��H;p�H;��H;#�H;!�H;��H;��H;��H;@I;�I;^I;"I;? I;�*I;�7I;FI;�VI;riI;Y~I;��I;�I;֗I;7yI;�8I;_�H;�2H;�dG;)gF;�EE;-D;��B;��A;��@;Gp@;      ��2;D%3;�U4;g16;��8;-7;;��=;Ӡ@;�C;IE;�F;��G;��H;a<I;فI;��I;�I;<�I;�pI;o[I;<II;�9I;,I;� I;!I;I;QI;�I;K�H;c�H;`�H;.�H;;�H;��H;��H;]�H;�H;`�H;��H;��H;=�H;-�H;c�H;d�H;G�H;�I;VI;I;I;� I;,I;�9I;;II;o[I;�pI;6�I;�I;��I;ցI;a<I;��H;��G;�F;IE;�C;͠@;��=; 7;;��8;{16;�U4;/%3;      Z�;ϻ;
;	�;��#;t);��.;�W4;.|9;@�=;1�A;�D;��F;rH;��H;_I;ƓI;X�I;P�I;�uI;r^I;�JI;%:I;#,I;> I;~I;NI;�I;%I;��H;�H;9�H;�H;m�H;d�H;��H;W�H;��H;`�H;j�H;�H;7�H;�H;��H;I;�I;TI;I;: I; ,I;%:I;�JI;r^I;�uI;Q�I;Q�I;ȓI;~_I;��H;pH;��F;ވD;4�A;>�=;)|9;�W4;��.;v);��#;�;
;��;      ���:m��:���:k
�:]+�:��;��;��;��&;T�/;D=7;[D=;��A;�E;G7G;b�H;n8I;�I;
�I;��I;xI;�_I;�JI;�9I;�*I;�I;5I;=I;�I;9I;�H;��H;�H;<�H;��H;�H;��H;�H;��H;;�H;�H;��H;�H;<I;I;<I;9I;�I;�*I;�9I;�JI;�_I;�wI;��I;
�I;�I;n8I;_�H;F7G;�E;��A;WD=;F=7;S�/;��&;��;��;��;�+�:U
�:���:W��:      0�x9���9���9p	:��^:� �:�ɼ:�P�:��;�h;ڣ#;�</;�;8;��>;�oC;�fF;>(H;NI;�I;ŜI;��I;�wI;n^I;;II;�7I;)I;I;�I;�I;GI;O I;L�H;T�H;=�H;��H;��H;��H;��H;��H;9�H;T�H;I�H;P I;JI;�I;�I;I;)I;�7I;;II;n^I;�wI;��I;ĜI;�I;JI;@(H;�fF;�oC;��>;�;8;�</;ۣ#;�h;��;�P�:�ɼ:� �:D�^:x	:��9@��9      ������J��:񳺠dt��F�`�8��&:0��:%��:�Z;KC;7�&;�'3;!<;��A;�E;p�G;AI;^|I;ȜI;��I;~uI;r[I;FI;�4I;(&I;�I;LI;�	I;�I;;�H;��H;8�H;t�H;z�H;�H;|�H;q�H;4�H;��H;:�H;�I;�	I;II;�I;.&I;�4I;FI;u[I;�uI;��I;ŜI;^|I;CI;n�G;�E;��A;<;�'3;5�&;HC;�Z;!��:&��:��&:@�8�F�xdt�P�L�ຨ���      N��;��b����g���7}�d�D����.x��(
�����9��:���:	;�;��.;��9;��@;�]E;m�G;CI;�I;	�I;M�I;�pI;�VI;�AI;z0I;�"I;�I;�I;�I;�I;��H;`�H;w�H;^�H;��H;^�H;t�H;]�H;��H;�I;�I;�I;�I;�"I;~0I;�AI;�VI;�pI;K�I;�I;�I;CI;m�G;�]E;��@;��9;��.;�;	;���:��:���90
��(x�����i�D��7}��g��f���8��      ��?��<<��1��h!��z��B�`���n����-�:��}��8�&:d��:4��:��;#�+;ۍ8;A�@;�]E;n�G;II;�I;S�I;8�I;riI;7PI;<I;�+I;�I;nI;TI;+I;sI;��H;��H;N�H;��H;Q�H;��H;��H;sI;+I;TI;oI;�I;�+I;<I;7PI;liI;8�I;Q�I;�I;FI;n�G;�]E;>�@;؍8;!�+;��;4��:d��:4�&:�}��@𳺃�-��n��`���B黴z��h!��1��<<�      b��R���I��{�������^��75��z���̻�눻�R�dt�P�x9B��:pm�:�h;c�*;ލ8;��@;�E;=(H;k8I;��I;�I;Q~I;�`I;�HI;�5I;_&I;rI;5I;�	I;�I;� I;��H;T�H;��H;T�H;��H;� I;�I;�	I;6I;tI;]&I;�5I;�HI;�`I;K~I;�I;��I;i8I;9(H;�E;��@;ۍ8;b�*;�h;lm�:D��:P�x9$dt��R��눻��̻�z��75��^����|����I��Q��      '��b��
����]��HC���t����|���?���	�$���V��������:��:�h;#�+;��9;��A;�fF;^�H;y_I;��I;��I;sI;�VI;s@I;�.I;� I;VI;I;�I;kI;O I;{�H;�H;|�H;J I;gI;�I;	I;VI;� I;�.I;u@I;�VI;�rI;��I;��I;x_I;[�H;zfF;��A;��9; �+;�h;��:��:@�����V�&����	���?���|��t��HC��^������
�b�      ��t��p�.�d� �Q�|�9�^*����a�ҼzI���o���'��ڻb6}�6���8���:fm�:��;��.;<;�oC;C7G;��H;ՁI;ٜI;҅I;fI;>LI;�7I;�'I;�I;tI;NI;JI;�I;� I;O I;� I;�I;HI;LI;qI;�I;�'I;�7I;?LI;fI;хI;՜I;ցI;��H;A7G;�oC;<;��.;��;hm�:��: 9�8��f6}��ڻ��'��o�zI��a�Ҽ���^*�}�9� �Q�.�d��p�      ��Ž4���̷�R���z����}��Q�T�'����'C��+\��,<<��>n��,��@�>��:4��:�;�'3;��>;�E;mH;d<I;ԗI;��I;�vI;�XI;�AI;v/I;�!I;�I;�I;Q	I;aI;!I;rI;#I;^I;S	I;�I;�I;�!I;y/I;�AI;�XI;�vI;��I;͗I;d<I;nH;�E;��>;�'3;�;6��:B��:@�8�ກn���>�-<<�+\��(C�����U�'��Q���}��z��R��̷�4���      c.��3�Ȥ�V����ΈŽ75�����YG�2��bkּG����xC��>�\6}����P�x9l��:	;6�&;�;8;��A;��F;��H;7yI;��I;�I;0fI;�KI;N7I;'I;�I;�I;ZI;I;�I;�I;�I;I;WI;�I;�I;}'I;O7I;�KI;1fI;�I;��I;0yI;��H;��F;��A;�;8;9�&;	;f��:P�x9���a6}��>��xC�H���bkּ2��YG����75��ΈŽ��V��Ȥ��3�      Hx��s���d�N�N�`�3�|I����H����z����\�B*�	�ݼH���,<<��ڻ�V�0dt�(�&:���:EC;�</;TD=;ڈD;��G;�8I;ȘI;��I;tI;(VI;Z?I;�-I;b I;�I;]I;�
I;�I;I;�I;�
I;ZI;�I;a I;�-I;\?I;,VI;tI;��I;ǘI;�8I;��G;ۈD;QD=;�</;FC;���:4�&:(dt��V��ڻ-<<�H���
�ݼC*���\��z��H������|I�`�3�N�N���d��s�      ,l¾(��T������������d���7�x��8Sؽ[���d�C*�bkּ+\����'�&���R�(~��~�:�Z;أ#;@=7;/�A;�F;[�H;q�I;�I;��I;�`I;�GI;�3I;'%I;tI;�I;TI;M
I;L	I;M
I;TI;�I;tI;$%I;�3I;�GI;�`I;��I;�I;o�I;W�H;�F;.�A;<=7;Σ#;�Z;|�:~���R�'����'�+\��bkּC*��d�[��8Sؽx����7��d���������T���(��      �V������������Ͼ�d���ǆ�D�N��3��c�[����\�2��(C���o���	��눻L����9!��:�h;T�/;=�=;JE;�2H;�WI;��I;��I;�kI;�OI;$:I;�)I;$I;�I;�I;�I;yI;�I;�I;�I;$I;�)I;":I;�OI;�kI;��I;��I;�WI;�2H;IE;>�=;R�/;�h;#��:���9L��눻��	��o�(C��2����\�[���c཰3�D�N��ǆ��d����Ͼ���������      �,b�ý\��>M���5�<��1r��%l¾青�"&W��3�8Sؽ�z��YG����zI����?���̻��-�`
�� ��:��;��&;|9;�C;�dG;KI;@�I;P�I;SvI;|WI;,@I;�.I;�!I;�I;UI;�I;�I;�I;VI;�I;�!I;�.I;)@I;{WI;RvI;Q�I;?�I;NI;�dG;�C;!|9;��&;��;"��:�
����-���̻��?�zI�����YG��z��8Sؽ�3�"&W�青�%l¾1r��<����5��>M�ý\�      ���$��Z���M䂿½\���1�����J˾青�D�N�x��H������U�'�b�Ҽ��|��z��n��8x����&:�P�:��;�W4;Ԡ@;(gF;`�H;�I;�I;1�I;_I;�EI;3I;!%I;DI;�I;�I;�I;�I;�I;DI;!%I;3I;�EI;!_I;1�I; �I;�I;e�H;%gF;Ӡ@;�W4;��;�P�:��&:Bx���n���z���|�c�ҼU�'����H���x��D�N�青��J˾�����1�½\�M䂿Z���$��      }߿�$ڿ.�ʿ����	����Ps�PX:����%l¾�ǆ���7����75���Q�����t���75�h�������8�ɼ:��;��.;��=;�EE;�YH;�hI;#�I;��I;)fI;KI;&7I;F(I;�I;�I;�I;wI;�I;�I;�I;H(I;&7I;KI;+fI;��I;&�I;�hI;�YH;�EE;��=;��.;��;�ɼ:��8���g���75��t������Q�75�������7��ǆ�%l¾���PX:��Ps�	�������.�ʿ�$ڿ      z�����p������ſ$���Ps���1�1r���d���d�|I�ΈŽ��}�_*�IC���^��B�u�D��F๚ �:��;r); 7;;)D;1�G;UHI;��I;��I;�lI;�OI;�:I;+I; I;�I;yI;/I;yI;�I; I;+I;�:I;�OI;�lI;��I;��I;THI;=�G;*D;!7;;p);��;� �:�F�w�D��B��^�IC��_*���}�ΈŽ|I��d��d��1r����1��Ps�$����ſ��꿃p����      ��7��3�ע%�z��<����ſ	���½\�<����Ͼ����`�3��轻z��|�9�^�Ἒ���z��7}�|dt�(�^:e+�:��#;��8;��B;	sG;o%I;��I;�I;	rI;TI;�=I;s-I;"I;HI;�I;}I;�I;KI;"I;s-I;�=I;TI;rI;�I;��I;r%I;sG;��B;��8;��#;g+�:�^:xdt��7}��z����^��|�9��z����`�3�������Ͼ<��½\�	�����ſ�<��z�ע%��3�      -�_��+Y��lG�f.�z���꿱���M䂿��5���󾍰��N�N�V��R�� �Q����|����h!��g��\񳺀	:]
�:��;]16;��A;8G;�I;8�I;x�I;lvI;NWI;l@I;m/I;�#I;�I;I;�I;
I;�I;�#I;o/I;o@I;KWI;rvI;x�I;9�I; I;CG;��A;_16;��;]
�:d	:Z񳺉g���h!�{������ �Q�R��V��N�N���������5�M䂿�������z�f.��lG��+Y�      Ѭ��#}�>tf��lG�ע%��p�.�ʿZ����>M����T�����d�Ȥ�̷�.�d��
��I���1�c���R��Ь�9���:;�U4;��@;ұF;2�H;ݎI;��I;�yI;�YI;<BI;�0I;�$I;�I;�I;�I;�I;�I;�$I;�0I;<BI;�YI;�yI;��I;��I;4�H;߱F;��@;�U4;;���:���9J��d����1��I���
�.�d�̷�Ȥ���d�T�������>M�Z���.�ʿ�p�ע%��lG�>tf�#}�      S���D���#}��+Y��3�����$ڿ%��ý\����(���s��3�5����p�b�S���<<�4���������9O��:һ;R%3;Ep@;�yF;��H;��I;�I;�{I;O[I;RCI;�1I;U%I;#I;ZI;I;WI;#I;U%I;�1I;SCI;K[I;�{I;�I;��I;��H;�yF;Gp@;Q%3;˻;I��:`��9����6���<<�S��b��p�5����3��s�(�����ý\�%���$ڿ����3��+Y�#}�D���      �Aq���i���U�F:�@�����<���v���{A�d5�� ��~^Z�����A���]�����d��H",��5����ѺP��9���: �;^Y4;H�@;JVF;��H;�GI;�bI;OI; :I;�)I;$I;�I;�I;�I;�I;�I;�I;�I;"I;�)I;:I;#OI;�bI;�GI;��H;ZVF;I�@;[Y4;�;���:(��9��Ѻ�5��H",��d������]��A�����~^Z�� ��d5�{A�v���<�������@�F:���U���i�      ��i���b�Z�O�.5�2i�������������q<�����e��`
V�GE	�!���IY�i9�C�����(��R����Ⱥh�:W��:�;A�4;>�@;hF;��H;II;ybI;�NI;�9I;�)I;�I;_I;�I;eI;`I;aI;�I;_I;�I;�)I;�9I;�NI;|bI;II;��H;(hF;?�@;?�4;ޔ;Q��:T�:��Ⱥ�R����(�C���i9��IY�!��GE	�`
V��e������q<������������2i�.5�Z�O���b�      ��U�Z�O�H-?�.�'���L�ῴ欿`�{�ea/���뾝���I����c���ZN�Z5������:H�` ��`�����":��:~�;��5;�`A;��F;K�H;MI;�aI;�MI;�8I;�(I;FI;�I;=I;I;I;I;>I;�I;FI;�(I;�8I;�MI;�aI;MI;N�H;��F;�`A;��5;v�;��:|�":X���b ��:H�����Z5���ZN�c������I�������ea/�`�{��欿L����.�'�H-?�Z�O�      F:�.5�.�'��������jȿ���k$_���W�Ҿە���6�����*���`=�<�漭)��GG�$6�����4�Q:��:�/";�7;^&B;��F;��H;�RI;�`I;yKI;7I;�'I;AI;I;�I;uI;t
I;oI;�I;I;AI;�'I;7I;KI;�`I;�RI;��H;��F;^&B;�7;�/";��:�Q:���$6��GG��)��<���`=��*������6�ە��W�Ҿ��k$_����jȿ�������.�'�.5�      @�2i�������I�ѿk��� ���q<��:��a����q����Wн潅���'�Tb̼�zl��.��F�X�T����:��;Ԏ&;ɫ9;$C;>MG;��H;8YI;�^I;�HI;�4I;�%I;�I;
I;�I;�
I;�	I;�
I;�I;
I;�I;�%I;�4I;�HI;�^I;<YI;��H;EMG;$C;ƫ9;ώ&;��;��:D��I�X��.���zl�Tb̼��'�潅��Wн����q��a���:��q<� ��k���I�ѿ������2i�      �������L��jȿk���������O���z]׾{����I�����A��=�d�m�}֮�RH��jλI�$��(�y��:JN;��+;�<;�3D;��G;�I;�^I;k[I;�DI;!2I;�#I;FI;�I;`I;�	I;�I;�	I;`I;�I;GI;�#I;!2I;�DI;n[I;�^I;�I;��G;�3D;�<;��+;JN;m��:`(�J�$��jλRH�}֮�m�=�d��A������I�{���z]׾����O�����k���jȿL�Ῡ��      <��������欿��� ����O��x����� ���l���"��ܽ���`=����u���k"�(R��2ۺ蓵9�?�:bL;��0;��>;�ME;M#H;�%I;�aI;�VI;�@I;�.I;?!I;AI;I;I;PI;�I;MI;I;I;@I;=!I;�.I;�@I; WI;�aI;�%I;Q#H;�ME;��>;��0;_L;�?�:�96ۺ(R���k"�v������`=����ܽ��"��l�� ����뾁x���O� ������欿����      v�������`�{�k$_��q<�������}��w��	�6�����!���h����෾�� d�y.���^e��H[���Z:h��:�, ;��5;�A;�VF;��H;�@I;pbI;�QI;�;I;=+I;nI;I;7I;	I;�I;/I;�I;�	I;:I;I;kI;;+I;�;I;�QI;vbI;�@I;��H;�VF;�A;��5;�, ;`��:��Z:�H[��^e�x.��� d�෾�����h�!������	�6�w���}��������q<�l$_�`�{�����      {A��q<�ea/����:�z]׾� ��w��>�CE	�����ڽ����3�]�꼘���
",��W��Y���
Q���:�M
;�f);��:;(@C;�?G;S�H;LTI;�_I;'KI;�6I;N'I;hI;�I;<I;�I;qI;�I;oI;�I;>I;�I;hI;O'I;�6I;*KI;�_I;HTI;S�H;�?G;(@C;��:;�f);�M
;���:�	Q�\���W��	",�����]�꼘�3�ڽ������DE	�>�w��� ��z]׾�:���ea/��q<�      d5�������W�Ҿ�a��{����l�	�6�DE	���Ƚk���aG����d֮��W����f�k� ���c,:���:�;��1;B�>;AE;#�G;I;*_I;AZI;6DI;�1I;0#I;CI;�I;
I;	I;�I;!I;�I;	I;
I;�I;BI;2#I;�1I;9DI;GZI;'_I;I;'�G;@E;E�>;��1;��;���:�c,:$��c�k�����W�d֮�����aG�k����ȽDE	�	�6��l�{����a��W�Ҿ������      � ���e�����ܕ����q��I���"���������k���ZN�[� ¼N�y��$��Q���� � HX���:0;*�&;�w8;o B;��F;ԐH;W@I;�aI;jRI;=I;,I;�I;�I;[I;�I;5I;I;cI;I;5I;�I;\I;�I;�I;,I;=I;pRI;�aI;V@I;ڐH;��F;s B;�w8;'�&;)0;��: LX��� ��Q���$�L�y� ¼Z��ZN�k������������"��I���q�ە������e��      ~^Z�`
V��I��6�������ܽ!��ڽ���aG�Z�	�ȼ�)��z�(�d��CG5������Z:'�:S;'1;��=;��D;1�G;��H;�XI;^I;II;�5I;�&I;�I;�I;�
I;�I;KI;` I;��H;` I;KI;�I;�
I;~I;�I;�&I;�5I;�II;^I;�XI;��H;1�G;��D;��=;'1;S;-�:��Z:���AG5�c��y�(��)���ȼZ��aG�ٽ��!���ܽ������6��I�`
V�      ���GE	��������Wн�A�����h���3���� ¼�)��0x/��һk�X�b#����9\��:�>;2f);j`9;a&B;��F;i}H;�6I;PaI;�UI;a@I;�.I;� I;GI;'I;�I;LI;P I;��H;��H;��H;O I;LI;�I;$I;KI;!I;�.I;d@I;�UI;OaI;�6I;j}H;��F;e&B;i`9;<f);�>;T��:��9\#��i�X�
�һ/x/��)�� ¼�����3��h��󑽡A���Wн��콺��FE	�      �A��!��c���*��潅�>�d��`=����]��d֮�L�y�{�(��һ�]e�ބ���f9���:>�;K1";�4;�m?;�E;��G;g�H;�WI;�^I;KI;r7I;�'I;�I;"I;�
I;#I;I;k�H;��H;:�H;��H;j�H;I; I;�
I;(I;�I;�'I;u7I;KI;}^I;�WI;h�H;��G;�E;�m?;$�4;N1";<�;���:�f9ք���]e��һz�(�K�y�c֮�\�꼖���`=�=�d�潅��*��c��!��      �]��IY��ZN��`=���'�m����߷�������W��$�f��n�X�℮��9���:g��:v�;��0;��<;U�C;#G;��H;�?I;&aI;�TI;?@I;/I;W!I;�I;I;xI;�I;��H;|�H;�H;��H;�H;z�H;��H;�I;uI;I;�I;Z!I;/I;B@I;�TI;-aI;�?I;��H;)G;W�C;��<;��0;p�;m��:���:�9ք��k�X�b���$��W�����߷�����l���'��`=��ZN��IY�      ���i9�Z5��:��Sb̼}֮�t��� d�	",�����Q��HG5�j#���f9���:��:�;��-;��:;�KB;<VF;KH;�I;�\I;\I;�HI;6I;'I;I;�I;
I;BI;��H;��H;��H;X�H;��H;W�H;��H;��H;��H;?I;
I;�I;I;"'I;	6I;�HI;$\I;�\I;�I;KH;BVF;�KB;��:;��-;�;��:���:�f9h#��AG5��Q�����	",�� d�u��|֮�Tb̼;��Z5��h9�      �d��B��������)���zl�RH��k"�t.���W��_�k�~� ������9���:s��:�;�-;ѫ9;HaA;��E;)�G;x�H;�RI;`I;�OI;�<I;�,I;�I;/I;I;zI;TI;��H;��H;��H;��H;`�H;��H;��H;��H;��H;TI;~I;I;/I;�I;�,I;�<I;�OI;`I;SI;}�H;,�G;��E;KaA;ͫ9;�-;�;u��:���:��9���{� �^�k��W��t.���k"�
RH��zl��)������@���      @",���(�9H�CG��.���jλ"R���^e�Y���� HX���Z:N��::�;t�;��-;ȫ9;|A;�cE; �G;��H;RGI;�`I;�UI;9BI;�1I;�#I;�I;�I;�I;�I;��H;H�H;��H;
�H;�H;��H;�H;�H;��H;G�H;�H;�I;�I;�I;�I;�#I;�1I;ABI;�UI;�`I;XGI;��H;'�G;�cE;{A;ϫ9;��-;t�;:�;P��:��Z: $X���O���^e�$R���jλ�.��DG�7H���(�      �5���R��` ��!6��I�X�8�$�"ۺ�H[��Q��c,:��:'�:�>;K1";��0;��:;HaA;�cE;��G;v�H;�=I;.`I;qYI;�FI;�5I;�'I;�I;�I;�
I;�I;��H;�H;�H;��H;�H;��H;<�H;��H;}�H;��H;�H;�H;��H;�I;�
I;�I;�I;�'I;�5I;�FI;qYI;2`I;�=I;|�H;��G;�cE;NaA;��:;��0;M1";�>;-�:��:�c,:�Q��H[�"ۺ>�$�F�X�&6��` ���R��      ��Ѻ��ȺB������L�� (�H��9��Z:���:���:,0;S;7f);�4;��<;�KB;��E;(�G;y�H;b:I;R_I;�[I;#JI;9I;�*I;�I;�I; I;]I;I;��H;��H;�H;/�H;��H;7�H;��H;3�H;��H;/�H;�H;��H;��H;I;]I;I;�I;�I;�*I;9I;%JI;�[I;X_I;c:I;}�H;%�G;��E;�KB;��<; �4;9f);S;,0;���:���:��Z:0��9�'�8�����X����Ⱥ      P��9,�:8�":�Q:��:w��:�?�:h��:�M
;�;(�&;'1;i`9;�m?;U�C;BVF;)�G;��H;�=I;R_I;\I;�KI;;I;�,I;� I;�I;�I;�I;JI;��H;6�H;x�H;5�H;��H;��H;��H;��H;��H;��H;��H;4�H;t�H;9�H;��H;HI;�I;�I;�I;� I;�,I;;I;�KI;\I;S_I;�=I;��H;,�G;DVF;X�C;�m?;j`9;'1;,�&;�;�M
;b��:�?�:k��:��:�Q:d�":@�:      ���:{��:��:��:��;NN;_L;�, ;�f);��1;�w8;��=;b&B;�E;)G;KH;}�H;YGI;3`I;�[I;�KI;�;I;�-I;3"I;0I;I;	I;dI;��H;��H;��H;l�H;y�H;�H;G�H;��H;g�H;��H;D�H;�H;y�H;h�H;��H;��H;��H;gI;	I;I;5I;3"I;�-I;�;I;�KI;�[I;5`I;VGI;�H;KH;)G;�E;d&B;��=;�w8;��1;�f);�, ;fL;FN;��;��:��:i��:      7�;�;x�;�/";ǎ&;��+;��0;��5;��:;I�>;| B;��D;��F;��G; �H;�I;SI;�`I;qYI;$JI;;I;�-I;�"I;I;�I;�	I;*I;I�H;r�H;Z�H;��H;��H;��H;��H;��H;��H;c�H;��H;��H;��H;��H;��H;��H;Z�H;n�H;O�H;,I;�	I;�I;I;�"I;�-I;;I;%JI;uYI;�`I;SI;�I; �H;��G;��F;��D;� B;E�>;��:;��5;��0;��+;֎&;�/";w�;є;      ^Y4;K�4;��5;	�7;��9;�<;��>;�A;!@C;AE;��F;1�G;g}H;k�H;�?I;�\I;`I;�UI;�FI;9I;�,I;+"I; I;&I;[
I;�I;��H;��H;��H;��H;��H;��H;��H;��H;��H;��H;i�H;��H;��H;��H;��H;��H;��H;��H;��H;��H;��H;�I;b
I;&I;�I;0"I;�,I;9I;�FI;�UI;`I;�\I;�?I;j�H;g}H;5�G;��F;@E;'@C;�A;��>;�<;ɫ9;�7;��5;A�4;      i�@;B�@;�`A;X&B;C;4D;�ME;�VF;�?G;)�G;ސH;��H;�6I;�WI;.aI;+\I;�OI;HBI;�5I;�*I;� I;4I;�I;f
I;�I; I;0�H;��H;$�H;��H;��H;��H;N�H;|�H;��H;��H;h�H;��H;��H;|�H;I�H;��H;�H;��H; �H;��H;.�H; I;�I;f
I;�I;:I;� I;�*I;�5I;EBI;�OI;0\I;1aI;�WI;�6I;��H;ސH;)�G;�?G;�VF;�ME;�3D;*C;^&B;�`A;A�@;      LVF;/hF;��F;��F;2MG;��G;Q#H;��H;R�H;!I;[@I;�XI;UaI;�^I;�TI;�HI;�<I;�1I;�'I;�I;�I;I;�	I;�I; I;>�H;�H;[�H;��H;��H;z�H;K�H;@�H;{�H;	�H;��H;~�H;��H;�H;{�H;?�H;G�H;z�H;��H;��H;[�H;�H;E�H; I;�I;�	I;I;�I;�I;�'I;�1I;�<I;�HI;�TI;�^I;UaI;�XI;d@I;!I;T�H;��H;R#H;��G;JMG;��F;��F;-hF;      ��H;��H;H�H;��H;��H;�I;�%I;�@I;JTI;)_I;�aI;^I;�UI;KI;A@I;	6I;�,I;�#I;�I;�I;�I;	I;-I;��H;,�H;�H;H�H;�H;.�H;p�H;)�H;�H;8�H;��H;:�H;��H;��H;��H;7�H;��H;9�H;�H;*�H;p�H;+�H;�H;G�H;�H;4�H;��H;0I;	I;�I;�I;�I;�#I;�,I;6I;A@I;
KI;�UI;!^I;�aI;'_I;JTI;�@I;�%I;�I;��H;��H;H�H;��H;      �GI;II;MI;�RI;+YI;�^I;�aI;rbI;�_I;GZI;qRI;�II;b@I;y7I;/I;!'I;�I;�I;�I;I;�I;aI;E�H;��H;��H;R�H;�H;�H;|�H;)�H;�H;�H;e�H;��H;v�H;B�H;7�H;>�H;u�H;��H;g�H;	�H;�H;(�H;|�H;	�H;�H;[�H;��H;��H;H�H;dI;�I; I;�I;�I;�I;%'I;/I;y7I;a@I;�II;wRI;KZI;�_I;rbI;�aI;z^I;9YI;�RI;MI;II;      �bI;ubI;�aI;�`I;�^I;n[I;WI;�QI;#KI;9DI;=I;�5I;�.I;�'I;[!I;I;8I;�I;�
I;cI;QI;��H;m�H;��H;�H;��H;'�H;}�H;!�H;��H;��H;;�H;��H;,�H;��H;��H;��H;��H;��H;-�H;��H;8�H;��H;��H;�H;}�H;'�H;��H;!�H;��H;q�H;��H;OI;_I;�
I;�I;9I;I;^!I;�'I;�.I;�5I;=I;:DI;'KI;�QI;WI;e[I;�^I;�`I;�aI;qbI;      OI;�NI;�MI;sKI;�HI;�DI;�@I;�;I;�6I;�1I;,I;�&I;!I;�I;�I;�I;I;�I;�I;I;��H;��H;V�H;��H;��H;��H;n�H;*�H;�H; �H;&�H;�H;��H;��H;D�H;!�H;�H;�H;C�H;��H;��H;}�H;&�H;��H;��H;)�H;l�H;��H;��H;��H;[�H;��H;��H;I;�I;�I;I;�I;�I;�I;!I;�&I;,I;�1I;�6I;�;I;�@I;�DI;�HI;|KI;�MI;�NI;      :I;�9I;�8I;&7I;�4I;$2I;�.I;H+I;S'I;9#I;�I;�I;OI;/I;I;!
I;�I;�I;��H;��H;A�H;��H;��H;��H;��H;w�H;)�H;�H;��H;,�H;��H;��H;\�H;�H;��H;��H;��H;��H;��H;�H;_�H;��H;��H;)�H;��H;�H;(�H;}�H;�H;��H;��H;��H;?�H;��H;��H;�I;�I;%
I;I;.I;RI;�I;�I;;#I;W'I;E+I;�.I;2I;�4I;)7I;�8I;�9I;      �)I;�)I;�(I;�'I;�%I;�#I;?!I;tI;nI;HI;�I;�I;)I;�
I;|I;II;^I;��H;�H;��H;��H;l�H;��H;��H;��H;B�H;�H;�H;<�H;��H;��H;w�H;��H;��H;w�H;N�H;9�H;N�H;s�H;��H;��H;w�H;��H;�H;8�H;�H;�H;H�H;��H;��H;��H;o�H;}�H;��H;�H;��H;_I;LI;}I;�
I;+I;�I;�I;JI;mI;rI;I!I;�#I;�%I;�'I;�(I;�)I;      (I;�I;PI;CI;�I;=I;@I;I;�I;�I;aI;�
I;�I;(I;�I; I;��H;N�H;&�H;�H;B�H;}�H;��H;��H;L�H;<�H;9�H;l�H;��H;��H;Y�H;��H;��H;U�H;�H;�H;�H;�H;�H;X�H;��H;��H;Y�H;��H;��H;i�H;9�H;=�H;O�H;��H;��H;}�H;?�H;�H;&�H;O�H;��H; I;�I;(I;�I;�
I;bI;�I;�I;I;DI;8I;�I;AI;WI;�I;      xI;\I;�I;I;I;�I;I;?I;?I;
I;�I;�I;WI;&I;��H;��H;��H;��H;��H;6�H;��H;�H;��H;��H;x�H;t�H;��H;��H;/�H;��H;	�H;��H;X�H;�H;��H;��H;��H;��H;��H;�H;Z�H;��H;	�H;��H;)�H;��H;��H;x�H;z�H;��H;��H;�H;��H;1�H;��H;��H;��H;��H;��H;$I;UI;�I;�I;
I;BI;<I;I;�I;I;I;�I;hI;      �I;�I;DI;�I;�I;ZI;I;�	I;�I;I;BI;\I;^ I;z�H;��H;��H;��H;�H;��H;��H;��H;D�H;��H;��H;��H; �H;4�H;u�H;��H;G�H;��H;x�H;�H;��H;��H;��H;��H;��H;��H;��H;�H;z�H;��H;A�H;��H;r�H;5�H;�H;��H;��H;��H;C�H;��H;��H;��H;�H;��H;��H;��H;x�H;^ I;YI;EI;I;�I;�	I;I;[I;�I;�I;BI;�I;      �I;hI;
I;uI;�
I;�	I;WI;�I;pI;�I;'I;i I;��H;��H;�H;[�H;��H;�H;��H;:�H;��H;��H;��H;{�H;��H;��H;��H;A�H;��H;%�H;��H;S�H;�H;��H;��H;}�H;|�H;��H;��H;��H;	�H;S�H;��H; �H;��H;>�H;��H;��H;��H;{�H;��H;��H;��H;4�H;��H;�H;��H;_�H;�H;��H;��H;h I;)I;�I;sI;�I;aI;�	I;�
I;rI;I;vI;      �I;\I;"I;w
I;�	I;�I;�I;6I;�I;#I;qI;��H;�H;F�H;��H;��H;n�H;��H;C�H;��H;��H;i�H;`�H;`�H;f�H;u�H;��H;:�H;��H;%�H;��H;;�H;�H;��H;��H;w�H;��H;w�H;��H;��H;�H;=�H;��H;�H;��H;6�H;��H;y�H;e�H;_�H;c�H;g�H;��H;��H;C�H;��H;n�H;��H;��H;F�H;�H;��H;vI;%I;�I;6I;�I;�I;�	I;z
I;!I;hI;      �I;iI;I;rI;�
I;�	I;VI;�I;pI;�I;%I;k I;��H;��H;�H;[�H;��H;�H;��H;;�H;��H;��H;��H;{�H;��H;��H;��H;A�H;��H;$�H;��H;S�H;	�H;��H;��H;}�H;|�H;��H;��H;��H;	�H;S�H;��H;�H;��H;=�H;��H;��H;��H;z�H;��H;��H;��H;4�H;��H;�H;��H;^�H;�H;��H;��H;h I;+I;�I;sI;�I;]I;�	I;�
I;vI;
I;pI;      �I;�I;>I;�I;�I;WI;I;�	I;�I;I;AI;\I;^ I;z�H;��H;��H;��H;�H;��H;��H;��H;F�H;��H;��H;��H;��H;4�H;u�H;��H;F�H;��H;x�H;�H;��H;��H;��H;��H;��H;��H;��H;�H;x�H;��H;@�H;��H;q�H;5�H;�H;��H;��H;��H;D�H;��H;��H;��H;�H;��H;��H;��H;z�H;` I;\I;FI;I;�I;�	I;I;WI;�I;�I;DI;�I;      xI;^I;�I;I;I;�I;I;AI;BI;
I;�I;�I;VI;&I;��H;��H;��H;��H;��H;6�H;��H;!�H;��H;��H;{�H;v�H;��H;��H;0�H;��H;�H;��H;X�H;�H;��H;��H;��H;��H;��H;�H;Z�H;��H;�H;��H;)�H;��H;��H;x�H;x�H;��H;��H;�H;��H;2�H;��H;��H;��H;��H;��H;&I;VI;�I;�I;
I;BI;@I;I;�I;I;I;�I;_I;      %I;�I;SI;BI;�I;@I;>I;I;�I;�I;_I;�
I;�I;(I;�I; I;��H;N�H;$�H;�H;D�H;�H;��H;��H;P�H;9�H;9�H;l�H;��H;��H;X�H;��H;��H;U�H;�H;�H;�H;�H;�H;W�H;��H;��H;Y�H;��H;��H;h�H;9�H;<�H;L�H;��H;��H;{�H;;�H;�H;$�H;L�H;��H; I;�I;*I;�I;�
I;cI;�I;�I;I;EI;<I;�I;HI;[I;�I;      �)I;�)I;�(I;�'I;�%I;�#I;F!I;pI;kI;HI;�I;�I;+I;�
I;I;II;^I;��H;�H;��H;��H;o�H;��H;��H;��H;D�H;�H;�H;?�H;�H;��H;w�H;��H;��H;z�H;J�H;9�H;N�H;s�H;��H;��H;w�H;��H;}�H;8�H;�H;�H;E�H;��H;��H;��H;o�H;|�H;��H;�H;��H;_I;LI;I;�
I;.I;�I;�I;JI;mI;pI;G!I;�#I;�%I;�'I;�(I;�)I;      :I;�9I;�8I;#7I;�4I;"2I;�.I;K+I;S'I;9#I;�I;�I;RI;/I;I;$
I;�I;�I;��H;��H;C�H;��H;��H;��H;�H;v�H;(�H;�H;��H;*�H;��H;��H;]�H;�H;��H;��H;��H;��H;��H;�H;_�H;��H;��H;'�H;��H;�H;)�H;z�H;��H;��H;��H;��H;<�H;��H;��H;�I;�I;"
I;I;0I;RI;�I;�I;7#I;U'I;I+I;�.I; 2I;�4I;-7I;�8I;�9I;      )OI;�NI;�MI;�KI;HI;�DI;�@I;�;I;�6I;�1I;,I;�&I;!I;�I;�I;�I;I;�I;�I;I;��H;��H;W�H;��H;��H;��H;n�H;*�H;�H;�H;&�H;��H;��H;��H;F�H; �H;�H;!�H;C�H;��H;��H;��H;&�H;��H;��H;(�H;n�H;��H;��H;��H;]�H;��H;��H;I;�I;�I;I;�I;�I;�I;!I;�&I;,I;�1I;�6I;�;I;�@I;�DI;�HI;�KI;�MI;�NI;      �bI;sbI;�aI;�`I;�^I;s[I;WI;�QI;-KI;7DI;=I;�5I;�.I;�'I;^!I;I;6I;�I;�
I;bI;TI;��H;n�H;��H;"�H;��H;'�H;~�H;%�H;��H;��H;<�H;��H;,�H;��H;��H;��H;��H;��H;,�H;��H;<�H;��H;��H;�H;z�H;'�H;��H;�H;��H;r�H;��H;NI;_I; I;�I;6I;I;^!I;�'I;�.I;�5I;=I;7DI;'KI;�QI;WI;k[I;�^I;�`I;�aI;lbI;      �GI;II;MI;�RI;*YI;�^I;�aI;zbI;�_I;HZI;qRI;�II;a@I;x7I;/I;#'I;�I;�I;�I;I;�I;eI;G�H;��H;��H;T�H;�H;	�H;��H;(�H;�H;�H;e�H;��H;x�H;>�H;7�H;A�H;t�H;��H;h�H;�H;�H;(�H;z�H;�H;�H;V�H;��H;��H;K�H;cI;�I; I;�I;�I;�I;%'I;/I;v7I;a@I;�II;tRI;KZI;�_I;sbI;�aI;�^I;8YI;�RI;MI;II;      ��H;ėH;G�H;��H;��H;�I;�%I;�@I;LTI;)_I;�aI;#^I;�UI;
KI;B@I;6I;�,I;�#I;�I;�I;�I;	I;*I;��H;3�H;�H;H�H;�H;0�H;p�H;(�H;�H;8�H;��H;;�H;��H;��H;��H;7�H;��H;9�H;�H;*�H;p�H;+�H;�H;J�H;�H;0�H;��H;1I;	I;�I;�I;�I;�#I;�,I;6I;B@I;
KI;�UI;^I;�aI;'_I;JTI;�@I;�%I;�I;��H;��H;H�H;��H;      BVF;+hF;��F;��F;9MG;��G;P#H;��H;T�H; I;^@I;�XI;WaI;�^I;�TI;�HI;�<I;�1I;�'I;�I;�I;I;�	I;�I; I;?�H;�H;_�H;��H;��H;y�H;K�H;=�H;{�H;�H;��H;��H;��H;�H;{�H;@�H;L�H;}�H;��H;��H;[�H;�H;A�H; I;�I;�	I;I;�I;�I;�'I;�1I;�<I;�HI;�TI;�^I;VaI;�XI;a@I; I;M�H;��H;P#H;��G;CMG;��F;��F;hF;      f�@;<�@;�`A;^&B;C;4D;�ME;�VF;�?G;*�G;ސH;��H;�6I;�WI;4aI;0\I;�OI;IBI;�5I;�*I;� I;;I;�I;g
I;�I; I;1�H;��H;%�H;��H;��H;��H;I�H;{�H;��H;��H;i�H;��H;��H;~�H;L�H;��H;�H;��H;!�H;��H;0�H; I;�I;b
I;�I;8I;� I;�*I;�5I;CBI;�OI;0\I;3aI;�WI;�6I;��H;ސH;*�G;�?G;�VF;�ME;�3D;&C;^&B;�`A;>�@;      ;Y4;3�4;��5;�7;��9;�<;��>;�A;+@C;@E;��F;3�G;g}H;h�H;�?I;�\I;`I;�UI;�FI;9I;�,I;/"I;�I;(I;b
I;�I;��H;��H;��H;��H;��H;��H;��H;��H;��H;��H;k�H;��H;��H;��H;��H;��H;��H;��H;��H;��H;��H;�I;\
I;$I; I;."I;�,I;9I;�FI;�UI;`I;�\I;�?I;h�H;g}H;2�G;��F;AE;$@C;�A;��>;�<;ͫ9;)�7;��5;�4;      %�;ޔ;j�;�/";Ď&;��+;��0;��5;��:;K�>;y B;��D;��F;��G;�H;�I;SI; aI;tYI;'JI;;I;�-I;�"I;I;�I;�	I;*I;N�H;r�H;V�H;��H;��H;��H;��H;��H;��H;e�H;��H;��H;��H;��H;��H;��H;[�H;n�H;K�H;.I;�	I;�I; I;�"I;�-I;;I;'JI;wYI;�`I;SI;�I;�H;��G;��F;��D;{ B;H�>;��:;��5;��0;��+;Ǝ&;�/";l�;ʔ;      ���:y��:��:��:��;TN;fL;�, ;�f);��1;�w8;��=;e&B;�E;-G; KH;�H;[GI;3`I;�[I;�KI;�;I;�-I;3"I;7I;I;	I;gI;��H;��H;��H;m�H;y�H;�H;F�H;��H;h�H;��H;B�H;�H;y�H;l�H;��H;��H;��H;dI;	I;I;1I;3"I;�-I;�;I;�KI;�[I;5`I;UGI;}�H;KH;)G;�E;e&B;��=;�w8;��1;�f);�, ;bL;<N;��;��:��:e��:      ��9��:h�":4�Q:��:��:�?�:l��:�M
;��;+�&;'1;i`9;�m?;[�C;FVF;-�G;��H;�=I;U_I;\I;�KI;;I;�,I;� I;�I;�I;�I;JI;��H;6�H;{�H;5�H;��H;��H;��H;��H;��H;��H;��H;5�H;x�H;7�H;��H;GI;�I;�I;�I;� I;�,I;;I;�KI;\I;U_I;�=I;��H;,�G;DVF;[�C;�m?;j`9;'1;.�&;�;�M
;n��:�?�:w��:��:0�Q:��":@�:      |�Ѻ��ȺP������T���'�0��9�Z:���:���:-0;S;9f);�4;��<;�KB;��E;(�G;z�H;e:I;X_I;�[I;#JI;9I;�*I;�I;�I; I;_I;I;��H;��H;�H;2�H;��H;3�H;��H;6�H;��H;-�H;�H;��H;��H;I;]I; I;�I;�I;�*I;9I;$JI;�[I;V_I;c:I;|�H;$�G;��E;�KB;��<;�4;7f);S;,0;���:���:��Z:��90(�0�����R����Ⱥ      �5���R��a �� 6��M�X�:�$�"ۺ�H[��Q��c,:��:/�:�>;J1";��0;��:;KaA;�cE;��G;|�H;�=I;3`I;rYI;�FI;�5I;�'I;�I;�I;�
I;�I;��H;�H;�H;��H;}�H;��H;;�H;��H;z�H;��H;�H;�H;��H;�I;�
I;�I;�I;�'I;�5I;�FI;rYI;/`I;�=I;|�H;��G;�cE;IaA;��:;��0;K1";�>;)�:��:�c,: 	Q��H[�$ۺ<�$�K�X� 6��d ���R��      E",���(�;H�CG��.���jλ"R��~^e�R���� 8X���Z:P��::�;w�;��-;ͫ9;{A;�cE;%�G;��H;VGI;�`I;�UI;ABI;�1I;�#I;�I;�I;�I;�I;��H;G�H;��H;	�H;�H;��H;�H;�H;��H;G�H;��H;�I;�I;�I;�I;�#I;�1I;;BI;�UI;�`I;UGI;��H;'�G;�cE;zA;ʫ9;��-;v�;8�;L��:��Z: 8X���U���^e�"R���jλ�.��DG�=H���(�      �d��B��������)���zl�
RH��k"�s.���W��^�k�}� ������9���:{��:�;�-;Ы9;IaA;��E;-�G;|�H;SI;`I;�OI;�<I;�,I;�I;1I;I;|I;TI;��H;��H;��H;��H;a�H;��H;��H;��H;��H;SI;|I;I;1I;�I;�,I;�<I;�OI;`I;SI;y�H;(�G;��E;HaA;̫9;�-;�;u��:���:��9���~� �`�k��W��t.���k"�
RH��zl��)������A���      ���h9�Z5��:��Sb̼|֮�t��� d�",�����Q��AG5�j#���f9���:��:�;��-;��:;�KB;DVF;KH;�I;�\I;$\I;�HI;6I;'I;I;�I;
I;BI;��H;��H;��H;W�H;��H;W�H;��H;��H;��H;AI;
I;�I;I;'I;6I;�HI;\I;�\I;�I;KH;<VF;�KB;��:;��-;�;��:���:дf9j#��GG5��Q�����	",�� d�u��|֮�Tb̼:��[5��i9�      �]��IY��ZN��`=���'�l����߷�������W��$�b��k�X�܄���9���:m��:s�;��0;��<;[�C;'G; �H;�?I;,aI;�TI;<@I;/I;X!I;�I;I;yI;�I;��H;|�H;�H;��H;�H;y�H;��H;�I;vI;I;�I;[!I;/I;<@I;�TI;'aI;�?I;��H;&G;R�C;��<;��0;p�;q��:���:`9؄��o�X�d���$��W�����߷�����l���'��`=��ZN��IY�      �A��!��c���*��潅�=�d��`=����\��c֮�L�y�y�(��һ�]e�Є�� �f9���::�;K1"; �4;�m?;�E;��G;k�H;�WI;�^I;
KI;q7I;�'I;�I;(I;�
I; I;I;k�H;��H;:�H;��H;i�H;I; I;�
I;%I;�I;�'I;r7I;
KI;~^I;�WI;k�H;��G;�E;�m?;!�4;H1";:�;���:дf9܄���]e��һz�(�L�y�d֮�\�꼖���`=�=�d�潅��*��c��!��      ���FE	��������Wн�A�����h���3����¼�)��.x/��һe�X�\#����9V��:�>;9f);n`9;d&B;��F;k}H;�6I;PaI;�UI;a@I;�.I;� I;JI;(I;�I;OI;P I;��H;��H;��H;O I;LI;�I;%I;HI; !I;�.I;`@I;�UI;OaI;�6I;i}H;��F;b&B;f`9;:f);�>;P��:��9`#��i�X��һ0x/��)�� ¼�����3��h��󑽡A���Wн��콺��FE	�      ~^Z�`
V��I��6�������ܽ!��ڽ���aG�Z��ȼ�)��z�(�a��AG5������Z:)�:S;'1;��=;��D;3�G;��H;�XI;^I;~II;�5I;�&I;�I;I;�
I;�I;KI;^ I;��H;` I;JI;�I;�
I;I;�I;�&I;�5I;~II;^I;�XI;��H;2�G;��D;��=;'1;S;%�:��Z:���DG5�c��z�(��)��	�ȼZ��aG�ڽ��!���ܽ������6��I�`
V�      � ���e�����ە����q��I���"���������k���ZN�Z� ¼M�y��$��Q���� � LX���:%0;/�&;�w8;u B;��F;ڐH;Y@I;�aI;oRI;=I;,I;�I;�I;[I;�I;3I;I;cI;I;3I;�I;[I;�I;�I;,I;=I;oRI;�aI;V@I;ԐH;��F;v B;�w8;#�&;%0;��: LX��� ��Q���$�M�y� ¼Z��ZN�k������������"��I���q�ە������e��      d5�������W�Ҿ�a��{����l�	�6�DE	���Ƚk���aG����d֮��W����e�k�&���c,:���:�;��1;D�>;CE;'�G;I;&_I;CZI;7DI;�1I;3#I;CI;�I;
I;I;�I;I;�I;I;
I;�I;BI;2#I;�1I;7DI;CZI;$_I;I;%�G;CE;H�>;��1;��;���:�c,:$��c�k�����W�d֮�����aG�k����ȽDE	�	�6��l�{����a��W�Ҿ������      {A��q<�ea/����:�z]׾� ��w��>�DE	�����ڽ����3�]�꼘���	",��W��\��@
Q����:�M
;�f);��:;(@C;�?G;P�H;HTI;�_I;)KI;�6I;P'I;gI;�I;>I;�I;oI;�I;mI;�I;;I;�I;gI;O'I;�6I;*KI;�_I;HTI;S�H;�?G;,@C;��:;�f);�M
;���:@Q�Y���W��
",�����]�꼘�3�ڽ������DE	�>�w��� ��z]׾�:���ea/��q<�      v�������`�{�k$_��q<�������}��w��	�6�����!���h����෾�� d�x.���^e��H[���Z:p��:�, ;��5;�A;�VF;��H;�@I;pbI;�QI;�;I;>+I;nI;I;9I;~	I;�I;.I;�I;	I;7I;I;kI;>+I;�;I;�QI;sbI;�@I;��H;�VF;�A;��5;�, ;^��:��Z:�H[��^e�x.��� d�෾�����h�!������	�6�w���}��������q<�l$_�`�{�����      <��������欿��� ����O��x����� ���l���"��ܽ���`=����u���k"�*R��2ۺ���9�?�:aL;��0;��>;�ME;H#H;�%I;�aI; WI;�@I;�.I;?!I;@I;I;
I;MI;�I;LI;I;I;@I;=!I;�.I;�@I;WI;�aI;�%I;R#H;�ME;��>;��0;aL;�?�:���98ۺ(R���k"�v������`=����ܽ��"��l�� ����뾁x���O� ������欿����      �������L��jȿk���������O���z]׾{����I�����A��=�d�m�}֮�RH��jλH�$�@(�y��:HN;��+;�<;�3D;��G;�I;�^I;l[I;�DI;%2I;�#I;DI;�I;^I;�	I;�I;�	I;^I;�I;FI;�#I;!2I;�DI;n[I;�^I;�I;��G;�3D;�<;��+;HN;q��:0(�L�$��jλRH�}֮�m�=�d��A������I�{���z]׾����O�����k���jȿL�Ῡ��      @�2i�������I�ѿk��� ���q<��:��a����q����Wн潅���'�Tb̼�zl��.��F�X�H����:��;ю&;ƫ9;&C;8MG;��H;8YI;�^I;�HI;�4I;�%I;�I;
I;�I;�
I;�	I;�
I;�I;I;�I;�%I;�4I;�HI;�^I;<YI;��H;CMG;&C;ɫ9;ώ&;��;��:<��I�X��.���zl�Tb̼��'�潅��Wн����q��a���:��q<� ��k���I�ѿ������2i�      F:�.5�.�'��������jȿ���l$_���W�Ҿە���6�����*���`=�<�漭)��GG�"6�����8�Q:��:�/";�7;^&B;��F;��H;�RI;�`I;xKI;7I;�'I;?I;I;�I;tI;u
I;qI;�I;I;BI;�'I;7I;�KI;�`I;�RI;��H;��F;_&B;�7;�/";��:(�Q:���$6��FG��)��<���`=��*������6�ە��W�Ҿ��k$_����jȿ�������.�'�.5�      ��U�Z�O�H-?�.�'���L�ῴ欿`�{�ea/���뾝���I����c���ZN�Z5������;H�` ��^�����":��:}�;��5;�`A;��F;J�H;MI;�aI;�MI;�8I;�(I;DI;�I;;I;I;I;I;>I;�I;GI;�(I;�8I;�MI;�aI;MI;N�H;��F;�`A;��5;w�;��:|�":V���b ��:H�����Z5���ZN�c������I�������ea/�`�{��欿L����.�'�H-?�Z�O�      ��i���b�Z�O�.5�2i�������������q<�����e��`
V�GE	�!���IY�i9�D�����(��R����Ⱥh�:W��:�;A�4;<�@;hF;��H;II;ybI;�NI;�9I;�)I;�I;_I;�I;dI;aI;`I;�I;_I;�I;�)I;�9I;�NI;|bI;II;��H;*hF;?�@;@�4;ޔ;Q��:T�:��Ⱥ�R����(�C���i9��IY�!��GE	�`
V��e������q<������������2i�.5�Z�O���b�      �>���8���*�O������˿p��E�b�C\�4m־^��Q�:��J�(��D�B�;��������./��J����>:ot�:p ;�J6;�DA;ZIF;�NH;��H;�!I;�I;�I;�I;SI;�I;P I;��H;�H;��H;M I;�I;SI;�I;�I;�I;�!I;��H;�NH;gIF;�DA;�J6;
p ;it�:�>:D���./���������;��E�B�(���J�Q�:�^��4m־C\�E�b�p���˿����O���*���8�      ��8��4��g&�6��<����<ƿ񲗿�>]����P�Ѿ�p���*7����%W��KR?��|�p8�������̅����G:y �:�!;�6;�kA;eYF;�TH;D�H;�!I;�I;�I;lI;-I;�I;A I;��H;��H;��H;A I;�I;-I;lI;�I;�I;�!I;I�H;�TH;rYF;�kA;�6;�!;s �:��G:ȅ�������p8���|�LR?�%W�����*7��p��P�Ѿ����>]�񲗿�<ƿ<���6���g&��4�      ��*��g&��#�t�U[�pL�������M�r5��>ľ����,��D�蒐��5�1�ݼ���q
��x�uk���b:1l�:�#;Ɨ7;S�A;��F;�dH;�I;#"I;�I;GI;I;�I;�I;��H;`�H;��H;Y�H;��H;�I;�I;I;DI;�I;&"I;�I;�dH;��F;T�A;7;�#;'l�:��b: uk��x��q
���0�ݼ�5�蒐��DὩ�,����>ľr5���M����pL��U[�t��#��g&�      O�6��t����˿@1��6�y�Î6��z �����1�l�+��ͽ#�����&���˼>�k� �����X�� �~��:;�;�&;�9;k�B;��F;�}H;�	I;2"I;I;�I;|I;YI;(I;��H;	�H;f�H;�H;��H;(I;VI;}I;�I; I;5"I;�	I;�}H;��F;k�B;~9;�&;8�;v��:ܙ ���X����>�k���˼��&�#����ͽ+�1�l������z �Î6�6�y�@1���˿���t�6��      ����<���U[忶˿�T���{�R�����E۾җ����M���	������j��3�d����O�7�׻��/�0��G��:� 
;�*;P;;�jC;�'G;؛H;�I;�!I;�I;xI;�
I;�I;�I;%�H;��H;��H;��H;&�H;�I;�I;�
I;vI;�I;�!I;�I;ڛH;�'G;�jC;O;;�*;� 
;=��:����/�7�׻��O�d���3���j������	���M�җ���E۾���{�R���T���˿U[�<���      �˿�<ƿpL��@1����>]���)��$��ֳ���{���,�q��'��P`I��J���,���3/��+��� �@-69�4�:ք;�o.;.=;?aD;��G;V�H;�I;!I;?I;*I;�	I;�I;� I;��H;��H;E�H;��H;��H;� I;�I;�	I;*I;FI;!I;�I;S�H;��G;@aD;.=;�o.;҄;�4�:`-69� ��+���3/��,���J��P`I�'��q�齤�,���{�ֳ��$����)��>]��@1��pL���<ƿ      p��񲗿���6�y�{�R���)�nv��>ľ^���I�Xl����������&�ӮҼ�}�/B�Ȯ�������!:�*�:&z;\3;Lj?;r\E;��G;��H;LI;I;kI;�I;XI;�I;��H;��H;F�H;��H;C�H;��H;��H;�I;VI;�I;tI;�I;KI;��H;��G;v\E;Lj?;\3;$z;�*�:��!:���ʮ��.B��}�ӮҼ��&��������Xl��I�^���>ľnv���)�{�R�6�y����񲗿      E�b��>]���M�Î6�����$���>ľ"q��y�Z�+�Q9ݽ W����L���� F���G�
�׻ ;�o칈Ȋ:�i;P$;��7;X�A;�IF;CH;��H;� I;DI;WI;�I;
I;�I;��H;��H;v�H;��H;u�H;��H;��H;I;I;�I;]I;EI;� I;��H;CH;�IF;T�A;��7;P$;�i;�Ȋ: o� ;�
�׻�G� F�������L� W��Q9ݽ+�y�Z�"q���>ľ�$�����Î6���M��>]�      C\����r5��z ��E۾ֳ�^��y�Z�K?#����A����j�%��Cϼ�����ǵ���lۺ�9�9h4�:E�;J�,;X�;;�C;G; �H;�I;�!I;�I;%I;I;tI;$I;��H;��H;��H;�H;��H;��H;��H;#I;sI;I;)I;�I;�!I;�I;#�H;�G; �C;[�;;K�,;@�;v4�:�9�9�lۺƵ����� ��Bϼ$����j��A�����K?#�y�Z�^��ֳ��E۾�z �r5����      4m־P�Ѿ�>ľ����җ����{��I�+�����V���{�>�/�$���,��==�@�һg�@�$� ���k:��:�a;��3;
j?;R2E;��G;B�H;I;N I;�I;�I;�I;�I;��H;��H;��H;��H;8�H;��H;��H;��H;��H;�I;�I;�I;�I;Q I;I;A�H;��G;R2E;j?;��3;�a;��:��k:,� �d�@�>�һ==��,��$��>�/��{��V�����+��I���{�ӗ�������>ľP�Ѿ      ^���p����1�l���M���,�Xl�Q9ݽ�A���{���5��J��;���T[� ?�����TP��@P�9��:��;*;�9;5kB;��F;WNH;W�H; I;hI;�I; I;�I;"I;F�H;��H;��H;��H;I�H;��H;��H;��H;D�H; I;�I;I;�I;lI;  I;V�H;[NH;��F;9kB;�9;*;��;��:8P�9HP������?��T[�;���J����5��{��A��Q9ݽXl���,���M�1�l����p��      Q�:��*7���,�+���	�q�齂��� W����j�>�/��J���I���k�k�.��^�����Ȋ:1o�:�;Fr3;�>;�D;P�G;'�H;�I;!I;�I;fI;b
I;�I;A I;��H;x�H;��H;��H;@�H;��H;��H;{�H;��H;? I;�I;g
I;mI;�I;!I;�I;)�H;P�G;�D;�>;Gr3;�;;o�:�Ȋ:� ��^��
.��i��k��I���J��>�/���j� W������q�齂�	�+���,��*7�      �J�����D��ͽ���'�������L�%��#��;���k����iI����/��/�4�>:)��:�B;A�,;��:;�B;kxF;x<H;��H;�I;sI;�I;I;�I;�I;n�H;W�H;�H;N�H;~�H;M�H;~�H;N�H;�H;U�H;m�H;�I;�I; I;�I;tI;�I;��H;x<H;nxF;�B;��:;M�,;�B;'��:L�>:x/���/�fI������k�;��#��$����L����'������ͽ�D����      (��$W��璐�#�����j�Q`I���&����Bϼ�,���T[�k�jI��`;��nk��:�4�:�;�&;��6;�!@;2E;��G;��H;�I;� I;3I;�I;�
I;I;Q I;��H;��H;��H;@�H;t�H;$�H;t�H;?�H;��H;��H;��H;V I;!I;�
I;�I;3I;� I;�I;��H;��G;2E;�!@;��6;�&;�; 5�:�:�nk�Z;�hI��i��T[��,��Bϼ�����&�P`I���j�$���璐�$W��      D�B�LR?��5���&��3��J��ҮҼF�� ��<=�?�.����/��nk���9.׳:��;$!;?3;��=;��C;��F;�cH;��H;nI;�I;�I;I;�I;�I;!�H;��H;r�H;_�H; �H;d�H;�H;b�H;�H;`�H;r�H;��H;$�H;�I;�I;	I;�I;�I;tI;��H;�cH;�F;��C;��=;C3;!;��;.׳:��9�nk���/�
.��?�<=� ��F��ҮҼ�J���3���&��5�LR?�      8���|�/�ݼ��˼d���,���}���G����?�һ����b���/��:.׳:�;Sb;��0;r<;��B;�IF;NH;�H;�I;M I;�I;I;9
I;�I; I;�H;5�H;��H;�H;�H;\�H;�H;Z�H;��H;�H;��H;5�H;�H; I;�I;?
I;I;�I;T I;�I;�H;SH;�IF;��B;u<;��0;Wb;��;4׳:�:�/�]������>�һ�����G��}��,��d����˼0�ݼ�|�      ~���o8����>�k���O��3/�,B��׻õ��`�@�DP�� ��D�>: 5�:��;Yb;��/;;; �A;j�E;��G;ԭH;�
I;E I;�I;�I;�I;�I;�I;h�H;�H;��H;x�H;��H;��H;O�H;�H;K�H;��H;��H;w�H;��H;�H;j�H;�I;�I;�I;�I;�I;J I;�
I;٭H;��G;t�E;$�A;;;��/;Zb;��;5�:D�>:� ��>P��_�@�õ���׻.B��3/���O�?�k���m8��      ������q
����1�׻�+��Į���;��lۺ� �HP�9�Ȋ:��:�; !;��0;;;��A;�pE;S�G;��H;��H;�I;I;/I;I;�I;UI;��H;%�H;Z�H;��H;��H;��H;��H;F�H;�H;C�H;��H;��H;��H;��H;]�H;*�H;��H;WI;�I;�I;7I;I;�I;��H;��H;X�G;�pE;��A;;;��0;$!;�;!��:�Ȋ:xP�9� ��lۺ�;�Ʈ���+��,�׻����q
���      !/��!����x���X���/�� ������n��9�9ĩk:��:/o�:�B;�&;C3;t<; �A;�pE;EtG;�|H;�H;I;RI;&I;�I;M
I;�I;3 I;-�H;�H;��H;^�H;��H;��H;��H;X�H;C�H;V�H;��H;��H;��H;]�H;��H;�H;.�H;7 I;�I;K
I;�I;*I;RI;I;�H;�|H;GtG;�pE;%�A;t<;G3;�&;�B;7o�:��:��k:�9�9�n����� ���/���X��x�!���      <���Ѕ���tk��� �8���-69��!:�Ȋ:z4�:��:��;�;J�,;��6;��=;��B;q�E;[�G;�|H;x�H;XI;�I;bI;<I;�I;I;iI;(�H;��H;�H;��H;��H;��H;��H;��H;o�H;V�H;k�H;��H;��H;��H;��H;��H;�H;��H;.�H;iI;I;�I;?I;cI;�I;_I;z�H;�|H;W�G;t�E;��B;��=;��6;M�,;�;��;��:|4�:�Ȋ:��!:�-69��̙ ��tk�����      p�>:\�G:��b:n��:)��:�4�:�*�:�i;B�;�a;*;Br3;��:;�!@;��C;�IF;��G;��H;�H;WI;�I;I;I;�I;�I;:I;��H;n�H;��H;[�H;-�H;��H;}�H;��H;��H;��H;f�H;��H;��H;��H;|�H;��H;0�H;_�H;��H;p�H;��H;<I;�I;�I;I;%I; I;ZI;�H;��H;��G;�IF;��C;�!@;��:;Gr3;*;�a;@�;�i;�*�:�4�:C��:t��:��b:d�G:      ot�:� �:Ol�:L�;� 
;؄;$z;P$;Q�,;��3;�9;�>;�B;2E;�F;SH;٭H;��H;I;�I;%I;^I;I;�I;�I;��H;�H;1�H;��H;{�H;��H;��H;r�H;��H;�H;��H;��H;��H;�H;��H;r�H;��H;��H;|�H;��H;4�H;�H;��H;�I;�I;I;cI;)I;�I;I;��H;ޭH;UH;�F;2E;�B;	�>;�9;��3;P�,;
P$;*z;҄;� 
;C�;;l�:� �:      *p ;�!;�#;�&;�*;�o.;g3;��7;b�;;j?;@kB;�D;qxF;��G;�cH;�H;�
I;�I;UI;cI;I;I;�I;=I;�H;q�H;p�H;�H;��H;��H;��H;e�H;u�H;��H;9�H;�H;��H;��H;8�H;��H;u�H;c�H;��H;��H;��H;�H;p�H;u�H;�H;;I;�I;I;!I;fI;VI;�I;�
I;�H;�cH;��G;rxF;�D;FkB;j?;c�;;��7;f3;�o.;�*;�&;�#;�!;      �J6; �6;7;~9;E;;.=;Ij?;V�A;�C;T2E;��F;P�G;v<H;��H;��H;�I;J I;!I;(I;9I;�I;�I;7I;2�H;��H;��H;C�H;�H;!�H;��H;j�H;V�H;w�H;�H;��H;V�H;-�H;P�H;��H;�H;w�H;T�H;m�H;��H; �H;�H;A�H;��H;��H;2�H;7I;�I;�I;9I;)I;I;L I;�I;��H;��H;v<H;S�G;��F;U2E; �C;^�A;Hj?;.=;U;;~9;ė7;�6;      EA;�kA;P�A;g�B;�jC;PaD;~\E;�IF;�G;��G;bNH;.�H;��H;�I;vI;[ I;�I;<I;�I;�I;�I;�I;�H;��H;��H;_�H;�H;2�H;��H;{�H;O�H;h�H;��H;C�H;��H;��H;��H;��H;��H;C�H;��H;b�H;R�H;{�H;��H;3�H;�H;c�H;��H;��H;�H;�I;�I;�I;�I;:I;�I;^ I;yI;�I;��H;3�H;dNH;��G;�G;�IF;~\E;FaD;�jC;m�B;Q�A;�kA;      ]IF;vYF;��F;��F;w'G;G;��G;CH; �H;H�H;Z�H;�I;�I;� I;�I;�I;�I;I;M
I;I;@I;��H;q�H;��H;]�H;:�H;D�H;��H;|�H;_�H;I�H;��H;�H;�H;9�H;�H;	�H;�H;6�H;�H;�H;��H;I�H;\�H;|�H;��H;D�H;A�H;c�H;��H;t�H;��H;CI;I;O
I;I;�I; I;�I;� I;�I;�I;b�H;I�H;$�H;CH;��G;��G;�'G;��F;��F;tYF;      �NH;�TH;�dH;�}H;ϛH;V�H;��H;��H;�I;I; I;!I;qI;3I;�I;I;�I;�I;�I;mI;�H;�H;r�H;J�H;�H;A�H;��H;��H;N�H;N�H;��H;��H;W�H;��H;��H;��H;z�H;��H;��H;��H;W�H;��H;��H;P�H;M�H;��H;��H;J�H;�H;H�H;u�H;�H;	�H;lI;�I;�I;�I;I;�I;0I;sI;!I; I;I;�I;��H;��H;Q�H;�H;�}H;�dH;{TH;      ��H;L�H;�I;�	I;�I;�I;WI;� I;�!I;W I;mI;�I;�I;�I;I;?
I;�I;UI;5 I;+�H;q�H;.�H;�H;�H;+�H;��H;}�H;_�H;D�H;v�H;��H;4�H;��H;t�H;3�H;�H;��H;�H;3�H;u�H;��H;2�H;��H;u�H;D�H;`�H;}�H;��H;2�H;�H;�H;4�H;t�H;+�H;4 I;SI;�I;A
I;I;�I;�I;�I;sI;X I;�!I;� I;WI;�I;�I;�	I;�I;@�H;      �!I;�!I;#"I;D"I;�!I;!I;�I;HI;�I;�I;�I;oI; I;�
I;�I;�I;�I;��H;4�H;��H;��H;��H;��H;!�H;��H;u�H;G�H;G�H;��H;��H;"�H;��H;@�H;��H;��H;��H;��H;��H;��H;��H;D�H;��H;%�H;��H;��H;G�H;F�H;y�H;��H;�H;��H;��H;��H;��H;4�H;��H;�I;�I;�I;�
I;!I;oI;�I;�I;�I;HI;�I;!I;�!I;J"I;"I;�!I;      �I;�I;�I;I;�I;?I;nI;]I;(I;�I;I;k
I;�I;#I;�I; I;p�H;%�H;�H;#�H;c�H;y�H;��H;��H;v�H;T�H;J�H;w�H;��H;�H;��H;?�H;��H;��H;b�H;C�H;2�H;B�H;_�H;��H;��H;<�H;��H;�H;��H;y�H;I�H;\�H;}�H;��H;��H;{�H;a�H;�H;�H;#�H;q�H;
 I;�I;I;�I;i
I;	I;�I;+I;[I;rI;?I;�I;I;�I;�I;      �I;�I;PI;�I;wI;-I;�I;�I;I;	I;�I;�I;�I;^ I;+�H;�H;(�H;a�H;��H;��H;9�H;��H;��H;m�H;O�H;F�H;��H;��H;)�H;��H;�H;��H;o�H;4�H;�H;��H;��H;��H;�H;6�H;p�H;��H;�H;��H;%�H;��H;��H;M�H;U�H;m�H;��H;��H;6�H;��H;��H;a�H;)�H;�H;,�H;] I;�I;�I;�I;	I;I;�I;�I;#I;�I;�I;OI;�I;      �I;sI;I;tI;�
I;�	I;[I;I;}I;�I;"I;F I;t�H;��H;��H;=�H;��H;��H;h�H; �H;��H;��H;d�H;U�H;f�H;��H;��H;6�H;��H;@�H;��H;P�H;�H;��H;��H;��H;��H;��H;��H;��H;�H;M�H;��H;=�H;��H;3�H;��H;��H;j�H;Q�H;k�H;��H;��H;��H;g�H;��H;��H;@�H;��H;��H;r�H;E I;)I;�I;xI;I;dI;�	I;�
I;|I;I;rI;      ZI;9I;�I;[I;�I;�I;�I;�I; I;��H;J�H;��H;\�H;��H;y�H;��H;��H;�H;��H;��H;��H;y�H;u�H;w�H;��H;�H;W�H;��H;H�H;��H;l�H;�H;��H;��H;��H;g�H;a�H;g�H;��H;��H;��H;�H;j�H;��H;D�H;��H;Y�H;�H;��H;x�H;|�H;x�H;��H;��H;��H;�H;��H;��H;y�H;��H;]�H;��H;M�H;��H;#I;~I;�I;�I;�I;XI;�I;6I;      �I;�I;�I; I;�I;� I;��H;��H;��H;��H;��H;��H;!�H;��H;j�H;�H;��H;��H;��H;��H;��H;��H;��H;�H;?�H;{�H;��H;x�H;��H;��H;/�H;��H;��H;h�H;S�H;C�H;7�H;C�H;Q�H;i�H;��H;��H;1�H;��H;��H;t�H;��H;|�H;A�H;�H;��H;��H;��H;��H;��H;��H;��H;�H;g�H;��H;�H;��H;��H;��H;�H;��H; I;� I;�I;!I;�I;�I;      H I;V I; I;��H;4�H;~�H;��H;��H;��H;��H;��H;��H;\�H;M�H;-�H;
�H; �H;��H;��H;��H;�H;�H;6�H;��H;��H;/�H;��H;5�H;��H;f�H;��H;��H;��H;Q�H;0�H; �H;%�H;"�H;,�H;S�H;��H;��H;��H;_�H;��H;0�H;��H;2�H;��H;��H;;�H;�H;��H;��H;��H;��H;�H;�H;*�H;K�H;\�H;��H;��H;��H;��H;��H;��H;~�H;3�H;��H; I;V I;      ��H;��H;\�H;�H;��H;��H;P�H;}�H;��H;��H;��H;��H;��H;}�H;i�H;^�H;V�H;F�H;^�H;r�H;��H;��H;��H;H�H;��H;�H;��H;�H;��H;I�H;��H;��H;l�H;E�H;&�H;�H;
�H;�H;"�H;I�H;o�H;��H;��H;C�H;��H;�H;��H;�H;��H;H�H;�H;��H;��H;k�H;]�H;L�H;X�H;a�H;i�H;~�H;��H;��H;��H;��H;��H;{�H;X�H;��H;��H;�H;X�H;��H;      �H;��H;��H;l�H;��H;B�H;��H;��H;�H;;�H;W�H;N�H;Y�H;4�H;#�H;"�H;�H; �H;L�H;^�H;r�H;��H;��H;&�H;��H; �H;w�H;��H;��H;8�H;��H;��H;d�H;4�H;&�H;�H;�H;
�H;#�H;5�H;h�H;��H;��H;2�H;��H;��H;z�H;�H;��H;%�H;��H;��H;j�H;Z�H;L�H;#�H;�H;%�H;#�H;4�H;Y�H;L�H;[�H;<�H;	�H;��H;��H;A�H;��H;p�H;��H;��H;      ��H;��H;V�H;�H;��H;��H;P�H;{�H;��H;��H;��H;��H;��H;~�H;i�H;^�H;V�H;F�H;^�H;r�H;��H;��H;��H;H�H;��H;�H;��H;�H;��H;G�H;��H;��H;n�H;F�H;&�H;�H;
�H;�H; �H;H�H;o�H;��H;��H;B�H;��H;��H;��H;�H;��H;F�H;�H;��H;��H;m�H;]�H;J�H;V�H;a�H;i�H;{�H;��H;��H;��H;��H;��H;}�H;V�H;��H;��H;	�H;Y�H;��H;      < I;V I;  I;��H;6�H;z�H;��H;��H;��H;��H;��H;��H;^�H;M�H;-�H;�H; �H;��H;��H;��H;�H; �H;8�H;��H;��H;-�H;��H;3�H;��H;e�H;��H;��H;��H;Q�H;.�H;"�H;%�H;#�H;-�H;S�H;��H;��H;��H;_�H;��H;/�H;��H;3�H;��H;��H;;�H;�H;��H;��H;��H;��H;�H;�H;*�H;M�H;\�H;��H;��H;��H;��H;��H;��H;{�H;9�H;��H; I;W I;      �I;�I;�I;"I;�I;� I;��H;��H;�H;��H;��H;��H;�H;��H;j�H;�H;��H;��H;��H;��H;��H;��H;��H;�H;C�H;{�H;��H;w�H;��H;��H;/�H;��H;��H;h�H;V�H;B�H;7�H;C�H;Q�H;i�H;��H;��H;/�H;��H;��H;t�H;��H;}�H;A�H;�H;��H;��H;��H;��H;��H;��H;��H;�H;j�H;��H; �H;��H;��H;��H;�H;��H; I;� I;�I;$I;�I;�I;      YI;=I;�I;XI;�I;�I;�I;�I;#I;��H;H�H;��H;\�H;��H;|�H;��H;��H;�H;��H;��H;��H;y�H;t�H;x�H;��H;�H;Y�H;��H;J�H;��H;i�H;�H;��H;��H;��H;h�H;a�H;h�H;��H;��H;��H; �H;j�H;��H;A�H;��H;Y�H;�H;��H;t�H;{�H;v�H;��H;��H;��H;�H;��H;��H;y�H;��H;`�H;��H;M�H;��H;$I;�I;�I;�I;�I;]I;�I;9I;      uI;sI;I;uI;�
I;�	I;aI;I;wI;�I;'I;H I;r�H;��H;��H;?�H;��H;��H;g�H;��H;��H;��H;g�H;U�H;j�H;��H;��H;7�H;��H;?�H;��H;M�H;�H;��H;��H;��H;��H;��H;��H;��H;�H;N�H;��H;=�H;��H;2�H;��H;��H;f�H;M�H;k�H;��H;��H;��H;e�H;��H;��H;?�H;��H;��H;u�H;H I;(I;�I;zI;I;aI;�	I;�
I;|I;I;nI;      �I;�I;LI;�I;}I;,I;�I; I;I;	I;�I;�I;�I;^ I;,�H;�H;)�H;a�H;��H;��H;;�H;��H;��H;n�H;T�H;F�H;��H;��H;,�H;��H;�H;��H;o�H;5�H;�H;��H;��H;��H;�H;8�H;p�H;��H;�H;��H;#�H;��H;��H;J�H;O�H;j�H;��H;��H;4�H;��H;��H;a�H;+�H;�H;.�H;^ I;�I;�I;�I;	I;I;I;�I;'I;�I;�I;SI;�I;      �I;�I;�I;!I;�I;JI;qI;dI;+I;�I;I;m
I;�I;!I;�I; I;p�H;(�H;�H;#�H;f�H;}�H;��H;��H;|�H;U�H;L�H;y�H;��H;�H;��H;?�H;��H;��H;e�H;B�H;2�H;D�H;a�H;��H;��H;@�H;��H;�H;��H;v�H;J�H;Y�H;{�H;��H;��H;{�H;_�H;�H;�H;#�H;p�H; I;�I;!I;�I;k
I;I;�I;)I;^I;uI;<I;�I;'I;�I;�I;      �!I;�!I;3"I;B"I;�!I;!I;�I;II;�I;�I;�I;pI;!I;�
I;�I;�I;�I;��H;3�H;��H;��H;��H;��H;"�H;��H;t�H;G�H;I�H;��H;��H;#�H;��H;A�H;��H;��H;��H;��H;��H;��H;��H;C�H;��H;%�H;��H;��H;C�H;G�H;x�H;��H;�H;��H;��H;��H;��H;5�H;��H;�I;�I;�I;�
I;!I;mI;�I;�I;�I;KI;�I;!I;�!I;B"I;3"I;�!I;      ��H;B�H;zI;�	I;�I;�I;YI;� I;�!I;X I;mI;�I;�I;�I;I;@
I;�I;WI;4 I;+�H;t�H;3�H;	�H;�H;3�H;��H;}�H;`�H;I�H;u�H;��H;4�H;��H;t�H;6�H;�H;��H;�H;3�H;u�H;��H;4�H;��H;v�H;C�H;\�H;}�H;��H;,�H;�H;�H;0�H;p�H;+�H;5 I;PI;�I;?
I;I;�I;�I;�I;rI;Y I;�!I;� I;YI;�I;�I;�	I;�I;B�H;      �NH;�TH;�dH;�}H;ޛH;X�H;��H;��H;�I;I; I;!I;pI;3I;�I;I;�I;�I;�I;lI;	�H;�H;o�H;M�H;�H;D�H;��H;��H;Q�H;N�H;��H;��H;V�H;��H;��H;��H;z�H;��H;��H;��H;W�H;��H;��H;N�H;K�H;�H;��H;H�H;�H;F�H;v�H;�H;�H;oI;�I;�I;�I;I;�I;0I;pI;!I; I;I;�I;��H;��H;T�H;�H;�}H;�dH;�TH;      SIF;rYF;��F;��F;~'G;̈G;��G;CH;$�H;F�H;a�H;�I;�I;� I;�I; I;�I;I;O
I;I;FI;��H;o�H;��H;c�H;;�H;D�H;��H;��H;\�H;I�H;��H;�H;��H;9�H;�H;�H;�H;6�H;�H;�H;��H;L�H;]�H;y�H;��H;G�H;;�H;`�H;��H;t�H;��H;AI;I;Q
I;I;�I; I;�I;� I;�I;�I;a�H;I�H;�H;CH;��G;��G;�'G;��F;��F;eYF;      EA;�kA;O�A;m�B;�jC;UaD;�\E;�IF;�G;��G;dNH;3�H;��H;�I;{I;^ I;�I;@I;�I;�I;�I;�I;�H;��H;��H;]�H;�H;3�H;��H;y�H;O�H;h�H;��H;C�H;��H;��H;��H;��H;��H;F�H;��H;i�H;T�H;|�H;��H;0�H;�H;b�H;��H;��H;�H;�I;�I;�I;�I;:I;�I;_ I;|I;�I;��H;0�H;bNH;��G;�G;�IF;�\E;GaD;�jC;k�B;J�A;�kA;      �J6;�6;��7;�9;@;; .=;Mj?;Z�A;$�C;R2E;��F;T�G;x<H;��H;��H;�I;L I;"I;)I;:I;�I;�I;7I;3�H;��H;��H;A�H;�H;"�H;��H;k�H;X�H;x�H;�H;��H;T�H;.�H;V�H;��H;�H;z�H;X�H;n�H;��H;�H;�H;D�H;��H;��H;0�H;9I;�I;�I;:I;*I;I;L I;�I;��H;��H;u<H;Q�G;��F;U2E;�C;T�A;Lj?;.=;W;;�9;��7;�6;      p ;�!;�#;�&;�*;�o.;c3;��7;h�;;j?;>kB;�D;qxF;��G;�cH;�H;�
I;�I;VI;fI;I;I;�I;>I;�H;n�H;o�H;�H;��H;��H;��H;h�H;t�H;��H;<�H;�H;��H;�H;6�H;��H;u�H;h�H;��H;��H;��H;�H;u�H;q�H;�H;:I;�I;I;I;fI;XI;�I;�
I;�H;�cH;��G;rxF;�D;>kB;j?;e�;;��7;c3;�o.;�*;�&;�#;�!;      gt�:� �:1l�:E�;� 
;��;,z;P$;R�,;��3;�9;�>;�B;2E;
�F;VH;ۭH;��H;I;�I;)I;cI;I;�I;�I;��H;�H;4�H;��H;y�H;��H;��H;r�H;��H;�H;��H;��H;��H;�H;��H;u�H;��H;��H;}�H;��H;1�H;�H;��H;�I;�I;I;aI;)I;�I;I;��H;ۭH;UH;�F;2E;�B;�>;�9;��3;R�,;P$;&z;Ȅ;� 
;7�;5l�:� �:      D�>:��G:��b:|��:/��:�4�:�*�:�i;E�;�a;*;Ir3;��:;�!@;��C;�IF;��G;��H;�H;[I; I;&I;I;�I;�I;9I;��H;n�H;��H;Z�H;,�H;��H;}�H;��H;��H;��H;f�H;��H;��H;��H;}�H;��H;0�H;^�H;��H;n�H;��H;9I;�I;�I;I;"I; I;[I;�H;��H;��G;�IF;��C;�!@;��:;Dr3;*;�a;A�;�i;�*�:�4�:S��:z��:��b:p�G:      ���ʅ���tk��� �8��.69��!:�Ȋ:�4�:��:��;�;K�,;��6;��=;��B;t�E;[�G;�|H;{�H;_I;�I;bI;:I;�I;I;eI;*�H;��H;�H;��H;��H;��H;��H;��H;k�H;V�H;m�H;��H;��H;��H;��H;��H;�H;��H;*�H;jI;I;�I;=I;fI;�I;]I;z�H;�|H;W�G;t�E;��B;��=;��6;J�,;�;��;��:z4�:�Ȋ:��!:�-69����� ��tk�҅��       /��!����x���X���/�� � ����n��9�9ĩk:��:;o�:�B;�&;H3;x<;#�A;�pE;FtG;�|H;�H;I;SI;&I;�I;K
I;�I;3 I;.�H;�H;��H;`�H;��H;��H;��H;V�H;C�H;W�H;��H;��H;��H;a�H;��H;�H;-�H;3 I;�I;K
I;�I;)I;SI;
I;�H;�|H;EtG;�pE;#�A;r<;G3;�&;�B;5o�:��:��k:�9�9�n� ���� ���/���X��x� ���      ������q
����/�׻�+��Į���;��lۺ� �`P�9�Ȋ:#��:�;$!;��0;;;��A;�pE;X�G;��H;��H;�I;I;5I;�I;�I;UI;��H;#�H;[�H;��H;��H;��H;��H;D�H;�H;F�H;��H;��H;��H;��H;]�H;%�H;��H;VI;�I;�I;0I;I;�I;��H;��H;X�G;�pE;��A;;;��0;$!;�;��:�Ȋ:pP�9� ��lۺ�;�Ů���+��.�׻����q
���      ���o8����<�k���O��3/�-B��׻ĵ��_�@�@P��� ��D�>:5�:��;]b;��/;;;#�A;q�E;��G;׭H;�
I;J I;�I;�I;�I;�I;�I;e�H;�H;��H;x�H;��H;��H;N�H;�H;N�H;��H;��H;w�H;��H;�H;h�H;�I;�I;�I;�I;�I;H I;�
I;ԭH;��G;r�E;!�A;;;��/;Zb;��; 5�:@�>:� ��>P��`�@�µ���׻.B��3/���O�>�k���n8��      8���|�0�ݼ��˼d���,���}���G����?�һ����]���/��:8׳:��;Tb;��0;t<;��B;�IF;RH;
�H;�I;T I;�I;I;7
I;�I;  I;�H;8�H;��H;�H;�H;Y�H;�H;Y�H;��H;�H;��H;6�H;�H; I;�I;9
I;I;�I;O I;�I;�H;PH;�IF;��B;q<;��0;Wb;�;0׳:�:�/�a������@�һ��� �G��}��,��d����˼1�ݼ�|�      D�B�KR?��5���&��3��J��ҮҼF�� ��<=�?�
.����/��nk�0��94׳:��;"!;C3;��=;��C;�F;�cH;��H;tI;�I;�I;I;�I;�I;$�H;��H;r�H;b�H; �H;b�H;�H;d�H;�H;`�H;r�H;��H;$�H;�I;�I;I;�I;�I;oI;��H;�cH;�F;��C;��=;?3;!;��;(׳:���9�nk���/�.��?�>=� ��F��ӮҼ�J���3���&��5�LR?�      (��$W��蒐�#�����j�P`I���&����Bϼ�,���T[�i�hI��[;��nk��: 5�:�;�&;��6;�!@;2E;��G;��H;�I;� I;0I;�I;�
I;I;V I;��H;��H;��H;?�H;s�H;&�H;v�H;:�H;��H;��H;��H;S I;I;�
I;�I;/I;� I;�I;��H;��G;2E;�!@;��6;�&;�;�4�:�:�nk�];�jI��j��T[��,��Bϼ�����&�P`I���j�#���璐�$W��      �J�����D��ͽ���'�������L�$��#��;���k����hI����/�|/�@�>:#��:�B;J�,;��:;�B;qxF;{<H;��H;�I;pI;�I;I;�I;�I;p�H;W�H;�H;N�H;~�H;M�H;~�H;L�H;�H;W�H;m�H;�I;�I;I;�I;qI;�I;��H;v<H;rxF;�B;��:;K�,;�B;!��:<�>:�/���/�iI������k�;��$��$����L����'������ͽ�D����      Q�:��*7���,�+���	�q�齂��� W����j�>�/��J���I���k�j�
.��]�� ���Ȋ:7o�:�;Nr3;�>;�D;S�G;+�H;�I;!I;�I;jI;`
I;�I;? I;��H;{�H;��H;��H;A�H;��H;��H;z�H;��H;? I;�I;d
I;mI;�I;!I;�I;$�H;S�G;�D;�>;Br3;�;1o�:�Ȋ:� ��_��.��k��k��I���J��>�/���j� W������q�齂�	�+���,��*7�      ^���p����1�l���M���,�Xl�Q9ݽ�A���{���5��J��;���T[�?�����RP��(P�9��:��;*;�9;;kB;��F;[NH;X�H;  I;iI;�I;I;�I;"I;F�H;��H;��H;��H;J�H;��H;��H;��H;F�H; I;�I;I;�I;kI;�I;W�H;YNH;��F;;kB;�9;	*;��;��:8P�9HP������ ?��T[�;���J����5��{��A��Q9ݽXl���,���M�1�l����p��      4m־P�Ѿ�>ľ����җ����{��I�+�����V���{�>�/�#���,��<=�>�һd�@�8� ���k:��:�a;��3;j?;U2E;��G;B�H;I;P I;�I;�I; 	I;�I;��H;��H;��H;��H;8�H;��H;��H;��H;��H;�I;�I;�I;�I;Q I;I;B�H;��G;R2E;j?;��3;�a;��:��k:,� �d�@�@�һ==��,��$��>�/��{��V�����+��I���{�җ�������>ľP�Ѿ      C\����r5��z ��E۾ֳ�^��y�Z�K?#����A����j�$��Cϼ �����ǵ���lۺ�9�9t4�:G�;H�,;Y�;; �C;�G; �H;�I;�!I;�I;%I;	I;tI;&I;��H;��H;��H;�H;��H;��H;��H;#I;vI;I;'I;�I;�!I;�I;#�H;�G;"�C;[�;;H�,;@�;v4�:�9�9�lۺǵ�������Cϼ%����j��A�����K?#�y�Z�^��ֳ��E۾�z �r5����      E�b��>]���M�Î6�����$���>ľ"q��y�Z�+�Q9ݽ W����L���� F���G�
�׻;��n칎Ȋ:�i;P$;��7;Z�A;�IF;CH;��H;� I;EI;WI;�I;
I;�I;��H;��H;t�H;��H;t�H;��H;��H;�I;	I;�I;]I;EI;� I;��H;CH;�IF;V�A;��7;P$;~i;�Ȋ:o� ;��׻�G� F�������L� W��Q9ݽ+�y�Z�"q���>ľ�$�����Î6���M��>]�      p��񲗿���6�y�{�R���)�nv��>ľ^���I�Xl����������&�ҮҼ�}�.B�ʮ�������!:�*�:&z;[3;Lj?;t\E;��G;��H;KI;I;mI;�I;XI;�I;��H;��H;C�H;��H;C�H;��H;��H;�I;ZI;�I;qI;�I;LI;��H;��G;s\E;Lj?;_3;$z;�*�:��!:���ʮ��.B��}�ӮҼ��&��������Xl��I�^���>ľnv���)�{�R�6�y����񲗿      �˿�<ƿpL��@1����>]���)��$��ֳ���{���,�q��'��P`I��J���,���3/��+��� ��-69�4�:҄;�o.;.=;?aD;��G;Q�H;�I;!I;BI;.I;�	I;�I;� I;��H;��H;E�H;��H;��H;� I;�I;�	I;*I;EI;!I;�I;T�H;��G;@aD;.=;�o.;҄;�4�:�-69� ��+���3/��,���J��P`I�'��q�齤�,���{�ֳ��$����)��>]��@1��pL���<ƿ      ����<���U[忶˿�T���{�R�����E۾җ����M���	������j��3�d����O�8�׻��/�(��G��:� 
;�*;O;;�jC;}'G;כH;�I;�!I;�I;xI;�
I;�I;�I;"�H;��H;��H;��H;%�H;�I;�I;�
I;vI;�I;�!I;�I;ۛH;�'G;�jC;R;;�*;� 
;=��: ����/�7�׻��O�d���3���j������	���M�җ���E۾���{�R���T���˿U[�<���      O�6��t����˿@1��6�y�Î6��z �����1�l�+��ͽ#�����&���˼>�k� �����X�ܙ ����::�;�&;}9;k�B;��F;�}H;�	I;2"I;I;�I;}I;VI;(I;��H;�H;f�H;�H;��H;%I;XI;I;�I;#I;5"I;�	I;�}H;��F;j�B;�9;�&;8�;z��:ؙ ���X����=�k���˼��&�#����ͽ+�1�l������z �Î6�6�y�@1���˿���t�6��      ��*��g&��#�t�U[�pL�������M�r5��>ľ����,��D�蒐��5�0�ݼ���q
��x�uk���b:+l�:�#;Ǘ7;V�A;��F;�dH;�I;#"I;�I;II;I;�I;�I;��H;]�H;��H;Y�H;��H;�I;�I;I;EI;�I;&"I;�I;�dH;��F;T�A;×7;�#;'l�:��b:�tk��x��q
���0�ݼ�5�蒐��DὩ�,����>ľr5���M����pL��U[�t��#��g&�      ��8��4��g&�6��<����<ƿ񲗿�>]����P�Ѿ�p���*7����%W��KR?��|�p8�������ʅ����G:y �:�!;�6;�kA;dYF;�TH;D�H;�!I;�I;�I;lI;-I;�I;A I;��H;��H;��H;A I;�I;-I;nI;�I;�I;�!I;I�H;�TH;rYF;�kA;�6;�!;s �:��G:ą�������p8���|�KR?�%W�����*7��p��P�Ѿ����>]�񲗿�<ƿ<���6���g&��4�      ��$������꿮�ſ�ޞ�%3s��2�=����� j���yHͽŸ����'�A<ͼo�n�b���;Q^��-.�r��:nW;_S%;fo8;��A;DF;�H;{�H;��H;��H;#�H;�H;&�H;��H;��H;��H;�H;��H;��H;��H;&�H;�H; �H;��H;��H;~�H;�H;DF;��A;co8;ZS%;lW;p��:�-.�<Q^�b���o�n�A<ͼ��'�Ÿ��yHͽ�� j���=����2�%3s��ޞ���ſ������$�      $�������忇�����cm�U�-�����Ph��Vde�!-�֪ɽ�v��'�$�~�ɼymj�5���X����ņ:hx;�%;2�8;EB;RF;�H;�H;�H;��H;F�H;�H;�H;{�H;��H;��H;�H;��H;��H;{�H;�H;�H;C�H;��H;�H;�H;�H;*RF;EB;0�8;�%;ex;�ņ:��X�4���ymj�~�ɼ'�$��v��֪ɽ!-�Vde�Ph������U�-�cm��������忝����      ����������ԿLw�����:�\�"����k��Y0X�����;����w����������]����F�����ɒ:��;�';��9;�oB;�zF;�!H;s�H;��H;�H;p�H;�H;�H;��H;��H;��H;��H;��H;��H;��H;�H;�H;n�H;�H;��H;t�H;�!H;�zF;�oB;��9;��';��;�ɒ:����F��黩�]����������w��;�����Y0X�k�����"�:�\����Lw���Կ��𿝏�      ������Կp���ޞ�_F�g�C�-E�!�;�I��D���"��e�c�|��֯���J��ѻʢ)��K�'��:�
;�M*;n�:;�C;ɸF;�8H;-�H;J�H;Z�H;��H;�H;�H;��H;��H;��H;��H;��H;��H;��H;�H;�H;��H;a�H;K�H;+�H;�8H;ӸF;�C;m�:;�M*;
�
;��:PK�̢)��ѻ��J��֯�{�e�c�"����D��I��!�;-E�g�C�_F��ޞ�p���Կ��      ��ſ���Lw���ޞ�����>�W�5�%�����hɰ��|x�f{+�ѱ����J��  �Ͷ��X�1�$���+�P 
9��:��;�-;��<;]�C;�G;�TH;$�H;��H;��H;��H;.�H;�H;g�H;��H;y�H;��H;u�H;��H;g�H;�H;,�H;��H;��H;��H;&�H;�TH;�G;^�C;��<;޷-;��;��:� 
9+�$���X�1�Ͷ���  ��J���ѱ�f{+��|x�hɰ�����5�%�>�W������ޞ�Lw�����      �ޞ�������_F�>�W�W�-���?Kɾ�G����O����ƽƸ��̈́-���ۼㄼ44�ǐ��ζ�,]:���:�;~�1;�c>;D�D;x\G;.sH;x�H;5�H;D�H;��H;K�H;�H;I�H;m�H;`�H;��H;\�H;k�H;G�H;�H;M�H;��H;K�H;5�H;x�H;-sH;�\G;E�D;�c>;z�1;�;��:0]:�ζ�ǐ�44�ㄼ��ۼ̈́-�Ƹ��ƽ�����O��G��?Kɾ��W�-�>�W�_F�������      %3s�cm�:�\�h�C�5�%����TҾj��	 j��C(����^P����[�{������Y�8��^X�P�<��k:>��:�� ;֟5;4R@;6uE;ϲG;�H;"�H;��H;��H;!�H;G�H;	�H;B�H;O�H;:�H;n�H;7�H;N�H;B�H;�H;D�H;�H;��H;��H; �H;�H;ֲG;9uE;2R@;ԟ5;�� ;0��:�k:T�<�_X�6����Y����{���[�^P����콪C(�	 j�j���TҾ��5�%�h�C�:�\�cm�      �2�U�-�"�-E�����?Kɾj����s�7�5���v㻽�v��	z0��;��+���*����+6� AS�OM�:R�	;r�(;�9;�/B;HDF; H;��H;]�H;��H;��H;L�H;d�H;��H;�H;�H;�H;9�H;�H;�H;�H;��H;b�H;J�H;��H;��H;]�H;��H;%H;MDF;�/B;�9;t�(;L�	;WM�:�@S�+6�����*��+���;�z0��v��v㻽��7�5���s�j��?Kɾ����-E�"�U�-�      =����������"�;hɰ��G��	 j�7�5��	�ΪɽY����J�r���沼��]�����	x�L	��,n:���:�v;��/;f-=;��C;�F;�HH;�H;��H;��H;�H;{�H;g�H;��H;��H;��H;��H;�H;��H;��H;��H;��H;g�H;{�H;�H;��H;�H;|�H;�HH;�F;��C;j-=;��/;�v;���:,n:N	���	x������]��沼r���J�Y���Ϊɽ�	�7�5�	 j��G��hɰ�!�;��徶���      ��Ph��k���I���|x���O��C(���Ϊɽ����QDX�H��&<ͼㄼ�X!��s���W��uK�!��:�y;�#;�H6;R@;�PE;h�G;\�H;��H;�H;��H;}�H;��H;U�H;��H;��H;��H;��H;��H;��H;��H;��H;��H;Q�H;��H;��H;��H;�H;��H;\�H;l�G;�PE;R@;�H6;��#;�y;!��:�uK��W��s���X!�ㄼ%<ͼH��QDX�����Ϊɽ���C(���O��|x��I��k��Ph��       j�Vde�Y0X�D�f{+�������u㻽Y���QDX������ۼʾ����;�D>ۻX�\�y��>":���:��;·-;��;;��B;ozF;�H;`�H;Z�H;��H;��H;��H;��H;N�H;��H;z�H;q�H;��H;[�H;��H;r�H;|�H;��H;J�H;��H;��H;��H;�H;Z�H;^�H;�H;mzF;��B;��;;��-;��;���:�>":D�y�X�B>ۻ��;�ʾ����ۼ���QDX�Y���u㻽��콂��g{+�D�Y0X�Vde�      ��"-������ѱ�ƽ^P���v���J�H����ۼ��b�J������+���rѺP(
9�M�:��;v $;��5;��?;\�D;A\G;�eH;��H;��H;��H;��H;��H;��H;3�H;R�H;9�H;2�H;D�H;�H;D�H;2�H;<�H;O�H;0�H;��H;�H;��H;��H;��H;��H;�eH;A\G;d�D;��?;��5;~ $;��;�M�:�(
9~rѺ�+������a�J�����ۼH���J��v��^P��ƽұ轃����!-�      yHͽ֪ɽ�;��"����Ƹ����[�z0�r��%<ͼʾ��b�J�����j��z*�`�:@b�:;�;��/;�L<;�C;mF;p�G;ݡH;��H;��H;��H;�H;1�H;��H;�H;�H;��H;��H;��H;��H;��H;��H;��H;�H;�H;��H;8�H;�H;��H;��H;��H;�H;p�G;mF;�C;�L<;��/;@�;:b�:���: �w*��j�����a�J�ɾ��%<ͼr��z0���[�Ƹ����"���;��֪ɽ      ĸ���v����w�f�c��J�΄-�{��;缄沼ㄼ��;������j���5�P��?Q:<��:Ri;�M*;h�8;g�@;�PE;�uG;iH;��H;��H;��H;��H;��H;U�H;��H;��H;��H;��H;��H;��H;~�H;��H;��H;��H;��H;��H;��H;^�H;��H;�H;��H;��H;��H;iH;�uG;�PE;h�@;p�8;�M*;Ri;F��:?Q:0�깞5��j��������;�ㄼ�沼�;�{�̈́-��J�f�c���w��v��      ��'�'�$����|��  ���ۼ����+����]��X!�B>ۻ�+��{*�P����>:���:��;%�%;ҟ5;y�>;�(D;��F;U!H;�H;*�H;��H;��H;��H;��H;L�H;��H;��H;i�H;m�H;I�H;4�H;N�H;2�H;G�H;p�H;i�H;��H;��H;S�H;��H;��H;��H;��H;0�H;�H;X!H;��F;�(D;��>;֟5;"�%;��;���:��>:0��w*��+��@>ۻ�X!���]��+�������ۼ�  �{����'�$�      ><ͼ}�ɼ�����֯�Ͷ��ㄼ��Y��*�����s��X��rѺp�?Q:���:��
;6�#;S�3;wc=;�#C;DF;��G;�H;��H;��H;�H;��H;5�H;��H;F�H;o�H;F�H;�H;1�H;��H;��H;��H;��H;��H;1�H;�H;C�H;s�H;J�H;�H;;�H;��H;�H;��H;��H;��H;��G;	DF;�#C;zc=;O�3;:�#;��
;���:?Q:`�|rѺX��s������*���Y�ㄼζ���֯�����|�ɼ      j�n�vmj���]���J�W�1�34�2������	x��W�4�y�`(
9���:F��:��;:�#;>�2;�<;OpB;�E;��G;�eH;��H;�H;��H;��H;��H;��H;�H;*�H;�H;��H;��H;��H;��H;��H;��H;��H;��H;��H;��H;��H;�H;-�H;�H;��H;��H;��H;��H;�H;��H;�eH;��G;�E;RpB;�<;B�2;=�#;�;J��:���:�(
9$�y��W��	x����4��24�X�1���J���]�tmj�      S���.������ѻ���ǐ�VX�$6�H	��@uK�?":�M�:4b�:Oi;"�%;L�3;�<;/0B;��E;U\G;�HH;$�H;y�H;@�H;��H;�H;�H;��H;��H;��H;��H;��H;��H;B�H;5�H;5�H;�H;4�H;4�H;C�H;��H;��H;��H;�H;��H;��H;�H;�H;��H;?�H;y�H;(�H;�HH;]\G;��E;,0B;�<;O�3;%�%;Pi;8b�:�M�: ?": uK�:	��$6�ZX�ǐ�����ѻ��/���      &Q^�X��F�Ƣ)�+��ζ�4�<��?S�<n:'��:ý�:��;=�;�M*;֟5;xc=;OpB;��E;�JG;/8H;K�H;g�H;��H;
�H;c�H;��H;s�H;��H;��H;��H;v�H;]�H;8�H;��H;��H;��H;��H;��H;��H;��H;7�H;Z�H;y�H;��H;��H;��H;s�H;��H;j�H;�H;��H;l�H;R�H;68H;�JG;��E;TpB;xc=;ڟ5;�M*;@�;��;˽�:)��:Hn:�?S�<�<��ζ�+�Т)��F�X�      �-.�$��X��0~K�@ 
9@]:D�k:OM�:���:�y;��;| $;��/;n�8;��>;�#C;�E;b\G;48H;��H;��H; �H;o�H;�H;h�H;3�H;��H;��H;��H;e�H;�H;��H;��H;��H;�H;x�H;^�H;r�H;|�H;��H;��H;��H;�H;e�H;��H;��H;��H;1�H;n�H;�H;o�H;�H;��H;��H;78H;]\G;�E;�#C;��>;n�8;��/;� $;��;�y;���:]M�:8�k:X]:� 
90K����H��      ���:�ņ:�ɒ:��:��:���:0��:O�	;�v;�#;·-;��5;~L<;g�@;�(D;DF;��G;�HH;P�H;��H;��H;*�H;��H;@�H;��H;n�H;��H;��H;B�H;�H;��H;��H;V�H;I�H;�H;�H;�H;
�H;�H;I�H;S�H;��H;��H;
�H;B�H;��H;��H;o�H;�H;>�H;��H;/�H;��H;��H;R�H;�HH;��G;DF;�(D;e�@;�L<;��5;Ʒ-;�#;�v;L�	;:��:��:��:��:�ɒ:�ņ:      pW;zx;��;�
;��;�;�� ;r�(;��/;�H6;��;;��?;�C;�PE;��F;��G;�eH;+�H;l�H;�H;/�H;��H;�H;��H;A�H;d�H;l�H;L�H;��H;��H;��H;0�H; �H;��H;��H;��H;��H;��H;��H;��H;��H;*�H;��H;��H;��H;O�H;i�H;h�H;F�H;��H;�H;��H;4�H;�H;n�H;*�H;�eH;��G;��F;�PE;�C;��?;��;;�H6;��/;x�(;�� ;;��;�
;��;ox;      zS%;	�%;��';�M*;۷-;��1;�5;��9;q-=;R@;��B;f�D;
mF;�uG;\!H;��H;��H;��H;��H;m�H;��H;�H;��H;J�H;a�H;X�H;�H;��H;��H;|�H;
�H;��H;��H;��H;p�H;[�H;<�H;U�H;n�H;��H;��H;��H;�H;{�H;��H;��H;�H;]�H;g�H;I�H;��H;�H;��H;p�H;��H;{�H;��H;��H;^!H;�uG;mF;j�D;��B;R@;r-=;��9;��5;��1;�-;�M*;��';��%;      fo8;<�8;��9;n�:;~�<;�c>;1R@;�/B;��C;�PE;lzF;@\G;o�G;iH;�H;��H;�H;E�H;�H;�H;>�H;��H;F�H;V�H;J�H;*�H;��H;��H;U�H;��H;��H;��H;G�H;�H;�H;�H;��H;�H;�H;�H;F�H;��H;��H;��H;S�H;��H;��H;0�H;P�H;V�H;F�H;��H;B�H;�H;�H;B�H;�H;��H;�H;iH;o�G;E\G;szF;�PE;��C;�/B;4R@;�c>;��<;m�:;��9;2�8;      ��A;HB;�oB;�C;V�C;V�D;CuE;MDF; �F;o�G;�H;�eH;�H;��H;2�H;��H;��H;��H;q�H;t�H;�H;H�H;g�H;V�H;�H;��H;��H;Z�H;��H;��H;b�H;3�H;��H;��H;��H;��H;��H;��H;��H;��H;��H;.�H;d�H;��H;��H;\�H;��H;��H;�H;V�H;i�H;L�H;�H;r�H;t�H;��H;��H;��H;7�H;��H;�H;�eH;�H;p�G;"�F;NDF;CuE;L�D;g�C;�C;�oB;HB;      DF;.RF;�zF;ȸF;�G;�\G;ֲG;.H;�HH;c�H;c�H;��H;��H;��H;��H;�H;��H;�H;��H;1�H;r�H;d�H;X�H;3�H;��H;u�H;I�H;��H;��H;U�H;	�H;��H;��H;��H;h�H;W�H;c�H;Q�H;e�H;��H;��H;��H;	�H;T�H;��H;��H;H�H;|�H;��H;1�H;[�H;h�H;u�H;3�H;��H;�H;��H;�H;��H;��H;��H;��H;k�H;d�H;�HH;.H;زG;{\G;�G;ӸF;�zF;-RF;      �H;H;�!H;�8H;�TH;0sH;%�H;��H;~�H;��H;Z�H;��H;��H;��H;��H;��H;��H; �H;w�H;��H;��H;k�H;�H;��H;��H;G�H;��H;z�H;=�H;�H;��H;��H;W�H;9�H;#�H;�H;�H;��H; �H;;�H;W�H;��H;��H;�H;9�H;z�H;��H;O�H;��H;��H; �H;o�H;��H;��H;y�H;�H;��H;��H;��H;��H;��H;��H;^�H;��H;~�H;��H;!�H;*sH;�TH;�8H;�!H;�H;      ��H;
�H;s�H;6�H;�H;~�H;.�H;_�H;�H;�H;�H;��H;��H;�H;��H;:�H;��H;��H;��H;��H;��H;I�H;��H;��H;S�H;��H;w�H;K�H;��H;��H;i�H;?�H;�H;��H;��H;��H;��H;��H;��H;��H;�H;;�H;i�H;��H;��H;K�H;u�H;��H;Y�H;��H;��H;M�H;��H;��H;��H;��H;��H;<�H;��H;�H;��H;��H;�H;�H;�H;c�H;0�H;q�H;*�H;8�H;s�H;��H;      ��H;�H;��H;]�H;��H;8�H;��H;��H;��H;��H;��H;��H;�H;��H;��H;�H;!�H;��H;��H;��H;J�H;��H;��H;U�H;��H;��H;6�H;��H;��H;b�H;+�H;��H;��H;��H;��H;��H;w�H;��H;��H;��H;��H;��H;-�H;a�H;��H;��H;5�H;��H;��H;R�H;��H;��H;I�H;��H;��H;��H;!�H;	�H;��H;��H;�H;��H;��H;��H;��H;��H;��H;1�H;��H;`�H;��H;�H;      ��H;��H;�H;T�H;��H;D�H;��H;��H;�H;��H;��H;�H;6�H;a�H;P�H;J�H;1�H;��H;��H;h�H;�H;��H;x�H;��H;��H;J�H;�H;��H;b�H;$�H;��H;��H;��H;��H;a�H;F�H;8�H;C�H;]�H;��H;��H;��H;��H;!�H;a�H;��H;�H;R�H;��H;��H;|�H;��H;
�H;e�H;��H;��H;4�H;N�H;P�H;^�H;8�H;�H;��H;��H;�H;��H;��H;D�H;��H;Z�H;�H;��H;      )�H;`�H;|�H;��H;��H;��H;'�H;U�H;��H;��H;��H;��H;��H;��H;��H;x�H;$�H;��H;}�H;'�H;��H;��H;
�H;��H;`�H;�H;��H;m�H;1�H;��H;��H;~�H;p�H;:�H;�H;"�H; �H;�H;�H;;�H;s�H;}�H;��H;��H;-�H;j�H;��H;�H;f�H;��H;�H;��H;��H;#�H;}�H;��H;&�H;{�H;��H;��H;��H;��H;��H;��H;��H;S�H;1�H;��H;��H;��H;|�H;^�H;      �H;�H;�H;�H;'�H;G�H;J�H;i�H;n�H;V�H;O�H;:�H;�H;��H;��H;L�H;��H;��H;b�H;�H;��H;2�H;��H;��H;0�H;��H;��H;@�H;��H;��H;w�H;]�H;;�H;�H;��H;��H;��H;��H;��H;�H;?�H;[�H;v�H;��H;��H;?�H;��H;��H;5�H;��H;��H;4�H;��H;��H;b�H;��H; �H;N�H;��H;��H;�H;7�H;T�H;X�H;m�H;i�H;R�H;H�H;5�H;�H;"�H;�H;      2�H;&�H;*�H;!�H;�H;�H;�H;��H;��H;��H;��H;[�H;�H;��H;p�H; �H;��H;��H;?�H;��H;c�H;�H;��H;G�H;��H;��H;W�H;�H;��H;��H;n�H;>�H;��H;��H;��H;��H;��H;��H;��H;��H;��H;?�H;l�H;��H;��H;�H;W�H;��H;�H;H�H;��H;�H;^�H;��H;?�H;��H;��H;#�H;o�H;��H;�H;Y�H;��H;��H;��H;��H;�H;��H;"�H;�H;3�H;%�H;      �H;x�H;��H;|�H;h�H;B�H;G�H;�H;��H;��H;��H;F�H;�H;��H;x�H;<�H;��H;J�H;��H;��H;S�H;��H;�H;�H;��H;��H;5�H;��H;��H;��H;4�H;�H;��H;��H;��H;��H;��H;��H;��H;��H;��H;
�H;4�H;~�H;��H;��H;6�H;��H;��H;�H;��H;��H;O�H;��H;��H;M�H;��H;<�H;w�H;��H;�H;C�H;��H;��H;��H;�H;L�H;>�H;n�H;|�H;��H;��H;      ��H;��H;��H;��H;��H;e�H;W�H;%�H;��H;��H;�H;C�H;�H;��H;U�H;��H;��H;;�H;��H;��H;"�H;��H;k�H;�H;��H;^�H;�H;��H;��H;d�H;�H;��H;��H;��H;��H;��H;��H;��H;��H;��H;��H;��H;�H;]�H;��H;��H;�H;a�H;��H;�H;q�H;��H;�H;�H;��H;>�H;��H;��H;U�H;��H;�H;C�H;��H;��H;��H;&�H;]�H;e�H;��H;��H;��H;��H;      ��H;��H;��H;��H;m�H;Z�H;E�H;#�H;��H;��H;��H;N�H;��H;��H;9�H;��H;��H;8�H;��H;y�H;�H;��H;R�H;�H;��H;J�H;��H;��H;��H;J�H;�H;��H;��H;��H;��H;��H;��H;��H;��H;��H;��H;��H;�H;E�H;��H;��H;��H;M�H;��H;�H;Y�H;��H;�H;u�H;��H;<�H;��H;��H;9�H;��H;��H;M�H;��H;��H;��H;#�H;L�H;Z�H;q�H;��H;��H;��H;      �H;�H;�H;��H;��H;��H;x�H;@�H;
�H;��H;i�H;'�H;��H;��H;\�H;��H;��H;�H;��H;h�H;�H;��H;<�H;��H;��H;\�H;�H;��H;}�H;A�H;�H;��H;��H;��H;��H;��H;{�H;��H;��H;��H;��H;��H;�H;;�H;w�H;��H;�H;_�H;��H;��H;@�H;��H;�H;d�H;��H;�H;��H;��H;[�H;��H;��H;%�H;k�H;��H;�H;A�H;}�H;��H;��H;��H;�H;�H;      ��H;��H;��H;��H;n�H;]�H;D�H;"�H;��H;��H;��H;N�H;��H;��H;9�H;��H;��H;8�H;��H;y�H;�H;��H;T�H;�H;��H;J�H;��H;��H;��H;I�H;�H;��H;��H;��H;��H;��H;��H;��H;��H;��H;��H;��H;�H;C�H;��H;��H;��H;N�H;��H;�H;X�H;��H;�H;u�H;��H;<�H;��H;��H;9�H;��H;��H;M�H;��H;��H;��H;%�H;I�H;Z�H;q�H;��H;��H;��H;      ��H;��H;��H;��H;��H;a�H;W�H;(�H;��H;��H;~�H;C�H;�H;��H;W�H;��H;��H;<�H;��H;��H;%�H;��H;m�H;�H;��H;^�H;�H;��H;��H;b�H;�H;��H;��H;��H;��H;��H;��H;��H;��H;��H;��H;��H;�H;]�H;��H;��H;�H;b�H;��H;�H;q�H;��H;�H;�H;��H;>�H;��H;��H;S�H;��H;�H;D�H;�H;��H;��H;,�H;^�H;a�H;��H;��H;��H;��H;      �H;x�H;��H;�H;h�H;D�H;E�H;�H;��H;��H;��H;D�H;�H;��H;z�H;<�H;��H;M�H;��H;��H;S�H;��H;��H;�H;��H;��H;6�H;��H;��H;��H;4�H;
�H;��H;��H;��H;��H;��H;��H;��H;��H;��H;�H;3�H;��H;��H;��H;6�H;��H;��H;�H;��H;��H;L�H;��H;��H;L�H;��H;=�H;z�H;��H;�H;D�H;��H;��H;��H;�H;N�H;A�H;o�H;�H;��H;y�H;      0�H;,�H;-�H;�H;�H;�H;�H;��H;��H;��H;��H;[�H;�H;��H;q�H;#�H;��H;��H;A�H;��H;c�H;�H;��H;H�H;�H;��H;U�H;�H;��H;��H;l�H;<�H;��H;��H;��H;��H;��H;��H;��H;��H;��H;?�H;l�H;��H;��H;�H;W�H;��H;��H;D�H;��H;�H;\�H;��H;A�H;��H;��H;#�H;p�H;��H;�H;Y�H;��H;��H;��H;��H;�H;�H;�H;%�H;6�H;&�H;      �H;�H;�H;�H;%�H;Q�H;O�H;g�H;j�H;U�H;Q�H;9�H;�H;��H;��H;N�H;��H;��H;b�H; �H;��H;4�H;��H;��H;5�H;��H;��H;@�H;��H;��H;v�H;Z�H;;�H;�H;��H;��H;��H;��H;��H;�H;>�H;[�H;u�H;��H;��H;=�H;��H;��H;0�H;��H;��H;4�H;��H;��H;b�H;��H; �H;M�H;��H;��H;�H;9�H;R�H;X�H;m�H;g�H;R�H;F�H;(�H;�H;�H;�H;      �H;^�H;y�H;��H;��H;��H;(�H;W�H;��H;��H;��H;��H;��H;��H;��H;{�H;&�H;��H;~�H;&�H;��H;��H;�H;��H;f�H;�H;��H;m�H;2�H;��H;��H;~�H;p�H;;�H;�H; �H; �H;"�H;�H;<�H;s�H;��H;��H;��H;+�H;j�H;��H;�H;b�H;��H;�H;��H;��H;%�H;~�H;��H;'�H;z�H;��H;��H;��H;��H;��H;��H;��H;X�H;-�H;��H;��H;��H;~�H;]�H;      ��H;��H;�H;a�H;��H;O�H;��H;��H;
�H;��H;��H;�H;9�H;_�H;S�H;L�H;2�H; �H;��H;i�H;�H;��H;x�H;��H;��H;K�H;�H;��H;e�H;&�H;��H;��H;��H;��H;a�H;E�H;8�H;F�H;^�H;��H;��H;��H;��H;#�H;_�H;��H;�H;Q�H;��H;��H;�H;��H;�H;e�H;��H;��H;2�H;M�H;Q�H;_�H;8�H;�H;��H;��H;�H;��H;��H;A�H;��H;f�H;�H;��H;      ��H;�H;�H;[�H;��H;<�H;��H;��H;��H;��H;��H;��H;�H;��H;��H;�H;!�H; �H;��H;��H;M�H;��H;��H;W�H;��H;��H;5�H;��H;��H;a�H;+�H;��H;��H;��H;��H;��H;w�H;��H;��H;��H;��H;��H;-�H;b�H;��H;��H;6�H;��H;��H;N�H;��H;��H;H�H;��H;��H;��H; �H;	�H;��H;��H;�H;��H;��H;��H;��H;��H;��H;5�H;��H;Y�H;�H;�H;      ��H;��H;f�H;8�H;�H;��H;0�H;h�H;�H;�H;�H;��H;��H;�H;��H;>�H;��H;��H;��H;��H;��H;M�H;��H;��H;\�H;��H;u�H;K�H;��H;��H;i�H;?�H;�H;��H;��H;��H;��H;��H;��H;��H;�H;?�H;j�H;��H;��H;H�H;w�H;��H;U�H;��H;��H;L�H;��H;��H;��H;��H;��H;<�H;��H;�H;��H;��H;�H;�H;�H;c�H;.�H;w�H;'�H;8�H;p�H;��H;      �H;H;�!H;�8H;�TH;4sH;%�H;��H;��H;��H;\�H;��H;��H;��H;��H;��H;��H;%�H;w�H;��H;��H;o�H;�H;��H;��H;G�H;��H;{�H;?�H;�H;��H;��H;U�H;9�H;$�H;��H;�H;��H; �H;;�H;W�H;��H;��H;�H;9�H;x�H;��H;N�H;��H;��H; �H;n�H;��H;��H;y�H;�H;��H;��H;��H;��H;��H;��H;[�H;��H;~�H;��H;&�H;.sH;�TH;�8H;�!H;�H;      DF;-RF;�zF;ɸF;�G;�\G;ղG;1H;�HH;b�H;h�H;��H;��H;��H;��H;�H;��H;�H;��H;3�H;w�H;h�H;Z�H;4�H;��H;v�H;H�H;��H;��H;T�H;	�H;��H;��H;��H;i�H;S�H;f�H;U�H;e�H;��H;��H;��H;�H;U�H;��H;��H;K�H;y�H;��H;0�H;[�H;g�H;s�H;3�H;��H;�H;��H;�H;��H;��H;��H;��H;g�H;c�H;�HH;)H;ҲG;{\G;�G;ɸF;zzF;RF;      ��A;CB;�oB;�C;Z�C;Z�D;DuE;PDF;#�F;r�G;�H;�eH;�H;��H;8�H;��H;��H;��H;t�H;t�H;�H;M�H;h�H;W�H;�H;��H;��H;\�H;��H;��H;b�H;3�H;��H;��H;��H;��H;��H;��H;��H;��H;��H;5�H;g�H;��H;��H;W�H;��H;��H;�H;S�H;i�H;L�H;
�H;t�H;u�H;��H;��H;��H;8�H;��H;�H;�eH;�H;p�G;�F;NDF;CuE;M�D;b�C;�C;�oB;CB;      Bo8;"�8;��9;z�:;x�<;�c>;7R@;�/B;��C;�PE;rzF;E\G;p�G;iH;�H;��H;�H;I�H;�H;�H;D�H;��H;F�H;W�H;Q�H;*�H;��H;��H;V�H;��H;��H;��H;G�H;�H;�H;�H;��H;�H;�H;�H;H�H;��H;��H;��H;S�H;��H;��H;,�H;M�H;T�H;F�H;��H;B�H;�H;�H;B�H;�H;��H;�H;iH;o�G;C\G;pzF;�PE;��C;�/B;5R@;�c>;��<;��:;��9;�8;      eS%;�%;��';�M*;ط-;��1;ܟ5;�9;x-=;R@;��B;j�D;mF;�uG;`!H;��H;��H;��H;��H;p�H;��H;�H;��H;L�H;h�H;W�H;�H;��H;��H;y�H;�H;��H;��H;��H;q�H;[�H;?�H;[�H;m�H;�H;��H;��H;�H;}�H;��H;��H;�H;X�H;d�H;H�H;��H;�H;��H;p�H;��H;{�H;��H;��H;_!H;�uG;mF;f�D;��B;R@;t-=;�9;ܟ5;��1;ط-;�M*;��';��%;      lW;zx;��;�
;��;�;�� ;z�(;��/;�H6;��;;��?;�C;�PE;��F;��G;�eH;,�H;l�H;�H;4�H;��H;�H;��H;I�H;b�H;l�H;O�H;��H;��H;��H;0�H;��H;��H;��H;��H;��H;��H;��H;��H;��H;2�H;��H;��H;��H;L�H;n�H;e�H;C�H;��H;�H;��H;2�H;�H;l�H;(�H;�eH;��G;��F;�PE;�C;��?;��;;�H6;��/;x�(;�� ;s;��;�
;��;qx;      ���:Ɔ:�ɒ:#��:��:��::��:R�	;�v;��#;ķ-;��5;�L<;g�@;�(D;DF;��G;�HH;Q�H;��H;��H;1�H;��H;A�H;�H;l�H;��H;��H;C�H;�H;��H;��H;U�H;K�H;�H;�H;�H;�H;�H;G�H;U�H;��H;��H;�H;A�H;��H;��H;l�H;��H;@�H;��H;,�H;��H;��H;Q�H;�HH;��G;DF;�(D;e�@;�L<;��5;Ƿ-;�#;�v;S�	;>��:���:�:��:�ɒ:�ņ:      �-.������ ~K�P 
9d]:D�k:iM�:���:�y;��;� $;��/;n�8;��>;�#C;�E;b\G;68H;��H;��H;�H;o�H;�H;o�H;1�H;��H;��H;��H;a�H;�H;��H;��H;��H;}�H;r�H;^�H;t�H;{�H;��H;��H;��H; �H;d�H;��H;��H;��H;1�H;j�H;�H;p�H;�H;��H;��H;68H;]\G;�E;�#C;��>;n�8;��/;� $;��;�y;���:[M�:4�k:4]:� 
9�~K���� ��      %Q^�X��F�â)�!+��ζ�8�<��>S�Pn:)��:ý�:��;@�;�M*;ܟ5;{c=;RpB;��E;�JG;68H;R�H;k�H;��H;�H;k�H;��H;r�H;��H;��H;��H;v�H;[�H;7�H;��H;��H;��H;��H;��H;��H;��H;5�H;]�H;y�H;��H;��H;��H;s�H;��H;f�H;�H;��H;j�H;Q�H;68H;�JG;��E;QpB;wc=;ڟ5;�M*;=�;��;ý�:%��:Dn:�>S�<�<��ζ�+�Ţ)��F�X�      Z���(������ѻ���ǐ�TX�6�>	��uK�?":�M�::b�:Pi;'�%;P�3;�<;/0B;��E;]\G;�HH;(�H;}�H;B�H;��H;�H;�H;��H;��H;��H;��H;��H;��H;C�H;5�H;4�H;�H;7�H;3�H;C�H;��H;��H;��H;��H;��H;��H;�H;�H;��H;?�H;{�H;$�H;�HH;]\G;��E;,0B;�<;O�3;%�%;Oi;2b�:�M�:?":@uK�>	��"6�WX�ǐ�����ѻ"��,���      j�n�vmj���]���J�V�1�24�2������	x��W�0�y��(
9���:J��:�;?�#;B�2;�<;QpB;�E;��G;�eH;��H;�H;��H;��H;��H;��H;�H;'�H;�H;��H;��H;��H;��H;��H;��H;��H;��H;��H;��H;��H;�H;+�H;�H;��H;��H;��H;��H;�H;��H;�eH;��G;�E;OpB;�<;?�2;=�#;�;F��:���:�(
9(�y��W��	x����5��24�X�1���J���]�tmj�      ><ͼ}�ɼ�����֯�Ͷ��ㄼ��Y��*�����s��X�xrѺP�?Q:���:��
;8�#;P�3;xc=;�#C;DF;��G;��H;��H;��H;�H;��H;5�H;�H;D�H;q�H;F�H;�H;5�H;��H;��H;��H;��H;��H;1�H;�H;F�H;q�H;G�H;��H;7�H;��H;�H;��H;��H;�H;��G;DF;�#C;uc=;L�3;9�#;��
;���:?Q:p�~rѺX��s������*���Y�ㄼζ���֯�����}�ɼ      ��'�'�$����{��  ���ۼ����+����]��X!�@>ۻ�+��w*�@����>:���:��;$�%;֟5;��>;�(D;��F;_!H;�H;.�H;��H;��H;��H;��H;L�H;��H;��H;i�H;p�H;I�H;1�H;N�H;2�H;G�H;p�H;h�H;��H;��H;M�H;��H;��H;��H;��H;+�H;�H;[!H;��F;�(D;��>;ҟ5;!�%;��;���:��>:H��z*��+��B>ۻ�X!���]��+�������ۼ�  �|����(�$�      ĸ���v����w�e�c��J�̈́-�{��;缄沼ㄼ��;������j���5���?Q:D��:Pi;�M*;n�8;n�@;�PE;�uG; iH;��H;��H;��H;��H;��H;W�H;��H;��H;��H;��H;��H;��H;�H;��H;��H;��H;��H;��H;��H;[�H;��H; �H;��H;��H;��H;iH;�uG;�PE;d�@;n�8;�M*;Pi;D��:?Q:H�깠5��j��������;�ㄼ�沼�;�{�̈́-��J�f�c���w��v��      yHͽ֪ɽ�;��"����Ƹ����[�z0�r��%<ͼɾ��a�J�����j��s*� ����::b�:=�;��/;�L<;�C;mF;u�G;�H;��H;��H;��H;�H;2�H;��H;�H;�H;��H;��H;��H;��H;��H;��H;��H;�H;�H;��H;6�H;�H;��H;��H;��H;ݡH;o�G;mF;�C;|L<;��/;;�;8b�:���:P�w*��j�����b�J�ʾ��&<ͼr��z0���[�Ƹ����"���;��֪ɽ      ��!-������ѱ�ƽ^P���v���J�H����ۼ��a�J������+��xrѺ�(
9�M�:��;~ $;��5;��?;f�D;D\G;�eH;��H;��H;��H;��H;��H;��H;2�H;U�H;<�H;2�H;A�H;�H;D�H;0�H;:�H;T�H;2�H;��H;�H;��H;��H;��H;��H;�eH;D\G;f�D;��?;��5;~ $;��;�M�:`(
9�rѺ�+������b�J�����ۼH���J��v��^P��ƽұ轃����!-�       j�Vde�Y0X�D�f{+�������u㻽Y���QDX������ۼʾ����;�A>ۻX�P�y��>":���:��;ɷ-;��;;��B;ozF;�H;a�H;X�H;��H;��H;��H;��H;N�H;��H;|�H;p�H;��H;[�H;��H;p�H;{�H;��H;K�H;��H;��H;��H;�H;W�H;^�H;�H;pzF;��B;��;;��-;��;���:�>":L�y�X�D>ۻ��;�ʾ����ۼ���QDX�Y���v㻽��콂��g{+�D�Z0X�Vde�      ��Ph��k���I���|x���O��C(���Ϊɽ����PDX�H��%<ͼㄼ�X!��s���W��uK�%��:�y;�#;�H6;R@;�PE;n�G;]�H;��H;�H;��H;~�H;��H;T�H;��H;��H;��H;��H;��H;��H;��H;��H;��H;R�H;��H;��H;��H;
�H;��H;\�H;i�G;�PE;R@;�H6;��#;�y;��:�uK��W��s���X!�ㄼ&<ͼH��QDX�����Ϊɽ���C(���O��|x��I��k��Ph��      =����������!�;hɰ��G��	 j�7�5��	�ΪɽY����J�r���沼��]�����	x�N	��<n:���:�v;��/;h-=;��C;�F;�HH;|�H;��H;��H;�H;~�H;g�H;��H;��H;��H;��H;�H;��H;��H;��H;��H;i�H;{�H;�H;��H;��H;~�H;�HH;�F;��C;k-=;��/;�v;���:(n:L	���	x������]��沼r���J�Y���Ϊɽ�	�7�5�	 j��G��hɰ�!�;��徶���      �2�U�-�"�-E�����?Kɾj����s�7�5���v㻽�v��z0��;��+���*����/6�@@S�QM�:S�	;t�(;��9;�/B;MDF;H;��H;\�H;��H;��H;M�H;d�H;��H;�H;�H;�H;9�H;�H;�H;�H;��H;c�H;L�H;��H;��H;]�H;��H;%H;JDF;�/B;��9;t�(;L�	;WM�: AS�+6�����*��+���;�	z0��v��v㻽��7�5���s�j��?Kɾ����-E�"�U�-�      %3s�cm�:�\�g�C�5�%����TҾj��	 j��C(����^P����[�{������Y�6��aX�T�<��k::��:�� ;ԟ5;2R@;8uE;ϲG;�H;�H;��H;��H;#�H;G�H;	�H;B�H;L�H;7�H;n�H;6�H;N�H;A�H;�H;G�H; �H;��H;��H;"�H;�H;ղG;6uE;4R@;؟5;�� ;0��:�k:X�<�_X�6����Y����{���[�^P����콪C(�	 j�j���TҾ��5�%�g�C�:�\�cm�      �ޞ�������_F�>�W�W�-���?Kɾ�G����O����ƽƸ��̈́-���ۼㄼ34�ǐ��ζ�4]:���:�;|�1;�c>;D�D;w\G;-sH;x�H;7�H;G�H; �H;N�H;�H;I�H;k�H;]�H;��H;]�H;j�H;H�H;�H;N�H;��H;K�H;8�H;{�H;0sH;�\G;E�D;�c>;|�1;;���:<]:�ζ�ǐ�34�ㄼ��ۼ̈́-�Ƹ��ƽ�����O��G��?Kɾ��W�-�>�W�_F�������      ��ſ���Lw���ޞ�����>�W�5�%�����hɰ��|x�f{+�ѱ����J��  �Ͷ��X�1�&���+�� 
9��:��;߷-;��<;]�C;�G;�TH;$�H;��H;��H;��H;,�H;�H;h�H;��H;x�H;��H;t�H;��H;d�H;�H;.�H;��H;��H;��H;(�H;�TH;�G;]�C;��<;޷-;��;��:� 
9+�$���X�1�Ͷ���  ��J���ѱ�f{+��|x�hɰ�����5�%�>�W������ޞ�Lw�����      ������Կp���ޞ�_F�g�C�-E�!�;�I��D���"��e�c�{��֯���J��ѻɢ)�pK�'��:
�
;�M*;l�:;�C;ƸF;�8H;-�H;H�H;X�H;��H;�H;�H;��H;��H;��H;��H;��H;��H;��H;�H;�H;��H;b�H;M�H;.�H;�8H;ѸF;�C;n�:;�M*;
�
;!��:K�̢)��ѻ��J��֯�|�e�c�"����D��I��!�;-E�g�C�_F��ޞ�p���Կ��      ����������ԿLw�����:�\�"����k��Y0X�����;����w����������]����F�����ɒ:��; �';��9;�oB;�zF;�!H;s�H;��H;�H;r�H;�H;�H;��H;��H;��H;��H;��H;��H;��H;�H;�H;o�H;�H;��H;w�H;�!H;�zF;�oB;��9;��';��;�ɒ:����F��黪�]����������w��;�����Y0X�k�����"�:�\����Lw���Կ��𿝏�      $�������忇�����cm�U�-�����Ph��Vde�!-�֪ɽ�v��'�$�~�ɼymj�6���X����ņ:hx;�%;2�8;CB;RF;�H;�H;�H;��H;H�H;�H;�H;{�H;��H;��H;�H;��H;��H;{�H;�H;�H;C�H;��H;�H;�H; H;-RF;CB;0�8;�%;ex;�ņ:��X�4���ymj�~�ɼ'�$��v��֪ɽ!-�Vde�Ph������U�-�cm��������忝����      dܿ3�ֿ�aǿ=^��/���Yo���7����iþ�(���-=��` �
A���_�/]�.p����I�O�ѻ~�)�`�R���:0�
;�*; �:;��B;�HF;'�G;�lH;�H;v�H;=�H;��H;��H;O�H;�H;�H;��H;	�H;}�H;P�H;��H;��H;<�H;��H;��H;�lH;+�G;IF;��B;�:;�*;.�
;��:�R��)�N�ѻ��I�.p��/]��_�
A���` ��-=��(���iþ����7�Yo�/���=^���aǿ3�ֿ      2�ֿCpѿ�¿������_Xi�Е3��
�UD��Fl��@�9��.���R�� \� �dx��.�E��ͻ�$� �ߍ�:?�;K�*;5�:;�B;�TF;��G;(nH;��H;��H;j�H;��H;��H;]�H;��H;!�H;��H;�H;��H;]�H;��H;��H;g�H;ɷH;��H;)nH;��G;�TF;�B;2�:;E�*;>�;ۍ�:� ��$��ͻ.�E�cx�� �\��R���.��@�9�Fl��UD���
�Е3�_Xi��������¿Cpѿ      �aǿ�¿����������"Y��f'�����6o���.}��k/����%ڟ� <Q�-#�ע��(;�,���2�� e7���:�;s,;��;;�C;�vF;�G;�rH;�H;��H;�H;��H;��H;��H;��H;P�H;��H;G�H;��H;��H;��H;��H;�H;��H;�H;�rH;�G;wF;�C;��;;n,;�;�: ^7�4��,����(;�ע�,#� <Q�%ڟ�����k/��.}�7o�������f'��"Y�����������¿      =^������k���Yo���@�)�#�޾����8ce�0����ڽ󻒽�f@������R���O*�FG������C^92��:;]d.;��<;��C;�F;��G;�yH;��H;�H;�H;��H;k�H;��H;��H;��H;�H;~�H;��H;��H;k�H;��H;�H;!�H;��H;�yH;��G;��F;��C;��<;Vd.;;.��:D^9���EG���O*��R�������f@�󻒽��ڽ/��8ce�����#�޾)���@�Yo�k�������      /����������Yo��!J�K�#��\��VD������zPH�����b��C��� +���ټ'����꿐����l�:(��:G�;�Y1;>;�0D;|�F;aH;C�H;ĨH;�H;Z�H;��H;�H;b�H;J�H;��H;_�H;��H;J�H;c�H;�H;��H;W�H;�H;ĨH;F�H;eH;��F;�0D;>;�Y1;G�;&��:��:
���鿐���'����ټ� +�C���b�����zPH�����VD���\��K�#��!J�Yo��������      Yo�_Xi��"Y���@�K�#��
��о�A���i���(�~��vr��
�_��5��ɺ�n�`��<��_�d�P�\�`�X:�P�:�`;ʱ4;��?;��D;u8G;m0H;��H;k�H;r�H;�H;��H;��H;��H;��H;�H;��H;�H;��H;��H;��H;��H; �H;{�H;m�H;��H;n0H;~8G;��D;��?;Ǳ4;�`;�P�:h�X:P�\�^�d��<��n�`��ɺ��5�
�_�vr��~����(��i��A���о�
�K�#���@��"Y�_Xi�      ��7�Е3��f'�)��\���о�����.}��-=�{
���Ľ[��+:�����������7�GĻ��$��N��ÿ�:�{;�D&;�+8;JA;�E;��G;}LH;�H;v�H;2�H;��H; �H;��H;��H;�H;��H;�H;�H;�H;��H;��H;��H;��H;9�H;x�H;�H;{LH;��G;�E;JA;�+8;�D&;�{;Ͽ�:�N����$�GĻ��7���������*:�[����Ľ{
��-=��.}������о�\��)��f'�Е3�      ���
�����#�޾VD���A���.}�(�D�ht���ڽ�!��\����Z�ļ�
v�;��ƿ���Iɺ S�9���:(;�-;��;;��B;hIF;��G;fH;��H;�H;,�H;��H;f�H;��H;\�H;��H;��H;e�H;��H;��H;]�H;��H;b�H;��H;4�H;�H;��H;fH;��G;jIF;��B;��;;�-;(;���:(S�9�Iɺƿ��:���
v�Y�ļ���\��!����ڽht�(�D��.}��A��VD��#�޾�����
�      �iþUD��6o�����������i��-=�ht�����R��gys�y +����x񗼒(;�'�ѻ�s@�ȅ!�4j:�P�:��;�D3;3�>;FD;��F;�	H;;|H;��H;s�H;3�H;��H;��H;��H;�H;,�H;n�H;��H;k�H;/�H;�H;��H;��H;��H;:�H;t�H;��H;<|H;�	H;��F;FD;5�>;�D3;��;�P�:4j:̅!��s@�&�ѻ�(;�x����y +�gys��R�����ht��-=��i���������6o��UD��      �(��Fl���.}�8ce�zPH���(�{
���ڽ�R����{�B�6�� �,p��\�`�˨��,��>IҺ�L^9���:ޣ;�~(;/�8;�IA;|E;jG;�=H;C�H;լH;�H;\�H;%�H;j�H;��H;��H;��H;��H;I�H;��H;��H;��H;��H;h�H;&�H;d�H; �H;֬H;C�H;�=H;jG;|E;�IA;3�8;�~(;�;���:�L^98IҺ�,��ʨ�\�`�+p��� �B�6���{��R����ڽ{
���(�zPH�8ce��.}�Fl��      �-=�@�9��k/�0�����~��Ľ�!��hys�B�6�$#��ɺ��vz����>^��b�$��~�T�r:��:��;�Y1;�H=;'xC;(wF;�G;�eH;I�H;��H;��H;��H;N�H;��H;��H;��H;c�H;v�H;��H;w�H;d�H;��H;��H;��H;N�H;��H;��H;��H;J�H;�eH;�G;'wF;+xC;I=;�Y1;��;��:X�r:x~�`�$�<^������vz��ɺ�$#�B�6�gys��!����Ľ~���0���k/�@�9�      �` ��.�����ڽ�b��vr��[��\�y +�� ��ɺ�?��O*�Dͻ�5R�ǅ�М:2��:��;�);�t8;d�@;X*E;n8G;>$H;>�H;D�H;�H;!�H;��H;k�H;a�H;�H;M�H;��H;��H;�H;��H;��H;O�H;��H;^�H;m�H;��H;)�H;��H;@�H;?�H;B$H;m8G;^*E;i�@;�t8;�);��;6��:�:ǅ��5R�Aͻ�O*�>��ɺ�� �y +�\�[��vr���b����ڽ��.��      
A���R��%ڟ�󻒽C��
�_�*:�������+p���vz��O*��4ֻ	k�$���`�096�:1;R� ;�D3;H�=;��C;�kF;��G;�\H;��H;O�H; �H;:�H;��H;v�H;��H;��H;�H;��H;T�H;��H;S�H;��H;	�H;��H;��H;x�H;��H;>�H;�H;L�H;��H;�\H;��G;�kF;��C;I�=;�D3;Y� ;1;B�:��09���k��4ֻ�O*��vz�+p����輣��*:�
�_�C��󻒽%ڟ��R��      �_�\� <Q� g@� +��5�����Y�ļx�[�`����Eͻk��Hɺ �6�H�:�P�:-�;�d.;G�:;%�A;*|E;xNG;F'H;��H;ǥH;^�H;��H;#�H;J�H;Y�H;3�H;��H;��H;�H;��H;��H;��H;	�H;��H;��H;0�H;\�H;T�H;*�H;��H;]�H;ƥH;�H;F'H;~NG;.|E;%�A;Q�:;�d.;,�;�P�:J�: �6��Hɺk�Bͻ���[�`�w�X�ļ�����5�� +� g@� <Q�\�      .]� �,#�������ټ�ɺ������
v��(;�˨�<^���5R�&��� �6����:���:��;,�*;�+8;�!@;Y�D;c�F;��G;�eH;�H;��H;��H;��H;��H;��H;�H;s�H;��H;b�H;x�H;)�H;V�H;(�H;w�H;d�H;��H;o�H;!�H;��H;��H;��H;��H;��H;��H;�eH;��G;g�F;\�D;�!@;�+8;'�*;��;���:���: �6�����5R�8^��ʨ��(;��
v������ɺ���ټ����-#� �      +p��cx��ע��R��'��o�`���7�9��'�ѻ�,��]�$�ǅ�`�09H�:���:�;�~(;�Z6;��>;̨C;�HF;ܠG;�DH;I�H;��H;��H;�H;)�H;�H;��H;��H;��H;��H;�H;��H;��H;��H;�H;��H;�H;��H;��H;��H;��H;�H;-�H;�H;��H;��H;I�H;�DH;�G;�HF;ըC;��>;�Z6;�~(;�;���:J�:��09�ƅ�Z�$��,��$�ѻ8����7�l�`�(���R��ע�bx��      �I�+�E��(;��O*����<��GĻÿ���s@�,IҺ`~�Ԝ:B�:�P�:��;�~(;�5;�>;:C;1�E;zcG;;$H;�{H;:�H;�H;��H;��H;;�H;��H;�H;V�H;��H;O�H;��H;@�H;��H;��H;��H;=�H;��H;L�H;��H;X�H;!�H;��H;=�H;��H;��H;�H;;�H;�{H;?$H;~cG;9�E;;C;�>;�5;�~(;�;�P�:D�:�:@~�(IҺ�s@�¿��GĻ�<�����O*��(;�)�E�      A�ѻ�ͻ*���@G��忐�]�d���$��Iɺą!��L^9`�r:(��:
1;,�;'�*;�Z6;�>;?�B;��E;�8G;�	H; nH;�H;I�H;��H;d�H;��H;��H;H�H;��H;��H;v�H;��H;��H;��H;�H;"�H;�H;��H;��H;��H;r�H;��H;�H;I�H;��H;��H;b�H;��H;J�H;�H;nH;�	H;�8G;��E;<�B;�>;�Z6;*�*;,�;1;2��:t�r: M^9��!��Iɺ��$�X�d�ῐ�BG��&����ͻ      e�)�#�$�2�� �������\��N��HS�9,4j:���:��:��;X� ;�d.;�+8;��>;:C;��E;�)G;��G;dH;��H;��H;_�H;��H;5�H;��H;��H;��H;��H;��H;I�H;{�H;`�H;��H;7�H;K�H;4�H;��H;_�H;x�H;F�H;��H;��H;��H;��H;��H;6�H;��H;b�H;��H;��H;dH;��G;�)G;��E;>C;��>;�+8;�d.;[� ;��;��:���:84j:HS�9�N��(�\�
������2��#�$�       �R�@ � V7�E^9l�:p�X:㿙:���:�P�:�;��;�);�D3;N�:;�!@;ӨC;8�E;�8G;��G;�`H;o�H;�H;�H;{�H;:�H;2�H;M�H;^�H;��H;��H;��H;�H;��H;��H;-�H;n�H;d�H;j�H;-�H;��H;��H;	�H;��H;��H;��H;b�H;M�H;3�H;A�H;|�H;�H;�H;v�H;�`H;��G;�8G;8�E;ըC;�!@;N�:;�D3;�);��;�;�P�:���:ۿ�:��X:��: D^9 ^7�� �      ��:���:��:��:��:�P�:�{;(;��;�~(;�Y1;�t8;F�=;$�A;[�D;�HF;{cG;�	H;dH;n�H;H�H;ֶH;3�H;��H;��H;;�H;I�H;��H;#�H;��H;~�H;��H;U�H;��H;H�H;��H;��H;��H;I�H;��H;T�H;��H;��H;��H;!�H;��H;G�H;;�H;��H;��H;0�H;ٶH;O�H;r�H;dH;�	H;~cG;�HF;]�D;#�A;I�=;�t8;�Y1;�~(;��;(;�{;�P�:(��: ��:��:���:      0�
;N�;�;;E�;�`;�D&;�-;�D3;6�8;	I=;f�@;��C;0|E;g�F;�G;A$H;nH;��H;�H;ٶH;��H;9�H; �H;i�H;��H;��H;u�H;j�H;�H; �H;��H;��H;!�H;g�H;��H;��H;��H;d�H;!�H;��H;��H;!�H;�H;j�H;v�H;��H;��H;m�H; �H;6�H;��H;߶H;�H;��H;nH;D$H;�G;k�F;-|E;��C;k�@;
I=;3�8;�D3;�-;�D&;�`;\�;;��;B�;      �*;N�*;o,;nd.;�Y1;ֱ4;�+8;��;;>�>;�IA;4xC;a*E;�kF;�NG;��G;�DH;�{H;�H;��H;�H;2�H;7�H;��H;��H;��H;_�H;
�H;��H;��H;��H;��H;p�H;��H;=�H;��H;��H;��H;��H;��H;>�H;��H;k�H;��H;��H;��H;��H;�H;b�H;��H;��H;��H;=�H;7�H;�H;��H;�H;�{H;�DH;��G;�NG;�kF;e*E;7xC;�IA;>�>;��;;�+8;ѱ4;�Y1;ld.;o,;7�*;      �:;?�:;��;;��<;>;��?;JA;��B;FD;|E;'wF;m8G;��G;G'H;�eH;M�H;<�H;N�H;b�H;x�H;��H;�H;��H;��H;�H;��H;��H;4�H;w�H;q�H;�H;��H;�H;^�H;��H;��H;��H;��H;}�H;`�H;�H;��H;�H;p�H;u�H;7�H;��H;��H;�H;��H;��H;�H;��H;y�H;`�H;J�H;>�H;O�H;�eH;F'H;��G;p8G;.wF;|E;FD;��B;JA;��?;>;��<;��;;4�:;      գB;�B;�C;��C;�0D;��D;��E;lIF;��F;jG;&�G;F$H;�\H;
�H;��H;��H;'�H;��H;��H;F�H;��H;m�H;��H;!�H;��H;q�H;��H;E�H;+�H;��H;��H;��H;/�H;t�H;��H;��H;��H;��H;��H;u�H;-�H;��H;��H;��H;(�H;E�H;��H;v�H;��H; �H;��H;r�H;��H;C�H;��H;��H;+�H;¨H;��H;�H;�\H;L$H;'�G;jG;��F;lIF; �E;��D;�0D;��C;�C;�B;      �HF;�TF;wF;�F;v�F;�8G;��G;��G;�	H;�=H;fH;E�H;��H;ϥH;��H;��H;��H;g�H;6�H;2�H;@�H;��H;^�H;��H;p�H;��H;#�H;�H;��H;F�H;��H;#�H;6�H;r�H;��H;��H;��H;��H;��H;r�H;6�H;�H;��H;D�H;��H;�H;"�H;��H;t�H;��H;^�H;��H;A�H;2�H;7�H;e�H;��H;��H;��H;˥H;��H;F�H;fH;�=H;�	H;��G;��G;w8G;��F;��F;wF;�TF;      <�G;��G;�G;��G;[H;p0H;�LH;fH;8|H;C�H;J�H;@�H;L�H;`�H;��H;�H;��H;��H;��H;O�H;O�H;��H;
�H;��H;��H;"�H;��H;��H;Q�H;��H;��H;2�H;O�H;u�H;��H;��H;��H;��H;��H;v�H;R�H;/�H;��H;��H;N�H;��H;��H;)�H;��H;��H;�H;��H;R�H;M�H;��H;��H;��H;�H;��H;]�H;L�H;D�H;M�H;B�H;8|H;fH;�LH;i0H;rH;��G;�G;��G;      �lH;-nH;�rH;�yH;<�H;��H;��H;��H;��H;ܬH;��H;��H; �H;��H;��H;-�H;>�H;��H;��H;`�H;��H;r�H;��H;7�H;A�H;�H;��H;6�H;��H;��H;�H;=�H;`�H;e�H;�H;��H;��H;��H;}�H;g�H;`�H;7�H;�H;��H;��H;3�H;��H;�H;E�H;6�H;��H;u�H;��H;^�H;��H;��H;@�H;0�H;��H;��H; �H;��H;��H;ݬH;��H;��H;��H;��H;I�H;�yH;�rH;nH;      �H;��H;�H;��H;��H;m�H;�H;�H;l�H;�H;��H;(�H;>�H;*�H;��H;�H;��H;P�H;��H;��H;+�H;i�H;��H;w�H;'�H;��H;H�H;��H;��H;�H;*�H;L�H;`�H;e�H;d�H;o�H;m�H;j�H;c�H;g�H;a�H;H�H;,�H;�H;��H;��H;G�H;��H;*�H;s�H;��H;i�H;*�H;��H;��H;N�H;��H;�H;��H;)�H;=�H;&�H;��H;!�H;p�H;�H;}�H;f�H;ĨH;��H;�H;��H;      |�H;��H;��H;�H;�H;r�H;5�H;.�H;7�H;b�H;��H;��H;��H;U�H;��H;��H;&�H;�H;��H;��H;��H;�H;��H;p�H;��H;<�H;��H;��H;�H;"�H;@�H;D�H;O�H;d�H;N�H;\�H;q�H;Y�H;I�H;c�H;P�H;@�H;@�H;!�H;�H;��H;��H;C�H;��H;m�H;��H;�H;��H;��H;��H;�H;'�H;�H;��H;Q�H;��H;��H;��H;f�H;9�H;0�H;8�H;q�H;�H;�H;��H;��H;      D�H;��H;�H;&�H;X�H;�H;��H;��H;��H;,�H;U�H;x�H;�H;c�H;(�H;��H;b�H;��H;��H;��H;��H;$�H;��H;�H;��H;��H;��H;�H;/�H;E�H;V�H;O�H;>�H;@�H;a�H;O�H;/�H;I�H;]�H;@�H;@�H;N�H;V�H;B�H;,�H;
�H;��H;��H;��H;�H;��H;$�H;��H;��H;��H;��H;e�H;��H;'�H;a�H;��H;x�H;W�H;-�H;��H;��H;��H;��H;e�H;%�H;�H;��H;      ��H;��H;��H;��H;��H;��H;�H;i�H;��H;j�H;��H;g�H;��H;>�H;w�H;��H;��H;}�H;Q�H;�H;��H;��H;n�H;��H;��H;�H;,�H;=�H;K�H;E�H;I�H;V�H;;�H;9�H;K�H;,�H;%�H;,�H;G�H;9�H;@�H;V�H;H�H;D�H;H�H;:�H;-�H;�H;��H;��H;u�H;��H;��H;�H;P�H;�H;��H;��H;v�H;:�H;��H;g�H;��H;m�H;��H;j�H;�H;��H;��H;��H;��H;��H;      ��H;��H;�H;n�H;�H;��H;��H;��H;��H;��H;��H;�H;�H;��H;��H;��H;X�H;�H;��H;��H;b�H;��H;��H;�H;/�H;2�H;O�H;g�H;e�H;U�H;;�H;@�H;D�H;>�H;�H;�H;L�H;�H;�H;>�H;D�H;@�H;:�H;O�H;a�H;c�H;P�H;4�H;2�H;�H;��H;��H;_�H;��H;��H;�H;Z�H;��H;��H;��H;�H;�H;��H;��H;��H;��H;��H;��H;�H;i�H;�H;��H;      I�H;[�H;��H;��H;f�H;��H;��H;^�H;�H;��H;��H;Y�H;�H;��H;n�H;�H;��H;�H;g�H;��H;��H;#�H;9�H;Y�H;r�H;m�H;q�H;g�H;e�H;g�H;:�H;;�H;>�H;)�H;�H;�H;&�H;�H;�H;)�H;A�H;:�H;:�H;c�H;c�H;c�H;r�H;o�H;u�H;W�H;A�H;"�H;��H;��H;f�H;�H;��H;�H;l�H;��H;�H;V�H;��H;��H;�H;^�H;��H;��H;o�H;��H;��H;e�H;      {�H;��H;��H;��H;Z�H;��H;$�H;��H;5�H;��H;o�H;��H;��H;�H;��H;��H;J�H;��H;�H;6�H;P�H;d�H;��H;t�H;��H;��H;��H;�H;e�H;P�H;Y�H;N�H;�H;�H;#�H;�H;��H;�H;!�H;�H;"�H;O�H;W�H;I�H;a�H;{�H;��H;��H;��H;u�H;��H;d�H;K�H;/�H; �H;��H;N�H;��H;��H;�H;��H;��H;r�H;��H;7�H;��H;+�H;��H;Z�H;��H;��H;��H;      	�H;$�H;N�H;��H;��H;�H;��H;��H;n�H;��H;��H;��H;\�H;��H;0�H;��H;��H;	�H;;�H;o�H;��H;��H;��H;��H;��H;��H;��H;��H;q�H;`�H;K�H;2�H;!�H;�H;�H;�H;�H;�H;�H;"�H;#�H;2�H;I�H;Z�H;m�H;��H;��H;��H;��H;��H;��H;��H;��H;k�H;:�H;�H;��H;��H;/�H;��H;Z�H;��H;��H;��H;q�H;��H;��H;	�H;��H;�H;L�H;/�H;      ��H;��H;��H;�H;]�H;��H;�H;m�H;��H;M�H;��H;+�H;��H;	�H;d�H;��H;��H;,�H;R�H;o�H;��H;��H;��H;��H;��H;��H;��H;��H;q�H;y�H;,�H;*�H;P�H;%�H;��H;�H; �H;�H;��H;&�H;U�H;,�H;,�H;t�H;m�H;��H;��H;��H;��H;��H;��H;��H;��H;h�H;R�H;-�H;��H;��H;c�H;	�H;��H;+�H;��H;O�H;��H;m�H;#�H;��H;`�H;�H;��H;��H;      	�H;&�H;J�H;��H;��H;�H;��H;��H;n�H;��H;~�H;��H;\�H;��H;0�H;��H;��H;�H;;�H;o�H;��H;��H;��H;��H;��H;��H;��H;��H;r�H;^�H;K�H;3�H;"�H;�H;�H;�H;�H;�H;�H;!�H;#�H;2�H;I�H;Z�H;m�H;��H;��H;��H;��H;��H;��H;��H;��H;k�H;:�H;�H;��H;��H;0�H;��H;Z�H;��H;��H;��H;o�H;��H;��H;	�H;��H;��H;P�H;-�H;      o�H;��H;��H;��H;[�H;��H;&�H;��H;3�H;��H;n�H;��H;��H;�H;��H;��H;J�H;��H;�H;6�H;R�H;h�H;��H;u�H;��H;��H;��H;�H;e�H;O�H;W�H;N�H;!�H;�H;%�H;�H;��H;�H;"�H;�H;#�H;N�H;W�H;I�H;a�H;{�H;��H;��H;��H;r�H;��H;e�H;K�H;0�H;�H;��H;M�H;��H;��H;�H;��H;��H;o�H;��H;5�H;��H;+�H;��H;`�H;��H;��H;��H;      J�H;[�H;��H;��H;h�H;��H;��H;a�H;�H;��H;��H;V�H;�H;��H;o�H;�H;��H;�H;i�H;��H;��H;&�H;=�H;]�H;v�H;m�H;r�H;g�H;g�H;g�H;:�H;;�H;>�H;)�H;�H;�H;&�H;�H;�H;)�H;A�H;;�H;9�H;c�H;a�H;d�H;r�H;o�H;r�H;U�H;A�H;%�H;��H;��H;g�H;�H;��H;�H;n�H;��H;�H;V�H;��H;��H;�H;c�H;��H;��H;o�H;��H;��H;]�H;      ��H;��H;�H;k�H;�H;��H;��H;��H;��H;��H;��H;�H;�H;�H;��H;��H;X�H;�H;��H;��H;b�H;��H;��H;�H;3�H;/�H;O�H;e�H;g�H;U�H;:�H;=�H;B�H;>�H;�H;�H;L�H;�H;�H;@�H;D�H;A�H;:�H;P�H;`�H;a�H;P�H;4�H;/�H;�H;��H;��H;[�H;��H;��H;�H;X�H;��H;��H;�H;�H;�H;��H;��H;��H;��H;��H;��H;�H;r�H;�H;��H;      |�H;��H;��H;��H;��H;��H;	�H;g�H;��H;j�H;��H;g�H;��H;:�H;z�H;��H;��H;�H;P�H;�H;��H;��H;p�H;��H;��H;�H;,�H;=�H;N�H;D�H;G�H;V�H;;�H;9�H;L�H;,�H;%�H;/�H;H�H;9�H;@�H;V�H;G�H;B�H;H�H;:�H;,�H;!�H;��H;��H;w�H;��H;��H;�H;P�H;}�H;��H;��H;w�H;;�H;��H;g�H;��H;l�H;��H;g�H;�H;��H;��H;��H;��H;��H;      :�H;��H;�H;"�H;_�H;�H;��H;��H;��H;,�H;W�H;x�H;��H;e�H;*�H;��H;d�H;��H;��H;��H;��H;&�H;��H;�H;��H;��H;��H;
�H;0�H;E�H;U�H;O�H;>�H;A�H;c�H;N�H;/�H;O�H;^�H;B�H;A�H;O�H;U�H;B�H;*�H;�H;��H;��H;��H;�H;��H;&�H;��H;��H;��H;��H;g�H;��H;(�H;c�H;�H;x�H;U�H;,�H;��H;��H;��H; �H;l�H;,�H;�H;��H;      ��H;��H;��H; �H;�H;~�H;8�H;7�H;;�H;d�H;��H;��H;��H;T�H;��H;��H;&�H;�H;��H;��H;��H;
�H;��H;o�H;��H;=�H;��H;��H;�H;#�H;@�H;B�H;L�H;d�H;N�H;Z�H;q�H;\�H;K�H;d�H;R�H;D�H;@�H;!�H;�H;��H;��H;C�H;��H;j�H;��H;�H;��H;��H;��H;�H;&�H; �H;��H;T�H;��H;��H;��H;d�H;7�H;4�H;9�H;n�H;�H;$�H;��H;��H;       �H;��H;-�H;��H;��H;t�H;}�H;�H;t�H;�H;��H;(�H;@�H;,�H;��H;�H;��H;S�H;��H;��H;.�H;k�H;��H;y�H;*�H;��H;H�H;��H;��H;�H;)�H;L�H;`�H;e�H;d�H;n�H;m�H;n�H;c�H;e�H;a�H;K�H;*�H;�H;��H;��H;J�H;��H;'�H;p�H;��H;j�H;*�H;��H;��H;N�H;��H;�H;��H;)�H;>�H;%�H;��H;�H;q�H;�H;��H;m�H;��H;��H;-�H;��H;      �lH;!nH;�rH;�yH;8�H;��H;��H;��H;��H;߬H;��H;��H;�H;��H;��H;/�H;@�H;��H;��H;`�H;��H;v�H;��H;:�H;E�H;�H;��H;3�H;��H;��H;	�H;:�H;]�H;e�H;�H;��H;��H;��H;}�H;g�H;c�H;;�H;	�H;��H;��H;2�H;��H;	�H;A�H;3�H;��H;s�H;��H;^�H;��H;��H;@�H;/�H;��H;��H;�H;��H;��H;ݬH;��H;��H;��H;��H;F�H;�yH;�rH;!nH;      /�G;��G;�G;��G;iH;t0H;�LH;#fH;<|H;E�H;M�H;E�H;K�H;^�H;��H;�H;��H;��H;��H;O�H;R�H;��H;�H;��H;��H;"�H;��H;��H;Q�H;��H;��H;2�H;N�H;u�H;��H;��H;��H;��H;��H;v�H;P�H;3�H;��H;��H;M�H;��H;��H;)�H;��H;��H;�H;��H;N�H;P�H;��H;��H;��H;�H;��H;]�H;L�H;D�H;L�H;C�H;:|H;%fH;�LH;m0H;rH;��G;�G;��G;      �HF;�TF;wF;�F;�F;�8G;��G;��G;�	H;�=H;fH;I�H;��H;ͥH;��H;��H;��H;k�H;7�H;2�H;D�H;��H;\�H;��H;v�H;��H;"�H;�H;��H;D�H;��H;#�H;4�H;r�H;��H;��H;��H;��H;��H;r�H;6�H;#�H;��H;F�H;��H;�H;#�H;��H;q�H;��H;_�H;��H;@�H;2�H;7�H;b�H;��H;��H;��H;ʥH;��H;E�H;fH;�=H;�	H;��G;��G;w8G;��F;�F;�vF;�TF;      УB;�B;�C;��C;�0D;��D; �E;oIF;��F;jG;&�G;N$H;�\H;�H;��H;ŨH;(�H;��H;��H;E�H;��H;q�H;��H;#�H;��H;o�H;��H;F�H;+�H;��H;��H;��H;,�H;u�H;��H;��H;��H;��H;��H;v�H;-�H;��H;��H;��H;(�H;B�H;��H;t�H;��H;�H;��H;p�H;��H;C�H;��H;��H;)�H;��H;��H;�H;�\H;H$H;$�G;jG;��F;jIF;��E;��D;�0D;��C;�C;�B;      ��:;&�:;|�;;	�<;�>;ɧ?;JA;��B;FD;|E;,wF;r8G;��G;F'H;�eH;R�H;>�H;Q�H;b�H;{�H;��H;�H;��H;��H;�H;��H;��H;7�H;w�H;o�H;�H;��H;�H;^�H;�H;��H;��H;��H;|�H;^�H;�H;��H;�H;q�H;w�H;4�H;��H;��H;�H;��H;��H;�H;��H;{�H;b�H;L�H;>�H;P�H;�eH;F'H;��G;n8G;+wF;|E;FD;��B;JA;��?;>;!�<;{�;;�:;      �*;D�*;d,;vd.;�Y1;α4;�+8;��;;D�>;�IA;0xC;c*E;�kF;�NG;��G;�DH;�{H;#�H;��H;�H;6�H;:�H;��H;��H;��H;\�H;�H;��H;��H;��H;��H;q�H;��H;=�H;��H;��H;��H;��H;��H;;�H;��H;q�H;��H;��H;��H;��H;�H;_�H;��H;��H;��H;9�H;5�H;�H;��H;�H;�{H;�DH;��G;�NG;�kF;a*E;1xC;�IA;A�>;��;;�+8;̱4;�Y1;vd.;d,;-�*;      .�
;N�;��;;J�;�`;�D&;�-;�D3;3�8;
I=;n�@;��C;.|E;k�F;�G;D$H;	nH;��H;�H;߶H;��H;7�H;!�H;p�H;��H;��H;w�H;k�H;�H; �H;��H;��H;!�H;d�H;��H;��H;��H;a�H;�H;��H;��H;#�H;�H;j�H;u�H;��H;��H;j�H;!�H;9�H;��H;ܶH;�H;��H;nH;B$H;�G;j�F;-|E;��C;i�@;	I=;0�8;�D3;�-;�D&;�`;]�;;��;F�;      ��:���:��:2��:��:�P�:�{;(;��;�~(;�Y1;�t8;K�=;$�A;`�D;�HF;~cG;�	H;dH;r�H;L�H;ڶH;2�H;��H;��H;9�H;G�H;��H;$�H;��H;��H;��H;T�H;��H;I�H;��H;��H;��H;G�H;��H;T�H;��H;��H;��H;!�H;��H;I�H;:�H;��H;��H;2�H;ֶH;L�H;q�H;dH;�	H;}cG;�HF;]�D;#�A;I�=;�t8;�Y1;�~(;��;(;�{;�P�:6��:,��:�:Ս�:      ��R�  � ^7�PE^9x�:��X:忙:���:�P�:�;��;�);�D3;N�:;�!@;רC;9�E;�8G;��G;�`H;v�H;�H;�H;|�H;B�H;0�H;J�H;`�H;��H;��H;��H;�H;��H;��H;/�H;j�H;d�H;k�H;,�H;��H;��H;�H;��H;��H;��H;^�H;M�H;0�H;<�H;�H;�H;�H;r�H;�`H;��G;�8G;9�E;֨C;�!@;L�:;�D3;�);��;�;�P�:���:ۿ�:h�X:��:�D^9 \7�0 �      d�)�!�$�4����������\��N��XS�9@4j:���:��:��;[� ;�d.;�+8;��>;=C;��E;�)G;��G;dH;��H;��H;`�H;��H;3�H;��H;��H;��H;��H;��H;I�H;{�H;`�H;��H;6�H;K�H;6�H;��H;`�H;{�H;I�H;��H;��H;��H;��H;��H;3�H;��H;b�H;��H;��H;dH;��G;�)G;��E;;C;��>;�+8;�d.;X� ;��;��:���:84j:`S�9�N��(�\��������9���$�      H�ѻ�ͻ.���>G��㿐�R�d���$��Iɺ��!��L^9h�r:2��:1;+�;,�*;�Z6;�>;?�B;��E;�8G;�	H;nH;�H;J�H;��H;d�H;��H;��H;I�H;��H;��H;v�H;��H;��H;��H;�H;"�H;�H;��H;��H;��H;v�H;��H;�H;I�H;��H;��H;a�H;��H;I�H;�H;nH;�	H;�8G;��E;<�B;�>;�Z6;*�*;)�;
1;,��:p�r:�L^9��!��Iɺ��$�[�d�㿐�AG��1����ͻ      �I�+�E��(;��O*����<��GĻ�����s@�(IҺP~��:D�:�P�:�;�~(;�5;�>;;C;5�E;�cG;>$H;�{H;:�H;!�H;��H;��H;9�H;��H;�H;X�H;��H;O�H;��H;A�H;��H;��H;��H;=�H;��H;L�H;��H;Z�H;�H;��H;:�H;��H;��H;�H;:�H;�{H;;$H;zcG;8�E;:C;�>;�5;�~(;�;�P�:B�:��:P~�.IҺ�s@�¿��GĻ�<�����O*��(;�*�E�      +p��bx��ע��R��'��l�`���7�8��&�ѻ�,��[�$��ƅ���09H�:���:�;�~(;�Z6;��>;ӨC;�HF;�G;�DH;K�H;��H;��H;�H;)�H;�H;��H;��H;��H;��H;�H;��H;�H;��H;�H;��H;�H;��H;��H;��H;��H;�H;*�H;�H;��H;��H;I�H;�DH;ޠG;�HF;ӨC;��>;�Z6;�~(;�;���:H�:`�09ǅ�\�$��,��&�ѻ8����7�l�`�(���R��ע�cx��      .]� �-#�������ټ�ɺ������
v��(;�ʨ�:^���5R���� �6����:���:��;)�*;�+8;�!@;`�D;g�F;��G;�eH;��H;��H;��H;��H;��H;��H;!�H;r�H;��H;e�H;z�H;'�H;V�H;(�H;w�H;e�H;��H;p�H; �H;��H;��H;��H;��H;��H;��H;�eH;��G;e�F;V�D;�!@;�+8;$�*;��;���:���: �6�&����5R�;^��˨��(;��
v������ɺ���ټ����-#� �      �_�\� <Q��f@� +��5�����X�ļw�[�`����@ͻk��Hɺ |6�R�:�P�:,�;�d.;L�:;+�A;-|E;�NG;G'H;�H;ʥH;]�H;��H;)�H;M�H;\�H;3�H;��H;��H;�H;��H;��H;��H;�H;��H;��H;2�H;Y�H;O�H;(�H;��H;[�H;ĥH;��H;G'H;�NG;)|E; �A;N�:;�d.;+�;�P�:H�: �6��Hɺk�Bͻ���\�`�w�X�ļ�����5�� +� g@� <Q�\�      
A���R��%ڟ�󻒽C��
�_�*:�������+p���vz��O*��4ֻk������09>�:1;V� ;�D3;O�=;��C;�kF;��G;�\H;��H;L�H; �H;>�H;��H;x�H;��H;��H;	�H;��H;S�H;��H;S�H;��H;�H;��H;��H;w�H;��H;>�H; �H;K�H;��H;�\H;��G;�kF;��C;E�=;�D3;T� ;
1;:�:`�09 ���k��4ֻ�O*��vz�+p����輣��*:�
�_�C��󻒽%ڟ��R��      �` ��.�����ڽ�b��vr��[��\�y +�� ��ɺ�>��O*�Bͻ�5R� ǅ���:,��:��;�);u8;i�@;a*E;p8G;D$H;B�H;A�H;�H;#�H;��H;o�H;`�H;�H;N�H;��H;��H;�H;��H;��H;N�H; �H;`�H;m�H;��H;&�H;�H;@�H;?�H;?$H;n8G;a*E;f�@;�t8;�);��;,��:ܜ:ǅ��5R�Cͻ�O*�>��ɺ�� �y +�\�[��vr���b����ڽ��.��      �-=�@�9��k/�0�����~��Ľ�!��hys�B�6�$#��ɺ��vz����:^��`�$��~�L�r:	��:��;�Y1;I=;0xC;)wF;�G; fH;H�H;��H;��H;��H;Q�H;��H;��H;��H;a�H;v�H;��H;v�H;a�H;��H;��H;��H;N�H;��H;��H;��H;H�H;�eH;�G;(wF;-xC;�H=;�Y1;��;��:L�r:�~�b�$�>^������vz��ɺ�$#�B�6�hys��!����Ľ~���0���k/�@�9�      �(��Fl���.}�8ce�zPH���(�{
���ڽ�R����{�B�6�� �+p��\�`�ʨ��,��6IҺ�L^9���:�;�~(;2�8;�IA;|E;jG;�=H;B�H;լH;�H;_�H;&�H;i�H;��H;��H;��H;��H;I�H;��H;��H;��H;��H;h�H;&�H;b�H; �H;֬H;B�H;�=H;jG;|E;�IA;/�8;�~(;�;���:pL^98IҺ�,��˨�\�`�,p��� �B�6���{��R����ڽ{
���(�zPH�8ce��.}�Fl��      �iþUD��6o�����������i��-=�ht�����R��gys�y +����x񗼒(;�&�ѻ�s@�̅!�$4j:�P�:��;�D3;7�>;FD;��F;�	H;;|H;��H;t�H;4�H;��H;��H;��H;�H;+�H;j�H;��H;j�H;,�H;�H;��H;��H;��H;6�H;t�H;��H;<|H;�	H;��F;FD;8�>;�D3;��;�P�:4j:̅!��s@�&�ѻ�(;�x����y +�hys��R�����ht��-=��i���������6o��UD��      ���
�����#�޾VD���A���.}�(�D�ht���ڽ�!��\����Z�ļ�
v�:��ƿ���Iɺ(S�9���: (;�-;��;;��B;jIF;��G;fH;��H;�H;,�H;��H;f�H;��H;\�H;��H;��H;e�H;��H;��H;Y�H;��H;c�H;��H;3�H;�H;��H;fH;��G;hIF;��B;��;;�-;(;���:S�9�Iɺƿ��;���
v�Y�ļ���\��!����ڽht�(�D��.}��A��VD��#�޾�����
�      ��7�Е3��f'�)��\���о�����.}��-=�{
���Ľ[��*:�����������7�GĻ��$��N��ɿ�:�{;�D&;�+8;JA;�E;��G;zLH;�H;x�H;2�H;��H; �H;��H;��H;�H;�H;�H;~�H;�H;��H;��H; �H;��H;8�H;x�H;�H;}LH;��G;�E;JA;�+8;�D&;�{;ѿ�: O����$�GĻ��7���������+:�[����Ľ{
��-=��.}������о�\��)��f'�Е3�      Yo�_Xi��"Y���@�K�#��
��о�A���i���(�~��vr��
�_��5��ɺ�n�`��<��a�d�P�\�h�X:�P�:�`;ȱ4;��?;��D;t8G;k0H;��H;m�H;w�H;�H;��H;��H;��H;��H;�H;��H;�H;��H;��H;��H;��H; �H;z�H;n�H;��H;p0H;~8G;��D;��?;ʱ4;�`;�P�:p�X:T�\�a�d��<��n�`��ɺ��5�
�_�vr��~����(��i��A���о�
�K�#���@��"Y�_Xi�      /����������Yo��!J�K�#��\��VD������zPH�����b��C��� +���ټ'����뿐����|�:,��:G�;�Y1;	>;�0D;y�F;`H;C�H;¨H;�H;Z�H;��H;�H;e�H;E�H;��H;]�H;��H;F�H;a�H;	�H;��H;X�H;�H;ŨH;F�H;hH;��F;�0D;	>;�Y1;G�;&��:��:
���运���'����ټ� +�C���b�����zPH�����VD���\��K�#��!J�Yo��������      =^������k���Yo���@�)�#�޾����8ce�0����ڽ󻒽�f@������R���O*�FG������C^94��:;Zd.;��<;��C;�F;��G;�yH;��H;�H; �H;��H;k�H;��H;��H;��H;�H;�H;��H;��H;l�H;��H;�H;"�H;��H;�yH;��G;��F;��C;��<;Yd.;;.��:@D^9���DG���O*��R�������f@�󻒽��ڽ/��8ce�����#�޾)���@�Yo�k�������      �aǿ�¿����������"Y��f'�����6o���.}��k/����%ڟ� <Q�,#�ע��(;�,���2�� d7��:�;q,;��;;�C;�vF;�G;�rH;�H;��H;�H;��H;��H;��H;��H;M�H;��H;I�H;��H;��H;��H;��H;�H;��H;�H;�rH;�G;wF;�C;��;;l,;�;�: ]7�4��,����(;�ע�,#� <Q�%ڟ�����k/��.}�6o�������f'��"Y�����������¿      3�ֿCpѿ�¿������_Xi�Е3��
�UD��Fl��@�9��.���R�� \� �dx��.�E��ͻ�$� �㍨:?�;K�*;5�:;�B;�TF;��G;(nH;��H;��H;j�H;��H;��H;]�H;��H; �H;��H;�H;��H;]�H;��H;��H;g�H;ɷH;��H;)nH;��G;�TF;�B;4�:;E�*;<�;ۍ�:� ��$��ͻ/�E�cx�� �\��R���.��@�9�Fl��UD���
�Е3�_Xi��������¿Cpѿ      �?��|h��=v��� ��7�X��O/�/y�@�;ఖ��+X��� �ѽ����^n;�Z�������B(�ؚ��N����e9"�:�;�Y.;T�<;eWC;�ZF;��G;0H;3jH;7�H;F�H;��H;)�H;��H;Z�H;��H;��H;��H;V�H;��H;(�H;�H;C�H;B�H;4jH;0H;��G;�ZF;bWC;S�<;�Y.;�;�:Пe9P��֚���B(�����Z��^n;����� �ѽ���+X�ఖ�@�;/y��O/�7�X�� ��=v��|h��      |h��/���a�����y�VvS�pM+��v�9ɾ�����T� ]�\ν����x\8�����x��%�L���l��h�9u-�:j�;��.;�<;�nC;�dF;�G;�1H;�jH;��H;��H;˵H;j�H;��H;e�H;��H;��H;��H;g�H;��H;i�H;˵H;��H;��H;�jH;�1H;�G;�dF;�nC;�<;��.;g�;o-�:��9l��J���%��x�����x\8�����\ν ]��T�����9ɾ�v�pM+�VvS���y�a���/���      =v��b���W ��`�h�6E�W��i���|㼾}���nH�ӈ�x�ý�Ȅ��s/��o��#�����!J�� к`	�9\g�:�l;$0;]=;ٲC;րF;n�G;6H;mH;%�H;��H;~�H;��H;@�H;��H;�H;��H; �H;��H;@�H;��H;�H;��H;/�H; mH;6H;t�G;�F;ٲC;]=;0;�l;\g�:�	�9$к!J������#���o��s/��Ȅ�x�ýӈ��nH�}��|㼾i���W��6E�`�h�W ��a���      � ����y�`�h���N��O/����B�߾B���*|��6�p}�䳽hSt�;�!�nrμ?F{��_��X��ē��L:0��:�Z;�2;�O>;mD;'�F;y�G;=H;�pH;��H;G�H;˷H;��H;��H;\�H;}�H;_�H;v�H;^�H;��H;��H;̷H;D�H;��H;�pH;=H;}�G;3�F;lD;�O>;�2;�Z;.��:h:ē���X���_�?F{�nrμ;�!�hSt�䳽p}��6��*|�B��B�߾����O/���N�`�h���y�      7�X�VvS�6E��O/��S�GW����������LS\��� ���9����Y�z��σ����]������b���Y�H�Y:��:f`;9�4;�?;9�D;��F;�G;FH;DuH;��H;��H;��H;�H;��H;�H;�H;��H;�H;�H;��H;�H;��H;��H;ƓH;GuH;FH;�G;��F;9�D;�?;5�4;f`;��:X�Y:��Y��b�������]�σ��z���Y�9����彑� �LS\���������GW���S��O/�6E�VvS�      �O/�pM+�W�����GW��9ɾA���Mw�� :�i��w�ý�L��[n;�\���rv���E<��˻��-���jy�:�^;�%;~�7;v�@;5E;�"G;
�G;7PH;�zH;��H;W�H;y�H;��H;��H;
�H;��H;��H;��H;	�H;��H;��H;{�H;T�H;H;�zH;:PH;�G;�"G;5E;u�@;��7;�%;�^;ry�:����-��˻�E<�rv��\���[n;��L��w�ýi��� :��Mw�A��9ɾGW�����W��pM+�      /y��v�i���B�߾����A��?����nH���C὜u����d�/O�hrμH"�����	����뺠r89\;�:b�;�+;R|:;{7B;��E;�aG;qH;�ZH;b�H;)�H;��H;�H;H�H;D�H;�H;��H;r�H;��H;�H;D�H;E�H;�H;��H;0�H;c�H;�ZH;rH;bG;��E;y7B;R|:;�+;`�;h;�:�r89���	�����H"��hrμ/O���d��u��C����nH�?���A������B�߾i����v�      @�;9ɾ|㼾B�������Mw��nH�����Z�䳽ʕ��q\8�m#������^N�J���b��Hx�H5:��:1�;��0;]=;A�C;�[F;ӞG;�)H;�eH;r�H;#�H;:�H;��H;�H;��H;(�H;��H;k�H;��H;*�H;��H;�H;��H;:�H;+�H;s�H;�eH;�)H;ٞG;�[F;=�C;]=;��0;-�;��:P5:�Hx��b�I��^N�����m#��p\8�ʕ��䳽�Z񽰯��nH��Mw�����B��|㼾9ɾ      ఖ�����}���*|�LS\�� :����Z�k$������ �K�u���Oļ����������=&����I/�:�^;��#;�G6;7�?;��D;E�F;��G;@H;�pH;ޏH;r�H;�H;K�H;0�H;j�H;n�H;��H;w�H;��H;p�H;j�H;*�H;K�H;�H;z�H;ޏH;�pH;@H;��G;I�F;��D;;�?;�G6;��#;�^;O/�:���<&������������Oļu�� �K�����k$���Z���� :�LS\��*|�}������      �+X��T��nH��6��� �i��C�
䳽�����mR����ټ�����E<��?ݻ2d\������ :�d�:��;)�,;z�:;V7B;��E;mLG;,H;ZSH;�{H;|�H;�H;�H;=�H;T�H;
�H;��H;��H;��H;��H;��H;
�H;O�H;9�H;�H;�H;��H;�{H;\SH;.H;rLG;��E;Y7B;}�:;&�,;��;�d�:� :����0d\��?ݻ�E<�����ټ����mR�����
䳽B�i���� ��6��nH��T�      �� ]�ӈ�p}���w�ý�u��ʕ�� �K�����o�iv���&R���S^��x�� �>����:_B;:";i�4;��>;=D;��F;�G;�)H;fdH;q�H;�H;^�H;%�H;-�H;��H;��H;�H;	�H;��H;
�H;�H;��H;}�H;(�H;(�H;f�H;�H;r�H;gdH;�)H;��G;��F;@D;��>;g�4;C";bB;���: |>�v��R^�����&R�hv���o���� �K�ʕ���u��w�ý��p}�ӈ�]�       �ѽ\νx�ý䳽9����L����d�q\8�u��ټgv����Y��_� ���9���[���Y:]��:Lm;�r-;�:;m�A;+oE;�"G;K�G;XGH;�sH;�H;��H;�H;"�H;�H;��H;u�H;{�H;%�H;��H;%�H;|�H;y�H;��H;�H;%�H;�H;��H;�H;�sH;YGH;N�G;�"G;/oE;p�A;�:;�r-;Om;_��:��Y:�[�6�������_���Y�gv��ټu��p\8���d��L��9���䳽y�ý\ν      ���������Ȅ�iSt��Y�[n;�/O�l#���Oļ�����&R��_������N3�ԅY��3:�:د;�?&;�G6;X?;�D;$xF;��G;-!H;�^H;��H;�H;íH;;�H;��H;��H;��H;�H;��H;M�H;�H;M�H;��H;�H;��H;��H; �H;E�H;ɭH;�H;��H;�^H;3!H;��G;'xF;�D;�X?;�G6;�?&;կ;�:4:ȅY��N3������_��&R������Oļl#��/O�[n;��Y�iSt��Ȅ�����      ]n;�w\8��s/�<�!�y��^���grμ��������E<��� ����N3�DHx���9��:�^;U ;,2;a�<;�B;��E;$5G;�G;*FH;xqH;��H;>�H;��H;D�H;��H;��H;��H;��H;�H;k�H; �H;k�H;�H;��H;��H;��H;��H;P�H;��H;B�H;��H;vqH;.FH;�G;)5G;��E;��B;k�<;02;T ;�^;��:��9,Hx��N3��������E<��������grμ\���z��<�!��s/�v\8�      X������o�nrμσ��qv��H"��
^N�����?ݻQ^��>��ԅY���9��:٦�:��;R�.;~|:;�>A;��D;#�F;��G;�)H;aH;�H;u�H;۬H;,�H;�H;.�H;V�H;��H;�H;N�H;��H;��H;��H;M�H;�H;��H;Q�H;0�H;�H;2�H;�H;u�H;�H;aH;�)H;��G;&�F;��D;�>A;�|:;N�.;��;ݦ�:��:��9ȅY�8��O^���?ݻ���
^N�H"��pv��у��nrμ�o����      �����x���#��=F{���]��E<����F�뻦���0d\�n�뺬[��3:��:ߦ�:z[;d�,;��8;!@;�0D;r[F;{G;�
H;=PH;vH;ېH;6�H;��H;�H;]�H;p�H;��H;��H;s�H;n�H;��H;��H;��H;k�H;s�H;��H;��H;s�H;c�H;#�H;��H;8�H;אH;vH;>PH;�
H;{G;s[F;�0D;!@;��8;i�,;|[;��:��:�3:�[�h��,d\�����E�뻠���E<���]�>F{��#���x��      �B(� %�����_�����˻�����b�5&����� l>���Y:�:�^;��;i�,;`8;c�?;��C;lF;�FG;B�G;�?H;kH;�H;��H;�H;L�H;��H;b�H;i�H;�H;s�H;��H;��H;}�H;��H;x�H;~�H;��H;p�H;�H;n�H;f�H;��H;O�H;�H;��H;��H;!kH;�?H;D�G;�FG;uF;³C;^�?;`8;k�,;��;�^;�:��Y: \>�����3&���b� 	���˻�����_�����%�      ɚ��E��� J���X���b���-�����Hx����!:��:Q��:ѯ;R ;N�.;��8;X�?;��C;��E;*#G;��G;�1H;�aH;A�H;k�H;o�H;��H;��H;S�H;�H;&�H;/�H;��H;�H;��H;3�H;��H;0�H;~�H;�H;��H;*�H;,�H;�H;U�H;��H;��H;m�H;r�H;A�H;�aH;�1H;��G;3#G;��E;��C;\�?;��8;Q�.;T ;ӯ;]��:��:!:@���Hx������-��b��X��J��E���      �����"к������Y����@s89d5:U/�:�d�:iB;Im;�?&;02;�|:;!@;��C;��E;rG;��G;N(H;�ZH;czH;0�H;ɤH;��H;\�H;��H;��H;U�H;��H;��H;B�H;$�H;C�H;��H;u�H;��H;@�H;$�H;@�H;��H;��H;Z�H;��H;��H;\�H;��H;ФH;3�H;`zH;�ZH;R(H;��G;uG;��E;ĳC;!@;�|:;12;�?&;Om;lB;�d�:[/�:l5:s89�����Y�ғ��"к���      ��e9P�9�	�9�:8�Y:xy�:~;�:��:�^;��;C";�r-;�G6;i�<;�>A;�0D;uF;7#G;��G;�$H;UWH;�vH;k�H;5�H;7�H;o�H;�H;��H;q�H;0�H;��H;w�H;��H;!�H;�H;��H;��H;��H;�H;!�H;��H;t�H;��H;0�H;o�H;��H;�H;o�H;>�H;8�H;i�H;�vH;YWH;�$H;��G;4#G;uF;�0D;�>A;f�<;�G6;�r-;H";��;�^;���:x;�:�y�:T�Y:L:x	�9��9      b�:[-�:(g�:��:��:�^;^�;-�;��#;)�,;j�4;�:;�X?;�B;��D;v[F;�FG;��G;Q(H;PWH;_uH;��H;�H;�H;�H;��H;��H;��H;��H;��H;��H;��H;��H;��H;��H;S�H;M�H;L�H;��H;��H;��H;��H;��H;��H;��H;��H;��H;��H;�H;�H;
�H;��H;cuH;UWH;R(H;��G;�FG;v[F;��D;�B;�X?;�:;m�4;)�,;��#;,�;d�;�^;��:��:@g�:S-�:      �;x�;�l;[;d`;�%;�+;��0;�G6;��:;��>;m�A;�D;��E;*�F;{G;G�G;�1H;�ZH;�vH;��H;A�H;��H;ƸH;~�H;J�H;��H;��H;��H;��H;3�H;4�H;��H;��H;e�H;��H;��H;��H;b�H;��H;��H;/�H;6�H;��H;��H;��H;��H;M�H;��H;ŸH;��H;C�H;��H;�vH;�ZH;�1H;I�G;{G;-�F;��E;�D;s�A;��>;}�:;�G6;��0;�+;�%;z`;�Z;�l;k�;      �Y.;��.;0;�2;1�4;��7;c|:;)]=;C�?;`7B;HD;2oE;*xF;55G;��G;�
H;�?H;�aH;dzH;g�H;
�H;��H;B�H;��H;\�H;��H;��H;��H;�H;��H;��H;X�H;R�H;A�H;��H;�H;@�H;�H;��H;B�H;O�H;T�H;��H;��H;�H;��H;��H;��H;b�H;��H;?�H;��H;�H;j�H;ezH;�aH;�?H;�
H;��G;25G;-xF;6oE;LD;]7B;C�?;(]=;b|:;��7;@�4;�2;0;��.;      T�<;'�<;]=;�O>;�?;}�@;|7B;@�C;�D;��E;��F;�"G;��G;�G;�)H;APH;"kH;J�H;3�H;4�H;�H;��H;��H;1�H;*�H;-�H;?�H;��H;�H;5�H;��H;
�H;�H;��H;@�H;}�H;��H;v�H;=�H;��H;�H;�H;��H;4�H;�H;��H;<�H;1�H;/�H;/�H;��H;øH;�H;4�H;2�H;C�H;"kH;DPH;�)H;�G;��G;�"G;��F;��E;��D;H�C;|7B;k�@;��?;�O>;]=;�<;      �WC;�nC;ֲC;lD;7�D;(5E;��E;�[F;N�F;uLG;��G;R�G;3!H;5FH;aH;vH;��H;{�H;פH;B�H; �H;��H;b�H;4�H;��H;��H;;�H;��H;��H;��H;��H;��H;��H;1�H;��H;��H;��H;��H;��H;4�H;��H;��H;��H;��H;��H;��H;7�H;�H;��H;3�H;b�H;��H; �H;?�H;ؤH;v�H; �H;vH;aH;4FH;5!H;X�G;��G;vLG;P�F;�[F;��E;5E;C�D;jD;زC;�nC;      �ZF;�dF;ހF;)�F;��F;�"G;bG;�G;��G;5H;�)H;`GH;�^H;�qH;�H;ߐH;��H;q�H;��H;l�H;��H;H�H;��H;1�H;��H;�H;��H;��H;h�H;��H;��H;��H;�H;t�H;��H;�H;�H;�H;��H;t�H; �H;��H;��H;��H;e�H;��H;��H;#�H;�H;0�H;��H;K�H;��H;n�H;��H;m�H;�H;ߐH;�H;}qH;�^H;_GH;�)H;6H;��G;�G;bG;�"G;��F;/�F;�F;�dF;      �G;�G;q�G;~�G;�G;
�G;~H;�)H;@H;]SH;hdH;�sH;��H;��H;u�H;;�H;�H;��H;^�H;�H;��H;��H;��H;C�H;9�H;��H;��H;;�H;~�H;��H;^�H;��H;p�H;��H;�H;6�H;Q�H;/�H;��H;��H;q�H;��H;]�H;��H;z�H;9�H;��H;��H;;�H;A�H;��H;��H;��H;�H;^�H;��H;�H;=�H;w�H;��H;��H;�sH;jdH;ZSH; @H;�)H;{H;�G;�G;p�G;p�G;ݪG;      0H;�1H;6H;=H;�EH;=PH;�ZH;�eH;�pH;�{H;r�H;�H;�H;F�H;ެH;��H;O�H;��H;��H;��H;��H;��H;��H;��H;��H;��H;9�H;u�H;\�H;H�H;��H;b�H;��H;	�H;A�H;V�H;A�H;Q�H;?�H;	�H;��H;^�H;��H;F�H;Y�H;r�H;6�H;��H;��H;��H;��H;��H;��H;��H;��H;��H;P�H;��H;ެH;E�H;�H;�H;w�H;�{H;�pH;�eH;�ZH;1PH;FH;=H;6H;�1H;      /jH;�jH;mH;�pH;6uH;�zH;j�H;r�H;ُH;}�H;�H;��H;ɭH;��H;2�H;&�H;��H;\�H;��H;u�H;��H;��H;�H;�H;��H;b�H;u�H;]�H;P�H;��H;M�H;��H;��H;0�H;`�H;f�H;V�H;b�H;\�H;0�H;��H;��H;N�H;��H;O�H;Z�H;r�H;b�H;��H;�H;�H;��H;��H;q�H;��H;Y�H;��H;'�H;2�H;��H;ɭH;��H;�H;��H;ُH;r�H;j�H;�zH;DuH;�pH;mH;�jH;      ;�H;��H;3�H;��H;ƓH;��H;-�H;&�H;x�H;�H;e�H;�H;B�H;P�H;�H;b�H;j�H;�H;U�H;1�H;��H;��H;��H;3�H;��H;��H;��H;I�H;��H;C�H;��H;��H;,�H;X�H;c�H;x�H;��H;w�H;`�H;V�H;.�H;��H;��H;@�H;��H;I�H;�H;��H;��H;1�H;��H;��H;��H;.�H;U�H;�H;j�H;d�H;�H;M�H;B�H;�H;e�H;�H;x�H;&�H;0�H;��H;ȓH;��H;6�H;��H;      P�H;��H;��H;L�H;��H;X�H;��H;>�H;�H;�H;/�H;-�H;�H;��H;9�H;z�H;w�H;3�H;��H;��H;��H;9�H;��H;��H;��H;��H;[�H;��H;P�H;��H;��H;"�H;V�H;g�H;��H;�H;z�H;|�H;~�H;i�H;[�H;!�H;��H;��H;M�H;��H;Z�H;��H;��H;��H;��H;9�H;��H;��H;��H;2�H;z�H;{�H;7�H;��H;	�H;/�H;/�H;�H;�H;@�H;��H;M�H;��H;I�H;��H;��H;      ��H;յH;�H;��H;~�H;q�H;��H;��H;P�H;?�H;.�H;�H;��H;��H;]�H;��H;�H;7�H;��H;�H;��H;6�H;V�H;
�H;��H;��H;��H;c�H;��H;��H;�H;<�H;`�H;�H;��H;��H;��H;��H;��H;��H;f�H;9�H;�H;��H;��H;a�H;��H;��H;��H;�H;\�H;8�H;��H;|�H;��H;9�H; �H;��H;[�H;��H;��H;�H;2�H;@�H;P�H;��H;��H;t�H;��H;ŷH;��H;յH;      /�H;u�H;�H;��H;�H;��H;I�H;�H;)�H;T�H;��H;��H;��H;��H;��H;��H;|�H;��H;L�H;��H;��H;��H;P�H;�H;��H;�H;o�H;��H;��H;3�H;V�H;f�H;u�H;��H;��H;��H;��H;��H;��H;��H;x�H;d�H;U�H;,�H;��H;��H;p�H;�H;��H;�H;V�H;��H;��H;��H;L�H;��H;��H;��H;��H;��H;��H;��H;��H;U�H;-�H;�H;J�H;|�H;!�H;��H;�H;t�H;      ��H;��H;D�H;��H;��H;��H;K�H;��H;n�H;�H;��H;��H;�H;��H;�H;}�H;��H;�H;+�H;+�H;��H;��H;>�H;��H;-�H;o�H;��H;�H;.�H;[�H;c�H;��H;��H;��H;��H;��H;��H;��H;��H;��H;��H;��H;c�H;X�H;,�H;�H;��H;p�H;/�H;��H;E�H;��H;��H;$�H;*�H;�H;��H;}�H;�H;��H;�H;�H;��H;�H;q�H;��H;N�H;��H;��H;��H;I�H;��H;      V�H;w�H;��H;b�H;.�H;�H;�H;.�H;u�H;��H;$�H;��H;��H;�H;[�H;v�H;��H;��H;H�H;�H;��H;e�H;��H;5�H;��H;��H;��H;@�H;b�H;g�H;{�H;��H;��H;��H;��H;��H;��H;��H;��H;��H;��H;��H;z�H;b�H;[�H;<�H;��H;��H;��H;5�H;��H;b�H;��H;�H;D�H;��H;��H;v�H;X�H;�H;��H;��H;'�H;��H;z�H;/�H;�H;�H;.�H;c�H;��H;y�H;      ��H;��H;�H;z�H;�H;��H;��H;��H;��H;��H;�H;.�H;T�H;w�H;��H;��H;��H;6�H;��H;��H;W�H;��H;�H;m�H;��H;�H;.�H;U�H;i�H;�H;~�H;��H;��H;��H;��H;��H;��H;��H;��H;��H;��H;��H;|�H;z�H;f�H;T�H;2�H;�H;��H;o�H;�H;��H;S�H;��H;��H;7�H;��H;��H;��H;t�H;U�H;-�H;�H;��H;��H;��H;��H;��H;�H;v�H;�H;��H;      ��H;��H;��H;a�H;��H;��H;|�H;o�H;~�H;��H;��H;��H;�H;�H;��H;��H;��H;��H;|�H;��H;X�H;��H;@�H;��H;��H;	�H;K�H;H�H;\�H;��H;w�H;��H;��H;��H;��H;��H;��H;��H;��H;��H;��H;��H;w�H;��H;X�H;F�H;O�H;�H;��H;��H;F�H;��H;S�H;��H;{�H;��H;��H;��H;��H;�H;�H;��H;��H;��H;�H;r�H;��H;��H;��H;b�H;��H;��H;      ��H;��H; �H;y�H;�H;��H;��H;��H;��H;��H;�H;.�H;T�H;u�H;��H;��H;��H;5�H;��H;��H;X�H;��H;�H;m�H;��H;	�H;.�H;U�H;j�H;~�H;~�H;��H;��H;��H;��H;��H;��H;��H;��H;��H;��H;��H;|�H;x�H;f�H;R�H;0�H;�H;��H;m�H;�H;��H;S�H;��H;��H;9�H;��H;��H;��H;r�H;T�H;-�H;�H;��H;��H;��H;��H;��H;�H;z�H;�H;��H;      I�H;z�H;��H;[�H;/�H; �H;�H;1�H;u�H;��H;$�H;��H;��H;�H;\�H;x�H;��H;��H;H�H;�H;��H;g�H;��H;5�H;��H;��H;��H;@�H;`�H;f�H;z�H;��H;��H;��H;��H;��H;��H;��H;��H;��H;��H;��H;z�H;`�H;]�H;<�H;��H;��H;��H;4�H;��H;d�H;��H;�H;F�H;��H;��H;x�H;V�H;�H;��H;��H;$�H;��H;w�H;6�H;�H; �H;5�H;_�H;��H;|�H;      ��H;��H;A�H;��H;��H;��H;H�H;��H;p�H;�H;��H;�H;�H;��H;�H;~�H;��H;�H;+�H;)�H;��H;��H;A�H;��H;/�H;p�H;��H;�H;0�H;[�H;c�H;��H;��H;��H;��H;��H;��H;��H;��H;��H;��H;��H;b�H;X�H;)�H;�H;��H;s�H;.�H;��H;E�H;��H;��H;%�H;+�H;�H;��H;~�H;�H;��H;�H;�H;��H;�H;p�H;��H;P�H;��H;��H;��H;I�H;��H;      /�H;x�H;
�H;��H;�H;��H;F�H;�H;*�H;V�H;��H;��H;��H;��H;��H;��H;~�H;��H;K�H;��H;��H;��H;P�H;�H;��H;�H;o�H;��H;��H;3�H;U�H;c�H;u�H;��H;��H;��H;��H;��H;��H;��H;w�H;f�H;U�H;.�H;��H;��H;p�H;�H;��H;�H;W�H;��H;��H;��H;I�H;��H;}�H;��H;��H;��H;��H;��H;��H;U�H;,�H;�H;O�H;��H;�H;��H;�H;r�H;      t�H;ҵH;u�H;ķH;}�H;��H;��H;��H;O�H;?�H;/�H;�H;��H;��H;`�H;��H;�H;9�H;��H;�H;��H;9�H;X�H;	�H;��H;��H;��H;c�H;��H;��H;�H;:�H;c�H;~�H;��H;��H;��H;��H;��H;��H;d�H;:�H;�H;��H;��H;a�H;��H;��H;��H; �H;]�H;8�H;��H;{�H;��H;6�H;�H;��H;[�H;��H;��H;�H;/�H;?�H;R�H;��H;��H;t�H;~�H;ƷH;{�H;͵H;      C�H;��H;��H;H�H;��H;X�H;��H;A�H;�H;�H;-�H;0�H;�H;��H;:�H;{�H;y�H;2�H;��H;��H;��H;:�H;��H;��H;��H;��H;Z�H;��H;S�H;��H;��H;"�H;V�H;g�H;��H;~�H;z�H;�H;~�H;i�H;[�H;$�H;��H;��H;L�H;��H;[�H;��H;��H;��H;��H;:�H;��H;��H;��H;2�H;|�H;{�H;9�H;��H;�H;/�H;-�H;�H;�H;D�H;��H;V�H;��H;R�H;��H;��H;      F�H;��H;.�H;��H;��H;ŗH;0�H;-�H;{�H;�H;e�H;�H;E�H;P�H;�H;c�H;i�H;�H;W�H;3�H;��H;��H;��H;3�H;��H;��H;��H;J�H;��H;C�H;��H;��H;)�H;X�H;c�H;w�H;��H;x�H;`�H;X�H;.�H;��H;��H;@�H;��H;F�H;��H;��H;��H;-�H;��H;��H;��H;.�H;W�H;�H;j�H;c�H;�H;P�H;B�H;�H;f�H;�H;x�H;*�H;1�H;��H;ȓH;��H;6�H;��H;      =jH;�jH;-mH;�pH;2uH;{H;j�H;s�H;��H;|�H;�H;��H;˭H;��H;3�H;'�H;��H;^�H;��H;t�H;��H;��H;�H;�H;��H;a�H;t�H;\�H;S�H;��H;M�H;��H;��H;/�H;]�H;d�H;V�H;d�H;\�H;/�H;��H;��H;N�H;��H;M�H;Y�H;t�H;e�H;��H;�H;�H;��H;��H;r�H;��H;Y�H;��H;(�H;3�H;��H;ʭH;��H;�H;|�H;ݏH;y�H;o�H;�zH;@uH;�pH;-mH;�jH;      0H;�1H;6H;=H;�EH;FPH;�ZH;�eH;�pH;�{H;w�H;�H;�H;F�H;�H;��H;P�H;��H;��H;��H;��H;��H;��H;��H;��H;��H;6�H;t�H;]�H;F�H;��H;b�H;��H;�H;?�H;R�H;A�H;T�H;=�H;	�H;��H;_�H;��H;H�H;Z�H;r�H;8�H;��H;��H;��H;��H;��H;��H;��H;��H;��H;P�H;��H;�H;C�H;�H;�H;x�H;�{H;�pH;�eH;�ZH;6PH;FH;=H;6H;�1H;      �G;��G;k�G;��G;�G;�G;~H;�)H;@H;]SH;jdH;�sH;��H;��H;w�H;<�H;�H;��H;`�H;�H;��H;��H;��H;F�H;;�H;��H;��H;;�H;~�H;��H;[�H;��H;o�H;��H;�H;2�H;O�H;0�H;��H;��H;p�H;��H;^�H;��H;z�H;8�H;��H;��H;9�H;?�H;��H;��H;��H;�H;`�H;��H;�H;=�H;x�H;��H;��H;�sH;hdH;\SH;@H;�)H;H;�G;�G;��G;p�G;�G;      �ZF;�dF;�F;'�F;��F;�"G; bG;�G;��G;3H;�)H;bGH;�^H;qH;�H;�H;��H;t�H;��H;n�H;��H;K�H;��H;4�H; �H;�H;��H;��H;i�H;��H;��H;��H;�H;t�H;��H;�H;�H;�H;��H;s�H;�H;��H;��H;��H;c�H;��H;��H;!�H;��H;.�H;��H;J�H;��H;n�H;��H;m�H;�H;�H;�H;}qH;�^H;_GH;�)H;5H;��G;ߞG;�aG;�"G;��F;&�F;ЀF;�dF;      �WC;�nC;ҲC;iD;9�D;+5E;��E;�[F;P�F;uLG;��G;U�G;3!H;4FH;aH;vH; �H;|�H;ڤH;B�H; �H;��H;b�H;7�H;��H;��H;9�H;��H;��H;��H;��H;��H;��H;1�H;��H;��H;��H;��H;��H;2�H;��H;��H;��H;��H;��H;��H;:�H; �H;��H;2�H;c�H;��H; �H;B�H;ڤH;v�H; �H;vH;aH;2FH;4!H;U�G;��G;vLG;L�F;�[F;��E;5E;?�D;jD;ҲC;�nC;      1�<;�<;]=;�O>;݁?;��@;7B;D�C;��D;��E;��F;�"G;��G;�G;�)H;EPH;$kH;K�H;3�H;5�H;�H;øH;��H;4�H;/�H;*�H;?�H;��H;�H;3�H;��H;�H;�H;��H;?�H;z�H;��H;{�H;=�H;��H;�H;
�H;��H;4�H;�H;��H;?�H;.�H;,�H;1�H;��H;¸H;�H;6�H;5�H;D�H;$kH;BPH;�)H;�G;��G;�"G;��F;��E;��D;@�C;|7B;v�@;�?;�O>;]=;��<;      �Y.;��.;0;�2;/�4;��7;\|:;+]=;G�?;_7B;ED;6oE;+xF;35G;��G;�
H;�?H;�aH;ezH;j�H;�H;��H;A�H;��H;b�H;��H;��H;��H;�H;��H;��H;X�H;O�H;A�H;��H;�H;C�H;�H;��H;?�H;P�H;X�H;��H;��H;�H;��H;��H;��H;^�H;��H;A�H;��H;�H;k�H;ezH;�aH;�?H;�
H;��G;/5G;+xF;3oE;GD;_7B;F�?;,]=;\|:;��7;.�4;�2;0;��.;      �;x�;�l;�Z;h`;�%;�+;��0;�G6;}�:;��>;u�A;�D;��E;-�F;!{G;I�G;�1H;�ZH;�vH;��H;D�H;��H;ƸH;��H;H�H;��H;��H;��H;��H;4�H;4�H;��H;��H;b�H;��H;��H;��H;b�H;��H;��H;2�H;7�H;��H;��H;��H;��H;K�H;�H;ǸH;��H;C�H;��H;�vH;�ZH;�1H;G�G;{G;,�F;��E;�D;s�A;��>;}�:;�G6;��0;�+;�%;|`;�Z;�l;n�;      N�:�-�:Jg�:.��:��:�^;d�;1�;��#;)�,;m�4;�:;�X?;�B;��D;y[F;�FG;��G;R(H;UWH;buH;��H;�H;��H;�H;��H;��H;��H;��H;��H;��H;��H;��H;��H;��H;M�H;O�H;O�H;��H;��H;��H;��H;��H;��H;��H;��H;��H;��H;�H;�H;
�H;��H;buH;VWH;R(H;��G;�FG;v[F;��D;�B;�X?;
�:;n�4;)�,;��#;3�;d�;�^;��:(��:dg�:g-�:      Рe9��9�	�9�:@�Y:�y�:�;�:���:�^;��;H";�r-;�G6;h�<;�>A;�0D;uF;7#G;��G;�$H;ZWH;�vH;k�H;8�H;>�H;n�H;�H;��H;r�H;,�H;��H;x�H;��H;"�H;�H;��H;��H;��H;�H;�H;��H;w�H;��H;.�H;q�H;��H;�H;o�H;8�H;;�H;j�H;�vH;WWH;�$H;��G;4#G;wF;�0D;�>A;h�<;�G6;�r-;H";��;�^;��:x;�:ry�:X�Y:t:�	�9`�9      �����"к������Y���� s89l5:W/�:�d�:hB;Om;�?&;.2;�|:;"!@;��C;��E;sG;��G;S(H;�ZH;ezH;2�H;ФH;��H;\�H;��H;��H;T�H;��H;��H;A�H;$�H;D�H;��H;u�H;��H;C�H;#�H;A�H;��H;��H;W�H;��H;��H;\�H;��H;ʤH;3�H;dzH;�ZH;Q(H;��G;rG;��E;³C;!@;�|:;-2;�?&;Lm;iB;�d�:[/�:t5:�r89�����Y�����,кv��      К��@���#J���X���b���-�����Hx�P��!:��:_��:կ;Q ;T�.;��8;\�?;��C;��E;1#G;��G;�1H;�aH;C�H;r�H;m�H;��H;��H;V�H;�H;*�H;-�H;��H;�H;�H;2�H;��H;3�H;}�H;�H;��H;-�H;*�H;�H;U�H;��H;��H;l�H;k�H;A�H;�aH;�1H;��G;1#G;��E;��C;Z�?;��8;R�.;P ;ѯ;Y��:��:!:`���Hx������-��b��X��(J��@���      �B(��%�����_�}����˻ 	����b�5&����� d>���Y:�:�^;��;m�,;`8;b�?;��C;tF;�FG;F�G;�?H;!kH;��H;��H;�H;J�H;��H;_�H;l�H;�H;s�H;��H;��H;{�H;��H;{�H;~�H;��H;p�H;�H;n�H;b�H;��H;J�H;�H;��H;�H;kH;�?H;@�G;�FG;sF;��C;^�?;`8;i�,;��;�^;�:��Y: d>�����3&���b�	���˻�����_�����%�      �����x���#��<F{���]��E<����D�뻤���.d\�h�뺌[� 4:��:��:~[;f�,;��8;!@;�0D;y[F;{G;�
H;>PH;vH;ݐH;5�H;��H;!�H;]�H;q�H;��H;��H;t�H;o�H;��H;��H;��H;k�H;q�H;��H;��H;q�H;`�H;!�H;��H;4�H;֐H;vH;;PH;�
H;{G;n[F;�0D;!@;��8;f�,;z[;��:��:�3:�[�l��/d\�����F�뻡���E<���]�=F{��#���x��      Y������o�mrμσ��pv��H"��
^N�����?ݻP^��8��ȅY���9 �:��:��;Q�.;�|:;�>A;��D;)�F;��G;�)H;aH;�H;t�H;ݬH;0�H;�H;0�H;V�H;��H;�H;N�H;��H;��H;��H;N�H;�H;��H;S�H;/�H;�H;2�H;ݬH;q�H;�H;aH;�)H;��G;&�F;��D;�>A;~|:;K�.;��;٦�:��:��9ԅY�:��P^���?ݻ���
^N�H"��qv��Ѓ��orμ�o����      ]n;�w\8��s/�<�!�y��\���grμ��������E<��������N3�,Hx��9�:�^;R ;.2;f�<;��B;��E;+5G;�G;0FH;}qH;��H;?�H;��H;I�H;��H;��H;��H;��H;�H;k�H; �H;m�H;�H;��H;��H;��H;��H;M�H;��H;A�H;��H;uqH;*FH;�G;/5G;��E;�B;h�<;*2;Q ;�^;��:��94Hx��N3��������E<��������hrμ]���z��<�!��s/�v\8�      ���������Ȅ�iSt��Y�[n;�.O�l#���Oļ�����&R��_������N3���Y�4:
�:֯;�?&;�G6;�X?;�D;-xF;��G;3!H;�^H;��H;�H;ʭH;?�H; �H;��H;��H;�H;��H;M�H;�H;M�H;��H;�H;��H;��H;��H;B�H;ɭH;�H;��H;�^H;-!H;��G;+xF;�D;{X?;�G6;�?&;ѯ;
�:�3:ȅY��N3������_��&R������Oļl#��/O�[n;��Y�iSt��Ȅ�����       �ѽ\νx�ý䳽9����L����d�p\8�u��ټgv����Y��_�����5���[���Y:W��:Om;�r-;�:;q�A;4oE;�"G;P�G;[GH;�sH;�H;��H;�H;&�H;�H;��H;x�H;|�H;#�H;��H;%�H;z�H;v�H;��H;�H;#�H;�H;��H;�H;�sH;WGH;J�G;�"G;3oE;m�A;�:;�r-;Jm;W��:��Y:�[�7�������_���Y�gv��ټu��p\8���d��L��9���䳽x�ý\ν      ��]�ӈ�p}���w�ý�u��ʕ�� �K�����o�hv���&R���P^��r�� �>����:aB;>";n�4;��>;ED;��F;��G;�)H;fdH;q�H;�H;a�H;(�H;+�H;��H;��H;�H;
�H;��H;
�H;�H;��H;}�H;(�H;%�H;e�H;�H;q�H;ddH;�)H;�G;��F;DD;��>;b�4;>";^B;���: �>�v��S^�����&R�hv���o���� �K�ʕ���u��w�ý��p}�ӈ� ]�      �+X��T��nH��6��� �i��C�
䳽�����mR����ټ�����E<��?ݻ0d\������ :�d�:��;.�,;|�:;_7B;��E;rLG;0H;ZSH;�{H;�H;�H;�H;<�H;T�H;�H;��H;��H;��H;��H;��H;
�H;O�H;9�H;�H;�H;�H;�{H;YSH;.H;nLG;��E;\7B;y�:;"�,;��;�d�:� :����2d\��?ݻ�E<�����ټ����mR�����
䳽C�i���� ��6��nH��T�      ఖ�����}���*|�LS\�� :����Z�k$������ �K�u���Oļ����������;&����M/�:�^;��#;�G6;<�?;��D;L�F;��G;@H;�pH;��H;u�H;�H;K�H;.�H;k�H;n�H;��H;w�H;��H;m�H;j�H;*�H;K�H;�H;x�H;ޏH;�pH;@H;��G;I�F;��D;>�?;�G6;��#;�^;G/�:���<&������������Oļu�� �K�����k$���Z���� :�LS\��*|�}������      @�;9ɾ|㼾B�������Mw��nH�����Z�䳽ʕ��q\8�m#������^N�I���b� Ix�T5:��:4�;��0;]=;@�C;�[F;֞G;�)H;�eH;r�H;#�H;=�H;��H;�H;��H;'�H;��H;k�H;��H;(�H;��H;�H;��H;:�H;*�H;u�H;�eH;�)H;؞G;�[F;?�C;]=;��0;,�;��:H5:�Hx��b�J��^N�����m#��q\8�ʕ��䳽�Z񽰯��nH��Mw�����B��|㼾9ɾ      /y��v�i���B�߾����A��?����nH���C὜u����d�/O�hrμH"�����	����뺐r89f;�:d�;�+;R|:;y7B;��E;�aG;pH;�ZH;e�H;,�H;��H;�H;F�H;D�H;�H;��H;r�H;��H;�H;B�H;C�H;�H;��H;1�H;f�H;�ZH;tH;bG;��E;{7B;W|:;�+;]�;j;�:�r89��� 	�����H"��hrμ/O���d��u��C����nH�?���A������B�߾i����v�      �O/�pM+�W�����GW��9ɾA���Mw�� :�i��w�ý�L��[n;�\���rv���E<��˻��-���py�:�^;�%;~�7;v�@;5E;�"G;	�G;7PH;�zH;��H;Z�H;|�H;��H;��H;
�H;��H;��H;��H;	�H;��H;��H;{�H;T�H;H;�zH;:PH;�G;�"G;5E;v�@;��7;�%;�^;vy�:����-��˻�E<�rv��\���[n;��L��w�ýi��� :��Mw�A��9ɾGW�����W��pM+�      7�X�VvS�6E��O/��S�GW����������LS\��� ���9����Y�z��σ����]����� �b���Y�T�Y:��:f`;6�4;�?;<�D;��F;�G;FH;FuH;��H;��H;��H;�H;��H;�H;�H;��H;�H;�H;��H;�H;��H;��H;ɓH;GuH;FH;�G;��F;;�D;�?;6�4;f`;��:X�Y:��Y��b�������]�σ��z���Y�9����彑� �LS\���������GW���S��O/�6E�VvS�      � ����y�`�h���N��O/����B�߾B���*|��6�p}�䳽hSt�;�!�nrμ?F{��_��X����X:4��:�Z;�2;�O>;mD;&�F;w�G;=H;�pH;��H;I�H;̷H;��H;��H;^�H;z�H;a�H;w�H;[�H;��H;��H;ͷH;G�H;��H;�pH;=H;}�G;3�F;lD;�O>;�2;�Z;.��:p:Ɠ���X���_�?F{�nrμ;�!�hSt�䳽p}��6��*|�B��B�߾����O/���N�`�h���y�      =v��b���W ��`�h�6E�W��j���|㼾}���nH�ӈ�x�ý�Ȅ��s/��o��#�����"J�� кh	�9^g�:�l;"0;]=;ڲC;րF;m�G;6H;mH;%�H;��H;��H;��H;>�H;��H;�H;��H;�H;��H;>�H;��H;�H;��H;/�H; mH;6H;t�G;�F;ٲC;]=;0;�l;Xg�:�	�9"к!J������#���o��s/��Ȅ�x�ýӈ��nH�}��|㼾j���W��6E�`�h�W ��b���      |h��/���b�����y�VvS�pM+��v�9ɾ�����T� ]�\ν����x\8�����x��%�K���h��x�9{-�:j�;��.;�<;�nC;�dF;�G;�1H;�jH;��H;��H;͵H;j�H;��H;g�H;��H;��H;��H;e�H;��H;i�H;͵H;��H;��H;�jH;�1H;�G;�dF;�nC;�<;��.;g�;o-�:��9n��J���%��x�����x\8�����\ν ]��T�����9ɾ�v�pM+�VvS���y�b���/���      EEb�`]��N��7����s� ���˾��(�j��!,�o���K��Bm�+��6,˼��x�Z���1�����`�:v�:�;�1;7,>;e�C;SwF;��G;m H;�>H;�hH;,�H;B�H;�H;��H;��H;�H;m�H;�H;��H;��H;�H;A�H;)�H;�hH;�>H;n H;�G;cwF;e�C;6,>;�1;�;t�:p�:����1��Z����x�6,˼+��Bm�K��o����!,�(�j�����˾s� �����7��N�`]�      `]�d�W��TI�v3��D�������Ǿv����f�7)�$��r;���Fi��k���Ǽ�[t�L�	�)Ȅ�X��ؠ:��:��;*J2;SZ>;'	D;;F;8�G;�H;�?H;viH;H;��H;S�H;�H;��H;7�H;��H;1�H;��H;�H;Q�H;��H;��H;~iH;�?H;�H;=�G;IF;'	D;SZ>;&J2;��;��:�:X��(Ȅ�L�	��[t���Ǽ�k��Fi�r;��$��7)��f�v�����Ǿ�����D�v3��TI�d�W�      �N��TI���;�/�'�l������x󐾲Z��K ��s�@����&^���"����g����̨u�� ���2<:��:�
;9g3;��>;UBD;u�F;ޔG;iH;BH;\kH;,�H;��H;	�H;��H;C�H;��H;$�H;��H;B�H;��H;�H;��H;(�H;ekH;BH;kH;�G;��F;WBD;��>;5g3;�
;��:�2<:� ��ʨu������g��"����&^�@����s潥K ��Z�x������l�/�'���;��TI�      �7�v3�/�'����s� ��{Ծ ���H���y�F�����ӽ���]�L�Iv��뮼PT����PV���=�`)i:z��:�z ;�$5;��?;�D;��F;�G;rH;dFH;rnH;a�H;K�H;K�H;��H;�H;1�H;��H;-�H;�H;��H;J�H;K�H;]�H;znH;fFH;rH;�G;��F;�D;��?;z$5;�z ;z��:t)i:��=��PV���OT��뮼Iv�]�L�����ӽ���y�F�H�������{Ծs� ����/�'�v3�      ����D�l�s� �V�ݾj���V͓��f��>/�����'���섽O�6�}t�w��]�:�%Tʻz.�۷�Bt�:�;��$;�Y7;R�@;�	E;��F;*�G;�H;LH;�rH;��H;��H;��H;��H;�H;$�H;��H; �H;�H;��H;��H;��H;��H;�rH;	LH;�H;.�G;��F;�	E;R�@;�Y7;��$;�;Nt�: ۷�x.�%Tʻ]�:�w��~t�O�6��섽�'������>/��f�V͓�j���V�ݾs� �l��D�      s� ��������{Ծj���v���Y�x��SC��^��޽?���x�e�'��B�Ѽ#G������R����� ޤ8Ň�:�Y;G�);��9;��A;��E;G;�G;@!H;	SH;�wH;I�H;Y�H;�H;��H;K�H;V�H;��H;P�H;I�H;��H;�H;Z�H;G�H;�wH;
SH;A!H;�G;�G;��E;��A;��9;G�);�Y;χ�:@ޤ8����R�����#G��B�Ѽ'��w�e�?����޽�^��SC�Z�x�v���j����{Ծ�쾠���      ��˾��Ǿ���� ���V͓�Y�x���J��K �m���������?����뮼)�[����3|��W����:=�:�';a/;=g<;�C;DF;�NG;��G;-H;;[H;�}H;��H;��H;��H;�H;��H;��H;��H;��H;��H;�H;��H;��H;��H;�}H;>[H;-H;��G;�NG;GF;�C;=g<;b/;�';I�:��:�W��3|����)�[��뮼���?������l����K ���J�Y�x�V͓� ���������Ǿ      ��v���x�G����f��SC��K �nn����Ž���
�Z��k�}ռ,X��`y-�*���n.�h��P�:�+�:~�;4;�>;�D;�wF;��G;��G;�9H;'dH;S�H;~�H;2�H;H�H;��H;~�H;+�H;E�H;(�H;�H;��H;E�H;/�H;}�H;[�H;)dH;�9H;��G;�G;�wF;�D;�>;4;{�;�+�:�P�:X��m.�)���_y-�,X��}ռ�k�
�Z������Žmn���K ��SC��f�G���x�v���      (�j��f��Z�y�F��>/��^�l�����ŽF ���Fi��Q+�zt�mT��l�W�����1��"Ⱥ0X�9wP�:�Y;��(;��8;�A;�E;��F;8�G;rH;�FH;�mH;j�H;��H;�H;H�H;��H;`�H;��H;��H;��H;`�H;��H;D�H;�H;��H;q�H;�mH;�FH;sH;9�G;��F;�E;�A;��8;��(;�Y;}P�:(X�9Ⱥ�1�����k�W�mT��zt�Q+��Fi�F ����Žl����^��>/�y�F��Z��f�      �!,�7)��K ��������޽������Fi��0����鷼��x�����.��O�(����+i:z��:%�;��0;8�<;oC;��E;�<G;��G;�$H;:TH;�wH;ȒH;�H;!�H;X�H;�H;c�H;q�H;M�H;p�H;d�H;�H;T�H;�H;�H;ΒH;�wH;>TH;�$H;��G;�<G;��E;rC;<�<;��0;.�;���:+i:���M�(��.�������x�鷼����0��Fi�������޽�������K �7)�      o���$��s��ӽ�'��?������
�Z��Q+�����"��G����0���׻ƕb�4W���X�9ԡ�: `;~*';�Y7;�#@;�D;�F;�G;��G;8H;�aH;́H;5�H;y�H;H�H;k�H;v�H;V�H;"�H;
�H;%�H;X�H;x�H;h�H;F�H;z�H;<�H;ҁH;�aH;8H;��G;��G;��F;�D;�#@;�Y7;�*';"`;ԡ�:Y�92W��ĕb���׻��0�G���"������Q+�
�Z����?����'���ӽ�s�$��      J��r;��@�������섽x�e��?��k�zt�鷼G���e7�����Ǆ�l0�@�t�u�:,�:n;l1;B�<;I�B; �E;�G;��G;0H;RJH;3oH;ҋH;��H;�H;m�H;��H;��H;i�H;��H;��H;��H;i�H;��H;��H;i�H;�H;��H;ڋH;6oH;QJH;2H;��G;�G;�E;N�B;E�<;x1;p;,�:(u�: �t�f0��Ǆ���껁e7�G��鷼zt��k��?�w�e��섽���@���r;��      Bm��Fi��&^�^�L�N�6�'����}ռmT����x���0����������ط��n`:��:�;�*;�8;��@;�D;D�F;�}G;z�G;k1H;�[H;E|H;��H;��H;W�H;��H;��H;]�H;e�H;��H;D�H;��H;e�H;]�H;��H;��H;]�H;��H;��H;F|H;�[H;k1H;��G;�}G;G�F;!�D;��@;'�8;�*;�;��:o`:xط��������껽�0���x�lT��}ռ��'��O�6�^�L��&^��Fi�      )���k��Jv�{t�C�Ѽ�뮼+X��l�W������׻�Ǆ��� ��5<:Y��:�Y;�t%;�$5;�Z>;�`C;��E;*G;B�G;�H;�GH;FlH;ɈH;ӞH;��H;��H;n�H;��H;��H;H�H;E�H; �H;C�H;G�H;��H;��H;j�H;��H;��H;ܞH;̈H;FlH;�GH;�H;B�G;*G;��E;�`C;�Z>;�$5;�t%;�Y;Y��:5<:������Ǆ���׻���j�W�+X���뮼B�Ѽ~t�Jv���k�      5,˼��Ǽ�"���뮼w��#G��)�[�]y-�����.��b�t0㺘ط�5<:�L�:�\;r�!;�J2;�g<;-0B;CE;�F;%�G;��G;_4H;v\H;�{H;~�H;v�H;/�H;��H;�H;h�H;#�H;#�H;��H;�H;��H;#�H;$�H;g�H;�H;��H;6�H;|�H;��H;�{H;s\H;c4H;��G;'�G;�F;CE;80B;�g<;�J2;z�!;�\;�L�:5<:�ط�j0㺾�b��.�����]y-�)�[�"G��w���뮼�"����Ǽ      ��x��[t���g�NT�]�:�������&����1��L�(�.W����t��n`:[��:�\;{ ;��0;R;;�<A;��D;�wF;�cG;-�G;�!H;�MH;WoH;J�H;Z�H;��H;e�H;7�H;��H;-�H;B�H;��H;k�H;��H;j�H;��H;B�H;*�H;��H;:�H;k�H;��H;^�H;J�H;SoH;�MH;�!H;.�G;�cG;�wF;��D;�<A;N;;��0;{ ;�\;[��:�n`:��t�&W��J�(��1��%���������_�:�NT���g��[t�      W��J�	������"Tʻ�R��3|�i.�Ⱥ���0Y�9 u�:��:�Y;v�!;��0;ו:;��@;�BD;e2F;X8G;��G;�H;@@H;�cH;��H;K�H;�H;�H;!�H;c�H;��H;��H;@�H;��H;��H;X�H;��H;�H;B�H;��H;��H;g�H;%�H;�H;�H;I�H;��H;�cH;C@H;�H;��G;[8G;l2F;�BD;��@;ٕ:;��0;z�!;�Y;��:(u�:PY�9���Ⱥg.�3|��R��%Tʻ�����H�	�      �1��$Ȅ�̨u��PV�l.����~W��8��@X�9+i:ܡ�:�+�:�;�t%;�J2;K;;��@;]D;�F;G;W�G;gH;X5H;VZH;xH;�H;��H;�H;�H;,�H;=�H;��H; �H;��H;�H;2�H;��H;/�H;�H;��H;��H;��H;C�H;4�H;�H;�H;��H;�H;
xH;VZH;U5H;jH;Z�G;	G;�F;\D;��@;J;;�J2;�t%;�;�+�:衼:+i:hX�9 ��W�����h.��PV�Ĩu�#Ȅ�      إ��.X��� ��|�=� ۷��ߤ8��:�P�:P�:���:)`;l;�*;�$5;�g<;�<A;�BD;�F;�G;V�G;@�G;y-H;�RH;-qH;��H;��H;S�H;�H;�H;��H;��H;��H;%�H;��H;r�H;j�H;��H;g�H;p�H;��H;"�H;��H;��H;��H;�H;�H;P�H;��H;��H;1qH;�RH;{-H;D�G;Z�G;�G;�F;�BD;�<A;�g<;�$5;�*;r;-`;���:�P�:�P�:��: ߤ8۷���=�� ��.X��      T�:Р:�2<:�)i:<t�:ч�:]�:�+�:�Y;.�;�*';v1;&�8;�Z>;:0B;��D;j2F;G;Z�G;��G;X)H;]NH;JlH; �H;8�H;W�H;q�H;�H;Z�H;��H;�H;��H;�H;/�H;��H;��H;��H;��H;��H;/�H;�H;��H;�H;��H;Z�H;�H;p�H;W�H;=�H;#�H;IlH;^NH;\)H;��G;]�G;G;l2F;��D;;0B;�Z>;&�8;x1;�*';/�;�Y;�+�:W�:߇�:Ht�:X)i:�2<:��:      ��:���:���:d��:�;�Y;�';{�;��(;��0;�Y7;@�<;��@;�`C;CE;�wF;Z8G;b�G;C�G;U)H;�LH;�iH;�H;/�H;x�H;��H;��H;7�H;��H;��H;��H;/�H;��H;r�H;��H;}�H;��H;w�H;��H;q�H;��H;(�H;��H;��H;��H;9�H;��H;��H;~�H;/�H;�H;�iH;�LH;W)H;D�G;\�G;[8G;�wF;CE;�`C;��@;D�<;�Y7;��0;��(;x�;�';�Y;�;d��:��:���:      �;��;;�z ;��$;H�);a/;4;��8;<�<;$@;I�B;!�D;��E;�F;�cG;��G;nH;}-H;^NH;�iH;�H;��H;��H;��H;��H;z�H;w�H;�H;��H;J�H;�H;�H;��H;��H;G�H;��H;A�H;��H;��H;�H;�H;K�H;��H;�H;w�H;w�H;��H;��H;��H;��H;�H;�iH;`NH;}-H;kH;��G;�cG;�F;��E;"�D;O�B;$@;:�<;��8;4;e/;A�);��$;�z ; ;��;      -�1;.J2;5g3;�$5;Y7;��9;Pg<;�>;�A;xC;�D;	�E;I�F;*G;*�G;3�G;�H;_5H;�RH;HlH;	�H;��H;��H;��H;]�H;>�H;3�H;	�H;��H;��H;a�H;��H;^�H;��H;��H;�H;L�H;�H;��H;��H;]�H;��H;d�H;��H;��H;�H;0�H;A�H;c�H;��H;��H;��H;�H;IlH;�RH;Z5H;�H;3�G;+�G;*G;K�F;�E;�D;uC;�A;�>;Ng<;��9;�Y7;�$5;4g3;J2;      6,>;^Z>;��>;��?;K�@;��A;�C;�D;�E;��E;�F;�G;�}G;G�G;��G;�!H;E@H;_ZH;/qH;�H;.�H;��H;��H;��H;��H;��H;�H;��H;��H;��H;<�H;�H;��H;{�H;@�H;��H;��H;��H;=�H;{�H;�H;�H;?�H;��H;��H;��H;�H;��H;��H;�H;��H;��H;/�H;�H;.qH;YZH;E@H;�!H;��G;D�G;�}G;�G;�F;��E;�E;�D;�C;��A;V�@;��?;��>;TZ>;      ��C;'	D;TBD;�D;�	E;��E;RF;�wF;��F;�<G;��G;��G;��G;�H;f4H;�MH;dH;xH;��H;C�H;��H;��H;a�H;��H;"�H;��H;��H;O�H;V�H;��H;��H;Z�H;x�H;3�H;��H;>�H;A�H;8�H;��H;4�H;w�H;T�H;��H;��H;S�H;O�H;��H;��H;%�H;��H;c�H;��H;��H;?�H;��H;xH;dH;�MH;h4H;�H;��G;��G;��G;�<G;��F;�wF;TF;��E;�	E;�D;UBD;'	D;      QwF;FF;}�F;��F;��F;�G;�NG;�G;;�G;��G;��G;7H;o1H;�GH;y\H;\oH;��H;�H;��H;U�H;��H;��H;:�H;��H;��H;A�H;�H;�H;��H;y�H;	�H;H�H;(�H;��H;h�H;��H;��H;��H;e�H;��H;)�H;C�H;�H;y�H;��H;�H;�H;E�H;��H;��H;<�H;��H;��H;T�H;��H;�H;��H;\oH;w\H;�GH;o1H;9H;��G;��G;;�G;�G;�NG;�G;��F;��F;��F;EF;      �G;A�G;�G;�G;#�G;�G;��G;��G;oH;�$H;8H;PJH;�[H;IlH;�{H;M�H;O�H;�H;U�H;r�H;��H;x�H;3�H; �H;��H;�H;��H;X�H;@�H;��H;(�H;�H;��H;~�H;��H; �H;	�H;��H;��H;��H;��H; �H;(�H;��H;=�H;W�H;��H;�H;��H;�H;6�H;{�H;��H;q�H;T�H;��H;P�H;O�H;�{H;FlH;�[H;TJH;8H;�$H;mH;��G;��G;�G;;�G;ߣG;�G;-�G;      n H;�H;hH;zH;�H;C!H;-H;�9H;�FH;BTH;�aH;:oH;E|H;͈H;��H;]�H;�H;�H;�H;�H;:�H;v�H;�H;��H;J�H;
�H;W�H;O�H;��H;��H;��H;��H;o�H;��H;�H;W�H;[�H;S�H;�H;��H;n�H;��H;��H;��H;��H;N�H;S�H;�H;O�H;��H;	�H;v�H;:�H;�H;�H;�H;�H;`�H;��H;͈H;E|H;;oH;�aH;BTH;�FH;�9H;-H;9!H;�H;wH;iH;�H;      �>H;|?H;BH;tFH;�KH;SH;D[H;&dH;�mH;�wH;ԁH;ڋH;��H;ٞH;{�H;��H;"�H;�H;�H;^�H;��H;�H;��H;��H;R�H;�H;9�H;��H;�H;��H;��H;b�H;��H;.�H;h�H;��H;��H;��H;f�H;/�H;��H;^�H;��H;��H;�H;��H;6�H;��H;S�H;��H;��H;�H;��H;Z�H;�H;�H;"�H;��H;{�H;؞H;��H;ًH;ՁH;�wH;�mH;&dH;A[H;SH;LH;tFH;BH;�?H;      �hH;piH;jkH;nnH;�rH;�wH;�}H;T�H;o�H;ΒH;<�H;��H;��H;��H;5�H;h�H;(�H;2�H;��H;��H;��H;��H;}�H;��H;��H;q�H;��H;��H;��H;��H;h�H;��H;�H;t�H;��H;��H;��H;��H;��H;t�H;�H;��H;h�H;��H;��H;��H;��H;u�H;��H;��H;��H;��H;��H;��H;��H;/�H;(�H;k�H;5�H;��H;��H;��H;=�H;ђH;o�H;X�H;�}H;�wH;�rH;pnH;jkH;oiH;      4�H;؈H;5�H;g�H;��H;K�H;��H;��H;��H;�H;��H;�H;c�H;��H;��H;A�H;p�H;H�H;��H;�H;��H;M�H;a�H;=�H;��H;�H;'�H;��H;��H;o�H;��H;'�H;~�H;��H;��H;��H;��H;��H;��H;��H;��H;&�H;��H;k�H;��H;��H;%�H;�H;��H;<�H;g�H;M�H;��H;�H;��H;F�H;r�H;C�H;��H;��H;d�H;�H;��H;��H;��H;��H;��H;A�H;��H;b�H;6�H;؈H;      B�H;��H;��H;C�H;��H;R�H;��H;3�H;�H;"�H;M�H;t�H;��H;x�H;�H;��H;��H;��H;��H;�H;4�H;	�H;��H;�H;X�H;A�H;�H;��H;b�H;��H;!�H;t�H;��H;��H;��H;��H;�H;��H;��H;��H;��H;s�H; �H;��H;`�H;��H; �H;D�H;[�H;�H;��H;�H;2�H;�H;��H;��H;��H;��H;�H;u�H;��H;r�H;Q�H;$�H;�H;7�H;��H;S�H;��H;D�H;��H;��H;      �H;`�H;�H;M�H;�H;�H;��H;E�H;A�H;Z�H;p�H;��H;��H;��H;n�H;6�H;��H;�H;.�H;�H;��H;"�H;^�H;~�H;z�H;%�H;��H;u�H;��H;�H;}�H;��H;��H;��H;�H;�H;��H;�H;�H;��H;��H;��H;{�H;�H;��H;p�H;��H;&�H;|�H;~�H;b�H;"�H;��H;�H;.�H;�H;��H;9�H;n�H;��H;��H;��H;r�H;[�H;F�H;E�H;��H;�H;�H;G�H;�H;^�H;      �H;�H;��H;��H;��H;��H;��H;��H;��H;�H;��H;��H;h�H;��H;-�H;L�H;J�H;�H;��H;7�H;y�H;��H;��H;r�H;0�H;��H;y�H;��H;.�H;x�H;��H;��H;��H;��H;'�H;2�H;�H;0�H;%�H;��H;��H;��H;��H;t�H;+�H;��H;z�H;��H;4�H;q�H;��H;��H;u�H;2�H;��H;�H;N�H;K�H;-�H;��H;g�H;��H;��H;�H;��H;��H;��H;��H;�H;��H;��H;�H;      ��H;��H;O�H;�H;�H;B�H;��H;��H;e�H;p�H;d�H;w�H;v�H;U�H;.�H;��H;��H;�H;w�H;��H;��H;��H;�H;2�H;��H;^�H;��H;�H;i�H;��H;��H;��H;�H;)�H;�H;'�H;F�H;(�H;	�H;+�H;�H;��H;��H;��H;f�H;�H;��H;`�H;��H;3�H;��H;��H;��H;��H;r�H;�H;��H;��H;.�H;T�H;v�H;x�H;g�H;q�H;i�H;��H;��H;D�H;�H;�H;P�H;��H;      �H;5�H;��H;/�H;!�H;L�H;��H;.�H;��H;{�H;/�H;��H;��H;M�H;��H;n�H;��H;3�H;n�H;��H;��H;F�H;��H;��H;7�H;��H;��H;X�H;��H;��H;��H;��H;�H;5�H;)�H;�H;2�H;�H;(�H;7�H;�H;��H;��H;��H;��H;W�H;��H;��H;8�H;��H;�H;C�H;}�H;��H;m�H;5�H;��H;q�H;��H;M�H;��H;��H;2�H;}�H;��H;2�H;��H;O�H;$�H;*�H;��H;C�H;      s�H;��H;=�H;��H;��H;��H;��H;H�H;��H;T�H;�H;��H;R�H;�H;��H;�H;e�H;��H;��H;��H;��H;��H;K�H;��H;?�H;��H;�H;c�H;��H;��H;��H;�H;�H;�H;G�H;0�H; �H;0�H;D�H;�H;�H;�H;��H;��H;��H;_�H;	�H;��H;B�H;��H;P�H;��H;��H;��H;��H;��H;e�H;�H;��H;�H;R�H;��H;�H;U�H;��H;K�H;��H;��H;��H;��H;<�H;��H;      �H;8�H;��H;.�H;!�H;R�H;��H;.�H;��H;{�H;-�H;��H;��H;O�H;��H;n�H;��H;3�H;n�H;��H;��H;G�H;��H;��H;7�H;��H;��H;X�H;��H;��H;��H;��H;�H;6�H;,�H;�H;2�H;�H;(�H;6�H;�H;��H;��H;��H;��H;U�H;��H;��H;8�H;��H;�H;A�H;}�H;��H;m�H;6�H;��H;q�H;��H;L�H;��H;��H;2�H;z�H;��H;2�H;��H;O�H;%�H;1�H;��H;?�H;      ��H;��H;I�H;�H;�H;A�H;��H;��H;e�H;p�H;d�H;w�H;u�H;U�H;0�H;��H;��H;�H;w�H;��H;��H;��H;�H;3�H;��H;]�H;��H;�H;i�H;��H;��H;��H;�H;)�H;�H;(�H;F�H;(�H;�H;+�H;�H;��H;��H;��H;f�H;�H;��H;a�H;��H;2�H;��H;��H;��H;��H;t�H;�H;��H;��H;-�H;T�H;v�H;x�H;d�H;p�H;g�H;��H;��H;A�H;�H;�H;O�H;��H;      �H;�H;��H;��H;��H;��H;��H;��H;��H;�H;��H;��H;g�H;��H;.�H;L�H;M�H;�H;��H;6�H;y�H;��H;��H;u�H;3�H;��H;z�H;��H;/�H;x�H;��H;��H;��H;��H;)�H;0�H;�H;0�H;'�H;��H;��H;��H;��H;t�H;*�H;��H;z�H;��H;2�H;m�H;��H;��H;q�H;2�H;��H;�H;M�H;L�H;-�H;��H;g�H;��H;��H;�H;��H;��H;��H;��H;�H;��H;��H;�H;       �H;d�H;�H;J�H;�H;�H;��H;H�H;C�H;[�H;p�H;��H;��H;��H;r�H;7�H;��H;�H;.�H;�H;��H;#�H;]�H;��H;|�H;#�H;��H;u�H;��H;!�H;}�H;��H;��H;��H;�H;	�H;��H;�H;�H;��H;��H;��H;}�H;�H;��H;o�H;��H;&�H;z�H;}�H;e�H;"�H;��H;
�H;.�H;�H;��H;7�H;n�H;��H;��H;��H;p�H;Z�H;F�H;H�H;��H;�H;�H;O�H;!�H;^�H;      7�H;��H;��H;D�H;��H;a�H;��H;5�H;�H;"�H;N�H;t�H;��H;w�H; �H;��H;��H;��H;��H;�H;7�H;�H;��H;�H;\�H;C�H; �H;��H;e�H;��H;!�H;s�H;��H;��H;��H;��H;�H;��H;��H;��H;��H;s�H;�H;��H;`�H;��H; �H;F�H;X�H;�H;��H;�H;/�H;�H;��H;��H;��H;��H;�H;u�H;��H;t�H;M�H;$�H;�H;6�H;��H;V�H;��H;F�H;��H;��H;      )�H;؈H;6�H;b�H;��H;L�H;��H;��H;��H;�H;��H;��H;c�H;��H;��H;C�H;q�H;H�H;��H;�H;��H;O�H;b�H;?�H;��H;�H;%�H;��H;��H;o�H;��H;'�H;�H;��H;��H;��H;��H;��H;��H;��H;��H;'�H;��H;l�H;��H;��H;%�H;�H;��H;9�H;h�H;N�H;��H;�H;��H;F�H;t�H;C�H;��H;��H;c�H;��H;��H;�H;��H;��H;��H;I�H;��H;l�H;<�H;׈H;      �hH;tiH;dkH;znH;�rH;�wH;�}H;]�H;r�H;ђH;<�H;��H;��H;��H;6�H;i�H;(�H;2�H;��H;��H;��H;��H;}�H;��H;��H;q�H;��H;��H;��H;��H;h�H;��H;�H;t�H;��H;��H;��H;��H;��H;t�H;�H;��H;h�H;��H;��H;��H;��H;x�H;��H;��H;��H;��H;��H;��H;��H;/�H;(�H;k�H;5�H;��H;��H;��H;=�H;ђH;o�H;[�H;�}H;�wH;�rH;~nH;nkH;piH;      �>H;|?H;#BH;rFH;�KH;SH;A[H;'dH;�mH;�wH;ҁH;ۋH;��H;ܞH;�H;��H;!�H;�H;�H;\�H;�H;�H;��H;��H;V�H;}�H;6�H;��H;�H;��H;��H;b�H;��H;.�H;h�H;��H;��H;��H;f�H;.�H;��H;a�H;��H;��H;�H;��H;7�H;��H;P�H;��H;��H;�H;��H;[�H;�H;�H;!�H;��H;|�H;؞H;��H;׋H;ԁH;�wH;�mH;,dH;E[H;SH;LH;pFH;#BH;z?H;      { H;�H;^H;yH;�H;N!H;-H;�9H;�FH;CTH;�aH;;oH;H|H;ΈH;��H;`�H;�H;�H;�H;�H;=�H;y�H;�H;��H;P�H;�H;T�H;N�H;��H;��H;��H;��H;k�H;��H;�H;T�H;\�H;U�H;�H;��H;o�H;��H;��H;��H;��H;K�H;U�H;�H;J�H;��H;�H;w�H;9�H;�H;�H;�H;�H;^�H;��H;̈H;E|H;:oH;�aH;BTH;�FH;�9H;-H;>!H;�H;wH;hH;�H;      ��G;K�G;ܔG;��G;2�G;�G;��G;��G;rH;�$H;8H;UJH;�[H;HlH;�{H;N�H;R�H;�H;W�H;q�H;��H;}�H;2�H;%�H;��H;�H;��H;X�H;@�H;��H;'�H;�H;��H;~�H;��H;��H;�H;��H;��H;~�H;��H;�H;(�H;��H;;�H;W�H;��H;�H;��H;�H;7�H;{�H;��H;t�H;U�H;��H;P�H;O�H;�{H;FlH;�[H;RJH;8H;�$H;oH;��G;��G;�G;9�G;�G;ߔG;6�G;      EwF;FF;��F;��F;��F;�G;�NG;�G;=�G;��G;��G;;H;p1H;�GH;z\H;^oH;��H;�H;��H;U�H;��H;��H;:�H;��H;��H;?�H;�H;�H;��H;x�H;	�H;G�H;&�H;��H;g�H;��H;��H;��H;b�H;��H;&�H;F�H;	�H;x�H;��H;�H;�H;E�H;��H;��H;<�H;��H;��H;U�H;��H;�H;��H;]oH;|\H;�GH;o1H;9H;��G;��G;5�G;
�G;�NG;�G;��F;��F;n�F;8F;      ��C;%	D;PBD;�D;�	E;��E;UF;�wF;��F;�<G;��G;��G;��G;�H;i4H;�MH;dH;xH;ÉH;B�H;��H;��H;a�H;��H;'�H;��H;��H;O�H;V�H;��H;��H;Z�H;u�H;3�H;��H;;�H;?�H;:�H;��H;3�H;w�H;X�H;��H;��H;R�H;L�H;��H;��H;"�H;��H;d�H;��H;��H;@�H;ÉH;xH;dH;�MH;j4H;�H;��G;��G;��G;�<G;��F;�wF;QF;��E;�	E;�D;PBD;$	D;      ,>;HZ>;��>;��?;D�@;��A;�C;�D;�E;��E;�F;�G;�}G;E�G;��G;�!H;F@H;`ZH;1qH;�H;2�H;��H;��H;��H;��H;��H;�H;��H;��H;��H;=�H;�H;��H;z�H;=�H;��H;��H;��H;:�H;w�H;��H;�H;@�H;��H;��H;��H;�H;��H;��H;��H;��H;��H;0�H; �H;1qH;[ZH;F@H;�!H;��G;E�G;�}G;�G;�F;��E;�E;�D;�C;��A;Z�@;ɯ?;��>;.Z>;      �1;(J2;)g3;�$5;|Y7;��9;Jg<; �>;�A;xC;�D;�E;I�F;*G;.�G;5�G;�H;a5H;�RH;IlH;�H;��H;��H;��H;c�H;:�H;3�H;�H;��H;}�H;b�H;��H;]�H;��H;��H;�H;N�H;�H;��H;��H;]�H;��H;e�H;��H;��H;�H;4�H;>�H;^�H;��H;��H;��H;�H;IlH;�RH;Z5H;�H;3�G;.�G;*G;I�F;	�E;�D;vC;�A; �>;Ig<;��9;|Y7;�$5;)g3;J2;      �;��;�
;�z ;��$;N�);g/;4;��8;:�<;$@;R�B;"�D;��E;�F;�cG;��G;oH;}-H;aNH;�iH;�H;��H;��H;��H;��H;z�H;w�H;�H;��H;J�H;�H;�H;��H;��H;C�H;��H;D�H;��H;��H;�H;�H;M�H;��H;�H;w�H;z�H;��H;��H;��H;��H;�H;�iH;aNH;}-H;kH;��G;�cG;�F;��E;!�D;N�B; $@;8�<;��8;4;`/;7�);��$;�z ; ;��;      ��:!��:��:v��:�;�Y;�';|�;��(;��0;�Y7;D�<;��@;�`C;CE;�wF;]8G;a�G;E�G;X)H;�LH;�iH;�H;0�H;~�H;��H;��H;7�H;��H;��H;��H;-�H;��H;q�H;��H;x�H;��H;z�H;��H;m�H;��H;*�H;��H;��H;��H;7�H;��H;��H;z�H;0�H;	�H;�iH;�LH;X)H;D�G;\�G;[8G;�wF;CE;�`C;��@;B�<;�Y7;��0;��(;�;�';�Y;�;n��:(��:���:      ��:�:�2<:�)i:Bt�:݇�:a�:�+�:�Y;0�;�*';x1;'�8;�Z>;;0B;�D;l2F;G;\�G;��G;^)H;aNH;JlH;!�H;=�H;U�H;p�H;�H;\�H;��H;�H;��H;�H;2�H;��H;��H;��H;��H;��H;,�H;�H;��H;�H;��H;[�H;�H;q�H;W�H;9�H;#�H;JlH;^NH;[)H;��G;\�G;
G;l2F;��D;;0B;�Z>;&�8;w1;�*';,�;�Y;�+�:Y�:ˇ�:Jt�:|)i:�2<:Р:      ֥��*X��� ��l�=�8۷��ߤ8��:�P�:�P�:���:)`;r; �*;�$5;�g<;�<A;�BD;�F;�G;Z�G;G�G;}-H;�RH;.qH;��H;��H;Q�H;�H;�H;��H;��H;��H;'�H;��H;r�H;h�H;��H;h�H;p�H;��H;$�H;��H;��H;��H;�H;�H;S�H;��H;��H;/qH;�RH;z-H;C�G;Z�G;�G;�F;�BD;�<A;�g<;�$5;�*;n;)`;~��:�P�:�P�:��:@ߤ8@۷�|�=�� �� X��      �1��Ȅ�Шu��PV�i.����|W�����hX�9+i:ࡼ:�+�:�;�t%;�J2;O;;��@;\D;�F;	G;\�G;jH;\5H;XZH;xH;�H;��H;�H;�H;,�H;A�H;��H; �H;��H;�H;0�H;��H;0�H;�H;��H; �H;��H;A�H;2�H;�H;�H;��H;�H;xH;VZH;[5H;hH;W�G;	G;�F;YD;��@;K;;�J2;�t%;�;�+�:桼:+i:`X�9��W�����l.��PV�٨u�Ȅ�      W��J�	������ Tʻ�R��3|�e.�Ⱥ���8Y�9,u�:��:�Y;|�!;��0;ٕ:;��@;�BD;j2F;_8G;��G;�H;C@H;�cH;��H;I�H;�H;�H; �H;g�H;��H;��H;B�H;��H;��H;Z�H;��H;�H;@�H;��H;��H;g�H;$�H;�H;�H;I�H;��H;�cH;B@H;�H;��G;W8G;j2F;�BD;��@;ؕ:;��0;z�!;�Y;��:&u�:8Y�9���Ⱥh.�3|��R��&Tʻ�����H�	�      ��x��[t���g�LT�]�:�������$����1��K�(�&W��@�t��n`:[��:�\;{ ;��0;O;;�<A;��D;�wF;�cG;3�G;�!H;�MH;ZoH;H�H;Z�H;��H;e�H;<�H;��H;-�H;E�H;��H;j�H;��H;j�H;��H;A�H;*�H;��H;:�H;h�H;��H;\�H;H�H;UoH;�MH;�!H;3�G;�cG;�wF;��D;�<A;K;;��0;{ ;�\;[��:�n`:��t�*W��L�(��1��&���������`�:�NT���g��[t�      5,˼��Ǽ�"���뮼w��"G��)�[�]y-�����.����b�l0㺀ط�5<:�L�:�\;x�!;�J2;�g<;40B;CE;�F;.�G;��G;e4H;y\H;�{H;��H;|�H;0�H;��H;�H;h�H;&�H;%�H;��H;�H;��H;#�H;$�H;g�H;�H;��H;2�H;|�H;��H;�{H;r\H;^4H;��G;+�G;�F;CE;60B;�g<;�J2;v�!;�\;�L�:5<:�ط�n0���b��.�����]y-�)�[�#G��w���뮼�"����Ǽ      *���k��Jv�|t�B�Ѽ�뮼+X��k�W������׻�Ǆ������5<:a��:�Y;�t%;�$5;�Z>;�`C;��E;*G;E�G;�H;�GH;FlH;ʈH;ٞH;��H;��H;n�H;��H;��H;J�H;B�H; �H;F�H;F�H;��H;��H;k�H;��H;��H;ٞH;ɈH;ClH;�GH;�H;E�G;*G;��E;�`C;�Z>;�$5;�t%;�Y;U��:5<:������Ǆ���׻���k�W�+X���뮼B�Ѽ}t�Jv���k�      Bm��Fi��&^�^�L�N�6�'����}ռmT����x���0���������`ط�o`:��:�;�*;#�8;�@;!�D;K�F;�}G;��G;n1H;�[H;E|H;��H;��H;\�H;��H;��H;`�H;h�H;��H;D�H;��H;e�H;]�H;��H;��H;Z�H;��H;��H;E|H;�[H;h1H;z�G;�}G;K�F;�D;��@;$�8;�*;�;��:�n`:�ط��������껽�0���x�lT��}ռ��'��P�6�^�L��&^��Fi�      K��r;��@�������섽w�e��?��k�zt�鷼G���e7�����Ǆ�d0㺀�t�$u�:�+�:n;t1;I�<;L�B;	�E;�G;��G;3H;QJH;3oH;׋H;��H;�H;k�H;��H;��H;j�H;��H;��H;��H;g�H;��H;��H;j�H;�H;��H;ًH;3oH;PJH;0H;��G;�G;
�E;K�B;>�<;v1;l;�+�: u�:��t�h0��Ǆ���껂e7�G��鷼zt��k��?�w�e��섽���@���r;��      n���$��s��ӽ�'��?������
�Z��Q+�����"��G����0���׻b�0W���X�9ԡ�: `;�*';�Y7;�#@;
�D;�F;��G;��G;8H;�aH;сH;6�H;}�H;J�H;k�H;y�H;W�H;%�H;�H;#�H;W�H;x�H;h�H;F�H;y�H;:�H;ҁH;�aH;8H;��G;�G;�F;
�D;�#@;�Y7;�*';`;Ρ�: Y�96W��ƕb���׻��0�G���"������Q+�
�Z����?����'���ӽ�s�$��      �!,�7)��K ��������޽������Fi��0����鷼��x�����.��L�(���� +i:~��:+�;��0;:�<;tC;��E;�<G;��G;�$H;:TH;�wH;ʒH;�H; �H;X�H;�H;d�H;p�H;M�H;o�H;c�H;�H;U�H;�H;�H;̒H;�wH;;TH;�$H;��G;�<G;��E;uC;6�<;��0;,�;x��:�*i:���O�(��.�������x�鷼����0��Fi�������޽�������K �7)�      (�j��f��Z�y�F��>/��^�m�����ŽF ���Fi��Q+�zt�lT��l�W�����1�� ȺX�9}P�:�Y;��(;��8;�A;�E;��F;9�G;sH;�FH;�mH;m�H;��H;�H;H�H;��H;^�H;��H;��H;��H;^�H;��H;D�H;�H;��H;n�H;�mH;�FH;sH;9�G;��F;�E;�A;��8;~�(;�Y;uP�:X�9"Ⱥ�1�����l�W�mT��zt�Q+��Fi�F ����Žm����^��>/�y�F��Z��f�      ��v���x�G����f��SC��K �mn����Ž���
�Z��k�}ռ,X��_y-�(���n.����P�:�+�:��;4;�>;�D;�wF;�G;��G;�9H;'dH;T�H;��H;3�H;H�H;��H;~�H;(�H;D�H;(�H;~�H;��H;E�H;/�H;��H;[�H;)dH;�9H;��G;�G;�wF;�D;�>;4;y�;�+�:�P�:`��m.�*���_y-�,X��}ռ�k�
�Z������Žmn���K ��SC��f�G���x�v���      ��˾��Ǿ���� ���V͓�Y�x���J��K �m���������?����뮼)�[����3|��W����:C�:�';d/;=g<;�C;GF;�NG;��G;-H;=[H;�}H;��H;��H;��H;�H;��H;��H;��H;��H;��H;�H;��H;��H;��H;�}H;>[H;
-H;��G;�NG;FF;�C;Bg<;a/;�';I�:��:�W��3|����)�[��뮼���?������l����K ���J�Z�x�V͓� ���������Ǿ      s� ��������{Ծj���v���Y�x��SC��^��޽?���w�e�'��B�Ѽ#G������R�����@ޤ8ˇ�:�Y;E�);��9;��A;��E;�G;�G;A!H;
SH;�wH;L�H;\�H;�H;��H;I�H;S�H;��H;S�H;I�H;��H;�H;Z�H;H�H;�wH;SH;C!H;�G;�G;��E;��A;��9;D�);�Y;χ�: ޤ8����R�����#G��B�Ѽ'��w�e�?����޽�^��SC�Y�x�v���j����{Ծ�쾠���      ����D�l�s� �V�ݾj���V͓��f��>/�����'���섽O�6�~t�w��\�:�$Tʻ|.� ۷�Ft�:�;��$;�Y7;R�@;�	E;��F;)�G;�H;	LH;�rH;��H;��H;��H;��H;�H;$�H;��H; �H;�H;�H;��H;��H;��H;�rH;
LH;�H;0�G;��F;�	E;S�@;�Y7;��$;�;Jt�:(۷�x.�%Tʻ]�:�w��~t�O�6��섽�'������>/��f�V͓�j���V�ݾs� �l��D�      �7�v3�/�'����s� ��{Ծ���H���y�F�����ӽ���]�L�Iv��뮼OT����PV���=�l)i:���:�z ;}$5;��?;�D;��F;�G;rH;eFH;rnH;d�H;M�H;K�H;��H;�H;1�H;��H;-�H;�H;��H;K�H;M�H;a�H;|nH;fFH;sH;�G;��F;�D;��?;{$5;�z ;v��:�)i:��=��PV���OT��뮼Iv�]�L�����ӽ���y�F�H��� ����{Ծs� ����/�'�v3�      �N��TI���;�/�'�l��쾀���x󐾲Z��K ��s�@����&^���"����g����̨u�� ���2<:"��:�
;8g3;��>;WBD;t�F;ߔG;kH;BH;^kH;/�H;��H;	�H;��H;B�H;��H;"�H;��H;B�H;��H;�H;��H;+�H;ekH;BH;lH;�G;��F;WBD;��>;4g3;�
;��:�2<:� ��̨u������g��"����&^�@����s潥K ��Z�x󐾀�����l�/�'���;��TI�      `]�d�W��TI�v3��D�������Ǿv����f�7)�$��r;���Fi��k���Ǽ�[t�L�	�)Ȅ�X��ܠ:��:��;,J2;SZ>;'	D;:F;8�G;�H;�?H;viH;ÈH;��H;S�H;�H;��H;5�H;��H;1�H;��H;�H;Q�H;��H;��H;~iH;�?H;�H;>�G;IF;%	D;SZ>;&J2;��;��:�:X��(Ȅ�L�	��[t���Ǽ�k��Fi�r;��$��7)��f�v�����Ǿ�����D�v3��TI�d�W�      1�$��� ����#��?��'�þ�*��0Dx���=�����Pν���#'K��c���n�V����E^���S��w[:���:e;)�4;E`?;�mD;R�F;LvG;�G;=H;aOH;�sH;��H;|�H;��H;�H;U�H;&�H;O�H;�H;��H;{�H;��H;�sH;mOH;=H;�G;QvG;a�F;�mD;D`?;%�4;e;���:�w[:��S�
E^����n�V����c�#'K�����Pν�����=�0Dx��*��'�þ?��#������� �      �� ����R��O��/������0��4�s�ր:�g9��ʽ1Z����G��8�
.���5S�����/X�p�D�rBd:�B�: ;��4;ʈ?;�~D;�F;yG;��G;M H;*PH;tH;�H;΢H;ưH;,�H;r�H;5�H;n�H;,�H;ưH;̢H;�H;tH;3PH;O H;��G;yG;�F;�~D;ʈ?;��4; ;�B�:�Bd:l�D��/X���껬5S�
.���8���G�0Z���ʽg9�ր:�4�s��0�����/��O��R�����      ���R��8�
������Yؾ���ޥ����f���0�Z[�N8��ΐ���>�����IȤ��6H�_�ܻrF�����}:��:d";/�5;��?;T�D;��F;	�G;��G;/#H;`RH;�uH;F�H;ģH;v�H;źH;�H;��H;�H;ĺH;v�H;��H;F�H;�uH;iRH;0#H;��G;�G;��F;V�D;��?;)�5;b";��:,�}:���rF�_�ܻ�6H�HȤ������>�ϐ��N8��Z[���0���f�ޥ������Yؾ����8�
�Q��      #��O������>I�(�þ�R��;���tS��Q"��s������}��0��켈�����6�D�ƻ6}*�������:}x;Z%;�l7;ڳ@;��D;��F;��G;��G;�'H;�UH;]xH;N�H;F�H;��H;��H;��H;z�H;��H;��H;��H;D�H;M�H;XxH;�UH;�'H;��G;��G;��F;��D;ܳ@;�l7;X%;}x;��:����4}*�D�ƻ��6��������0���}�����s��Q"�tS�;����R��(�þ=Iᾣ���O��      ?��/�待Yؾ(�þĪ�|쏾�k�ր:�~�z�ؽ�����c�\y���Ҽ����B� �h�(�� #(7E�:��
;��(;�_9;��A;h\E;l�F;��G;��G;�.H;�ZH;�{H;�H;I�H;P�H;�H;��H;x�H;��H;�H;Q�H;H�H;�H;�{H;�ZH;�.H;��G;��G;x�F;j\E;��A;}_9;��(;��
;S�: #(7(��h�B� �������Ҽ\y��c�����{�ؽ~�ր:��k�|쏾Ī�(�þ�Yؾ/��      '�þ��� ����R��|쏾4�s��H�����������ΐ����D��c�����:�f�R,�����P��X�9˳�:�;"j-;M�;;u�B;��E;[G;��G;��G;�6H;�`H;W�H;L�H;թH;N�H;��H;R�H;��H;N�H;��H;M�H;ҩH;L�H;V�H;�`H;�6H;��G;��G;dG;��E;s�B;L�;;"j-;�;ճ�:`�9�P�����R,�:�f������c���D�ΐ�������������H�4�s�|쏾�R�� ������      �*���0��ޥ��;����k��H��#%�Z[��Pνt��`�f�2/%���伅���s�=��?ػ�FL���D�l�R:��:4�;42;��=;��C;f0F;FGG;��G;#H;�?H;�gH;��H;,�H;��H;��H;��H;��H;r�H;��H;��H;��H;��H;*�H;��H;�gH;�?H;#H;��G;MGG;i0F;��C;��=;62;2�;��:l�R:��D��FL��?ػs�=��������1/%�`�f�t���PνZ[��#%��H��k�;���ޥ���0��      0Dx�4�s���f�tS�ր:����Z[��7ս�榽��}���;��8�T�����r����8G�����̬�)��:	�;�}$;Ä6;�?;��D;ƔF;�pG;��G;�H; JH;>oH;;�H;v�H;��H;6�H;��H;��H;&�H;��H;��H;9�H;��H;s�H;9�H;GoH;$JH;�H;��G;�pG;ʔF;��D;�?;Ƅ6;�}$;�;)��:�̬���8G�������r�T����8���;���}��榽�7սZ[����׀:�sS���f�4�s�      ��=�ր:���0��Q"�~������Pν�榽?����G�1����Ҽ ��GE:�:�ܻ�D^�����li:A��:�;8|,;��:;K�A;AiE;��F;�G;�G;�(H;2UH;{wH;o�H;!�H;��H;�H;��H;��H;�H;��H;��H;�H;��H;#�H;o�H;�wH;5UH;�(H;��G;�G;��F;?iE;N�A;��:;8|,;�;G��:hi:�����D^�8�ܻGE:� ����Ҽ1����G�?���榽�Pν����~��Q"���0�ր:�      ���g9�Z[��s�z�ؽ���t����}���G�����0c��V�V�D,��*����������:��:Q ;c�3;�0>;ÚC;�F;�8G;*�G;kH;�7H;�`H;�H;�H;��H;K�H;��H;G�H;��H;�H;��H;G�H;��H;G�H;��H;�H;�H;�`H;�7H;lH;*�G;�8G;�F;ƚC;�0>;b�3;X ;��:��:�������*��D,�U�V�/c��������G���}�t�����{�ؽ�s�Z[�g9�      �Pν�ʽN8���������ΐ��`�f���;�1����BȤ�2�f�(��Jߵ�Ro5���D�<�-:H��:�>;�+;�_9;�A;c�D; �F;�vG;��G;H;uGH;ZlH;��H;��H;��H;,�H;��H;��H;�H;"�H;�H;��H;��H;*�H;�H;��H;ǈH;`lH;yGH;!H;��G;�vG; �F;h�D;�A;�_9;�+;�>;F��:L�-:��D�Po5�Hߵ�'��1�f�AȤ���1����;�`�f�ΐ���������N8���ʽ      ���1Z��ΐ����}��c���D�1/%��8���Ҽ/c��1�f�����ƻ|/X�V������9�:=�;�";��3;=>;?YC;r�E;�G;�G;c�G;�,H;WH;xH;��H;/�H;�H;�H;��H;0�H;D�H;-�H;B�H;0�H;��H;�H;�H;2�H;��H;xH;WH;�,H;c�G;�G;�G;y�E;FYC;?>;��3;�";=�;�:���9R���x/X��ƻ���0�f�0c����Ҽ�8�1/%���D��c���}�ϐ��0Z��      #'K���G��>��0�\y��c����S��� ��U�V�'���ƻ�od�~�º (7�4�:���:��;�P.;ҡ:;zA;,�D;ƨF;MnG;8�G;�H;�@H;$fH;]�H;.�H;��H;ԸH;��H;��H;��H;{�H;6�H;z�H;��H;��H;��H;иH;��H;5�H;c�H;%fH;�@H;�H;?�G;NnG;ʨF;0�D;zA;ݡ:;�P.;��;���:�4�: �(7t�º�od��ƻ'��U�V� ��S�����伔c�]y��0��>���G�      �c��8���������Ҽ����������r�GE:�C,�Hߵ�~/X���º�Ƭ�p�}:�:�;K�);%m7;�?;��C;F;U)G;�G;E�G;�)H;�SH;�tH;\�H;|�H;�H;��H;��H;��H;�H;��H;J�H;��H;�H;��H;��H;��H;�H;��H;f�H;�tH;�SH;�)H;L�G;�G;\)G;
F;��C;�?;(m7;H�);�;�:|�}:@Ƭ�~�ºx/X�Fߵ�C,�EE:���r�����������Ҽ�켶����8�      ��
.��JȤ���������:�f�s�=����:�ܻ�*��Mo5�`��� ~(7x�}:�n�:-�;�>&;��4;��=;��B;�E;�F;��G;��G;+H;�AH;�eH;<�H;јH;Y�H;ڷH;i�H;�H;��H;j�H;��H;N�H;��H;h�H;��H;�H;c�H;ݷH;_�H;ؘH;A�H;�eH;~AH;/H;��G;��G;�F;�E;��B;��=;��4;�>&;,�;�n�:��}: �(7T���Jo5��*��6�ܻ���s�=�8�f���������JȤ�
.��      h�V��5S��6H���6�B� �S,��?ػ6G���D^������D����9�4�:�:,�;�%;��3; �<;XB;�E;��F;�XG;��G;E H;h0H;LWH;YvH;�H;{�H;��H;��H;��H;o�H;M�H;��H;��H;7�H;��H;��H;N�H;l�H;��H;��H;ñH;�H;�H;[vH;GWH;l0H;F H; �G;�XG;�F;�E;YB;�<;��3;�%;.�;�:�4�:���9��D�����D^�4G���?ػP,�E� ���6��6H��5S�      ��ﻪ��d�ܻF�ƻd󩻶���FL�������@��X�-:	�:���:�;�>&;��3;T9<;�A;۰D;AZF;5G;��G;��G;i!H;,JH;/kH;��H;��H;c�H;��H;��H;��H;��H;��H;��H;c�H;��H;_�H;��H;��H;��H;��H;��H;��H;g�H;��H;��H;*kH;2JH;l!H;��G;��G;!5G;HZF;ްD;�A;W9<;��3;�>&;�;���:�:d�-:@����������FL����h�I�ƻi�ܻ���      �D^��/X�rF�*}*����P��|�D� ̬�ti:��:P��:7�;��;H�);��4;�<;�A;&�D;v9F;�G;m�G;C�G;=H;?H;ZaH;}H;|�H;v�H;��H;�H;��H;b�H;�H;�H;��H;(�H;��H;%�H;��H;�H;{�H;]�H;��H;�H;��H;v�H;{�H;}H;_aH;?H;:H;F�G;q�G;�G;w9F;#�D;�A;�<;��4;H�);��;:�;^��:��:�i:�ˬ���D��P����2}*��qF��/X�      0�S���D����Ȇ�� $(7��9��R:3��:I��: ��:�>;�";�P.;*m7;��=;YB;ݰD;~9F;G;�G;R�G;�H;�6H;iYH;�uH;�H;�H;��H;��H;��H;�H;��H;�H;8�H;a�H;��H;��H;��H;^�H;6�H;�H;��H; �H;��H;��H;��H;�H;�H;�uH;lYH;�6H;�H;W�G;�G; G;y9F;�D;VB;��=;*m7;�P.;�";�>;��:O��:3��:��R:��9 &(70��������D�      �w[:nBd:<�}:��:=�:ճ�:�:�;�;Z ;�+;��3;ܡ:;�?;��B;�E;HZF;�G;�G;o�G;>H;S1H;�SH;`pH;ׇH;H�H;�H;{�H;��H;��H;��H;��H;r�H;"�H;��H;�H;\�H;�H;��H;!�H;p�H;��H;��H;��H;��H;|�H;�H;G�H;ۇH;bpH;�SH;U1H;DH;r�G; �G;�G;HZF;�E;��B;�?;ܡ:;��3;�+;Z ;�;�;�:��:I�:��:�}:2Bd:      *��:�B�:���:ox;��
;�;3�;�}$;8|,;e�3;�_9;:>;zA;��C;�E;�F;5G;x�G;W�G;=H;�/H;�PH;mH;H�H;��H;��H;n�H;��H;��H;�H;\�H;��H;��H;��H;k�H;L�H;��H;D�H;j�H;��H;��H;��H;^�H;�H;��H;��H;i�H;��H;��H;H�H;�lH;�PH;�/H;?H;X�G;t�G;"5G;�F;�E;��C;zA;?>;�_9;e�3;6|,;�}$;9�;�;��
;px;ֆ�:�B�:      
e; ;q";h%;��(;$j-;42;Ä6;��:;�0>;�A;AYC;0�D;F;�F;�XG;��G;L�G;�H;T1H;�PH;�kH;t�H;{�H;1�H;,�H;׼H;��H;��H;�H;m�H;��H;v�H;p�H;��H;a�H;��H;[�H;��H;p�H;u�H;��H;n�H;�H;��H;��H;ӼH;.�H;5�H;{�H;p�H;�kH;�PH;U1H;�H;I�G;��G;�XG;�F;
F;1�D;HYC;�A;�0>;��:;ʄ6;82;j-; �(;\%;g"; ;      B�4;��4;(�5;�l7;{_9;W�;;��=;�?;X�A;͚C;q�D;{�E;ͨF;b)G;��G;�G;��G;EH;�6H;�SH;�lH;r�H;��H;�H;��H;O�H;#�H;2�H;��H;��H;�H;��H;2�H;��H;��H;b�H;��H;[�H;��H;��H;2�H;��H;�H;�H;��H;3�H;�H;P�H;��H;�H;��H;u�H;mH;�SH;�6H;?H;��G;�G;��G;])G;ͨF;��E;t�D;ʚC;X�A;�?;��=;S�;;�_9;�l7;(�5;��4;      E`?;Ԉ?;��?;ֳ@;��A;w�B;��C;�D;8iE;�F;#�F;�G;NnG;�G;��G;I H;l!H;?H;lYH;[pH;E�H;w�H;�H;C�H;��H;%�H;C�H;�H;��H;s�H;S�H;��H;��H;��H;��H;<�H;M�H;5�H;��H;��H;��H;��H;V�H;r�H;��H;�H;?�H;(�H;��H;A�H;�H;z�H;F�H;]pH;jYH;?H;l!H;K H;��G;�G;KnG;�G;&�F;�F;?iE;��D;��C;h�B;��A;ӳ@;��?;ˈ?;      �mD;�~D;S�D;��D;a\E;��E;r0F;ǔF;��F;�8G;�vG;�G;@�G;Q�G;2H;r0H;7JH;haH;�uH;��H;��H;5�H;��H;��H;��H;��H;j�H;�H;��H;��H;\�H;A�H;��H;��H;��H;��H;)�H;��H;��H;��H;��H;;�H;_�H;��H;��H;�H;d�H;��H;��H;��H;��H;6�H;��H;އH;�uH;eaH;9JH;u0H;2H;M�G;@�G;��G;�vG;�8G;��F;ʔF;u0F;��E;o\E;��D;V�D;�~D;      M�F;�F;��F;��F;l�F;dG;PGG;�pG;�G;4�G;��G;i�G;�H;*H;�AH;PWH;2kH;}H;�H;D�H;��H;(�H;K�H;%�H;��H;/�H;��H;�H;��H;�H;�H;��H;��H;��H;:�H;��H;��H;��H;7�H;��H;��H;��H;�H;�H;��H;�H;��H;3�H;��H;"�H;L�H;)�H;��H;D�H;�H;}H;3kH;NWH;�AH;*H;�H;j�G;��G;2�G;�G;�pG;QGG;[G;��F;��F;��F;�F;      dvG;yG;
�G;��G;��G;��G;��G;��G;~�G;lH;!H;�,H;�@H;�SH;�eH;]vH;��H;��H;�H;�H;p�H;ּH;#�H;D�H;g�H;��H;c�H;]�H;��H;��H;^�H;��H;��H;@�H;��H;&�H;#�H;�H;��H;B�H;��H;��H;`�H;��H;��H;\�H;^�H;��H;k�H;@�H;#�H;׼H;r�H;�H;�H;|�H;��H;]vH;�eH;�SH;�@H;�,H;!H;kH;}�G;��G;��G;��G;˝G;��G;�G; yG;      �G;��G;��G;��G;��G;��G;1H;�H;�(H;�7H;yGH;WH;$fH;�tH;=�H;�H;��H;v�H;��H;y�H;��H;��H;-�H;�H;�H;}�H;]�H;��H;��H;d�H;��H;��H;U�H;��H;O�H;��H;��H;��H;M�H;��H;W�H;��H;��H;e�H;��H;��H;X�H;�H;�H;�H;0�H;��H;��H;y�H;��H;t�H;��H;�H;<�H;�tH;$fH;
WH;|GH;�7H;�(H;�H;3H;��G;��G;��G;��G;��G;      :H;E H;,#H;(H;w.H;�6H;�?H; JH;.UH;�`H;alH;xH;a�H;b�H;֘H;�H;j�H;��H;�H;��H;��H;��H;��H;��H;��H;��H;��H;��H;1�H;��H;��H;O�H;��H;s�H;��H;��H;��H;��H;��H;u�H;��H;I�H;��H;��H;3�H;��H;��H;��H;��H;��H;��H;��H;��H;��H;�H;��H;j�H;��H;֘H;`�H;`�H;xH;blH;�`H;.UH; JH;�?H;6H;�.H; (H;-#H;I H;      cOH;%PH;kRH;�UH;�ZH;�`H;�gH;@oH;�wH;�H;ǈH;��H;3�H;��H;[�H;��H;��H;�H;��H;��H;�H;	�H;z�H;n�H;��H;	�H;��H;d�H;��H;��H;I�H;��H;e�H;��H;��H;�H;4�H;�H;��H;��H;g�H;��H;H�H;��H;��H;d�H;��H;�H;��H;k�H;~�H;�H;�H;��H;��H;�H;��H;��H;Y�H;��H;3�H;��H;ǈH;�H;wH;EoH;�gH;�`H;�ZH;�UH;nRH;"PH;      �sH;-tH;�uH;`xH;�{H;X�H;��H;;�H;s�H;�H;��H;9�H;��H;��H;�H;��H;��H;��H;&�H;�H;d�H;p�H;�H;S�H;\�H;�H;`�H;��H;��H;O�H;��H;k�H;��H;�H;X�H;c�H;[�H;_�H;U�H;�H;��H;h�H;��H;L�H;��H;��H;[�H;�H;a�H;R�H;�H;n�H;a�H;��H;%�H;��H;��H;��H;�H;��H;��H;;�H;��H;�H;t�H;@�H;��H;P�H;�{H;^xH;�uH;.tH;      ��H;�H;F�H;D�H;�H;B�H;4�H;w�H;(�H;��H;��H;�H;۸H;��H;i�H;��H;��H;g�H;��H;��H;��H;��H;��H;��H;@�H;��H;��H;��H;L�H;��H;e�H;��H;�H;Z�H;��H;�H;��H;�H;��H;[�H;�H;��H;d�H;��H;K�H;��H;��H;��H;B�H;��H;��H;��H;��H;��H;��H;i�H;��H;��H;i�H;��H;ڸH;�H;��H;��H;(�H;|�H;:�H;E�H;��H;G�H;O�H;�H;      ��H;ڢH;̣H;G�H;R�H;ҩH;��H;��H;��H;N�H;4�H;�H;��H;��H;$�H;v�H;��H;��H;�H;z�H;��H;z�H;/�H;��H;��H;��H;��H;Z�H;��H;l�H;��H;�H;Q�H;��H;��H;��H;��H;��H;��H;��H;S�H;�H;��H;g�H;��H;Y�H;��H;��H;��H;��H;6�H;w�H;��H;u�H;�H;��H;��H;w�H;%�H;��H;��H;�H;4�H;O�H;��H;��H;��H;ʩH;U�H;B�H;٣H;ڢH;      |�H;°H;x�H;��H;S�H;F�H;��H;;�H;��H;��H;�H;��H;��H;��H;��H;V�H;��H;"�H;=�H;)�H;��H;q�H;��H;��H;��H;��H;=�H;��H;p�H;��H;	�H;Z�H;��H;��H;��H;��H;��H;��H;��H;��H;��H;Z�H;	�H;��H;n�H;��H;>�H;��H;��H;��H;��H;p�H;��H;�H;<�H;#�H;��H;V�H;��H;��H;��H;��H;�H;��H;��H;@�H;��H;C�H;[�H;��H;��H;ͰH;      �H;=�H;ӺH;��H;�H;��H;��H;��H;��H;R�H;��H;<�H;��H;�H;t�H;��H;��H;��H;c�H;��H;q�H;��H;��H;��H;��H;2�H;��H;P�H;��H;�H;T�H;��H;��H;��H;��H;��H;��H;��H;��H;��H;��H;��H;Q�H;��H;��H;L�H;��H;3�H;��H;��H;��H;��H;k�H;��H;`�H;��H;��H;��H;t�H;�H;��H;>�H;��H;S�H;��H;��H;��H;��H;�H;��H;ҺH;A�H;      N�H;o�H;�H;��H;��H;H�H; �H;��H;��H;��H;�H;L�H;��H;��H;��H;��H;f�H;(�H;��H;�H;P�H;`�H;Z�H;,�H;��H;��H;"�H;��H;��H;$�H;a�H;��H;��H;��H;��H;��H;��H;��H;��H;��H;��H;��H;_�H;�H;��H;��H;#�H;��H;��H;.�H;a�H;]�H;K�H;�H;��H;)�H;i�H;��H;��H;��H;��H;L�H;�H;��H;��H;��H;�H;I�H;��H;��H;�H;}�H;      +�H;4�H;��H;x�H;u�H;��H;|�H;*�H;�H;�H;5�H;?�H;D�H;[�H;[�H;?�H;��H;��H;��H;d�H;��H;��H;��H;D�H;*�H;��H;�H;��H;��H;=�H;X�H;��H;��H;��H;��H;��H;��H;��H;��H;��H;��H;��H;X�H;8�H;��H;��H;#�H;��H;*�H;F�H;��H;��H;��H;]�H;��H;��H;��H;B�H;[�H;[�H;F�H;>�H;6�H;�H;�H;-�H;��H;��H;v�H;x�H;��H;=�H;      O�H;r�H;�H;��H;��H;N�H;��H;��H;��H;��H;�H;L�H;��H;��H;��H;��H;e�H;(�H;��H;�H;R�H;a�H;Z�H;,�H;��H;��H;"�H;��H;��H;#�H;a�H;��H;��H;��H;��H;��H;��H;��H;��H;��H;��H;��H;_�H;�H;��H;��H;"�H;��H;��H;,�H;a�H;[�H;K�H;�H;��H;)�H;h�H;��H;��H;��H;��H;L�H;�H;��H;��H;��H;�H;I�H;��H;��H;�H;{�H;      ߹H;@�H;̺H;��H;�H;��H;��H;��H;��H;S�H;��H;<�H;��H;�H;u�H;��H;��H;��H;c�H;��H;r�H;��H;��H;��H;��H;2�H;��H;Q�H;��H;�H;S�H;��H;��H;��H;��H;��H;��H;��H;��H;��H;��H;��H;Q�H;��H;��H;J�H;��H;4�H;��H;��H;��H;��H;j�H;��H;`�H;��H;��H;��H;r�H;�H;��H;?�H;��H;S�H;��H;��H;��H;��H;!�H;��H;ѺH;A�H;      ~�H;��H;w�H;��H;V�H;J�H;��H;>�H;��H;��H;�H;��H;��H;��H;��H;V�H;��H;%�H;=�H;&�H;��H;t�H;��H;��H;��H;��H;=�H;��H;r�H;��H;	�H;Z�H;��H;��H;��H;��H;��H;��H;��H;��H;��H;Z�H;�H;��H;l�H;��H;=�H;��H;��H;��H;��H;q�H;��H;!�H;=�H;"�H;��H;X�H;��H;��H;��H;��H; �H;��H;��H;A�H;��H;G�H;]�H;��H;��H;ðH;      ��H;�H;УH;D�H;N�H;թH;��H;��H;��H;O�H;3�H;�H;��H;��H;'�H;w�H;��H;��H;�H;z�H;��H;z�H;/�H;��H;��H;��H;��H;]�H;��H;l�H;��H;�H;P�H;��H;��H;��H;��H;��H;��H;��H;P�H;�H;��H;g�H;��H;W�H;��H;��H;��H;��H;7�H;y�H;��H;w�H;�H;��H;��H;w�H;%�H;��H;��H;�H;3�H;N�H;��H; �H;��H;ѩH;S�H;L�H;ڣH;ڢH;      ��H;�H;8�H;G�H;�H;S�H;8�H;|�H;&�H;��H;��H;�H;ڸH;��H;k�H;��H;��H;i�H;��H;��H;��H;��H;��H;��H;B�H;��H;��H;��H;P�H;��H;d�H;��H;�H;X�H;��H;��H;��H;��H;��H;Z�H;�H;��H;b�H;��H;K�H;��H;��H;��H;@�H;��H;��H;��H;��H;��H;��H;f�H;��H;��H;i�H;��H;ڸH;�H;��H;��H;+�H;|�H;;�H;I�H;�H;F�H;A�H;	�H;      �sH;,tH;�uH;]xH;�{H;[�H;��H;=�H;v�H;�H;��H;<�H;��H;��H;�H;��H;��H;��H;&�H; �H;e�H;q�H;�H;V�H;b�H;�H;[�H;��H;��H;N�H;��H;i�H;��H;�H;Z�H;b�H;[�H;c�H;W�H;�H;��H;i�H;��H;K�H;��H;��H;]�H;�H;\�H;O�H;�H;q�H;`�H; �H;%�H;��H;��H;��H;�H;��H;��H;<�H;��H;��H;t�H;B�H;��H;X�H;�{H;hxH;�uH;-tH;      mOH;)PH;fRH;�UH;�ZH;�`H;�gH;GoH;�wH;�H;ǈH;��H;6�H;��H;]�H;��H;��H;�H;��H;��H;�H;�H;{�H;o�H;��H;�H;��H;g�H;��H;��H;I�H;��H;d�H;��H;��H;�H;4�H;�H;��H;��H;g�H;��H;H�H;�H;��H;a�H;��H;�H;��H;h�H;��H;�H;�H;��H;��H;�H;��H;��H;[�H;��H;5�H;��H;ɈH;�H;�wH;GoH;�gH;�`H;�ZH;�UH;qRH;#PH;      EH;E H;@#H; (H;p.H;�6H;�?H; JH;5UH;�`H;`lH;xH;a�H;c�H;ژH;��H;j�H;��H;�H;��H;��H;��H;��H;��H;��H;��H;��H;��H;5�H;��H;��H;O�H;��H;s�H;��H;��H;��H;��H;��H;s�H;��H;L�H;��H;��H;.�H;��H;��H;��H;��H;��H;��H;��H;��H;��H;�H;��H;h�H;��H;טH;`�H;a�H;xH;alH;�`H;4UH;%JH;�?H;�6H;.H;�'H;@#H;E H;      !�G;��G;��G;��G;��G;��G;3H;�H;�(H;�7H;|GH;	WH;%fH;�tH;A�H;�H;��H;x�H;��H;x�H;��H;��H;/�H;�H;�H;y�H;Y�H;��H;��H;d�H;��H;��H;U�H;��H;O�H;��H;��H;��H;O�H;��H;W�H;��H;��H;d�H;��H;��H;Y�H;��H;�H;�H;3�H;��H;��H;x�H;��H;s�H;��H;�H;?�H;�tH;$fH;	WH;{GH;�7H;�(H;�H;1H;��G;��G;��G;��G;��G;      SvG;"yG;	�G;��G;ÝG;��G;��G;��G;��G;mH;"H;�,H;�@H;�SH;�eH;_vH;��H;��H;�H;�H;s�H;ؼH; �H;H�H;j�H;��H;`�H;]�H;��H;��H;^�H;��H;��H;A�H;��H; �H;#�H; �H;��H;A�H;��H;��H;`�H;��H;��H;[�H;`�H;��H;h�H;@�H;&�H;ּH;o�H;�H;�H;|�H;��H;_vH;�eH;�SH;�@H;�,H;H;kH;~�G;��G;��G;��G;˝G;��G;
�G;
yG;      C�F;�F;��F;��F;p�F;lG;JGG;�pG;�G;2�G;��G;l�G;�H;*H;�AH;RWH;2kH;}H;�H;D�H;��H;,�H;L�H;(�H;��H;-�H;��H;��H;��H;�H;�H;��H;��H;��H;9�H;��H;��H;��H;7�H;��H;��H;��H;�H;�H;��H;�H;��H;3�H;��H;"�H;N�H;)�H;��H;D�H;�H;}H;2kH;OWH;�AH;*H;�H;i�G;��G;4�G;�G;�pG;IGG;[G;x�F;��F;��F;	�F;      �mD;�~D;P�D;��D;d\E;��E;u0F;ȔF;��F;�8G;�vG;��G;>�G;O�G;5H;w0H;9JH;jaH;�uH;��H;��H;;�H;��H;��H;��H;��H;g�H;�H;��H;��H;^�H;A�H;��H;��H;��H;��H;)�H;��H;��H;��H;��H;>�H;a�H;��H;��H;�H;g�H;��H;��H;��H;��H;8�H;��H;��H;�uH;baH;7JH;s0H;4H;M�G;@�G;��G;�vG;�8G;��F;ȔF;p0F;��E;k\E;��D;R�D;�~D;      &`?;��?;��?;�@;��A;|�B;C;��D;FiE;�F;(�F;�G;NnG;�G;��G;L H;m!H;!?H;lYH;^pH;J�H;z�H;�H;H�H;��H;!�H;@�H;�H;��H;p�H;U�H;��H;��H;��H;��H;9�H;N�H;:�H;��H;��H;��H;��H;W�H;s�H;��H;�H;A�H;(�H;��H;E�H;�H;w�H;F�H;^pH;jYH;?H;l!H;K H;��G;�G;MnG;�G;$�F;�F;>iE;��D;��C;r�B;��A;��@;��?;��?;      1�4;��4;�5;�l7;y_9;R�;;��=;�?;]�A;˚C;m�D;~�E;̨F;`)G;��G;�G;��G;HH;�6H;�SH;mH;u�H;��H;�H;��H;I�H; �H;2�H;��H;}�H;�H;��H;2�H;��H;��H;a�H;��H;_�H;��H;��H;0�H;��H;�H;��H;��H;2�H;#�H;P�H;��H;�H;��H;r�H;mH;�SH;�6H;>H;��G;�G;��G;[)G;ʨF;|�E;m�D;ʚC;Y�A;�?;��=;P�;;y_9;�l7;�5;��4;      e; ;d";^%;��(;)j-;:2;Ƅ6;��:;�0>;�A;HYC;1�D;
F;�F;�XG;��G;M�G;�H;W1H;�PH;�kH;t�H;}�H;8�H;(�H;ԼH;��H;��H;�H;n�H;��H;u�H;p�H;��H;]�H;��H;^�H;��H;n�H;v�H;��H;r�H;�H;��H;��H;׼H;,�H;4�H;}�H;r�H;�kH;�PH;U1H;�H;F�G;��G;�XG;�F;F;1�D;FYC;�A;�0>;��:;Ʉ6;42;j-;�(;R%;f"; ;      ��:�B�:��:zx;��
;�;7�;�}$;:|,;c�3;�_9;>>;zA;��C;�E;�F;"5G;x�G;Z�G;AH;�/H;�PH;mH;J�H;��H;��H;i�H;��H;��H;�H;]�H;��H;��H;��H;j�H;H�H;��H;I�H;j�H;��H;��H;��H;^�H;�H;��H;��H;l�H;��H;��H;I�H;mH;�PH;�/H;?H;W�G;t�G;"5G;�F;�E;��C;zA;=>;�_9;e�3;8|,;�}$;9�;�;��
;tx;���:�B�:      �w[:�Bd:�}:��:E�:��:�:�;�;Z ;�+;��3;ܡ:;�?;��B;�E;IZF;�G;�G;s�G;FH;Z1H;�SH;apH;އH;E�H;�H;y�H;��H;��H;��H;��H;s�H;#�H;��H;�H;\�H;�H;��H;�H;p�H;��H;��H;��H;��H;y�H;�H;H�H;هH;dpH;�SH;S1H;?H;p�G;�G;�G;IZF;�E;��B;�?;ܡ:;��3;�+;Z ;�;�;�:ѳ�:K�:��:$�}:jBd:      4�S���D�������� !(7��9��R:3��:O��:��:�>;�";�P.;(m7;��=;[B;ްD;{9F; G;�G;[�G;�H;�6H;iYH;�uH;�H;�H;��H; �H;��H;�H;��H;�H;9�H;a�H;��H;��H;��H;^�H;6�H;�H;��H;"�H;��H;��H;��H;�H;�H;�uH;mYH;�6H;�H;T�G;�G; G;w9F;ްD;VB;��=;(m7;�P.;�";�>;��:M��:9��:��R:��9 (7І��Ԗ���D�      �D^��/X�rF�(}*����P��|�D�@ˬ��i:��:R��::�;��;H�);��4;�<;�A;&�D;y9F;�G;r�G;G�G;AH;?H;aaH;}H;x�H;v�H;��H;�H;��H;b�H;�H;�H;��H;&�H;��H;&�H;��H;�H;|�H;`�H;��H;�H;��H;v�H;|�H;}H;ZaH;?H;>H;C�G;m�G;�G;t9F;#�D;�A;�<;��4;F�);��;9�;X��:��:�i:�ˬ���D��P����0}*�rF��/X�      ��ﻩ��c�ܻB�ƻb󩻴���FL� ������@��`�-:�:���:�;�>&;��3;W9<;�A;ްD;FZF;$5G;��G;��G;l!H;5JH;-kH;��H;��H;j�H;��H;��H;��H;��H;��H;��H;c�H;��H;b�H;��H;��H;��H;��H;��H;��H;g�H;��H;��H;,kH;,JH;j!H;��G;��G;5G;FZF;ݰD;�A;U9<;��3;�>&;�;���:�:X�-:`������ ���FL����i�H�ƻh�ܻ���      i�V��5S��6H���6�B� �P,��?ػ4G���D^������D����9�4�:�:0�;�%;��3;�<;XB;�E;�F;�XG;�G;H H;n0H;NWH;YvH;�H;�H;��H;��H;��H;p�H;T�H;��H;��H;7�H;��H;��H;K�H;m�H;��H;��H;��H;|�H;�H;XvH;HWH;g0H;E H;�G;�XG;��F;�E;VB;�<;��3;�%;-�;
�:�4�:���9��D�����D^�4G���?ػQ,�E� ���6��6H��5S�      ��
.��KȤ���������8�f�s�=����9�ܻ�*��Lo5�V��� �(7��}:�n�:0�;�>&;��4;��=;��B;�E;�F;��G;��G;/H;�AH;�eH;?�H;ؘH;[�H;ݷH;f�H;!�H;��H;j�H;��H;N�H;��H;h�H;��H;�H;c�H;۷H;\�H;ؘH;<�H;�eH;}AH;*H;��G;��G;�F;�E;��B;��=;��4;�>&;*�;�n�:|�}: ~(7Z���Mo5��*��8�ܻ���s�=�9�f���������KȤ�
.��      �c��8���������Ҽ����������r�FE:�C,�Fߵ�y/X�|�º@Ƭ���}:�:�;H�);'m7;�?;��C;	F;])G;�G;L�G;*H;�SH;�tH;c�H;�H;�H;��H;��H;��H;�H;��H;J�H;��H;�H;��H;��H;��H;�H;��H;c�H;�tH;�SH;�)H;E�G;�G;\)G;F;��C;�?;$m7;F�);�;�:x�}:@Ƭ���ºz/X�Gߵ�D,�FE:���r�����������Ҽ�켴����8�      #'K���G��>��0�\y��c����S��� ��U�V�&���ƻ�od�t�º �(7�4�:���:��;�P.;ء:;zA;.�D;ΨF;QnG;?�G;�H;�@H;$fH;d�H;0�H;��H;ָH;��H;��H;��H;{�H;6�H;{�H;��H;��H;��H;ѸH;��H;2�H;c�H;!fH;�@H;�H;8�G;MnG;ʨF;-�D;zA;ڡ:;�P.;��;���:�4�: �(7z�º�od��ƻ'��U�V� ��S�����伔c�^y��0��>���G�      ���0Z��ΐ����}��c���D�1/%��8���Ҽ/c��0�f�����ƻz/X�N������9�:9�;�";��3;E>;DYC;|�E;�G;�G;f�G;�,H;WH;xH;��H;4�H;�H;�H;��H;0�H;B�H;.�H;D�H;-�H;��H;�H;�H;1�H;��H;xH;WH;�,H;`�G;�G;�G;|�E;BYC;;>;��3;�";:�;�:���9T���{/X��ƻ���1�f�/c����Ҽ�8�2/%���D��c���}�ϐ��0Z��      �Pν�ʽN8���������ΐ��`�f���;�1����AȤ�1�f�'��Iߵ�No5���D�@�-:H��:�>;�+;�_9;�A;j�D;#�F;�vG;��G;H;xGH;`lH;H;��H;��H;,�H;��H;��H;�H;$�H;�H;��H;��H;)�H;�H;��H;ňH;`lH;uGH;H;��G;�vG;!�F;j�D;�A;�_9;�+;�>;@��:@�-:��D�Ro5�Jߵ�(��2�f�AȤ����1����;�`�f�ΐ���������N8���ʽ      ���g9�Z[��s�z�ؽ���t����}���G�����/c��U�V�D,��*����������:��:W ;i�3;�0>;ʚC;�F;�8G;-�G;kH;�7H;�`H;
�H;�H;��H;K�H;��H;G�H;��H;�H;��H;E�H;��H;H�H;��H;�H;�H;�`H;�7H;iH;)�G;�8G;�F;ʚC;�0>;^�3;W ;��:��:�������*��D,�V�V�/c��������G���}�t�����{�ؽ�s�Z[�g9�      ��=�ր:���0��Q"�~������Pν�榽?����G�1����Ҽ ��GE:�9�ܻ�D^�����`i:I��:�;<|,;��:;O�A;BiE;��F;�G;�G;�(H;5UH;|wH;q�H;#�H;��H;�H;��H;��H;�H;��H;��H;�H;��H;!�H;p�H;�wH;5UH;�(H;��G;�G;��F;CiE;O�A;��:;6|,;�;A��:`i:�����D^�:�ܻGE:� ����Ҽ1����G�?���榽�Pν����~��Q"���0�ր:�      0Dx�4�s���f�sS�ր:����Z[��7ս�榽��}���;��8�T�����r����8G����@ͬ�-��:�;�}$;Ƅ6;�?;��D;ʔF;�pG;��G;�H;"JH;@oH;=�H;y�H;��H;7�H;��H;��H;%�H;��H;��H;6�H;��H;r�H;:�H;GoH;"JH;�H;��G;�pG;ȔF;�D;�?;6;�}$;�;%��:�̬���9G�������r�T����8���;���}��榽�7սZ[����ր:�sS���f�4�s�      �*���0��ޥ��;����k��H��#%�Z[��Pνt��`�f�2/%���伅���s�=��?ػ�FL���D�p�R:��:7�;82;��=;��C;h0F;IGG;��G;#H;�?H;�gH;��H;-�H;��H;��H;}�H;��H;r�H;��H;��H;��H;��H;*�H;��H;�gH;�?H;&H;��G;MGG;h0F;��C;��=;22;0�;��:d�R:��D��FL��?ػs�=��������2/%�`�f�t���PνZ[��#%��H��k�;���ޥ���0��      '�þ��� ����R��|쏾5�s��H�����������ΐ����D��c�����:�f�R,�����P��`�9ӳ�:�;"j-;M�;;u�B;��E;\G;��G;��G;�6H;�`H;[�H;O�H;թH;N�H;��H;O�H;��H;O�H;��H;M�H;ҩH;L�H;W�H;�`H;�6H;��G;��G;bG;��E;v�B;M�;;j-;�;׳�:P�9�P�����R,�:�f������c���D�ΐ�������������H�5�s�|쏾�R�� ������      @��/�待Yؾ(�þĪ�|쏾�k�ր:�~�z�ؽ�����c�\y���Ҽ����B� �g�+�� #(7K�:��
;��(;~_9;��A;j\E;l�F;��G;��G;�.H;�ZH;�{H;�H;I�H;P�H;�H;��H;u�H;��H;�H;M�H;H�H;�H;�{H;�ZH;�.H;��G;ÝG;v�F;g\E;��A;~_9;��(;��
;O�: "(7(��h�B� �������Ҽ]y��c�����z�ؽ~�ր:��k�|쏾Ī�(�þ�Yؾ/��      #��N������>I�(�þ�R��;���tS��Q"��s������}��0��켇�����6�D�ƻ6}*�������:�x;X%;�l7;ڳ@;��D;��F;��G;��G;�'H;�UH;`xH;N�H;F�H;��H;��H;��H;{�H;��H;��H;��H;F�H;N�H;]xH;�UH;�'H;��G;��G;��F;��D;ܳ@;�l7;X%;}x;��: ���3}*�D�ƻ��6��������0���}�����s��Q"�tS�;����R��(�þ>Iᾣ���O��      ���R��8�
������Yؾ���ޥ����f���0�Z[�N8��ϐ���>�����IȤ��6H�_�ܻrF�����}:���:c";-�5;��?;Y�D;��F;	�G;��G;/#H;`RH;�uH;H�H;£H;v�H;ĺH;�H;��H;�H;ĺH;v�H;��H;F�H;�uH;iRH;0#H;��G;�G;��F;T�D;��?;+�5;b";��:0�}:���rF�`�ܻ�6H�IȤ������>�ϐ��N8��Z[���0���f�ޥ������Yؾ����8�
�R��      �� ����R��N��/������0��4�s�ր:�g9��ʽ0Z����G��8�
.���5S�����/X�h�D�zBd:�B�: ;��4;ʈ?;�~D;�F;yG;��G;M H;*PH;tH;�H;΢H;ǰH;.�H;q�H;6�H;n�H;.�H;ǰH;̢H;�H;tH;3PH;P H;��G;yG;�F;�~D;Ȉ?;��4; ;�B�:�Bd:p�D��/X���껬5S�
.���8���G�1Z���ʽg9�ր:�4�s��0�����/��N��R�����      GF�Wh����VVھ7�������~���S��#��o��8S��p₽1�6�n���hy��UFB��Eֻ�A?�ľ	�oY�:���:g�";h46;\@;b�D;��F;�nG;��G;�H;@H;�fH;B�H;/�H;��H;гH;͹H;��H;ʹH;ϳH;��H;,�H;?�H;�fH;@H;�H;��G;�nG;��F;_�D;[@;b46;g�";���:wY�:ľ	��A?��EֻUFB�gy��n���1�6�p₽8S���o���#��S��~������7��VVھ��Wh��      Vh���b���쾧*־�v��(���*��'�O�U� �s��r���؀�F�3���>ݜ�;�>�R�ѻܡ9�����#o�:>% ;tM#;C�6;LA@;��D;��F;qG;L�G;H;�@H;ggH;��H;��H;ީH;�H;��H;޻H;��H;�H;ީH;��H;��H;cgH;�@H;H;L�G;qG;��F;��D;LA@;?�6;pM#;=% ;)o�:����ܡ9�Q�ѻ;�>�>ݜ���F�3��؀��r��s�U� �'�O�*��(����v���*־���b��      ���쾳�޾/5ʾL;���:��(�v��E�_'����q����u���+��W��A����4���Ļ9)�`j��{W�:b�;	%;�k7;$�@;��D;��F;�wG;T�G;2H;=CH;(iH;�H;��H;��H;��H;��H;r�H;��H;��H;��H;��H;�H;$iH;DCH;4H;U�G;�wG;��F;��D;"�@;�k7;%;d�;�W�:pj��9)���Ļ��4��A���W缃�+���u�q�����_'��E�(�v��:��L;��/5ʾ��޾��      VVھ�*־/5ʾr��������M���9b��5�����ս����Xc���ʖռ�I��U�$�kT���Z�@\���:��;k�';�8;RA;�9E;��F;ÂG;��G;@H;GH;lH;C�H;;�H;�H;��H;��H;Q�H;��H;ĵH;�H;8�H;B�H;lH;GH;CH;��G;łG;��F;�9E;RA;�8;k�';��;�:@\���Z�jT��T�$��I��ʖռ���Xc������ս���5��9b��M������r���/5ʾ�*־      7���v��M;������RP��E�r�z�H�U� ���5@��ѓ����K�`��վ���s�r���񕻛ܺ5u9&�:"�;-�+;~�:;�"B;o�E;��F;ԐG;��G;/H;5LH;�oH;;�H;t�H;��H;4�H;ؼH;��H;ԼH;7�H;��H;r�H;9�H;�oH;<LH;.H;��G;ՐG;��F;q�E;�"B;|�:;/�+;"�;&�:�4u9�ܺ��r����s��վ�`���K�ѓ��5@����U� �z�H�E�r�RP������M;���v��      ����(����:���M��E�r�&�O�#,�X�
��gٽpĥ���u�x1�h���)Ϥ���P�[�.o�np��@:c��:�P;>�/;9�<;C;�E;k!G;5�G;�G;�%H;�RH;�tH;��H;F�H;֯H;�H;[�H;�H;V�H;�H;ԯH;D�H;��H;�tH;�RH;�%H;�G;7�G;u!G;�E;C;7�<;>�/;�P;k��:D:hp���.o�[򻩎P�)Ϥ�g���w1���u�pĥ��gٽX�
�#,�&�O�E�r��M���:��(���      �~��*��(�v��9b�z�H�#,�MZ����7S��x^����N������μ�I���%+����ڝ.�p����j~:I��:-m;��3;�>;;�C;=PF;}FG;Q�G;��G;v/H;�YH;tzH;E�H;��H;\�H;�H;)�H;��H;&�H;�H;]�H;��H;D�H;rzH;ZH;y/H;��G;S�G;�FG;>PF;;�C;�>;��3;,m;W��:�j~:p���֝.�����%+��I����μ�����N�x^��7S�����MZ�#,�z�H��9b�(�v�*��      �S�'�O��E��5�U� �X�
���罤9��'l���Xc���(��������[�����ݎ�@ܺ�;9%��:/�	;Ed';e 8;<�@;�D;�F;jG;��G;NH;p:H;AbH;��H;�H;1�H;B�H;}�H;6�H;��H;5�H;��H;D�H;/�H;�H;��H;HbH;q:H;OH;��G;jG;�F;{�D;>�@;h 8;Ed';6�	;'��:�;9<ܺ�ݎ������[��������(��Xc�'l���9�����X�
�U� ��5��E�'�O�      �#�U� �_'������gٽ7S��'l��N�j�C�3��i��վ�y���(���Ļ^A?���B��@:�[�:
Q;�.;��;;{tB;�E;�F;%�G;��G;�H;TFH;%kH;��H;�H;�H;g�H;
�H;s�H;��H;o�H;�H;h�H;�H;�H;��H;*kH;VFH;�H;��G;(�G;��F;�E;~tB;��;;�.;Q;�[�:�@:��B�\A?���Ļ(�y����վ��i�C�3�M�j�'l��7S���gٽ����_'�U� �      �o��s��罫�ս4@��pĥ�x^���Xc�D�3���	�Ɍ˼�]��QFB��Z򻬜��hӺ ��8��:ܛ;�M#;u=5;?;K�C;|@F;:G;�G; �G;0'H;�RH;ztH;��H;{�H;+�H;��H;��H;��H;?�H;��H;��H;��H;(�H;x�H;��H;�tH;�RH;2'H; �G;�G;:G;{@F;O�C;?;w=5;�M#;ߛ;��:���8dӺ�����Z�QFB��]��Ɍ˼��	�C�3��Xc�x^��pĥ�5@����ս���s�      8S���r��q�����Г����u���N���(��i�ʌ˼�A����P�fs��8|�8����\:5�:r�;xn-;�:;�A;z,E;j�F;)oG;��G;�H;�7H;:_H;~H;�H;�H;t�H;�H;x�H;;�H;��H;;�H;x�H;�H;s�H;��H;�H;~H;@_H;�7H;�H;��G;/oG;k�F;~,E;��A;�:;�n-;u�;5�:�\:0���4|��fs���P��A��Ɍ˼�i���(���N���u�ѓ�����r���r��      o₽�؀���u��Xc���K�x1�������վ��]����P����?T����9���o��3�9z&�:a�	;\%;F�5;��>;��C;�F;�!G;��G;��G;DH;`HH;�kH;��H;J�H;��H;��H;t�H;J�H;��H;��H;��H;I�H;w�H;��H;��H;M�H;��H;�kH;bHH;EH;��G;��G;�!G;�F;��C;��>;T�5;`%;`�	;�&�:�3�9��o���9�>T�������P��]���վ�ߤ���v1���K��Xc���u��؀�      1�6�F�3���+���`�h�����μ���y���QFB�es�@T��&�D��{���:u9�q�:}��:�Y;�t0;��;;�B;�9E;�F;hG;ٿG;�G;z0H;�XH;'xH; �H;v�H;�H;��H;��H;�H;.�H;2�H;.�H;�H;��H;��H;��H;y�H;*�H;-xH;�XH;|0H;�G;޿G;hG;�F;�9E;�B;��;;�t0;}Y;���:�q�:�:u9�{��$�D�=T��es�QFB�x��������μh���a�����+�F�3�      l�����W�˖ռ�վ�*Ϥ��I����[�(��Z����9��{���;9SX�:`X�:=Q;B,;��8;�A@;BD;�@F;�,G;��G;��G;gH;�DH;hH;-�H;T�H;e�H;`�H;"�H;�H;��H;��H;c�H;��H;��H;�H; �H;[�H;j�H;\�H;7�H; hH;�DH;bH;��G;��G;�,G;�@F;BD;�A@;��8;@,;BQ;^X�:]X�:�;9�{����9���Z�(���[��I��)Ϥ��վ�˖ռ�W���      fy��?ݜ��A���I����s���P��%+������Ļ����2|��o��:u9YX�:�+�:Z;�);ׄ6;x�>;�PC;d�E;��F;�xG;+�G;zH;e1H;XH;wH;��H;�H;�H;~�H;�H;?�H;��H;��H;��H;��H;��H;B�H;�H;z�H;�H;�H;��H;wH;XH;a1H;}H;/�G;�xG;��F;h�E;�PC;}�>;ф6;�);Z;�+�:aX�:�:u9��o�.|�������Ļ����%+���P���s��I���A��>ݜ�      OFB�:�>���4�S�$�q��
[�����ݎ�bA?�cӺ(����3�9�q�:`X�:Z;��';�=5;��=;�B;GE;K�F;�UG; �G;��G;UH;�HH;jH;��H;u�H;H�H;1�H;J�H;��H;A�H;�H;�H;��H;�H;�H;@�H;��H;F�H;5�H;N�H;|�H;��H;jH;�HH;WH;��G;$�G;�UG;O�F;!GE;�B;|�=;�=5;��';\;`X�:�q�:�3�9���^ӺZA?��ݎ����[�t��T�$���4�7�>�      �EֻN�ѻ��ĻnT���񕻶.o�ҝ.�5ܺ|�B� ��8�\:|&�:���:AQ;�);�=5;�:=;,#B;��D;�uF;�6G;ÚG;]�G;tH;�:H;^H;�zH;��H;a�H;ŲH;�H;��H;\�H;�H;m�H;2�H;��H;-�H;j�H;�H;X�H;��H;�H;ȲH;e�H;��H;�zH;^H;�:H;vH;\�G;ǚG;�6G;�uF;��D;(#B;�:=;�=5;�);BQ;���:�&�:�\:`��8x�B�1ܺ֝.��.o���pT����ĻI�ѻ      oA?�ա9�9)��Z�ܺdp��(����;9�@:��:=�:\�	;yY;@,;Є6;y�=;!#B;��D;`XF;�!G;|�G;�G;�H;�.H;ySH;cqH;߉H;��H;c�H;��H;o�H;��H;��H;��H;��H;�H;��H;�H;�H;��H;��H;��H;r�H;ĹH;h�H;��H;މH;^qH;SH;�.H;�H; �G;��G;�!G;eXF;��D;%#B;v�=;ӄ6;>,;zY;]�	;G�:��:�@: <9X���`p��zܺ�Z�9)�ҡ9�      d�	� ���hj���[��5u9t:�j~:3��:�[�:�;|�;[%;�t0;��8;}�>;�B;��D;hXF;7G;_�G;��G;��G;�%H;KH;�iH;�H;��H;8�H;v�H;
�H;]�H;��H;��H;3�H;��H;��H;S�H;��H;}�H;2�H;��H;��H;`�H;�H;v�H;8�H;��H;�H;�iH;
KH;�%H;��G;��G;e�G;;G;eXF;��D;�B;~�>;��8;�t0;_%;}�;��;�[�:7��:�j~:\: 5u9 ]��pj�� ���      eY�:!o�:�W�:1�:&�:o��:k��:0�	;Q;�M#;�n-;Q�5;��;;�A@;�PC;"GE;�uF;�!G;b�G;��G;�G;H H;EH;�cH;8}H;u�H;��H;��H;��H;��H;��H;+�H;T�H;S�H;N�H;|�H;��H;u�H;K�H;S�H;R�H;(�H;��H;��H;��H;��H;��H;t�H;<}H;�cH;EH;J H;�G;��G;f�G;�!G;�uF;!GE;�PC;�A@;��;;R�5;�n-;�M#;Q;9�	;g��:{��:&�:�:uW�:�n�:      ���:/% ;H�;��;�;�P;-m;Cd';�.;x=5;�:;��>;�B;BD;f�E;P�F;�6G;��G;��G;�G;tH;�AH;
`H;LyH;~�H;"�H;Q�H;�H;K�H;��H;��H;2�H;��H;B�H;��H;��H;F�H;��H;��H;A�H;��H;-�H;��H;��H;K�H;�H;M�H;�H;��H;LyH;`H;�AH;zH;�G;��G;��G;�6G;P�F;i�E;BD;�B;��>;�:;w=5;�.;@d';3m;�P;$�;��;R�;+% ;      _�";xM#;%;x�';-�+;>�/;��3;d 8;��;;?;�A;��C;�9E;�@F;��F;�UG;ĚG;$�G;��G;I H;�AH;�^H;GwH;�H;��H;�H;��H;.�H;��H;%�H;�H;��H;��H;��H;m�H;L�H;|�H;D�H;j�H;��H;��H;��H;�H;(�H;��H;-�H;��H;ݫH;��H;�H;BwH;�^H;�AH;L H;��G;#�G;ʚG;�UG;��F;�@F;�9E;��C;�A;?;��;;m 8;��3;8�/;A�+;m�';	%;nM#;      46;B�6;�k7;*�8;v�:;@�<;+�>;H�@;�tB;U�C;�,E;�F;�F;�,G;�xG;(�G;b�G;�H;�%H;EH;`H;DwH;2�H;5�H;G�H;�H;��H;n�H;��H;��H;(�H;@�H;��H;]�H;��H;p�H;��H;k�H;��H;_�H;��H;<�H;*�H;��H;��H;n�H;��H;�H;K�H;3�H;-�H;HwH;`H;EH;�%H;�H;b�G;(�G;�xG;�,G;�F;�F;�,E;P�C;�tB;J�@;+�>;>�<;��:;*�8;�k7;&�6;      ^@;UA@;�@;RA;�"B;C;?�C;�D;�E;�@F;o�F;�!G;hG;��G;/�G;��G;vH;�.H;KH;�cH;IyH;�H;3�H;éH;�H;|�H;w�H;��H;�H;N�H;��H;J�H;9�H;��H;��H;_�H;��H;Z�H;��H;��H;9�H;I�H;��H;M�H;�H;��H;r�H;�H;	�H;��H;.�H;�H;JyH;�cH;KH;�.H;xH;��G;-�G;��G;hG;�!G;t�F;�@F;�E;��D;?�C;�
C;�"B;RA;�@;NA@;      ��D;��D;��D;�9E;h�E;)�E;FPF;�F;��F;:G;7oG;��G;ݿG;��G;H;]H;�:H;�SH;�iH;B}H;��H;��H;J�H;�H;=�H;��H;.�H;m�H;��H;(�H;��H;	�H;��H;��H;��H;%�H;c�H; �H;��H;��H;��H;�H;��H;+�H;��H;m�H;'�H;��H;?�H;	�H;J�H;��H;��H;?}H;�iH;�SH;�:H;]H;H;��G;޿G;��G;9oG;:G;��F;�F;HPF;!�E;r�E;�9E;��D;��D;      ��F;��F;��F;��F;��F;x!G;�FG;#jG;)�G;��G;��G;��G;�G;oH;e1H;�HH;^H;eqH;�H;p�H; �H;ګH;�H;|�H;��H;�H;�H;[�H;��H;��H;��H;��H;��H;��H;x�H;��H;	�H;��H;w�H;��H;��H;}�H;��H;��H;��H;Z�H;�H;�H;��H;z�H;�H;۫H; �H;q�H;�H;aqH;^H;�HH;e1H;iH;�G;��G;��G;�G;)�G;&jG;�FG;m!G;��F;��F;��F;��F;      �nG;qG;�wG;ǂG;̐G;1�G;_�G;��G;��G;"�G;�H;BH;y0H;�DH;XH;jH;�zH;�H;��H;��H;U�H;��H;��H;x�H;,�H;�H;=�H;��H;\�H;{�H;I�H;��H;��H;��H;6�H;��H;��H;��H;2�H;��H;��H;��H;K�H;z�H;\�H;��H;6�H;�H;-�H;t�H;��H;��H;T�H;��H;��H;߉H;�zH;jH;XH;�DH;y0H;EH;�H;�G;��G;��G;Z�G;0�G;�G;��G;�wG;qG;      ��G;I�G;N�G;��G;��G;��G;��G;LH;�H;7'H;�7H;gHH;�XH;"hH;wH;��H;��H;��H;8�H;��H;�H;*�H;j�H;��H;j�H;X�H;��H;9�H;v�H;@�H;��H;��H;��H;a�H;��H;�H;�H;��H;��H;c�H;��H;��H;��H;@�H;w�H;9�H;��H;[�H;o�H;��H;m�H;+�H;�H;��H;8�H;��H;��H;��H;wH;"hH;�XH;hHH;�7H;7'H;�H;NH;��G;��G;��G;��G;P�G;?�G;      �H;H;1H;OH;H;�%H;}/H;m:H;MFH;�RH;A_H;�kH;-xH;3�H;��H;z�H;g�H;j�H;z�H;¼H;N�H;��H;��H;�H;��H;��H;W�H;v�H;!�H;��H;��H;��H;S�H;��H;C�H;v�H;��H;r�H;C�H;��H;W�H;��H;��H;��H;"�H;v�H;S�H;��H;��H;	�H;��H;��H;K�H;��H;x�H;h�H;g�H;{�H;��H;1�H;*xH;�kH;D_H;�RH;OFH;m:H;}/H;�%H;+H;MH;1H;	H;      @H;�@H;HCH;GH;>LH;�RH;ZH;@bH;)kH;�tH;~H;��H;(�H;]�H;�H;H�H;ʲH;��H;�H;��H;��H;!�H;��H;H�H;*�H;��H;w�H;>�H;��H;��H;��H;g�H;��H;M�H;��H;��H;��H;��H;��H;M�H;��H;c�H;��H;��H;��H;>�H;t�H;��H;+�H;G�H;��H;"�H;��H;��H;�H;��H;ʲH;I�H;�H;[�H;'�H;��H;~H;�tH;(kH;FbH;ZH;�RH;>LH;GH;ICH;�@H;      �fH;{gH;.iH;lH;�oH;�tH;|zH;��H;��H;��H;��H;T�H;~�H;q�H;�H;:�H;�H;v�H;b�H;��H;��H; �H;&�H;��H;��H;��H;K�H;��H;��H;��H;g�H;�H;]�H;��H;��H;�H;'�H;�H;��H;��H;`�H; �H;g�H;��H;��H;��H;H�H;��H;��H;��H;,�H;�H;��H;��H;a�H;u�H;�H;8�H;�H;o�H;��H;U�H;�H;��H;��H;��H;�zH;�tH; pH;lH;/iH;}gH;      A�H;��H;�H;;�H;:�H;�H;L�H;�H;$�H;~�H;�H;��H;
�H;i�H;��H;M�H;��H;��H;��H;2�H;6�H;��H;=�H;H�H;	�H;}�H;��H;��H;��H;h�H;��H;s�H;��H;��H;&�H;@�H;@�H;@�H;$�H;��H;��H;o�H;��H;g�H;��H;��H;��H;�H;�H;B�H;A�H;��H;2�H;.�H;��H;��H;��H;O�H;��H;g�H;	�H;��H;�H;�H;#�H;�H;U�H;�H;E�H;<�H;�H;��H;      2�H;��H;��H;;�H;|�H;D�H;��H;.�H;�H;1�H;{�H;��H;�H;+�H;�H;��H;a�H;��H;��H;X�H;��H;��H;��H;6�H;��H;��H;��H;��H;Y�H;��H;[�H;��H;�H;5�H;T�H;v�H;}�H;v�H;Q�H;6�H;�H;��H;Z�H;��H;W�H;��H;��H;��H;��H;6�H;��H;��H;��H;U�H;��H;��H;b�H;��H;�H;+�H;�H;��H;}�H;2�H;�H;/�H;��H;=�H;��H;5�H;��H;��H;      ��H;ةH;��H;٫H;��H;ͯH;g�H;F�H;n�H;��H;�H;��H;��H;(�H;I�H;H�H;"�H;��H;7�H;W�H;G�H;��H;Y�H;��H;��H;��H;��H;d�H;��H;P�H;��H;��H;2�H;p�H;�H;��H;��H;��H;~�H;q�H;5�H;��H;��H;L�H;��H;`�H;��H;��H;��H;��H;`�H;��H;A�H;Q�H;6�H;��H;'�H;H�H;I�H;'�H;��H;��H;�H;��H;p�H;L�H;j�H;˯H;��H;ګH;��H;�H;      ̳H;#�H;ôH;ƵH;E�H;��H;*�H;~�H;�H;��H;��H;V�H;!�H;��H;��H;�H;q�H;��H;��H;R�H;��H;k�H;��H;��H;��H;p�H;-�H;��H;C�H;��H;��H;'�H;S�H;��H;��H;��H;��H;��H;��H;��H;W�H;'�H;��H;��H;?�H;��H;-�H;q�H;��H;��H;��H;j�H;��H;I�H;~�H;��H;v�H;�H;��H;��H;!�H;X�H;��H;��H;�H;��H;-�H;��H;E�H;ǵH;ŴH;'�H;      ͹H;��H;��H;��H;׼H;O�H;8�H;:�H;v�H;��H;F�H;��H;5�H;��H;��H;!�H;4�H;�H;��H;y�H;��H;I�H;h�H;P�H; �H;��H;��H;�H;y�H;��H;�H;D�H;{�H;��H;��H;��H;��H;��H;��H;��H;~�H;D�H;�H;��H;v�H;��H;��H;��H;!�H;Q�H;o�H;G�H;��H;u�H;��H; �H;6�H;#�H;��H;��H;5�H;��H;I�H;��H;y�H;?�H;<�H;R�H;ؼH;��H;��H;�H;      ȻH;ۻH;��H;N�H;�H;�H;��H;��H;��H;H�H;��H;��H;B�H;s�H;��H;��H;��H;��H;Y�H;��H;O�H;��H;��H;��H;d�H;�H;��H;�H;��H;��H;$�H;D�H;~�H;��H;��H;��H;��H;��H;��H;��H;��H;C�H;$�H;��H;��H;�H;��H;�H;d�H;��H;��H;��H;J�H;��H;W�H;��H;��H;��H;��H;s�H;A�H;��H;��H;J�H;�H;��H;��H;�H;��H;M�H;��H;�H;      ιH;��H;��H;��H;׼H;U�H;7�H;:�H;v�H;��H;D�H;��H;6�H;��H;��H;!�H;3�H;�H;��H;y�H;��H;K�H;h�H;P�H;!�H;��H;��H;�H;z�H;��H;�H;F�H;}�H;��H;��H;��H;��H;��H;��H;��H;~�H;D�H;�H;��H;v�H;��H;��H;��H;!�H;Q�H;o�H;E�H;��H;u�H;��H;!�H;4�H;$�H;��H;��H;5�H;��H;I�H;��H;y�H;@�H;:�H;R�H;ۼH;��H;��H;�H;      ĳH;&�H;��H;��H;H�H;��H;,�H;��H;�H;��H;��H;V�H;"�H;��H;��H;�H;q�H;��H;��H;R�H;��H;n�H;��H;��H;��H;n�H;/�H;��H;E�H;��H;��H;'�H;T�H;��H;��H;��H;��H;��H;��H;��H;W�H;&�H;��H;��H;?�H;��H;-�H;q�H;��H;��H;��H;k�H;��H;I�H;~�H;��H;v�H;�H;��H;��H;!�H;Z�H;��H;��H;�H;��H;2�H;��H;I�H;��H;´H;)�H;      ��H;٩H;��H;ݫH;��H;ЯH;d�H;J�H;o�H;��H;�H;�H;��H;(�H;J�H;G�H;%�H;��H;9�H;X�H;H�H;��H;[�H;��H;��H;��H;��H;d�H;��H;Q�H;��H;��H;2�H;p�H;�H;��H;��H;��H;~�H;p�H;5�H;��H;��H;L�H;��H;`�H;��H;��H;��H;��H;`�H;��H;@�H;S�H;6�H;��H;%�H;I�H;J�H;'�H;��H;��H;�H;��H;p�H;N�H;k�H;ϯH;��H;ګH;��H;۩H;      2�H;��H;��H;9�H;y�H;F�H;��H;1�H;�H;1�H;{�H;��H;�H;+�H;�H;��H;b�H;��H;��H;[�H;��H;��H;��H;6�H;��H;��H;��H;��H;\�H;��H;[�H;��H;�H;5�H;S�H;x�H;}�H;v�H;S�H;5�H;�H;��H;Z�H;��H;S�H;��H;��H;��H;��H;3�H;��H;��H;��H;V�H;��H;��H;b�H;��H;�H;+�H;�H;��H;{�H;1�H;�H;4�H;��H;C�H;|�H;=�H;��H;��H;      3�H;��H;��H;:�H;6�H;��H;P�H;�H;#�H;~�H;�H;��H;�H;g�H;��H;O�H;��H;��H;��H;0�H;;�H;��H;@�H;H�H;�H;�H;��H;��H;��H;g�H;��H;p�H;��H;��H;'�H;?�H;@�H;?�H;#�H;��H;��H;o�H;��H;e�H;��H;��H;��H;��H;	�H;?�H;D�H;��H;/�H;,�H;��H;��H;��H;N�H;��H;g�H;
�H;��H;�H;�H;'�H;
�H;S�H;�H;7�H;:�H;�H;��H;      �fH;ygH;1iH;lH;�oH;�tH;|zH;��H;��H;��H;��H;U�H;~�H;o�H;	�H;;�H;�H;x�H;d�H;��H;��H;#�H;)�H;��H;��H;��H;G�H;��H;��H;��H;g�H;�H;^�H;��H;��H;�H;&�H;�H;��H;��H;`�H;�H;e�H;��H;��H;��H;E�H;��H;��H;��H;-�H; �H;��H;��H;b�H;t�H;�H;8�H;�H;q�H;��H;W�H;��H;��H;��H;��H;�zH;�tH;pH;lH;6iH;{gH;      @H;�@H;BCH;GH;5LH;�RH;ZH;HbH;*kH;�tH;~H;��H;(�H;\�H;�H;K�H;˲H;��H;�H;��H;��H;&�H;��H;J�H;-�H;��H;w�H;@�H;��H;��H;��H;g�H;��H;O�H;��H;��H;��H;��H;��H;M�H;��H;e�H;��H;��H;��H;;�H;t�H;��H;(�H;C�H;��H;"�H;��H;��H;�H;��H;ʲH;K�H;�H;\�H;*�H;��H;~H;�tH;)kH;HbH;	ZH;�RH;>LH;GH;OCH;�@H;       H;H;BH;KH;H;�%H;{/H;m:H;UFH;�RH;A_H;�kH;-xH;4�H;��H;~�H;g�H;m�H;x�H;��H;P�H;��H;��H;�H;��H;��H;U�H;w�H;#�H;��H;��H;��H;U�H;��H;C�H;s�H;��H;s�H;C�H;��H;V�H;��H;��H;��H;�H;q�H;U�H;��H;��H;�H;��H;��H;K�H;��H;z�H;f�H;d�H;|�H;��H;3�H;,xH;�kH;B_H;�RH;TFH;q:H;/H;�%H;'H;HH;BH;H;      ��G;<�G;B�G;��G;��G;
�G;��G;RH;�H;7'H;�7H;gHH;�XH;#hH;wH;��H;��H;��H;8�H;��H;�H;/�H;j�H;��H;o�H;T�H;��H;9�H;z�H;>�H;��H;��H;��H;a�H;��H;��H;�H;��H;��H;c�H;��H;��H;��H;=�H;t�H;4�H;��H;[�H;j�H;��H;o�H;+�H;�H;��H;8�H;��H;��H;��H;wH;"hH;�XH;gHH;�7H;6'H;�H;NH;��G;��G;��G;��G;P�G;<�G;      �nG;$qG;�wG;΂G;ېG;9�G;_�G;��G;��G;"�G;�H;EH;v0H;�DH;XH;jH;�zH;�H;��H;��H;X�H;��H;��H;~�H;,�H;�H;9�H;��H;^�H;x�H;H�H;��H;��H;��H;4�H;��H;��H;��H;2�H;��H;��H;��H;K�H;x�H;Y�H;��H;9�H; �H;-�H;u�H;��H;��H;T�H;��H;��H;��H;�zH;jH;XH;�DH;w0H;GH;�H; �G;��G;��G;^�G;5�G;ߐG;ʂG;�wG;qG;      �F;��F;��F;��F;��F;!G;�FG;'jG;-�G;�G;��G;��G;�G;lH;i1H;�HH;^H;hqH;�H;q�H;%�H;ݫH;�H;�H;��H;�H;�H;Z�H;��H;��H;��H;��H;��H;��H;x�H;��H;
�H;��H;u�H;��H;��H;��H;��H;��H;��H;X�H;�H;�H;��H;{�H;�H;۫H; �H;q�H;�H;bqH;^H;�HH;j1H;kH;�G;��G;��G;��G;%�G;"jG;�FG;m!G;��F;��F;��F;��F;      ��D;��D;��D;�9E;j�E;,�E;KPF;�F;��F;:G;9oG;��G;޿G;��G;�H;`H;�:H;�SH;�iH;B}H;��H;��H;J�H;�H;A�H;��H;)�H;m�H;��H;'�H;��H;�H;��H;��H;��H;"�H;c�H;!�H;��H;��H;��H;�H;��H;*�H;��H;j�H;,�H;��H;=�H;�H;M�H;��H;��H;C}H;�iH;�SH;�:H;^H;�H;��G;�G;��G;6oG;:G;��F;�F;FPF;!�E;o�E;�9E;��D;��D;      ?@;@A@;�@;"RA;�"B;C;B�C;��D;#�E;@F;t�F;�!G;hG;��G;0�G;��G;yH;�.H;	KH;�cH;MyH;�H;1�H;ƩH;�H;x�H;u�H;��H;�H;K�H;��H;M�H;:�H;��H;��H;[�H;��H;\�H;��H;��H;<�H;J�H;��H;N�H;�H;��H;u�H;�H;�H;éH;3�H;�H;JyH;�cH;KH;�.H;vH;��G;-�G;��G;�gG;�!G;q�F;~@F;�E;{�D;?�C; C;�"B;4RA;�@;(A@;      q46;A�6;�k7;4�8;v�:;=�<;%�>;H�@;�tB;S�C;�,E;�F;�F;�,G;�xG;+�G;c�G;�H;�%H;EH;`H;IwH;0�H;7�H;M�H;�H;��H;m�H;��H;��H;)�H;A�H;��H;]�H;��H;p�H;��H;n�H;��H;\�H;��H;A�H;,�H;��H;��H;k�H;��H;�H;H�H;5�H;/�H;EwH;`H;EH;�%H;�H;b�G;'�G;�xG;�,G;�F;�F;�,E;R�C;�tB;J�@;$�>;;�<;r�:;0�8;�k7;*�6;      c�";zM#;%;o�';-�+;D�/;��3;h 8;��;;?;�A;��C;�9E;�@F;��F;�UG;ǚG;'�G;��G;M H;�AH;�^H;EwH;�H;��H;٫H;��H;-�H;��H;#�H;�H;��H;��H;��H;j�H;G�H;|�H;H�H;i�H;��H;��H;��H;#�H;(�H;��H;+�H;��H;ޫH;��H;�H;EwH;�^H;�AH;L H;��G; �G;ŚG;�UG;��F;�@F;�9E;��C;��A;?;��;;k 8;��3;-�/;D�+;a�';%;lM#;      ���:H% ;Z�;��;�;Q;0m;Cd';�.;u=5;�:;��>;�B;BD;l�E;S�F;�6G;��G;��G;�G;zH;�AH;
`H;MyH;��H;�H;M�H;�H;K�H;��H;��H;2�H;��H;E�H;��H;��H;G�H;��H;��H;@�H;��H;/�H;��H;��H;I�H;�H;Q�H; �H;�H;MyH;`H;�AH;wH;�G;��G;��G;�6G;P�F;k�E;BD;�B;��>;�:;x=5;�.;Gd';4m;�P;%�;��;h�;4% ;      �Y�:)o�:�W�:/�:
&�:{��:o��::�	;Q;�M#;�n-;Q�5;��;;�A@;�PC;$GE;�uF;�!G;f�G;��G;�G;L H;EH;�cH;?}H;r�H;��H;��H;üH;��H;��H;,�H;U�H;U�H;N�H;w�H;��H;w�H;K�H;P�H;R�H;)�H;��H;��H;¼H;��H;��H;u�H;9}H;�cH;EH;I H;�G;��G;c�G;�!G;�uF;!GE;�PC;�A@;��;;Q�5;�n-;�M#;Q;3�	;g��:i��:&�:�:�W�:o�:      d�	����pj��@[���4u9p:�j~:1��:�[�:��;|�;^%;�t0;��8;�>;�B;��D;hXF;:G;c�G;��G;��G;�%H;KH;�iH;�H;��H;7�H;w�H;�H;^�H;��H;��H;3�H;�H;��H;S�H;��H;~�H;2�H;��H;��H;`�H;�H;v�H;7�H;��H;�H;�iH;	KH;�%H;��G;��G;c�G;8G;dXF;��D;�B;�>;��8;�t0;\%;|�;��;�[�:7��:�j~:l:�4u9�[���j������      |A?�̡9�"9)��Z�zܺRp��0���0<9$�@:��:C�:]�	;zY;>,;Ԅ6;|�=;%#B;��D;dXF;�!G;��G;#�G;�H;�.H;SH;_qH;܉H;��H;h�H;��H;r�H;��H;��H;��H;��H;�H;��H;�H;|�H;��H;��H;��H;t�H;��H;f�H;��H;߉H;_qH;xSH;�.H;�H;�G;|�G;�!G;cXF;��D;!#B;x�=;Ԅ6;>,;xY;\�	;G�:��: �@:<98���`p���ܺ�Z�+9)�ˡ9�      �EֻN�ѻ��ĻjT���񕻲.o�ԝ.�2ܺ��B�@��8�\:�&�:���:AQ;�);�=5;�:=;+#B;��D;�uF;�6G;ǚG;b�G;vH;�:H;^H;�zH;��H;g�H;ĲH;	�H;��H;\�H;�H;m�H;0�H;��H;0�H;j�H;�H;X�H;��H;�H;ǲH;d�H;��H;�zH;^H;�:H;vH;`�G;ÚG;�6G;�uF;��D;%#B;�:=;�=5;�);AQ;���:�&�:�\: ��8x�B�1ܺ؝.��.o���nT����ĻJ�ѻ      OFB�:�>���4�R�$�q��[�����ݎ�^A?�aӺ����3�9�q�:bX�:^;��';�=5;�=;�B;GE;S�F;�UG;'�G;��G;ZH;�HH;jH;��H;|�H;H�H;4�H;H�H;��H;D�H;�H;�H;��H;�H;
�H;>�H;��H;F�H;4�H;K�H;z�H;��H;jH;�HH;UH;��G;%�G;�UG;H�F;GE;�B;{�=;�=5;��';\;`X�:�q�:�3�9���aӺ^A?��ݎ����[�t��S�$���4�9�>�      gy��>ݜ��A���I����s���P��%+������Ļ����0|���o��:u9aX�:�+�:^;�);ӄ6;{�>;�PC;k�E;��F;�xG;-�G;~H;f1H;XH;wH;��H;�H;�H;~�H;�H;C�H;��H;��H;��H;��H;��H;A�H;�H;z�H;�H;�H;��H; wH;XH;b1H;zH;-�G;�xG;��F;a�E;�PC;x�>;Є6;�);V;�+�:YX�:�:u9�o�2|�������Ļ����%+���P���s��I���A��>ݜ�      l�����W�˖ռ�վ�)Ϥ��I����[�(��Z����9��{�� <9aX�:hX�:AQ;>,;��8;�A@;BD;�@F;�,G;��G;��G;hH;�DH;hH;4�H;V�H;j�H;`�H;"�H;�H;��H;��H;c�H;��H;��H;�H;�H;[�H;g�H;Y�H;3�H;hH;�DH;dH;��G;��G;�,G;�@F;BD;�A@;��8;<,;AQ;ZX�:YX�:�;9�{����9���Z�(���[��I��)Ϥ��վ�˖ռ�W���      1�6�F�3���+���`�h�����μ���y���PFB�es�=T��"�D��{��;u9�q�:���:}Y;�t0;��;;�B;�9E;�F;hG;ݿG;�G;y0H;�XH;.xH;$�H;y�H;�H;��H;��H;�H;.�H;2�H;.�H;�H;��H;��H;��H;w�H;'�H;-xH;�XH;y0H;��G;׿G;hG;�F;�9E;�B;��;;�t0;xY;���:�q�:�:u9�{��'�D�>T��es�QFB�y��������μh���b�����+�F�3�      o₽�؀���u��Xc���K�w1����ߤ��վ��]����P����>T����9���o��3�9�&�:]�	;_%;N�5;��>;��C;�F;�!G;��G;��G;DH;`HH;�kH;��H;N�H;��H;��H;w�H;J�H;��H;��H;��H;H�H;u�H;��H;��H;L�H;��H;�kH;^HH;BH;��G;��G;�!G;�F;��C;��>;N�5;[%;]�	;~&�:�3�9��o���9�?T�������P��]���վ�ߤ���v1���K��Xc���u��؀�      8S���r��r�����Г����u���N���(��i�Ɍ˼�A����P�es��2|� ����\:1�:s�;~n-;�:;��A;�,E;k�F;-oG;��G;�H;�7H;>_H;~H;�H;�H;v�H;�H;x�H;;�H;��H;<�H;w�H;�H;q�H;��H;�H;~H;@_H;�7H;�H;��G;)oG;m�F;�,E;��A;ޞ:;~n-;o�;-�:�\:@���6|��fs���P��A��ʌ˼�i���(���N���u�ѓ�����r���r��      �o��s��罫�ս4@��pĥ�x^���Xc�C�3���	�Ɍ˼�]��QFB��Z򻪜��aӺ���8��:ߛ;�M#;{=5;?;O�C;~@F;	:G;�G;�G;0'H;�RH;|tH;��H;{�H;-�H;��H;��H;��H;?�H;��H;��H;��H;(�H;w�H;��H;}tH;�RH;0'H;�G;�G;:G;~@F;R�C;?;p=5;�M#;ܛ;��:���8gӺ�����Z�RFB��]��Ɍ˼��	�C�3��Xc�x^��pĥ�5@����ս���s�      �#�U� �_'������gٽ7S��'l��M�j�C�3��i��վ�y���(���ĻZA?���B� �@:�[�:Q;
�.;��;;tB;�E;��F;&�G;��G;�H;VFH;&kH;��H;�H;�H;h�H;�H;p�H;��H;o�H;
�H;g�H;�H;�H;��H;(kH;UFH;�H;��G;(�G;��F;�E;tB;��;;�.;Q;�[�: �@:��B�^A?���Ļ(�y����վ��i�C�3�M�j�'l��7S���gٽ����_'�U� �      �S�&�O��E��5�U� �X�
���罤9��'l���Xc���(��������[�����ݎ�<ܺ@;9+��:3�	;Hd';h 8;@�@;��D;�F;jG;��G;LH;q:H;AbH;��H;�H;4�H;C�H;{�H;6�H;��H;5�H;}�H;C�H;.�H;�H;��H;HbH;q:H;NH;��G;jG;�F;�D;@�@;e 8;Cd';4�	;#��:p;9;ܺ�ݎ������[��������(��Xc�'l���9�����X�
�U� ��5��E�&�O�      �~��*��(�v��9b�z�H�#,�LZ����7S��x^����N������μ�I���%+����֝.������j~:O��:/m;��3;�>;>�C;=PF;�FG;P�G;��G;y/H;ZH;wzH;G�H;��H;]�H;�H;)�H;��H;&�H;�H;]�H;��H;E�H;tzH;ZH;{/H;��G;S�G;�FG;=PF;?�C;�>;��3;)m;Y��:�j~:����ם.�����%+��I����μ�����N�x^��7S�����MZ�#,�z�H��9b�(�v�*��      ����(����:���M��E�r�&�O�#,�X�
��gٽpĥ���u�w1�h���)Ϥ���P�[�.o�pp��H:k��:�P;=�/;:�<;C;�E;n!G;4�G;�G;�%H;�RH;�tH;��H;F�H;ׯH; �H;X�H;�H;X�H;�H;ׯH;D�H;��H;�tH;�RH;�%H;�G;5�G;u!G;�E;C;9�<;:�/;�P;m��:<:np���.o�[򻩎P�)Ϥ�h���w1���u�pĥ��gٽX�
�#,�&�O�E�r��M���:��(���      8���v��M;������RP��E�r�z�H�T� ���5@��Г����K�`��վ���s�q���񕻠ܺ 5u9&�:$�;/�+;|�:;�"B;o�E;��F;ԐG;��G;/H;5LH;�oH;:�H;r�H;��H;2�H;׼H;��H;ӼH;4�H;��H;r�H;9�H;�oH;<LH;/H;��G;ڐG;��F;n�E;�"B;|�:;-�+;!�;&�:�4u9�ܺ��q����s��վ�a���K�ѓ��5@����U� �z�H�E�r�RP������M;���v��      VVھ�*־/5ʾr��������M���9b��5�����ս����Xc���ʖռ�I��T�$�jT���Z� \���:�;j�';�8;RA;�9E;��F;ÂG;��G;AH;GH;lH;C�H;9�H;�H;��H;��H;Q�H;��H;õH;�H;9�H;C�H;lH;GH;CH;��G;ƂG;��F;�9E;RA;�8;h�';��;�:`\���Z�jT��T�$��I��ʖռ���Xc������ս���5��9b��M������r���/5ʾ�*־      ���쾳�޾/5ʾL;���:��(�v��E�_'����q����u���+��W��A����4���Ļ9)�`j���W�:d�;%;�k7;$�@;��D;��F;�wG;T�G;4H;>CH;*iH;�H;��H;��H;��H;��H;r�H;��H;��H;��H;��H;�H;&iH;DCH;5H;U�G;�wG;��F;��D;$�@;�k7;%;b�;�W�:`j��9)���Ļ��4��A���W缂�+���u�q�����_'��E�(�v��:��L;��/5ʾ��޾��      Vh���b���쾧*־�v��(���*��'�O�U� �s��r���؀�G�3���>ݜ�;�>�Q�ѻޡ9�����'o�:A% ;tM#;C�6;LA@;��D;��F;qG;L�G;H;�@H;hgH;��H;��H;ީH;�H;��H;�H;��H;�H;ߩH;��H;��H;cgH;�@H;H;L�G;qG;��F;��D;LA@;?�6;pM#;<% ;-o�:����ܡ9�R�ѻ;�>�>ݜ���F�3��؀��r��s�U� �'�O�*��(����v���*־���b��      ���^�T_ݾ��ɾj*��쫖�{x�&G�P,�����b��]@{���/�����䙼�J;�M�ͻ��4� W���:6;��#;�6;[@;3�D;��F;�lG;��G;7H;�:H;�bH;߀H;,�H;/�H;ٱH;��H;ܹH;�H;رH;/�H;*�H;ۀH;�bH;�:H;6H;��G;�lG;��F;3�D;[@;�6;��#;4;��:W���4�L�ͻ�J;��䙼����/�]@{��b�����P,�&G�{x�쫖�i*����ɾT_ݾ^�      ^�3���:پ{�žg�����9t�p�C�������㪫�W`w�F-����)`����7�4Sɻ�K/��xƹ���:�/;�f$;�7;�~@;K�D;\�F;�nG;��G;"H;�;H;jcH;p�H;��H;q�H;�H;.�H;"�H;*�H;	�H;o�H;��H;m�H;dcH;�;H;#H;��G;�nG;f�F;K�D;�~@;�7;�f$;�/;���:�xƹ�K/�4Sɻ��7�)`�����E-�W`w�㪫�������p�C�9t���g���{�ž�:پ3��      U_ݾ�:پ�V;+���Ƥ�La����g��$:��Z�oݽ�ƣ�zl�e.%��߼g���9.�ʴ��JV�`1p��@�:x;N(&;4�7;:�@;�
E;��F;huG;$�G;OH;�=H;MeH;ĂH;u�H;M�H;��H;��H;��H;��H;��H;M�H;r�H;ÂH;GeH;�=H;OH;&�G;kuG;��F;�
E;6�@;.�7;L(&;x;�@�:�1p�JV�ʴ���9.�f���߼e.%�zl��ƣ�oݽ�Z��$:���g�La���Ƥ�+���V;�:پ      ��ɾ{�ž+��qת�쫖�!�����T��J+�:��2̽�s���yZ����Mμfy����[Ϩ�N,� �6��:��
;_�(;WN9;�A;|NE;0�F;�G;��G;|H;�AH;1hH;�H;A�H;թH;ͳH;��H;x�H;��H;ϳH;ԩH;=�H;�H;-hH;�AH;|H;��G;�G;9�F;~NE;��A;RN9;\�(;��
;��: �6J,�[Ϩ���ey��Mμ����yZ��s���2̽:��J+���T�!���쫖�qת�+��|�ž      j*��g����Ƥ�쫖��/��>�c��G=�����zｐж��ɇ�Q�C�
��""��p;k��&��-��l�˺8Y�9v��:9;�h,;�	;;�PB;b�E;� G;܌G;��G;hH;GH;OlH; �H;��H;��H;;�H;�H;ּH;�H;<�H;��H;��H;��H;JlH;GH;hH;��G;ߌG;� G;d�E;�PB;�	;;�h,;9;���:0Y�9j�˺�-���&�o;k�""��
��Q�C��ɇ��ж��z�����G=�>�c��/��쫖��Ƥ�g���      쫖���La��!���>�c�p�C�z#���RvϽ����zl�dg*����
���I���軼\c�퀺�t,:���:��;�_0;f�<;�1C;��E;t#G;S�G;	�G; H;�MH;6qH;��H;}�H;ޭH;*�H;��H;_�H;��H;,�H;ۭH;{�H;��H;5qH;�MH; H;�G;S�G;|#G;��E;�1C;c�<;�_0;�;���:�t,:퀺�\c�����I��
�����dg*�zl�����RvϽ��z#�p�C�>�c�!���La����      {x�9t���g���T��G=�z#�6�oݽ�b������AG����ލǼgy��I�$�c����$��uƹQ��:�&�:�� ;L4;t�>;ND;�[F;�FG;��G;�G;�)H;\UH;�vH;��H;�H;��H;j�H;��H;,�H;��H;l�H;��H;�H;��H;�vH;fUH;�)H;�G;~�G;�FG;�[F;ND;q�>;M4;�� ;�&�:Q��:�uƹ�$�d���I�$�gy��ލǼ���AG������b��nݽ6�z#��G=���T���g�9t�      %G�p�C��$:��J+������oݽ]���.I���yZ��"����ҫ��bT��� �M����˺�m9=ٶ:g�;`(;�8;d�@;��D;ޱF;>hG;��G;�H;/5H;�]H;e}H;�H;��H;S�H;ƻH;��H;5�H;��H;̻H;V�H;��H;�H;c}H;�]H;15H;�H;��G;DhG;�F;��D;d�@;�8;	`(;o�;=ٶ:�m9��˺M���� �bT�ҫ������"��yZ�-I��]���oݽ������J+��$:�p�C�      P,�����Z�:��z�RvϽ�b��-I��f]a�F-�g� � "��v�{�D�!�������4��P(�oQ:�L�:��;֊/;�'<;ڟB;��E;��F;��G;��G;4H;<AH;gH;M�H;3�H;ϪH;��H;~�H;��H;Q�H;��H;��H;��H;̪H;3�H;O�H;gH;@AH;6H;��G;��G;��F;��E;ݟB;�'<;֊/;�;�L�:�nQ:�P(���4�����C�!�u�{� "��g� �F-�f]a�-I���b��RvϽ�z�:��Z����      ������oݽ�2̽�ж����������yZ�F-�շ�-aļXO���J;����x�|���º�N@9ǂ�:>�;�f$;��5;�N?;:D;�LF;�:G;��G;��G;�!H;�MH;�pH;��H;ПH;/�H;�H;?�H;s�H;��H;q�H;B�H;�H;-�H;͟H;��H;�pH;�MH;�!H;��G;��G;�:G;�LF;;D;�N?;��5;�f$;@�;ǂ�:�N@9��ºt�|���軾J;�XO��-aļշ�F-��yZ����������ж��2̽oݽ���      �b��㪫��ƣ��s���ɇ�zl�BG��"�h� �-aļa���I��C��ۙ�@�uƹV�k:���:�;>>.;
;;��A;�AE;^�F;mG;��G;��G;U2H;�ZH;�zH;֒H;��H;��H;X�H;*�H;��H;�H;��H;,�H;[�H;��H;��H;ؒH;�zH;�ZH;X2H;��G;��G;mG;\�F;�AE;��A;
;;J>.;�;���:n�k:uƹ<��ۙ��C��I�a��-aļg� ��"�BG�zl��ɇ��s���ƣ�㪫�      \@{�W`w�zl��yZ�Q�C�dg*�������!"��XO���I�=|�7Ϩ�jK/�l$T�<Q:X��:��;�(&;�#6;�%?;��C;r#F;�#G;�G;��G;�H;)CH;�gH;}�H;X�H;k�H;�H;��H;�H;��H;��H;��H;�H;��H;�H;g�H;[�H;��H;�gH;*CH;�H;��G;"�G;�#G;w#F;��C;�%?;�#6;�(&;��;f��:HQ:d$T�fK/�6Ϩ�;|��I�XO�� "����鼮��cg*�R�C��yZ�zl�V`w�      ��/�E-�e.%����	�����ލǼѫ��v�{��J;��C�8Ϩ�FO:�����X[�9���:r;��;;.1;�'<;�5B;�NE;�F;1fG;�G;.�G;�*H;�SH;�tH; �H;��H; �H;L�H;w�H;��H; �H;�H; �H;��H;y�H;J�H;�H;��H;(�H;�tH;�SH;�*H;*�G;�G;1fG;�F;�NE;�5B;(<;D.1;��;x;���:x[�9����CO:�5Ϩ��C��J;�t�{�ѫ��ލǼ��������e.%�E-�      ������߼Nμ "���
��gy��aT�D�!���軺ۙ�lK/����� m9�A�:���:0�;D�,;�N9;@@;�^D;�LF;T.G;�G;��G;�H;�?H;dH;�H;n�H;�H;��H;��H;��H;��H;��H;v�H;��H;��H;��H;��H;��H;	�H;v�H;�H;dH;�?H;�H;��G;�G;Z.G;�LF;�^D;I@;�N9;C�,;9�;���:�A�:0m9����gK/��ۙ����B�!�_T�gy���
��""��Nμ�߼���      �䙼*`��h��fy��n;k��I�I�$��� �����t�|�;��$T�P[�9�A�:j��:"�;�);+7;��>;�tC;�E;��F;�uG;�G;��G;�+H;�SH;�sH;��H;a�H;�H;̻H;��H;4�H;n�H;��H;��H;��H;n�H;7�H;��H;ȻH;�H;g�H;��H;�sH;�SH;�+H;��G;�G;�uG;��F;�E;�tC;��>;'7; �);$�;l��:�A�:h[�9l$T�8�s�|������� �I�$��I�r;k�fy��h��)`��      �J;���7��9.����&����^���M����4���º uƹ8Q:���:���:"�;��(;��5;��=;��B;�[E;C�F;�TG;��G;��G;�H;�CH;fH;ɁH;u�H;��H;��H;��H;��H;U�H;��H;>�H;�H;<�H;��H;T�H;��H;��H;��H;��H;y�H;ˁH;fH;�CH;�H;��G;��G;�TG;G�F;�[E;��B;��=;��5;��(;&�;���:���:HQ:�tƹ��º��4�M��_�����軩&����9.���7�      F�ͻ1Sɻδ��^Ϩ��-���\c��$���˺�P(�O@9r�k:Z��:v;5�;�);��5;L�=;*QB;kE;�F;%8G;C�G;C�G;�	H;U5H;�YH;AwH;؎H;��H;ӰH;��H;��H;T�H;!�H;��H;u�H;�H;q�H;~�H;#�H;P�H;��H;��H;ְH;��H;َH;BwH;�YH;[5H;�	H;C�G;E�G;'8G;�F;oE;$QB;N�=;��5; �);7�;v;`��:z�k: O@9xP(���˺�$��\c��-��aϨ�Ӵ��,Sɻ      ��4��K/�NV�@,�N�˺�쀺puƹ�m9oQ:ӂ�:���:��;|�;A�,;$7;��=;QB;��D;�cF;$G;̇G;��G;��G;x)H;�NH;�mH;܆H;ŚH;%�H;�H;�H;��H;��H;��H;��H;w�H;�H;u�H;��H;��H;��H;��H;�H;�H;(�H;ŚH;܆H;�mH;�NH;x)H;��G;��G;ЇG;!$G;�cF;��D;#QB;��=;'7;A�,;�;��;���:т�:oQ:0m9�uƹ�쀺H�˺H,�FV��K/�      0V�(yƹ�1p� *�68Y�9�t,:i��:Iٶ:�L�:C�;�;�(&;?.1;�N9;��>;��B;lE;�cF;�G;*�G;��G;��G;V H;�EH;�eH;�H;��H;ҥH;��H;��H;�H;��H;��H;R�H;��H;J�H;��H;G�H;��H;Q�H;��H;��H;�H;��H;��H;ԥH;��H;�H;�eH;�EH;S H;��G;¿G;0�G;�G;�cF;qE;��B;��>;�N9;A.1;�(&;�;D�;�L�:Kٶ:c��:�t,:@Y�9 �6�1p�yƹ      ���:���: A�:5��:t��:���:�&�:g�;��;�f$;H>.;�#6;(<;G@;�tC;�[E;�F;&$G;-�G;��G;�G;�H;�?H;�_H;�yH;^�H;�H;��H;0�H;v�H;��H;N�H;q�H;��H;��H;�H;g�H;��H;��H;��H;p�H;J�H;��H;v�H;0�H;��H;�H;Z�H;�yH;�_H;�?H;�H;�G;��G;1�G;#$G;�F;�[E;�tC;F@;(<;�#6;L>.;�f$;�;p�;�&�:��:|��:��:�@�:���:      Z;�/;�w;�
;9;��;�� ;`(;Պ/;��5;
;;�%?;�5B;�^D;�E;G�F;%8G;؇G;��G;�G;�H;�<H;�[H;�uH;��H;U�H;:�H;>�H;��H;��H;��H;i�H;�H;��H;|�H;�H;��H;x�H;|�H;��H;�H;d�H;��H;��H;��H;>�H;7�H;T�H;��H;�uH;�[H;�<H;�H;�G;¿G;ՇG;)8G;I�F;�E;�^D;�5B;�%?; 
;;��5;ӊ/;`(;�� ;�;9;�
;x;�/;      ��#;�f$;Z(&;i�(;�h,;�_0;J4;�8;�'<;�N?;��A;��C;�NE;�LF;��F;�TG;D�G;��G;��G;�H;�<H;nZH;�sH;��H;��H;��H;ԵH;ɿH;��H;�H;:�H;3�H;T�H;v�H;��H;��H;�H;��H;��H;v�H;Q�H;/�H;>�H;�H;��H;˿H;еH;��H;��H;��H;�sH;pZH;�<H;�H;��G;��G;G�G;�TG;��F;�LF;�NE;��C;��A;�N?;�'<;�8;P4;�_0;�h,;^�(;N(&;�f$;      /�6;�7;.�7;dN9;�	;;m�<;��>;p�@;�B;BD;�AE;y#F;�F;b.G;�uG;��G;G�G;��G;V H;�?H;�[H;�sH;7�H;X�H;�H;*�H;��H;%�H;��H;$�H;N�H;��H;B�H;.�H;=�H;��H;0�H;��H;:�H;/�H;?�H;��H;R�H;$�H;��H;(�H;��H;*�H;�H;W�H;4�H;�sH;�[H;�?H;X H;��G;H�G;��G;�uG;^.G;�F;}#F;�AE;=D;�B;q�@;��>;j�<;�	;;cN9;+�7;�7;      [@;�~@;,�@;��A;�PB;�1C;RD;��D;��E;�LF;b�F;�#G;1fG;�G;�G;��G;�	H;)H;�EH;�_H;�uH;�H;U�H;d�H;;�H;�H;(�H;��H;Q�H;��H;�H;��H;��H;j�H;i�H; �H;B�H;��H;g�H;j�H;��H;��H;�H;��H;Q�H;��H;$�H;�H;>�H;c�H;S�H;��H;�uH;�_H;�EH;x)H;�	H;��G;�G;�G;1fG; $G;e�F;�LF;��E;��D;SD;�1C;�PB;��A;/�@;�~@;      V�D;I�D;�
E;uNE;`�E;��E;�[F;ޱF;��F;�:G;mG;%�G;�G;��G;��G;�H;_5H;�NH;�eH;�yH;��H;��H;�H;B�H;��H;��H;)�H;��H;��H;y�H;P�H;��H;R�H;z�H;z�H;��H;�H;��H;x�H;|�H;O�H;��H;U�H;z�H;��H;��H;#�H;��H;��H;@�H;��H;��H;��H;�yH;�eH;�NH;a5H;�H;��G;��G;�G;+�G;mG;;G;��F;�F;�[F;��E;h�E;pNE;�
E;I�D;      ��F;a�F;��F;/�F;� G;#G;�FG;NhG;��G;��G;��G;��G;1�G;�H;�+H;�CH;�YH;�mH;�H;Y�H;T�H;��H;%�H;�H;��H;��H;4�H;��H;�H;�H;[�H;�H;��H;~�H;]�H;��H;��H;��H;[�H;~�H;��H;�H;[�H;�H;�H;��H;.�H;��H;��H;�H;%�H;��H;T�H;V�H;�H;�mH;�YH;�CH;�+H;�H;1�G;��G;��G;��G;��G;PhG;�FG;t#G;� G;:�F;��F;d�F;      �lG;�nG;juG;�G;ՌG;P�G;��G;~�G;��G;��G;��G;�H;�*H;�?H;�SH;fH;EwH;�H;��H;�H;>�H;ѵH;�H;+�H;(�H;4�H;T�H;��H;��H;(�H;�H;h�H;��H;m�H;��H;\�H;x�H;U�H;��H;n�H;��H;d�H;�H;(�H;��H;��H;M�H;7�H;*�H;&�H;�H;ҵH;>�H;�H;��H;چH;EwH;fH;�SH;�?H;�*H;�H;��G;��G;��G;��G;��G;L�G;�G;�G;kuG;�nG;      ��G;��G;�G;��G;��G;�G;�G;�H;8H;�!H;[2H;0CH;�SH;dH;�sH;ʁH;؎H;ŚH;ԥH;��H;A�H;ȿH;!�H;��H;��H;��H;��H;��H;�H;��H;d�H;��H;t�H;6�H;|�H;��H;�H;��H;|�H;9�H;t�H;��H;d�H;��H;�H;��H;��H;��H;��H;��H;"�H;ȿH;>�H;��H;ѥH;��H;؎H;ˁH;�sH;dH;�SH;0CH;_2H;�!H;8H;�H;�G;��G;��G;��G; �G;��G;      3H;H;LH;�H;ZH; H;*H;+5H;6AH;�MH;�ZH;�gH;�tH;�H;��H;x�H;��H;,�H;��H;0�H;��H;��H;��H;P�H;��H;�H;��H;�H;��H;L�H;q�H;��H;3�H;��H;�H;L�H;V�H;F�H;�H;��H;6�H;��H;s�H;J�H;��H;�H;��H;�H;��H;L�H;��H;��H;��H;-�H;��H;(�H;��H;y�H;��H;�H;�tH;�gH;�ZH;�MH;9AH;+5H;*H; H;dH;�H;LH;H;      �:H;|;H;�=H;�AH;GH;�MH;cUH;�]H;gH;�pH;�zH;��H;'�H;x�H;d�H;��H;װH;�H;��H;s�H;��H;�H;�H;��H;y�H;�H;&�H;��H;J�H;��H;j�H;)�H;��H;1�H;��H;��H;��H;��H;��H;1�H;��H;%�H;j�H;��H;J�H;��H;!�H;�H;z�H;��H;"�H;�H;��H;p�H;��H;�H;װH;��H;d�H;u�H;'�H;��H;�zH;�pH;gH;�]H;cUH;�MH;GH;�AH;�=H;{;H;      �bH;{cH;QeH;3hH;MlH;9qH; wH;f}H;P�H;��H;��H;b�H;ǡH;�H;�H;��H;��H;�H;�H;��H;��H;>�H;O�H;�H;S�H;[�H;�H;h�H;t�H;p�H;;�H;��H;'�H;��H;��H;��H;�H;��H;��H;��H;*�H;��H;;�H;m�H;s�H;d�H;�H;^�H;V�H;�H;T�H;>�H;��H;��H;�H;�H;��H;��H;�H;�H;ɡH;d�H;��H;��H;S�H;i}H;	wH;/qH;WlH;1hH;SeH;}cH;      ހH;t�H;ĂH;߄H;��H;��H;�H;�H;9�H;ӟH;��H;r�H;&�H;��H;ϻH;��H;��H;��H;��H;S�H;o�H;4�H;��H;��H;��H;�H;d�H;��H;��H;*�H;��H;<�H;��H;��H;�H;9�H;-�H;9�H;�H;��H;��H;:�H;��H;)�H;��H;��H;b�H;�H;��H;��H;��H;6�H;i�H;N�H;��H;��H;��H;��H;һH;��H;&�H;r�H;��H;ӟH;9�H;�H;�H;��H;�H;�H;̂H;{�H;      ,�H;��H;��H;A�H;��H;{�H;�H;��H;˪H;2�H;��H;�H;V�H;��H;��H;��H;X�H;��H;��H;w�H;�H;U�H;?�H;��H;S�H;��H;��H;z�H;9�H;��H;&�H;��H;��H;�H;Q�H;b�H;/�H;b�H;N�H;�H;��H;��H;%�H;��H;7�H;w�H;��H;��H;V�H;��H;C�H;T�H;�H;s�H;��H;��H;Z�H;��H;��H;��H;V�H;�H;��H;3�H;ΪH;��H;�H;u�H;��H;:�H;��H;��H;      -�H;k�H;O�H;ͩH;��H;ҭH;��H;W�H;��H;��H;h�H;��H;��H;��H;>�H;\�H;(�H;��H;V�H;��H;��H;y�H;+�H;a�H;w�H;z�H;i�H;9�H;��H;4�H;��H;��H;�H;I�H;h�H;o�H;��H;m�H;e�H;I�H;�H;��H;��H;0�H;��H;4�H;g�H;{�H;z�H;`�H;0�H;w�H;��H;��H;U�H;��H;-�H;\�H;>�H;��H;��H;��H;i�H;��H;��H;\�H;��H;ҭH;��H;ͩH;X�H;x�H;      ձH;�H;��H;гH;L�H;%�H;w�H;˻H;��H;M�H;7�H;)�H;��H;��H;x�H;��H;��H;��H;��H;��H;��H;��H;6�H;[�H;t�H;T�H;��H;{�H;�H;��H;��H;�H;Q�H;i�H;p�H;��H;��H;��H;m�H;i�H;S�H;�H;��H;��H;�H;v�H;��H;U�H;v�H;[�H;;�H;��H;z�H;��H;��H;��H;��H;�H;v�H;��H;��H;*�H;;�H;M�H;��H;ϻH;z�H;(�H;J�H;ӳH;��H;�H;      ��H;,�H;��H;��H;�H;��H;��H;��H;��H;�H;
�H;��H;�H;��H;��H;>�H;w�H;v�H;K�H; �H;��H;��H;��H;��H;��H;��H;W�H;��H;O�H;��H;��H;?�H;h�H;s�H;��H;��H;��H;��H;��H;w�H;j�H;=�H;��H;��H;L�H;��H;Y�H;��H;��H;��H;��H;��H;}�H;��H;J�H;y�H;{�H;A�H;��H;��H;�H;��H;�H;��H;�H;��H;��H;��H;�H;��H;��H;:�H;      �H;�H;κH;u�H;мH;`�H;3�H;9�H;Z�H;��H; �H;��H;,�H;��H;��H;&�H;)�H;�H;��H;l�H;��H;�H;.�H;8�H;�H;��H;u�H;�H;Z�H;��H;�H;1�H;1�H;��H;��H;��H;��H;��H;��H;��H;5�H;/�H;�H;��H;V�H;�H;u�H;��H;�H;8�H;3�H;�H;��H;h�H;��H;�H;)�H;'�H;��H;��H;,�H;��H;!�H;��H;^�H;=�H;5�H;_�H;ѼH;r�H;ϺH;(�H;      ��H;-�H;��H;��H;�H;��H;��H;��H;��H;�H;�H;��H;	�H;��H;��H;>�H;w�H;v�H;K�H; �H;��H;��H;��H;��H;��H;��H;W�H;��H;P�H;��H;��H;?�H;i�H;t�H;��H;��H;��H;��H;��H;v�H;j�H;=�H;��H;��H;L�H;��H;W�H;��H;��H;��H;��H;��H;}�H;��H;J�H;y�H;z�H;A�H;��H;��H;�H;��H;�H;�H;�H;��H;��H;��H;	�H;��H;��H;5�H;      ͱH;�H;��H;ȳH;L�H;#�H;x�H;ͻH;��H;M�H;8�H;)�H;��H;��H;y�H;��H;��H;��H;��H;��H;��H;��H;6�H;[�H;v�H;T�H;��H;{�H;�H;��H;��H;�H;P�H;i�H;p�H;��H;��H;��H;o�H;i�H;U�H;�H;��H;��H;�H;u�H;��H;X�H;s�H;Z�H;;�H;��H;y�H;��H;��H;��H;��H;�H;v�H;��H;��H;,�H;8�H;M�H;��H;ԻH;~�H;"�H;M�H;ȳH;��H;�H;      ,�H;j�H;O�H;ѩH;��H;׭H;��H;Z�H;��H;��H;i�H;��H;��H;��H;@�H;[�H;+�H;��H;V�H;��H;��H;|�H;+�H;c�H;|�H;z�H;j�H;9�H;��H;4�H;��H;��H;�H;I�H;f�H;m�H;��H;o�H;e�H;G�H;�H;��H;��H;0�H;��H;4�H;g�H;}�H;w�H;]�H;0�H;y�H;��H;��H;V�H;��H;+�H;]�H;@�H;��H;��H;��H;h�H;��H;��H;^�H;��H;ԭH;��H;˩H;W�H;k�H;      -�H;��H;~�H;=�H;��H;|�H;�H;��H;˪H;3�H;��H;�H;V�H;��H;��H;��H;W�H;��H;��H;w�H;�H;X�H;?�H;��H;W�H;��H;��H;z�H;;�H;��H;%�H;��H;��H;�H;P�H;c�H;/�H;b�H;P�H;�H;��H;��H;%�H;��H;3�H;u�H;��H;��H;R�H;��H;F�H;T�H;
�H;t�H;��H;��H;Z�H;��H;��H;��H;W�H;�H;��H;3�H;ϪH;��H;�H;y�H;��H;D�H;��H;��H;      ΀H;z�H;��H;݄H;��H;��H;�H;�H;6�H;ҟH;��H;q�H;$�H;��H;һH;��H;��H;��H;��H;S�H;p�H;9�H;��H;��H;��H;�H;b�H;��H;��H;)�H;��H;;�H;��H;��H;�H;6�H;-�H;8�H;�H;��H;��H;8�H;��H;(�H;��H;��H;`�H;�H;��H;��H;��H;6�H;h�H;N�H;��H;��H;��H;��H;лH;��H;&�H;r�H;��H;ԟH;<�H;�H;
�H;��H;��H;ބH;��H;q�H;      �bH;{cH;TeH;.hH;SlH;9qH;�vH;e}H;Q�H;��H;ߒH;d�H;ǡH;�H;�H;��H;��H;�H;�H;��H;��H;B�H;O�H;�H;V�H;X�H;�H;e�H;w�H;n�H;;�H;��H;'�H;��H;��H;��H;�H;��H;��H;��H;*�H;��H;:�H;k�H;p�H;b�H;�H;\�H;R�H;�H;U�H;@�H;��H;��H;�H;�H;��H;��H;�H;�H;ǡH;f�H;ߒH;��H;Q�H;l}H;wH;6qH;]lH;;hH;[eH;|cH;      �:H;�;H;�=H;�AH;
GH;�MH;bUH;�]H;gH;�pH;�zH;��H;'�H;v�H;g�H;��H;ְH;�H;��H;u�H;��H;�H;�H;��H;|�H;�H;$�H;��H;M�H;��H;j�H;)�H;��H;1�H;��H;��H;��H;��H;��H;1�H;��H;(�H;j�H;��H;H�H;��H;!�H;�H;w�H;��H;%�H;�H;��H;p�H;��H;�H;װH;��H;g�H;v�H;'�H;��H;�zH;�pH;gH;^H;fUH;�MH;GH;�AH;�=H;{;H;      >H;H;]H;�H;PH; H;*H;+5H;?AH;�MH;�ZH;�gH;�tH;�H;��H;y�H;��H;-�H;��H;0�H;��H;��H;��H;P�H;��H;�H;��H;�H;��H;I�H;q�H;��H;4�H;��H;�H;J�H;V�H;I�H;�H;��H;6�H;��H;s�H;J�H;��H;	�H;��H;�H;��H;I�H;��H;��H;��H;/�H;��H;(�H;��H;y�H;��H;�H;�tH;�gH;�ZH;�MH;=AH;15H;*H; H;cH;�H;]H;H;      ��G;��G;�G;��G;��G;�G;�G;�H;6H;�!H;[2H;-CH;�SH;dH;�sH;ˁH;؎H;ȚH;ҥH;��H;C�H;̿H;!�H;��H;��H;��H;��H;��H;�H;��H;e�H;��H;r�H;7�H;{�H;��H;�H;��H;{�H;7�H;u�H;��H;d�H;��H;�H;��H;��H;��H;��H;��H;'�H;ȿH;<�H;��H;ҥH;��H;َH;ˁH;�sH;dH;�SH;/CH;\2H;�!H;8H;�H;�G;�G;��G;��G; �G;��G;      �lG;�nG;euG;�G;�G;Y�G;��G;��G;��G;��G;��G;�H;�*H;�?H;�SH;fH;GwH;�H;��H;�H;A�H;յH;��H;.�H;*�H;1�H;Q�H;��H;��H;'�H;�H;i�H;��H;m�H;��H;W�H;x�H;W�H;��H;n�H;��H;g�H;�H;'�H;��H;��H;P�H;8�H;)�H;'�H;�H;ԵH;<�H; �H;��H;܆H;EwH;fH;�SH;�?H;�*H;�H;��G;��G;��G;��G;��G;S�G;�G;�G;kuG;�nG;      ��F;c�F;��F;/�F;� G;�#G;�FG;PhG;��G;��G;��G;��G;4�G;�H; ,H;�CH;�YH;�mH;�H;W�H;X�H;��H;%�H;�H;��H;��H;1�H;��H;�H;�H;Z�H;�H;��H;~�H;\�H;��H;��H;��H;[�H;~�H;��H;�H;^�H;�H;�H;��H;1�H;��H;��H;�H;'�H;��H;T�H;Y�H;�H;�mH;�YH;�CH;,H;�H;3�G;��G;��G;��G;��G;LhG;�FG;u#G;� G;-�F;��F;R�F;      U�D;F�D;�
E;wNE;^�E;��E;�[F;߱F;��F;;G;mG;)�G;�G;��G;��G;�H;_5H;�NH;�eH;�yH;��H;��H;�H;D�H;��H;��H;%�H;��H;��H;v�H;S�H;��H;O�H;z�H;z�H;��H;�H;��H;x�H;|�H;R�H;��H;V�H;y�H;��H;��H;&�H;��H;��H;@�H;��H;��H;��H;�yH;�eH;�NH;a5H;�H;��G;��G;�G;(�G;mG;�:G;��F;߱F;�[F;��E;g�E;qNE;�
E;F�D;      �Z@;�~@;)�@;�A;�PB;�1C;UD;��D;�E;�LF;f�F;$G;1fG;�G;�G;��G;�	H;)H;�EH;�_H;�uH;��H;S�H;e�H;A�H;�H;&�H;��H;S�H;��H;	�H;��H;��H;j�H;h�H;��H;B�H;��H;g�H;h�H;��H;��H;�H;��H;S�H;��H;'�H;�H;=�H;e�H;U�H;��H;�uH;�_H;�EH;z)H;�	H;��G;�G;�G;0fG;�#G;c�F;�LF;��E;��D;RD;�1C;QB;�A;(�@;�~@;      $�6;�7;�7;lN9;�	;;k�<;��>;p�@;�B;AD;�AE;}#F;�F;b.G;�uG;��G;J�G;��G;X H;�?H;�[H;�sH;5�H;Z�H;��H;%�H;��H;%�H;��H; �H;Q�H;��H;A�H;.�H;=�H;��H;3�H;��H;:�H;,�H;A�H;��H;T�H;%�H;��H;$�H;�H;*�H;�H;W�H;5�H;�sH;�[H;�?H;X H;��G;H�G;��G;�uG;].G;�F;y#F;�AE;?D;�B;q�@;�>;h�<;�	;;gN9;�7;�7;      ��#;�f$;P(&;_�(;�h,;�_0;Q4;�8;�'<;�N?;��A;��C;�NE;�LF;��F;�TG;G�G;��G;��G;�H;�<H;qZH;�sH;��H;��H;��H;ѵH;˿H;��H;�H;>�H;4�H;R�H;w�H;��H;��H;�H;��H;��H;u�H;T�H;2�H;@�H;�H;��H;ɿH;ҵH;��H;��H;��H;�sH;pZH;�<H;�H;��G;��G;C�G;�TG;��F;�LF;�NE;��C;��A;�N?;�'<;�8;I4;�_0;�h,;T�(;P(&;�f$;      P;�/;x;��
;9;��;�� ;`(;ي/;��5;
;;�%?;�5B;�^D;�E;K�F;)8G;؇G;¿G;�G;�H;�<H;�[H;�uH;��H;T�H;5�H;<�H;��H;��H;��H;i�H;
�H;��H;|�H;{�H;��H;}�H;z�H;��H;�H;h�H;��H;��H;��H;<�H;:�H;U�H;��H;�uH;�[H;�<H;�H;�G;��G;чG;%8G;G�F;�E;�^D;�5B;�%?;
;;��5;֊/;`(;�� ;��;9;��
;x;�/;      /��:���:�@�:3��:x��:��:�&�:r�;�;�f$;N>.;�#6;(<;G@;�tC;�[E;�F;($G;0�G;��G;�G;�H;�?H;�_H;�yH;Z�H;�H;��H;2�H;r�H;��H;N�H;t�H;��H;��H;��H;h�H;��H;��H;��H;q�H;M�H;��H;u�H;0�H;��H; �H;\�H;�yH;�_H;�?H;�H;�G;��G;.�G;!$G;�F;�[E;�tC;E@;(<;�#6;J>.;�f$;�;i�;�&�:���:���:��:�@�:���:      @V�yƹ�1p� *�6 Y�9�t,:c��:Kٶ:�L�:D�;�;�(&;A.1;�N9;��>;��B;nE;�cF;�G;.�G;ÿG;��G;X H;�EH;�eH;�H;��H;ѥH;��H;��H;�H;��H;��H;T�H;��H;H�H;��H;H�H;��H;Q�H;��H;��H;�H;��H;��H;ѥH;��H;�H;�eH;�EH;V H;��G;��G;.�G;�G;�cF;lE;��B;��>;�N9;>.1;�(&;�;A�;�L�:Oٶ:e��:�t,:Y�9 &�6�1p��xƹ      ��4��K/�RV�B,�G�˺�쀺xuƹpm9 oQ:т�:���:��;��;C�,;*7;��=;!QB;��D;�cF;$G;ЇG;��G;��G;z)H;�NH;�mH;؆H;ĚH;)�H;�H;�H;��H;��H;��H;��H;v�H;�H;w�H;��H;��H;��H;��H;�H;�H;(�H;ĚH;܆H;�mH;�NH;x)H;��G;��G;̇G;$G;�cF;��D;QB;��=;)7;>�,;|�;��;���:т�:oQ:Pm9xuƹ�쀺P�˺H,�ZV��K/�      F�ͻ1Sɻδ��\Ϩ��-���\c��$���˺�P(� O@9z�k:d��:x;6�;"�);��5;P�=;'QB;lE;�F;,8G;G�G;G�G;�	H;\5H;�YH;AwH;ՎH;��H;ѰH;��H;��H;T�H;$�H;��H;u�H;!�H;u�H;~�H;!�H;Q�H;��H;��H;԰H;��H;ՎH;BwH;�YH;W5H;�	H;G�G;D�G;"8G;�F;kE;#QB;L�=;��5; �);5�;v;^��:v�k: O@9�P(���˺�$��\c��-��_Ϩ�Ҵ��.Sɻ      �J;���7��9.����&����^���M����4���º�tƹLQ:���:���:(�;��(;��5;��=;��B;�[E;K�F;�TG;��G;��G;�H;�CH;fH;ɁH;y�H;��H;��H;��H;��H;V�H;��H;<�H;�H;<�H;��H;R�H;��H;��H;��H;��H;x�H;ɁH;fH;�CH;�H;��G;��G;�TG;@�F;�[E;��B;��=;��5;��(;$�;���:���:8Q:�tƹ��º��4�M��b�����軪&����9.���7�      �䙼)`��i��ey��n;k��I�H�$��� �����r�|�8�p$T�h[�9�A�:t��:&�;�);*7;��>;�tC;�E;��F;�uG;�G;��G;�+H;�SH;�sH;��H;b�H;�H;̻H;��H;9�H;o�H;��H;��H;��H;k�H;6�H;��H;ȻH;�H;b�H;��H;�sH;�SH;�+H;��G;�G;�uG;��F;�E;�tC;��>;$7;�);"�;l��:�A�:P[�9x$T�;�v�|������� �I�$��I�r;k�gy��h��)`��      ������߼Nμ "���
��gy��`T�C�!���軸ۙ�hK/�����@m9�A�:���:6�;A�,;�N9;C@;�^D;�LF;Z.G;�G;��G;�H;�?H;dH;�H;q�H;	�H;��H;��H;��H;��H;��H;w�H;��H;��H;��H;��H;��H;�H;u�H;�H;dH;�?H;�H;��G;�G;^.G;�LF;�^D;F@;�N9;@�,;3�;���:�A�:m9����hK/��ۙ����C�!�`T�gy���
��""��Nμ�߼���      ��/�E-�e.%����	�����ލǼѫ��u�{��J;��C�6Ϩ�CO:������[�9���:t;��;>.1;(<;�5B;�NE;�F;4fG;�G;.�G;�*H;�SH;�tH;"�H;��H; �H;M�H;|�H;��H; �H;�H; �H;��H;w�H;I�H;�H;��H;%�H;�tH;�SH;�*H;,�G;�G;1fG;�F;�NE;�5B;(<;;.1;}�;t;���:�[�9����FO:�7Ϩ��C��J;�u�{�ѫ��ލǼ��������f.%�E-�      \@{�W`w�zl��yZ�Q�C�dg*������� "��XO���I�<|�7Ϩ�gK/�`$T�LQ:`��:��;�(&;�#6;�%?;��C;y#F;�#G;$�G;��G;�H;)CH;�gH;~�H;\�H;j�H;�H;��H;�H;�H;��H;��H;�H;��H;�H;h�H;Y�H;��H;�gH;(CH;�H;��G;�G;�#G;y#F;��C;�%?;�#6;�(&;��;\��:4Q:d$T�jK/�7Ϩ�<|��I�XO�� "����鼮��cg*�R�C��yZ�zl�V`w�      �b��㪫��ƣ��s���ɇ�zl�BG��"�h� �-aļa���I��C��ۙ�;�uƹ^�k:���:�;D>.;
;;��A;�AE;_�F;mG;��G;��G;Y2H;�ZH;�zH;ْH;��H;��H;[�H;*�H;��H;�H;��H;*�H;Z�H;��H;��H;֒H;�zH;�ZH;X2H;��G;��G;mG;_�F;�AE;��A;
;;F>.;�;���:b�k: uƹ>��ۙ��C��I�a��-aļh� ��"�BG�zl��ɇ��s���ƣ�㪫�      ������oݽ�2̽�ж����������yZ�F-�շ�,aļXO���J;����t�|���º�N@9ł�:@�;�f$;��5;�N?;;D;�LF;�:G;��G;��G;�!H;�MH;�pH;��H;ϟH;0�H;�H;?�H;s�H;��H;s�H;?�H;�H;,�H;͟H;��H;�pH;�MH;�!H;��G;��G;�:G;�LF;?D;�N?;��5;�f$;=�;���:�N@9��ºu�|���軿J;�XO��-aļշ�F-��yZ����������ж��2̽oݽ���      P,�����Z�:��z�RvϽ�b��-I��f]a�F-�g� � "��u�{�D�!�������4��P(��nQ:�L�:�;ڊ/;�'<;ߟB;��E;��F;��G;��G;5H;?AH;gH;P�H;5�H;ѪH;��H;~�H;��H;S�H;��H;�H;��H;̪H;3�H;O�H;gH;@AH;5H;��G;��G;��F; �E;��B;�'<;ӊ/;�;�L�:�nQ:�P(���4�����D�!�v�{� "��h� �F-�f]a�-I���b��RvϽ�z�:��Z����      %G�p�C��$:��J+������oݽ]���-I���yZ��"����ҫ��bT��� �M����˺�m9Aٶ:i�;`(;�8;i�@;��D;�F;AhG;�G;�H;/5H;�]H;f}H;�H;��H;V�H;ƻH;��H;5�H;��H;ɻH;U�H;��H;�H;e}H;�]H;15H;�H;�G;BhG;߱F;��D;g�@;�8;`(;l�;;ٶ:�m9��˺M���� �bT�ҫ������"��yZ�-I��]���oݽ������J+��$:�p�C�      {x�9t���g���T��G=�z#�6�oݽ�b������AG����ލǼgy��I�$�c����$��uƹS��:�&�:�� ;O4;v�>;OD;�[F;�FG;~�G;�G;�)H;_UH;�vH;��H;�H;��H;i�H;��H;*�H;��H;l�H;��H;�H;��H;�vH;eUH;*H;�G;��G;�FG;�[F;RD;w�>;L4;�� ;�&�:M��:�uƹ�$�d���I�$�gy��ލǼ���AG������b��nݽ6�z#��G=���T���g�9t�      뫖���La��!���>�c�p�C�z#���RvϽ����zl�dg*����
���I���軺\c�퀺�t,:���:��;�_0;h�<;�1C;��E;t#G;S�G;�G; H;�MH;;qH;��H;|�H;ޭH;,�H;��H;_�H;��H;,�H;ܭH;{�H;��H;6qH;�MH; H;�G;S�G;|#G;��E;�1C;f�<;�_0;�;���:�t,:퀺�\c�����I��
�����dg*�zl�����RvϽ��z#�p�C�>�c�!���La����      j*��g����Ƥ�쫖��/��>�c��G=�����zｐж��ɇ�Q�C�
��""��p;k��&��-��q�˺8Y�9|��:9;�h,;�	;;�PB;g�E;� G;܌G;��G;hH;GH;OlH;��H;��H;��H;8�H;�H;ּH;�H;;�H;��H;��H;��H;LlH;GH;jH;��G;�G;� G;e�E;�PB;�	;;�h,;9;���:0Y�9h�˺�-���&�p;k�""��
��Q�C��ɇ��ж��z�����G=�>�c��/��쫖��Ƥ�g���      ��ɾ{�ž+��qת�쫖�!�����T��J+�:��2̽�s���yZ����Mμfy����[Ϩ�N,� "�6��: �
;^�(;VN9;�A;NE;/�F;�G;��G;|H;�AH;3hH;�H;?�H;ԩH;ͳH;��H;y�H;��H;ͳH;ҩH;?�H;�H;0hH;�AH;|H;��G;�G;9�F;~NE;�A;RN9;\�(;��
;��: �6J,�ZϨ���ey��Mμ����yZ��s���2̽:��J+���T�!���쫖�qת�+��|�ž      U_ݾ�:پ�V;+���Ƥ�La����g��$:��Z�oݽ�ƣ�zl�e.%��߼g���9.�ɴ��KV�P1p��@�:x;L(&;4�7;:�@;�
E;��F;juG;$�G;OH;�=H;NeH;ĂH;s�H;L�H;��H;��H;��H;��H;��H;L�H;r�H;ÂH;IeH;�=H;OH;'�G;luG;��F;�
E;9�@;.�7;L(&;x;�@�:�1p�JV�ʴ���9.�g���߼e.%�zl��ƣ�oݽ�Z��$:���g�La���Ƥ�+���V;�:پ      ^�3���:پ{�žg�����9t�p�C�������㪫�W`w�F-����)`����7�4Sɻ�K/��xƹ���:�/;�f$;�7;�~@;K�D;Z�F;�nG;��G;"H;�;H;jcH;o�H;��H;q�H;	�H;-�H;$�H;*�H;	�H;q�H;��H;o�H;dcH;�;H;#H;��G;�nG;g�F;J�D;�~@;�7;�f$;�/;���:�xƹ�K/�5Sɻ��7�)`�����F-�W`w�㪫�������p�C�9t���g���{�ž�:پ4��      GF�Wh����UVھ7�������~���S��#��o��7S��p₽1�6�n���hy��VFB��Eֻ�A?�о	�nY�:���:g�";h46;^@;_�D;��F;�nG;��G;�H;@H;�fH;?�H;,�H;��H;ϳH;ιH;��H;˹H;ҳH;��H;.�H;A�H;�fH;@H;�H;��G;�nG;��F;_�D;Y@;_46;g�";���:rY�:Ծ	��A?��EֻUFB�gy��n���1�6�p₽7S���o���#��S��~������7��UVھ��Wh��      Vh���b���쾧*־�v��(���*��'�O�U� �s��r���؀�F�3���>ݜ�<�>�Q�ѻޡ9�����#o�:<% ;rM#;B�6;NA@;��D;��F;qG;J�G;H;�@H;ggH;��H;��H;ܩH;�H;��H;޻H;��H;�H;ܩH;��H;��H;cgH;�@H;H;M�G;qG;��F;��D;JA@;<�6;nM#;<% ;)o�:����ܡ9�P�ѻ<�>�>ݜ���F�3��؀��r��s�U� �'�O�*��)����v���*־���b��      ���쾳�޾/5ʾL;���:��(�v��E�_'����q����u���+��W��A����4���Ļ9)�pj��{W�:`�;	%;�k7;$�@;��D;��F;�wG;T�G;1H;;CH;(iH;�H;��H;��H;��H;��H;p�H;��H;��H;��H;��H;�H;#iH;DCH;4H;W�G;�wG;��F;��D; �@;�k7;%;`�;�W�:�j��9)���Ļ��4��A���W缃�+���u�p�����_'��E�(�v��:��L;��/5ʾ��޾��      UVھ�*־/5ʾr��������M���9b��5�����ս����Xc���ʖռ�I��U�$�kT���Z��\���:�;k�';�8;RA;�9E;��F;łG;��G;@H;	GH;lH;B�H;9�H;�H;��H;��H;N�H;��H;ĵH;�H;8�H;A�H;lH;GH;CH;��G;łG;��F;�9E;RA;�8;h�';��;�:�\���Z�jT��U�$��I��ʖռ���Xc������ս���5��9b��M������r���/5ʾ�*־      7���v��L;������RP��D�r�z�H�U� ���5@��ѓ����K�a��վ���s�q���񕻝ܺ�4u9&�:!�;-�+;~�:;�"B;m�E;��F;ԐG;��G;-H;4LH;�oH;:�H;t�H;��H;3�H;׼H;��H;ӼH;7�H;��H;q�H;9�H;�oH;<LH;.H;��G;ՐG;��F;n�E;�"B;z�:;,�+; �;&�:�4u9�ܺ��r����s��վ�`���K�ѓ��5@����U� �z�H�D�r�SP������L;���v��      ����)����:���M��D�r�&�O�#,�X�
��gٽpĥ���u�v1�h���)Ϥ���P�[�.o�pp��<:c��:�P;=�/;:�<;C;�E;m!G;5�G;��G;�%H;�RH;�tH;��H;F�H;֯H;�H;Y�H;�H;U�H;�H;ԯH;C�H;�H;�tH;�RH;�%H;�G;5�G;t!G;�E;C;6�<;;�/;�P;m��:@:lp���.o�[򻨎P�)Ϥ�g���v1���u�pĥ��gٽX�
�#,�&�O�D�r��M���:��)���      �~��*��(�v��9b�z�H�#,�MZ����6S��x^����N������μ�I���%+����ܝ.�x����j~:G��:,m;��3;�>;=�C;;PF;~FG;Q�G;��G;u/H;�YH;tzH;D�H;��H;\�H;�H;)�H;��H;&�H;�H;]�H;��H;B�H;rzH;ZH;{/H;��G;P�G;�FG;>PF;;�C;�>;��3;+m;U��:�j~:����؝.�����%+��I����μ�����N�x^��6S�����MZ�#,�z�H��9b�(�v�*��      �S�'�O��E��5�U� �X�
���罤9��(l���Xc���(��������[�����ݎ�Cܺp;9$��:/�	;Ed';d 8;<�@;�D;�F;jG;��G;NH;n:H;?bH;��H;�H;1�H;@�H;{�H;6�H;��H;5�H;~�H;B�H;/�H; �H;��H;HbH;r:H;PH;��G;jG;�F;z�D;>�@;e 8;Cd';6�	;&��:�;9?ܺ�ݎ������[��������(��Xc�'l���9�����X�
�U� ��5��E�'�O�      �#�U� �`'������gٽ6S��'l��O�j�B�3��i��վ�y���(���Ļ^A?���B��@:�[�:
Q;�.;��;;~tB;�E;�F;%�G;��G;�H;QFH;"kH;��H;�H;�H;e�H;�H;r�H;��H;o�H;
�H;h�H;�H;�H;��H;*kH;VFH;�H;��G;(�G;��F;�E;tB;��;;�.;Q;�[�: �@:��B�\A?���Ļ(�y����վ��i�B�3�N�j�'l��6S���gٽ����_'�U� �      �o��s��罫�ս4@��pĥ�x^���Xc�B�3���	�Ɍ˼�]��RFB��Z򻬜��jӺ ��8��:ܛ;�M#;u=5;?;L�C;|@F;:G;�G;�G;0'H;�RH;ytH;��H;{�H;+�H;��H;��H;��H;?�H;��H;��H;��H;(�H;x�H;��H;�tH;�RH;2'H;�G;�G;
:G;{@F;P�C;?;t=5;�M#;ޛ;��:���8hӺ�����Z�QFB��]��Ɍ˼��	�B�3��Xc�x^��pĥ�5@����ս���s�      7S���r��r�����Г����u���N���(��i�Ɍ˼�A����P�fs��8|�8����\:4�:p�;xn-;�:;��A;|,E;j�F;,oG;��G;�H;�7H;:_H;	~H;�H;�H;s�H;�H;w�H;9�H;�H;;�H;x�H;�H;s�H; �H;�H;~H;@_H;�7H;�H;��G;/oG;h�F;�,E;��A;�:;�n-;u�;4�:�\:0���6|��fs���P��A��Ɍ˼�i���(���N���u�ѓ�����r���r��      o₽�؀���u��Xc���K�v1�������վ��]����P����@T����9���o��3�9x&�:`�	;\%;F�5;��>;��C;�F;�!G;��G;��G;EH;`HH;�kH;��H;I�H;��H;��H;t�H;I�H;��H;��H;��H;I�H;x�H;��H;��H;M�H;��H;�kH;bHH;EH;��G;��G;�!G;�F;��C;��>;Q�5;_%;^�	;�&�:�3�9��o���9�>T�������P��]���վ�ߤ���v1���K��Xc���u��؀�      2�6�E�3���+���`�h�����μ���y���QFB�es�@T��)�D��{���:u9�q�:}��:�Y;�t0;��;;�B;�9E;�F;hG;ٿG;�G;z0H;�XH;'xH;�H;u�H;�H;��H;��H;�H;.�H;2�H;.�H;�H;��H;��H;��H;z�H;(�H;.xH;�XH;|0H;��G;޿G;hG;�F;�9E;�B;��;;�t0;|Y;���:�q�:�:u9�{��'�D�=T��es�QFB�x��������μh���a�����+�E�3�      k�����W�˖ռ�վ�*Ϥ��I����[�(��Z����9��{���;9SX�:ZX�:;Q;B,;��8;�A@;BD;�@F;�,G;��G;��G;gH;�DH;hH;,�H;Q�H;d�H;]�H;"�H;�H;��H;��H;c�H;��H;��H;�H; �H;[�H;j�H;\�H;5�H; hH;�DH;bH;��G;��G;�,G;�@F;BD;�A@;��8;>,;DQ;\X�:]X�:�;9�{����9���Z�(���[��I��)Ϥ��վ�˖ռ�W���      fy��>ݜ��A���I����s���P��%+������Ļ����4|��o��:u9WX�:�+�:X;�);Մ6;w�>;�PC;d�E;��F;�xG;+�G;zH;e1H;XH;�vH;��H;�H;��H;}�H;�H;?�H;��H;��H;��H;��H;��H;B�H;�H;z�H;�H;�H;��H;wH;XH;a1H;~H;,�G;�xG;��F;h�E;�PC;z�>;Є6;�);X;�+�:]X�:�:u9 �o�2|�������Ļ����%+���P���s��I���A��>ݜ�      OFB�:�>���4�S�$�q��
[�����ݎ�aA?�cӺ(����3�9�q�:\X�:X;��';�=5;��=;�B;GE;K�F;�UG;!�G;��G;SH;�HH;jH;��H;t�H;G�H;.�H;G�H;��H;>�H;�H; �H;��H;�H;�H;>�H;��H;D�H;5�H;L�H;{�H;��H;jH;�HH;YH;��G;$�G;�UG;O�F;!GE;�B;|�=;�=5;��';\;\X�:�q�:�3�9 ���`ӺZA?��ݎ����[�t��T�$���4�7�>�      �EֻM�ѻ��ĻlT���񕻶.o�ԝ.�;ܺ��B�@��8�\:z&�:���:AQ;�);�=5;�:=;,#B;��D;�uF;�6G;ĚG;\�G;uH;�:H;^H;�zH;��H;^�H;ĲH;�H;��H;\�H;�H;m�H;2�H;��H;-�H;j�H;�H;X�H;��H;�H;ǲH;e�H;��H;�zH;^H;�:H;uH;]�G;ǚG;�6G;�uF;��D;%#B;�:=;�=5;�);BQ;���:�&�:�\:@��8x�B�5ܺ؝.��.o���pT����ĻH�ѻ      oA?�ס9� 9)��Z��ܺjp��8����;9�@:��::�:Y�	;yY;<,;΄6;x�=;!#B;��D;aXF;�!G;|�G;�G;�H;�.H;xSH;bqH;މH;��H;b�H;��H;o�H;��H;��H;��H;��H;�H;��H;�H;�H;��H;��H;��H;t�H;ùH;f�H;��H;߉H;^qH;}SH;�.H;�H;!�G;��G;�!G;dXF;��D;$#B;u�=;ф6;<,;yY;\�	;F�:��: �@: <9X���dp��{ܺ�Z�9)�ԡ9�      l�	����xj���[���4u9t:�j~:0��:�[�:ߛ;z�;\%;�t0;��8;{�>;	�B;��D;jXF;7G;a�G;��G;��G;�%H;KH;�iH;�H;��H;8�H;v�H;�H;[�H;��H;��H;3�H;�H;��H;S�H;��H;~�H;2�H;��H;��H;^�H;�H;v�H;8�H;��H;�H;�iH;	KH;�%H;��G;��G;e�G;:G;dXF;��D;�B;~�>;��8;�t0;_%;}�;��;�[�:4��:�j~:`:5u9 ]��xj�����      dY�:#o�:�W�:1�:
&�:m��:i��:/�	;Q;�M#;�n-;O�5;��;;�A@;�PC;!GE;�uF;�!G;c�G;��G;�G;H H;EH;�cH;8}H;t�H;��H;��H;��H;��H;��H;,�H;T�H;S�H;N�H;z�H;��H;u�H;K�H;Q�H;R�H;)�H;��H;��H;��H;��H;��H;r�H;=}H;�cH;EH;J H;�G;��G;h�G;�!G;�uF;GE;�PC;�A@;��;;Q�5;�n-;�M#;Q;9�	;c��:{��:&�:�:wW�:o�:      ���:0% ;F�;��;�;�P;,m;@d';�.;w=5;�:;��>;�B;BD;f�E;O�F;�6G;��G;��G;�G;wH;�AH;`H;LyH;{�H;"�H;Q�H;�H;K�H;��H;��H;1�H;��H;@�H;��H;��H;D�H;��H;��H;A�H;��H;+�H;��H;��H;K�H;�H;N�H;�H;�H;LyH;`H;�AH;zH;�G;��G;��G;�6G;M�F;h�E;BD;�B;��>;�:;u=5; �.;>d';3m;�P;"�;��;R�;.% ;      `�";xM#;%;v�';,�+;=�/;��3;a 8;��;;?;��A;��C;�9E;�@F;��F;�UG;ŚG;$�G;��G;J H;�AH;�^H;HwH;�H;��H;�H;��H;.�H;��H;%�H;�H;��H;��H;��H;n�H;L�H;y�H;G�H;m�H;��H;��H;��H;�H;&�H;��H;-�H;��H;ޫH;��H;�H;BwH;�^H;�AH;L H;��G;!�G;ǚG;�UG;��F;�@F;�9E;��C;�A;?;��;;i 8;��3;7�/;?�+;k�';%;nM#;      }46;B�6;�k7;*�8;x�:;@�<;,�>;H�@;�tB;S�C;�,E;�F;�F;�,G;�xG;'�G;`�G;�H;�%H;EH;`H;GwH;2�H;5�H;G�H;�H;��H;n�H;��H;��H;(�H;?�H;��H;]�H;��H;o�H;��H;i�H;��H;_�H;��H;<�H;*�H;��H;��H;n�H;��H;�H;K�H;4�H;-�H;HwH;`H;EH;�%H;�H;b�G;$�G;�xG;�,G;�F;�F;�,E;O�C;�tB;J�@;(�>;>�<;��:;)�8;�k7;&�6;      _@;VA@;�@;RA;�"B;C;?�C;|�D;�E;@F;n�F;�!G;hG;��G;,�G;��G;vH;�.H;KH;�cH;JyH;�H;3�H;ĩH;�H;~�H;x�H;��H;�H;N�H;��H;J�H;:�H;��H;��H;^�H;��H;X�H;��H;��H;7�H;H�H;��H;M�H;�H;��H;r�H;�H;�H;��H;0�H;�H;JyH;�cH;KH;�.H;vH;��G;-�G;��G;�gG;�!G;q�F;@F;�E;��D;?�C;�
C;�"B;RA;�@;OA@;      ��D;��D;��D;�9E;h�E;'�E;FPF;�F;��F;:G;6oG;��G;ݿG;��G;~H;]H;�:H;�SH;�iH;B}H;��H;��H;K�H;�H;=�H;��H;-�H;m�H;��H;*�H;��H;	�H;��H;��H;��H;%�H;c�H;�H;��H;��H;��H;�H;��H;+�H;��H;m�H;&�H;��H;@�H;�H;K�H;��H;��H;@}H;�iH;�SH;�:H;\H;H;��G;޿G;��G;9oG;:G;��F;�F;HPF;!�E;r�E;�9E;��D;��D;      ��F;��F;��F;��F;��F;t!G;�FG;#jG;)�G;�G;��G;��G;�G;oH;e1H;�HH;^H;fqH;�H;q�H; �H;ګH;�H;~�H;��H;
�H;�H;[�H;��H;��H;��H;��H;��H;��H;x�H;��H;�H;��H;u�H;��H;��H;}�H;��H;��H;��H;Z�H;�H;�H;��H;{�H;�H;ݫH; �H;q�H;�H;aqH;^H;�HH;e1H;iH;�G;��G;��G;�G;,�G;'jG;�FG;j!G;��F;��F;��F;��F;      �nG;qG;�wG;ƂG;̐G;1�G;^�G;��G;��G;"�G;�H;AH;w0H;�DH;XH;jH;�zH;�H;��H;��H;V�H;��H;��H;{�H;,�H;�H;=�H;��H;]�H;{�H;I�H;��H;��H;��H;4�H;��H;��H;��H;2�H;��H;��H;��H;I�H;{�H;Z�H;��H;8�H;�H;.�H;u�H;��H;��H;V�H;��H;��H;މH;�zH;jH;XH;�DH;w0H;EH;�H;�G;��G;��G;W�G;.�G;�G;��G;�wG;qG;      ��G;H�G;P�G;��G;��G;��G;��G;LH;�H;7'H;�7H;gHH;�XH;#hH; wH;��H;��H;��H;:�H;��H;�H;*�H;k�H;��H;l�H;Z�H;��H;;�H;w�H;>�H;��H;��H;��H;a�H;��H; �H;�H;��H;��H;c�H;��H;��H;��H;A�H;v�H;9�H;��H;[�H;o�H;��H;m�H;+�H;�H;��H;8�H;��H;��H;��H;wH; hH;�XH;gHH;�7H;6'H;�H;NH;��G;��G;��G;��G;N�G;?�G;      �H;H;1H;OH;H;�%H;|/H;j:H;KFH;�RH;@_H;�kH;-xH;1�H;��H;z�H;e�H;l�H;{�H;¼H;N�H;��H;��H;�H;��H;��H;Y�H;w�H;!�H;��H;��H;��H;U�H;��H;C�H;u�H;��H;p�H;C�H;��H;V�H;��H;��H;��H;"�H;v�H;S�H;��H;��H;	�H;��H;��H;K�H;��H;x�H;h�H;g�H;z�H;��H;1�H;*xH;�kH;B_H;�RH;OFH;m:H;|/H;�%H;+H;KH;/H;H;      @H;�@H;ICH;	GH;?LH;�RH;ZH;=bH;&kH;~tH;~H;��H;&�H;\�H;�H;I�H;ʲH;��H;�H;��H;��H;"�H;��H;J�H;*�H;��H;z�H;A�H;��H;��H;��H;g�H;��H;M�H;��H;��H;��H;��H;��H;M�H;��H;d�H;��H;��H;��H;>�H;t�H;��H;-�H;G�H;��H;#�H;��H;��H;�H;��H;ȲH;K�H;�H;Y�H;(�H;��H;~H;�tH;(kH;FbH;ZH;�RH;>LH;	GH;KCH;�@H;      �fH;ygH;.iH;lH;�oH;�tH;~zH;��H;��H;��H;�H;S�H;}�H;o�H;�H;8�H;�H;x�H;b�H;��H;��H;�H;(�H;��H;��H;��H;K�H;��H;��H;��H;g�H;�H;^�H;��H;��H;�H;'�H;�H;��H;��H;`�H;�H;g�H;��H;��H;��H;H�H;��H;��H;��H;,�H;�H;��H;��H;a�H;u�H;�H;8�H;�H;n�H;��H;T�H;�H;��H;��H;��H;�zH;�tH;pH;lH;/iH;|gH;      C�H;��H;�H;>�H;:�H;�H;N�H;�H;$�H;~�H;�H;��H;�H;g�H;~�H;M�H;��H;��H;��H;/�H;8�H;��H;?�H;H�H;	�H;�H;��H;��H;��H;h�H;��H;u�H;��H;��H;&�H;@�H;@�H;@�H;#�H;��H;��H;o�H;��H;j�H;��H;��H;��H;��H;�H;B�H;A�H;��H;2�H;,�H;��H;��H;��H;N�H;��H;e�H;�H;��H;
�H;|�H;#�H;�H;S�H;�H;E�H;>�H;�H;��H;      0�H;��H;��H;;�H;}�H;C�H;��H;.�H;�H;/�H;z�H;��H;��H;)�H;�H;��H;a�H;��H;��H;Y�H;��H;��H;��H;6�H;��H;��H;��H;��H;Z�H;��H;[�H;��H;�H;5�H;T�H;w�H;}�H;w�H;Q�H;6�H;�H;��H;Z�H;��H;W�H;��H;��H;��H;��H;6�H;��H;��H;��H;U�H;��H;��H;b�H;��H;�H;)�H;�H;��H;{�H;1�H;�H;/�H;��H;=�H;��H;5�H;��H;��H;      ��H;٩H;��H;ګH;��H;̯H;g�H;F�H;n�H;��H;�H;��H;��H;'�H;H�H;G�H;!�H;��H;7�H;W�H;G�H;��H;[�H;��H;��H;��H;��H;c�H;��H;P�H;��H;��H;2�H;p�H;�H;��H;��H;��H;~�H;q�H;5�H;��H;��H;M�H;��H;`�H;��H;��H;��H;��H;`�H;��H;@�H;Q�H;6�H;��H;'�H;H�H;H�H;'�H;��H;~�H;�H;��H;r�H;L�H;k�H;̯H;��H;٫H;��H;�H;      ̳H;%�H;ôH;ǵH;E�H;��H;*�H;~�H;�H;��H;��H;V�H;�H;��H;��H;�H;q�H;��H;�H;O�H;��H;k�H;��H;��H;��H;p�H;/�H;��H;E�H;��H;��H;'�H;T�H;��H;��H;��H;��H;��H;��H;��H;U�H;'�H;��H;��H;?�H;��H;/�H;r�H;��H;��H;��H;i�H;��H;I�H;~�H;��H;v�H;�H;��H;��H;�H;W�H;��H;��H;�H;��H;,�H;��H;E�H;ɵH;ƴH;&�H;      ͹H;��H;��H;��H;׼H;Q�H;8�H;:�H;u�H;��H;F�H;��H;5�H;��H;��H;!�H;2�H;�H;��H;z�H;��H;H�H;h�H;Q�H;!�H;��H;��H;�H;y�H;��H;�H;D�H;}�H;��H;��H;��H;��H;��H;��H;��H;�H;D�H;�H;��H;u�H;��H;��H;��H; �H;Q�H;n�H;G�H;��H;u�H;��H; �H;6�H;#�H;��H;��H;3�H;��H;G�H;��H;y�H;?�H;<�H;R�H;ڼH;��H;��H;�H;      ȻH;ۻH;��H;P�H;�H;�H;��H;��H;��H;H�H;��H;��H;A�H;q�H;��H;��H;��H;��H;W�H;��H;O�H;��H;��H;��H;d�H;�H;��H;�H;��H;��H;$�H;D�H;��H;��H;��H;��H;��H;��H;��H;��H;��H;D�H;$�H;��H;��H;�H;��H;�H;d�H;��H;��H;�H;H�H;��H;W�H;��H;��H;��H;��H;s�H;@�H;��H;��H;I�H;�H;��H;��H;�H;��H;N�H;��H;�H;      ͹H;��H;��H;��H;ؼH;U�H;5�H;9�H;u�H;��H;D�H;��H;6�H;��H;��H;!�H;2�H;�H;��H;z�H;��H;I�H;h�H;Q�H;!�H;��H;��H;�H;|�H;��H;�H;G�H;�H;��H;��H;��H;��H;��H;��H;��H;�H;D�H;�H;��H;u�H;��H;��H;��H;�H;P�H;n�H;E�H;��H;u�H;��H;!�H;3�H;#�H;��H;��H;3�H;��H;G�H;��H;y�H;?�H;:�H;R�H;ݼH;��H;��H;�H;      ĳH;)�H;��H;��H;G�H;��H;,�H;��H;�H;��H;��H;V�H;!�H;��H;��H;�H;q�H;��H;�H;O�H;��H;m�H;��H;��H;��H;n�H;0�H;��H;F�H;��H;��H;(�H;T�H;��H;��H;��H;��H;��H;��H;��H;W�H;'�H;��H;��H;?�H;��H;,�H;r�H;��H;��H;��H;j�H;��H;I�H;~�H;��H;t�H;�H;��H;��H;�H;X�H;��H;��H;�H;��H;2�H;��H;H�H;��H;´H;'�H;      ��H;ةH;��H;ݫH;��H;ЯH;d�H;J�H;o�H;��H;�H;�H;��H;'�H;J�H;G�H;$�H;��H;7�H;W�H;H�H;��H;[�H;��H;��H;��H;��H;e�H;��H;Q�H;��H;��H;4�H;p�H;�H;��H;��H;��H;~�H;o�H;4�H;��H;��H;L�H;��H;^�H;��H;��H;��H;��H;`�H;��H;>�H;S�H;6�H;��H;$�H;G�H;I�H;&�H;��H;~�H;�H;��H;r�H;M�H;k�H;ͯH;��H;٫H;��H;۩H;      2�H;��H;��H;8�H;x�H;D�H;��H;1�H;�H;1�H;z�H;��H;�H;+�H;�H;��H;a�H;��H;��H;Y�H;��H;��H;��H;6�H;��H;��H;��H;��H;]�H; �H;[�H;��H;�H;5�H;T�H;x�H;}�H;v�H;S�H;4�H;�H;��H;Z�H;��H;S�H;��H;��H;��H;��H;2�H;��H;��H;��H;V�H;��H;��H;_�H;��H;�H;)�H;�H;��H;z�H;.�H;�H;4�H;��H;@�H;|�H;=�H;��H;��H;      3�H;��H;��H;:�H;6�H;��H;P�H;�H;!�H;|�H;�H;��H;�H;g�H;��H;N�H;��H;��H;��H;/�H;9�H;��H;=�H;F�H;�H;�H;��H;��H;��H;h�H;��H;r�H;��H;��H;'�H;?�H;@�H;@�H;$�H;��H;��H;p�H;��H;e�H;��H;��H;��H;��H;�H;>�H;D�H;��H;/�H;,�H;��H;��H;��H;M�H;�H;e�H;	�H;��H;�H;~�H;&�H;
�H;S�H;�H;:�H;;�H;�H;��H;      �fH;xgH;/iH;lH;�oH;�tH;|zH;��H;��H;��H;��H;U�H;~�H;o�H;�H;8�H;�H;x�H;b�H;��H;��H;"�H;(�H;��H;��H;��H;H�H;��H;��H;��H;g�H;�H;^�H;��H;��H;�H;'�H;�H;��H;��H;`�H;�H;e�H;��H;��H;��H;E�H;��H;��H;��H;-�H;�H;��H;��H;a�H;t�H;�H;7�H;�H;n�H;}�H;U�H;�H;��H;��H;��H;�zH;�tH;pH;lH;6iH;ygH;      @H;�@H;BCH;GH;3LH;�RH;ZH;HbH;,kH;�tH;~H;��H;*�H;]�H;�H;I�H;ʲH;��H;�H;��H;��H;%�H;��H;H�H;+�H;��H;w�H;A�H;��H;��H;��H;g�H;��H;M�H;��H;��H;��H;��H;��H;M�H;��H;e�H;��H;��H;��H;;�H;s�H;��H;(�H;D�H;��H;#�H;��H;��H;�H;��H;ȲH;H�H;�H;[�H;'�H;��H;~H;�tH;(kH;GbH;ZH;�RH;>LH;GH;SCH;�@H;      H;H;CH;JH;H;�%H;{/H;n:H;VFH;�RH;A_H;�kH;.xH;4�H;��H;|�H;e�H;m�H;z�H;¼H;P�H;��H;��H;�H;��H;��H;U�H;w�H;#�H;��H;��H;��H;V�H;��H;C�H;s�H;��H;s�H;C�H;��H;W�H;��H;��H;��H;�H;q�H;R�H;��H;��H;�H;��H;��H;K�H;��H;x�H;e�H;b�H;{�H;��H;1�H;,xH;�kH;B_H;�RH;TFH;p:H;}/H;�%H;&H;FH;BH;�H;      ��G;>�G;B�G;��G;��G;�G;��G;PH;�H;9'H;�7H;gHH;�XH;%hH;wH;��H;��H;��H;8�H;��H;�H;.�H;j�H;��H;o�H;T�H;��H;9�H;z�H;>�H;��H;��H;��H;a�H;��H;��H;�H;��H;��H;c�H;��H;��H;��H;>�H;t�H;4�H;��H;X�H;l�H;��H;o�H;+�H;޹H;��H;8�H;��H;��H;��H;wH; hH;�XH;dHH;�7H;4'H;�H;LH;��G;��G;��G;��G;P�G;>�G;      �nG;"qG;�wG;ЂG;ؐG;9�G;\�G;��G;��G;�G;�H;EH;w0H;�DH;XH;jH;�zH;�H;��H;��H;Y�H;��H;��H;~�H;-�H;�H;9�H;��H;^�H;z�H;H�H;��H;��H;��H;4�H;��H;��H;��H;2�H;��H;��H;��H;K�H;z�H;Y�H;��H;9�H;�H;-�H;w�H;��H;��H;T�H;��H;��H;މH;�zH;jH;XH;�DH;v0H;DH;�H;�G;��G;��G;a�G;5�G;ߐG;͂G;�wG;qG;      ��F;��F;��F;��F;��F;|!G;�FG;'jG;-�G;�G;��G;��G;�G;lH;f1H;�HH;^H;fqH;�H;q�H;%�H;ݫH;�H;~�H;��H;�H;�H;Z�H;��H;��H;��H;��H;��H;��H;x�H;��H;
�H;��H;u�H;��H;��H;��H;��H;��H;��H;X�H;�H;�H;��H;{�H;�H;ګH; �H;p�H;�H;_qH;^H;�HH;i1H;iH;�G;��G;��G;��G;&�G;"jG;�FG;m!G;��F;��F;��F;�F;      �D;��D;��D;�9E;h�E;,�E;FPF;�F;��F;:G;7oG;��G;ݿG;��G;�H;^H;�:H;�SH;�iH;@}H;��H;��H;J�H;�H;A�H;��H;)�H;m�H;��H;'�H;��H;	�H;��H;��H;��H;"�H;c�H;"�H;��H;��H;��H;�H;��H;(�H;��H;i�H;*�H;��H;=�H;�H;N�H;��H;��H;B}H;�iH;�SH;�:H;\H;�H;��G;ݿG;��G;4oG;:G;��F;�F;HPF; �E;o�E;�9E;��D;��D;      @@;>A@;�@;"RA;�"B;C;A�C;��D;!�E;~@F;q�F;�!G;�gG;��G;/�G;��G;vH;�.H;KH;�cH;MyH;�H;1�H;ƩH;�H;z�H;u�H;��H;�H;J�H;��H;L�H;9�H;��H;��H;\�H;��H;^�H;��H;��H;<�H;J�H;��H;K�H;�H;��H;w�H;~�H;�H;ƩH;1�H;�H;IyH;�cH;KH;�.H;uH;��G;-�G;��G;�gG;�!G;q�F;|@F;�E;z�D;>�C; C;�"B;1RA;�@;(A@;      p46;>�6;�k7;4�8;v�:;;�<;%�>;F�@;�tB;R�C;�,E;�F;�F;�,G;�xG;(�G;`�G;�H;�%H;EH;
`H;HwH;/�H;8�H;M�H;�H;��H;n�H;��H;��H;*�H;C�H;��H;]�H;��H;p�H;��H;n�H;��H;[�H;��H;@�H;-�H;��H;��H;m�H;��H;�H;H�H;4�H;/�H;GwH;`H;EH;�%H;�H;b�G;'�G;�xG;�,G;�F;�F;�,E;R�C;�tB;H�@;$�>;;�<;t�:;/�8;�k7;)�6;      c�";xM#;%;m�';,�+;D�/;��3;e 8;��;;?;�A;��C;�9E;�@F;��F;�UG;ȚG;&�G;��G;L H;�AH;�^H;DwH;�H;��H;۫H;��H;-�H;��H;#�H;�H;��H;��H;��H;k�H;H�H;{�H;H�H;j�H;��H;��H;��H; �H;&�H;��H;*�H;��H;ݫH;��H;�H;EwH;�^H;�AH;L H;��G;!�G;ĚG;�UG;��F;�@F;�9E;��C;��A;?;��;;i 8;��3;/�/;B�+;a�';%;jM#;      ���:F% ;X�;��;�;Q;/m;Ad';�.;t=5;�:;��>;�B;BD;k�E;R�F;�6G;��G;��G;�G;wH;�AH;
`H;NyH;��H;�H;M�H;߹H;K�H;��H;��H;2�H;��H;E�H;��H;��H;F�H;��H;��H;@�H;��H;/�H;��H;��H;H�H;޹H;O�H;�H;|�H;MyH;`H;�AH;uH;�G;��G;��G;�6G;M�F;i�E;BD;�B;��>;�:;u=5;�.;Ed';3m;�P;$�;��;f�;2% ;      �Y�:)o�:�W�:+�:
&�:w��:i��:9�	;Q;�M#;�n-;O�5;��;;�A@;�PC;$GE;�uF;�!G;f�G;��G;�G;L H;EH;�cH;?}H;r�H;��H;��H;üH;��H;��H;+�H;U�H;U�H;N�H;v�H;��H;w�H;K�H;P�H;T�H;+�H;��H;��H;��H;��H;��H;r�H;8}H;�cH;EH;I H;�G;��G;c�G;�!G;�uF;GE;�PC;�A@;��;;O�5;�n-;�M#;Q;2�	;c��:e��:&�:�:�W�:o�:      h�	����pj���[���4u9p:�j~:2��:�[�:ߛ;y�;^%;�t0;��8;�>;	�B;��D;hXF;:G;e�G;��G;��G;�%H;KH;�iH;�H;��H;5�H;w�H;�H;^�H;��H;��H;3�H;��H;��H;S�H;��H;~�H;2�H;��H;��H;^�H;�H;t�H;4�H;��H;�H;�iH;	KH;�%H;��G;��G;c�G;7G;cXF;��D;�B;~�>;��8;�t0;\%;z�;ޛ;�[�:4��:�j~:h:�4u9�[���j������      ~A?�С9�#9)��Z�wܺVp��@���@<9$�@:��:@�:]�	;yY;<,;ӄ6;{�=;$#B;��D;cXF;�!G;��G;#�G;�H;�.H;SH;_qH;ىH;��H;h�H;��H;r�H;��H;��H;��H;��H;�H;��H;�H;}�H;��H;��H;��H;r�H;��H;e�H;��H;މH;^qH;xSH;�.H;�H; �G;|�G;�!G;aXF;��D;!#B;v�=;ӄ6;<,;xY;Z�	;B�:��:�@:<9H���`p���ܺ�Z�-9)�С9�      �EֻN�ѻ��ĻkT���񕻵.o�֝.�6ܺ��B�`��8�\:�&�:���:AQ;�);�=5;�:=;(#B;��D;�uF;�6G;ǚG;`�G;xH;�:H;^H;�zH;��H;e�H;ĲH;	�H;��H;\�H;�H;m�H;0�H;��H;0�H;j�H;�H;W�H;��H;	�H;ŲH;b�H;��H;�zH;^H;�:H;vH;`�G;ĚG;�6G;�uF;��D;%#B;�:=;�=5;�);AQ;���:~&�:�\: ��8|�B�6ܺڝ.��.o���nT����ĻJ�ѻ      PFB�:�>���4�S�$�r��[�����ݎ�_A?�cӺ����3�9�q�:`X�:^;��';�=5;}�=;�B;GE;P�F;�UG;(�G;��G;YH;�HH;jH;��H;{�H;I�H;4�H;J�H;��H;B�H;�H; �H;��H;�H;�H;=�H;��H;D�H;1�H;H�H;x�H;�H;jH;�HH;SH;��G;'�G;�UG;H�F;GE;�B;{�=;�=5;��';\;ZX�:�q�:�3�9 ���dӺ`A?��ݎ����[�t��S�$���4�:�>�      fy��>ݜ��A���I����s���P��%+������Ļ����2|� �o��:u9_X�:�+�:\;�);ӄ6;z�>;�PC;k�E;��F;�xG;/�G;H;f1H;XH;wH;��H;�H;�H;}�H;�H;C�H;��H;��H;��H;��H;��H;A�H;�H;z�H;�H;�H;��H;�vH;XH;b1H;zH;/�G;�xG;��F;b�E;�PC;w�>;΄6;�);V;�+�:WX�:�:u9�o�5|�������Ļ����%+���P���s��I���A��>ݜ�      l�����W�˖ռ�վ�)Ϥ��I����[�(��Z����9��{�� <9aX�:dX�:@Q;<,;��8;�A@;BD;�@F;�,G;��G;��G;hH;�DH;hH;3�H;V�H;j�H;`�H;"�H;�H;��H;��H;c�H;��H;��H;�H;�H;Z�H;e�H;Y�H;4�H;hH;�DH;dH;��G;��G;�,G;�@F;
BD;�A@;��8;<,;@Q;ZX�:WX�:�;9�{����9���Z�(���[��I��)Ϥ��վ�˖ռ�W���      1�6�E�3���+���`�h�����μ���y���PFB�es�>T��&�D��{�� ;u9�q�:���:}Y;�t0;��;;�B;�9E;�F;hG;޿G;�G;y0H;�XH;-xH;$�H;y�H; �H;��H;��H;�H;.�H;2�H;.�H;�H;��H;��H;��H;v�H;'�H;-xH;�XH;w0H;�G;ٿG;hG;�F;�9E;�B;��;;�t0;yY;���:�q�:�:u9�{��*�D�?T��es�QFB�y��������μh���a�����+�E�3�      o₽�؀���u��Xc���K�v1����ߤ��վ��]����P����>T����9���o��3�9~&�:Z�	;^%;M�5;��>;��C;�F;�!G;��G;��G;BH;`HH;�kH;��H;M�H;��H;��H;w�H;I�H;��H;��H;��H;I�H;u�H;��H;��H;J�H;��H;�kH;`HH;AH;��G;��G;�!G;�F;��C;��>;N�5;[%;]�	;~&�:�3�9��o���9�?T�������P��]���վ�ߤ���v1���K��Xc���u��؀�      7S���r��r�����Г����u���N���(��i�Ɍ˼�A����P�fs��5|�0����\:0�:r�;~n-;�:;��A;�,E;m�F;/oG;��G;�H;�7H;>_H;~H;�H;�H;s�H;�H;w�H;<�H;��H;;�H;w�H;�H;p�H; �H;�H;~H;A_H;�7H;�H;��G;)oG;m�F;�,E;��A;ޞ:;n-;p�;.�:�\:@���8|��fs���P��A��Ɍ˼�i���(���N���u�ѓ�����r���r��      �o��s��罫�ս4@��pĥ�x^���Xc�B�3���	�Ȍ˼�]��QFB��Z򻪜��dӺ���8��:ܛ;�M#;x=5;?;P�C;~@F;
:G;�G;�G;2'H;�RH;}tH;��H;x�H;+�H;��H;��H;��H;?�H;��H;��H;��H;(�H;w�H;��H;~tH;�RH;/'H;�G;�G;:G;~@F;P�C;?;p=5;�M#;ٛ;��:���8jӺ�����Z�RFB��]��Ɍ˼��	�B�3��Xc�x^��pĥ�5@����ս���s�      �#�U� �_'������gٽ6S��'l��N�j�B�3��i��վ�y���(���ĻZA?���B���@:�[�:Q;�.;��;;tB;�E;��F;(�G;��G;�H;VFH;&kH;��H;�H;�H;h�H;�H;r�H;��H;p�H;
�H;g�H;�H;�H;��H;(kH;VFH;�H;��G;(�G;��F;�E;tB;��;;�.;Q;�[�: �@:��B�^A?���Ļ(�y����վ��i�B�3�N�j�'l��6S���gٽ����_'�U� �      �S�'�O��E��5�U� �X�
���罤9��(l���Xc���(��������[�����ݎ�?ܺ@;9(��:2�	;Gd';e 8;@�@;��D;�F;jG;��G;LH;p:H;?bH;��H;�H;1�H;C�H;{�H;6�H;��H;6�H;}�H;C�H;-�H; �H;��H;FbH;r:H;NH;��G;jG;�F;�D;>�@;d 8;Cd';6�	;"��:�;9=ܺ�ݎ������[��������(��Xc�'l���9�����X�
�U� ��5��E�'�O�      �~��*��(�v��9b�z�H�#,�MZ����6S��x^����N������μ�I���%+����؝.������j~:O��:/m;��3;�>;=�C;=PF;�FG;N�G;��G;y/H;ZH;uzH;D�H;��H;]�H;�H;)�H;��H;&�H;�H;\�H;��H;B�H;rzH;ZH;{/H;��G;P�G;�FG;;PF;=�C;�>;��3;+m;W��:�j~:����؝.�����%+��I����μ�����N�x^��6S�����MZ�#,�z�H��9b�(�v�*��      ����(����:���M��D�r�'�O�#,�X�
��gٽpĥ���u�v1�g���)Ϥ���P�[�.o�rp��D:i��:�P;=�/;:�<;C;�E;k!G;4�G;�G;�%H;�RH;�tH;��H;D�H;֯H; �H;Y�H;�H;Y�H;�H;֯H;C�H;��H;�tH;�RH;�%H;�G;4�G;t!G;�E;C;9�<;:�/;�P;m��:<:rp���.o�[򻨎P�)Ϥ�h���v1���u�pĥ��gٽX�
�#,�&�O�D�r��M���:��)���      7���v��L;������RP��D�r�z�H�T� ���5@��Г����K�`��վ���s�q���񕻡ܺ�4u9&�:$�;,�+;~�:;�"B;n�E;��F;ӐG;��G;.H;3LH;�oH;9�H;r�H;��H;2�H;ؼH;��H;ӼH;4�H;��H;q�H;:�H;�oH;<LH;1H;��G;אG;��F;m�E;�"B;z�:;,�+;!�;&�:�4u9�ܺ��r����s��վ�a���K�ѓ��5@����U� �z�H�D�r�RP������L;���v��      UVھ�*־/5ʾr��������M���9b��5�����ս����Xc���ʖռ�I��U�$�jT���Z�@\���:�;j�';�8;RA;�9E;��F;��G;��G;@H;GH;lH;B�H;6�H;�H;��H;��H;Q�H;��H;õH;ޫH;9�H;B�H;lH;GH;DH;��G;łG;��F;�9E;RA;�8;h�';��;�:�\���Z�jT��U�$��I��ʖռ���Xc������ս���5��9b��M������r���/5ʾ�*־      ���쾳�޾/5ʾL;���:��(�v��E�_'����q����u���+��W��A����4���Ļ9)�hj��W�:b�;%;�k7;$�@;��D;��F;�wG;U�G;1H;;CH;'iH;�H;��H;��H;��H;��H;r�H;��H;��H;��H;��H;�H;$iH;DCH;4H;W�G;�wG;��F;��D;$�@;�k7;%;`�;�W�:pj��9)���Ļ��4��A���W缃�+���u�q�����`'��E�(�v��:��L;��/5ʾ��޾��      Vh���b���쾦*־�v��(���*��'�O�U� �s��r���؀�F�3���>ݜ�<�>�P�ѻߡ9�����%o�:>% ;rM#;B�6;NA@;��D;��F;qG;J�G;H;�@H;egH;��H;��H;ܩH;�H;��H;�H;��H;�H;ީH;��H;��H;cgH;�@H;H;M�G;qG;��F;��D;KA@;<�6;nM#;<% ;+o�:����ܡ9�R�ѻ<�>�>ݜ���F�3��؀��r��s�U� �'�O�*��(����v���*־���b��      1�$��� ����#��@��'�þ�*��1Dx���=�����Pν���"'K��c���o�V����E^���S��w[:���:e;*�4;G`?;�mD;R�F;LvG;�G;=H;`OH;�sH;��H;z�H;~�H;�H;S�H;&�H;O�H;�H;��H;x�H;��H;�sH;kOH;=H;�G;PvG;^�F;�mD;B`?;"�4;e;���:�w[:��S�E^����o�V����c�!'K�����Pν�����=�0Dx��*��'�þ@��#������� �      �� ����R��O��/������0��4�s�׀:�g9��ʽ1Z����G��8�
.���5S�����/X���D�jBd:�B�: ;��4;ʈ?;�~D;�F;yG;��G;O H;)PH;tH;�H;ˢH;ŰH;)�H;o�H;4�H;m�H;,�H;ưH;ˢH;�H;tH;3PH;Q H;��G;yG;�F;�~D;ǈ?;��4; ;�B�:zBd:��D��/X���껭5S�	.���8���G�1Z���ʽg9�׀:�4�s��0�����/��O��R�����      ���R��8�
������Yؾ���ޥ����f���0�Z[�N8��ϐ���>�����IȤ��6H�a�ܻrF�Ȗ��}:��:c";0�5;��?;S�D;��F;�G;��G;0#H;`RH;�uH;E�H;��H;v�H;úH;�H;��H;�H;úH;v�H;��H;E�H;�uH;gRH;2#H;��G;	�G;��F;T�D;��?;)�5;`";��: �}:Ԗ�rF�a�ܻ�6H�HȤ������>�ΐ��N8��Z[���0���f�ޥ������Yؾ����8�
�R��      #��N������<I�(�þ�R��;���tS��Q"��s������}��0��켈�����6�G�ƻ8}*������:{x;X%;�l7;ܳ@;��D;��F;��G;��G;�'H;�UH;]xH;K�H;D�H;��H;��H;��H;w�H;��H;��H;��H;C�H;K�H;ZxH;�UH;�'H;��G;��G;��F;��D;س@;�l7;X%;zx;��: ���6}*�F�ƻ��6��������0���}�����s��Q"�tS�;����R��(�þ<Iᾣ���O��      @��/�待Yؾ(�þ
Ī�|쏾�k�׀:�~�z�ؽ�����c�\y���Ҽ����C� �i�*�� !(7E�:��
;��(;�_9;��A;g\E;n�F;��G;��G;�.H;�ZH;�{H;�H;H�H;P�H;	�H;��H;v�H;��H;�H;P�H;G�H;�H;�{H;�ZH;�.H;��G;��G;s�F;f\E;��A;{_9;��(;��
;M�:  (7)��h�C� �������Ҽ\y��c�����{�ؽ~�׀:��k�|쏾
Ī�(�þ�Yؾ/��      '�þ�������R��|쏾4�s��H�����������ΐ����D��c�����<�f�S,�����P��@�9˳�:�;!j-;P�;;s�B;��E;\G;��G;��G;�6H;�`H;W�H;J�H;ҩH;M�H;��H;R�H;��H;O�H;��H;K�H;ѩH;J�H;V�H;�`H;�6H;��G;��G;`G;��E;p�B;K�;;!j-;�;ѳ�:8�9�P�����S,�;�f������c���D�ΐ�������������H�4�s�|쏾�R��������      �*���0��ޥ��;����k��H��#%�Z[��Pνt��`�f�2/%���伅���t�=��?ػ�FL���D�d�R:��:3�;42;��=;��C;f0F;FGG;��G;#H;�?H;�gH;��H;)�H;��H;��H;~�H;��H;r�H;��H;��H;��H;��H;'�H;��H;�gH;�?H;#H;��G;JGG;f0F;��C;��=;42;0�;��:d�R:��D��FL��?ػs�=��������1/%�`�f�t���PνZ[��#%��H��k�;���ޥ���0��      0Dx�4�s���f�tS�׀:����Z[��7ս�榽��}���;��8�T�����r����:G���� ͬ�!��:
�;�}$;6;�?;�D;ǔF;�pG;��G;�H; JH;>oH;9�H;u�H;��H;6�H;��H;��H;&�H;��H;��H;9�H;��H;s�H;:�H;GoH;$JH;�H;��G;�pG;ǔF;�D;�?;ń6;�}$;�;%��: ͬ���:G�������r�T����8���;���}��榽�7սZ[����׀:�tS���f�4�s�      ��=�ր:���0��Q"�~������Pν�榽?����G�1����Ҽ ��HE:�<�ܻ�D^�����`i:=��:�;6|,;��:;L�A;AiE;��F;�G;�G;�(H;1UH;ywH;o�H;!�H;��H;�H;��H;��H;�H;��H;��H;�H;��H;!�H;o�H;�wH;5UH;�(H;~�G;�G;��F;<iE;N�A;��:;6|,;�;A��:`i:�����D^�:�ܻGE:� ����Ҽ1����G�?���榽�Pν����~��Q"���0�ր:�      ���g9�Z[��s�z�ؽ���t����}���G�����0c��V�V�E,��*����� ����:��:S ;c�3;�0>;ĚC;�F;�8G;+�G;kH;�7H;�`H;�H;�H;��H;I�H;��H;E�H;��H;�H;��H;I�H;��H;H�H;��H;�H;�H;�`H;�7H;iH;*�G;�8G;�F;ƚC;�0>;b�3;W ;��:��:�������*��D,�U�V�/c��������G���}�t�����{�ؽ�s�Z[�g9�      �Pν�ʽN8���������ΐ��`�f���;�1�����BȤ�3�f�)��Lߵ�So5���D�(�-:F��:�>;�+;�_9;�A;f�D;!�F;�vG;��G;H;tGH;WlH;��H;��H;��H;,�H;��H;��H;�H;$�H;�H;��H;��H;*�H;�H;��H;ǈH;alH;vGH;H;��G;�vG;�F;h�D;�A;�_9;�+;�>;D��:H�-:��D�Po5�Jߵ�(��2�f�AȤ����1����;�`�f�ΐ���������N8���ʽ      ���1Z��ΐ����}��c���D�1/%��8���Ҽ/c��2�f�����ƻ|/X�V������9�:=�;�";��3;=>;AYC;t�E;�G;�G;c�G;�,H;�VH;xH;��H;.�H;�H;�H;��H;0�H;D�H;.�H;E�H;1�H;��H;�H;�H;2�H;��H;xH;WH;�,H;b�G;�G;�G;x�E;FYC;>>;��3;�";=�;�:���9R���x/X��ƻ���1�f�0c����Ҽ�8�1/%���D��c���}�ΐ��1Z��      "'K���G��>��0�[y��c����S��� ��U�V�(���ƻ�od���º }(7�4�:���:��;�P.;ѡ:;zA;,�D;ǨF;MnG;8�G;�H;�@H;"fH;\�H;+�H;��H;ӸH;��H;��H;��H;z�H;7�H;{�H;��H;��H;��H;ѸH;��H;3�H;d�H;$fH;�@H;�H;>�G;MnG;ɨF;.�D;zA;ܡ:;�P.;��;���:�4�: �(7v�º�od��ƻ'��U�V� ��R�����伔c�\y��0��>���G�      �c��8���������Ҽ����������r�HE:�D,�Jߵ�~/X���º Ǭ�h�}:�:�;I�);$m7;�?;��C;F;U)G;�G;E�G;�)H;�SH;�tH;[�H;z�H;�H;��H;��H;��H;�H;��H;L�H;��H;�H;��H;��H;��H;�H;��H;f�H;�tH;�SH;�)H;J�G;�G;\)G;
F;��C;�?;'m7;H�);�;�:t�}:�Ƭ���ºz/X�Hߵ�D,�EE:���r�����������Ҽ�켶����8�      ��
.��IȤ���������;�f�s�=����<�ܻ�*��Oo5�`��� {(7p�}:�n�:,�;�>&;��4;��=;��B;�E;�F;��G;��G;*H;AH;�eH;:�H;ИH;V�H;ڷH;g�H; �H;��H;k�H;��H;Q�H;��H;j�H;��H;�H;d�H;ݷH;]�H;ؘH;@�H;�eH;}AH;1H;��G;��G;�F;�E;��B;��=;��4;�>&;,�;�n�:|�}: (7V���Lo5��*��8�ܻ���s�=�8�f���������JȤ�
.��      i�V��5S��6H���6�B� �S,��?ػ6G���D^������D����9�4�:�:,�;�%;��3;�<;VB;�E;��F;�XG;��G;E H;g0H;KWH;XvH;�H;x�H;��H;��H;��H;p�H;N�H;��H;��H;8�H;��H;��H;N�H;m�H;��H;��H;��H;�H;�H;\vH;GWH;l0H;E H; �G;�XG;�F;�E;XB;�<;��3;�%;0�;	�:�4�:���9��D�����D^�5G���?ػQ,�E� ���6��6H��5S�      ��ﻪ��e�ܻG�ƻd󩻶���FL�������`��H�-:�:���:�;�>&;��3;R9<;�A;ڰD;AZF;5G;��G;��G;i!H;)JH;-kH;��H;��H;a�H;��H;��H;��H;��H;��H;��H;c�H;��H;^�H;��H;��H;��H;��H;��H;��H;g�H;��H;��H;*kH;2JH;j!H;��G;��G;5G;HZF;ݰD;�A;U9<;��3;�>&;�;���:�:X�-:������� ���FL����g�J�ƻi�ܻ���      �D^��/X�rF�*}*����P����D�@̬�hi:��:J��:7�;��;F�);��4;�<;�A;&�D;t9F;�G;n�G;C�G;=H;?H;XaH;}H;{�H;t�H;��H;�H;��H;b�H;�H;�H;��H;%�H;��H;#�H;��H;�H;{�H;_�H;��H;�H;��H;v�H;|�H;}H;^aH;?H;:H;G�G;q�G;�G;w9F;#�D;�A;�<;��4;F�);��;9�;X��:��:ti:�ˬ���D��P����0}*��qF��/X�      <�S���D�Ȗ�Ȇ�� "(7��9��R:1��:E��:��:�>;�";�P.;(m7;��=;YB;۰D;~9F;G;�G;R�G;�H;�6H;hYH;�uH;�H;�H;��H;��H;��H;�H;��H;�H;5�H;^�H;��H;��H;��H;]�H;4�H;�H;��H; �H;��H;��H;��H;�H;�H;�uH;lYH;�6H;�H;W�G;�G; G;v9F;߰D;UB;��=;(m7;�P.;�";�>;��:M��:3��:��R:��9 $(70���Ȗ���D�      jw[:nBd:4�}:��:E�:ճ�:�:�;�;X ;�+;��3;ء:;�?;��B;�E;FZF;�G;�G;p�G;>H;T1H;�SH;^pH;ׇH;G�H;�H;x�H;��H;��H;��H;��H;o�H;!�H;��H;�H;X�H;�H;��H;�H;o�H;��H;��H;��H;��H;|�H;�H;E�H;ۇH;apH;�SH;U1H;DH;p�G;�G;�G;FZF;�E;��B;�?;١:;��3;�+;W ;�;�;�:��:I�:��:�}:BBd:      &��:�B�:���:px;��
;�;2�;�}$;6|,;c�3;�_9;8>;zA;��C;�E;�F;5G;v�G;U�G;>H;�/H;�PH;mH;F�H;��H;��H;n�H;��H;��H;�H;Z�H;��H;��H;��H;i�H;K�H;��H;D�H;j�H;��H;��H;��H;\�H;�H;��H;��H;k�H;��H;��H;F�H;�lH;�PH;�/H;>H;W�G;r�G;5G;�F;�E;��C;zA;;>;�_9;c�3;4|,;�}$;7�;�;��
;px;ֆ�:�B�:      e; ;r";h%;��(;"j-;42;��6;��:;�0>;�A;AYC;.�D;F;�F;�XG;��G;I�G;�H;U1H;�PH;�kH;u�H;{�H;1�H;.�H;ּH;��H;��H;�H;j�H;��H;u�H;n�H;��H;`�H;��H;Z�H;��H;m�H;s�H;��H;m�H;�H;��H;��H;ѼH;,�H;5�H;z�H;n�H;�kH;�PH;U1H;�H;F�G;��G;�XG;�F;F;.�D;DYC;�A;�0>;��:;Ʉ6;82;j-;��(;Z%;f"; ;      ?�4;��4;)�5;�l7;}_9;V�;;��=;
�?;U�A;ʚC;p�D;{�E;̨F;`)G;��G;�G;��G;DH;�6H;�SH; mH;r�H;��H;
�H;��H;P�H;"�H;2�H;��H;�H;�H;��H;2�H;��H;��H;a�H;��H;[�H;��H;��H;.�H;��H;�H;~�H;��H;4�H;�H;P�H;��H;�H;��H;u�H;mH;�SH;�6H;=H;��G;�G;��G;])G;̨F;~�E;p�D;ƚC;V�A;�?;��=;S�;;�_9;�l7;&�5;��4;      H`?;Ԉ?;��?;ٳ@;��A;v�B;��C;�D;5iE;�F;#�F;�G;MnG;�G;��G;H H;i!H;?H;lYH;^pH;H�H;v�H;�H;E�H;��H;&�H;A�H;�H;��H;r�H;R�H;��H;��H;��H;��H;<�H;M�H;6�H;��H;��H;��H;��H;S�H;p�H;��H;�H;=�H;(�H;��H;B�H;�H;x�H;F�H;]pH;iYH;?H;l!H;H H;��G;�G;KnG;�G;&�F;�F;>iE;��D;��C;d�B;��A;ӳ@;��?;ˈ?;      �mD;�~D;R�D;��D;a\E;��E;s0F;ƔF;��F;�8G;�vG;�G;<�G;O�G;/H;s0H;6JH;haH;�uH;�H;��H;6�H;��H;��H;��H;��H;j�H;�H;��H;��H;\�H;@�H;��H;��H;��H;��H;)�H;��H;��H;��H;��H;:�H;^�H;��H;��H;�H;e�H;��H;��H;��H;��H;8�H;��H;��H;�uH;caH;6JH;r0H;1H;L�G;>�G;�G;�vG;�8G;��F;ȔF;s0F;��E;m\E;��D;P�D;�~D;      J�F;�F;��F;��F;h�F;`G;PGG;�pG;�G;0�G;��G;f�G;�H;*H;AH;OWH;0kH;}H;�H;E�H;��H;(�H;N�H;(�H;��H;0�H;��H;��H;��H;�H;�H;��H;��H;��H;:�H;��H;��H;��H;7�H;��H;��H;��H;�H;�H;��H;��H;��H;3�H;��H;%�H;L�H;)�H;��H;B�H;�H;}H;2kH;NWH;AH;*H;�H;g�G;��G;1�G;�G;�pG;NGG;XG;}�F;��F;��F;�F;      avG;yG;�G;��G;��G;��G;��G;��G;{�G;iH;H;�,H;�@H;�SH;�eH;\vH;��H;��H;�H;�H;r�H;ԼH;%�H;G�H;h�H;��H;c�H;]�H;��H;��H;^�H;��H;��H;@�H;��H;%�H;#�H;�H;��H;A�H;��H;��H;^�H;��H;��H;\�H;^�H;��H;k�H;A�H;#�H;ּH;p�H;�H;�H;y�H;��H;[vH;�eH;�SH;�@H;�,H;H;iH;}�G;��G;��G;��G;ǝG;��G;�G;�xG;      �G;��G;��G;��G;��G;��G;1H;�H;�(H;�7H;vGH;WH;"fH;�tH;<�H;�H;��H;v�H;��H;x�H;��H;��H;0�H;�H;�H;�H;]�H;��H;��H;e�H;��H;��H;V�H;��H;O�H;��H;��H;��H;M�H;��H;V�H;��H;��H;d�H;��H;��H;X�H;��H;�H;�H;0�H;��H;��H;v�H;��H;q�H;��H;�H;9�H;�tH;$fH;WH;|GH;�7H;�(H;�H;0H;��G;��G;��G;��G;��G;      :H;F H;0#H;(H;u.H;�6H;�?H;JH;*UH;�`H;^lH;xH;`�H;`�H;ԘH;�H;j�H;��H;�H;��H;��H;��H;��H;��H;��H;��H;��H;��H;4�H;��H;��H;O�H;��H;r�H;��H;��H;��H;��H;��H;s�H;��H;I�H;��H;��H;1�H;��H;��H;��H;��H;��H;��H;��H;��H;��H;�H;��H;g�H;�H;ԘH;_�H;^�H;xH;blH;�`H;.UH;JH;�?H;6H;�.H; (H;-#H;I H;      aOH;"PH;nRH;�UH;�ZH;�`H;�gH;=oH;}wH;�H;ňH;��H;2�H;��H;X�H;��H;��H;�H;��H;��H;�H;	�H;}�H;p�H;��H;	�H;��H;g�H;��H;��H;H�H;��H;g�H;��H;��H;�H;4�H;�H;��H;��H;g�H;��H;H�H;��H;��H;d�H;��H;�H;��H;l�H;~�H;�H;�H;��H;��H;�H;��H;��H;X�H;��H;2�H;��H;ƈH;�H;wH;BoH;�gH;�`H;�ZH;�UH;mRH;#PH;      �sH;)tH;�uH;`xH;�{H;X�H;��H;=�H;s�H;�H;��H;6�H;��H;��H;�H;��H;��H;��H;#�H;�H;d�H;p�H;�H;U�H;_�H;�H;`�H;��H;��H;O�H;��H;k�H;��H;�H;X�H;c�H;[�H;a�H;W�H;�H;��H;h�H;��H;N�H;��H;��H;]�H;�H;c�H;S�H;�H;n�H;`�H;��H;#�H;��H;��H;��H;�H;��H;��H;9�H;��H;�H;s�H;@�H;��H;M�H;�{H;^xH;�uH;,tH;      ��H;
�H;F�H;J�H;�H;B�H;3�H;v�H;(�H;��H;��H;�H;ڸH;��H;f�H;��H;��H;f�H;��H;��H;��H;��H;��H;��H;@�H;��H;��H;��H;O�H;��H;d�H;��H;�H;Z�H;��H;�H;��H;��H;��H;[�H;�H;��H;b�H;��H;L�H;��H;��H;��H;B�H;��H;��H;��H;��H;��H;��H;g�H;��H;��H;g�H;��H;ظH;�H;��H;��H;'�H;w�H;8�H;C�H;��H;J�H;P�H;�H;      ��H;٢H;ϣH;F�H;P�H;ѩH;��H;��H;��H;N�H;2�H;�H;��H;��H;"�H;s�H;��H;��H;�H;v�H;��H;y�H;0�H;��H;��H;��H;��H;]�H;��H;n�H;��H;�H;S�H;��H;��H;��H;��H;��H;��H;��H;S�H;�H;��H;i�H;��H;W�H;��H;��H;��H;��H;5�H;w�H;��H;u�H;�H;��H;��H;v�H;"�H;��H;��H;�H;3�H;N�H;��H;��H;��H;˩H;V�H;@�H;٣H;٢H;      }�H;��H;w�H;��H;T�H;D�H;��H;;�H;��H;��H; �H;��H;��H;��H;��H;U�H;��H;!�H;<�H;&�H;��H;q�H;��H;��H;��H;��H;=�H;��H;r�H;��H;	�H;[�H;��H;��H;��H;��H;��H;��H;��H;��H;��H;Z�H;�H;��H;n�H;��H;;�H;��H;��H;��H;��H;p�H;��H;�H;;�H;"�H;��H;V�H;��H;��H;��H;��H;�H;��H;��H;>�H;��H;C�H;[�H;��H;��H;ͰH;      �H;@�H;ѺH;��H;�H;��H;��H;��H;��H;R�H;��H;<�H;��H;�H;r�H;��H;��H;��H;a�H;��H;p�H;��H;��H;��H;��H;3�H;��H;O�H;��H;�H;T�H;��H;��H;��H;��H;��H;��H;��H;��H;��H;��H;��H;P�H;��H;��H;J�H;��H;3�H;��H;��H;��H;��H;i�H;��H;^�H;��H;��H;��H;q�H;�H;��H;<�H;��H;S�H;��H;��H;��H;��H;�H;��H;ҺH;?�H;      O�H;m�H;�H;��H;��H;G�H; �H;��H;��H;��H;�H;L�H;��H;��H;��H;��H;e�H;#�H;��H;�H;O�H;^�H;[�H;.�H;��H;��H;"�H;��H;��H;$�H;a�H;��H;��H;��H;��H;��H;��H;��H;��H;��H;��H;��H;_�H;�H;��H;��H; �H;��H;��H;/�H;_�H;[�H;H�H;�H;��H;)�H;f�H;��H;��H;��H;�H;K�H;�H;��H;��H;��H;�H;I�H;��H;��H;�H;|�H;      +�H;2�H;��H;w�H;r�H;��H;z�H;)�H;�H;�H;3�H;<�H;D�H;Z�H;[�H;?�H;��H;��H;��H;b�H;��H;��H;��H;F�H;)�H;��H;"�H;��H;��H;?�H;X�H;��H;��H;��H;��H;��H;��H;��H;��H;��H;��H;��H;W�H;8�H;��H;��H; �H;��H;(�H;D�H;��H;��H;��H;]�H;��H;��H;��H;?�H;Y�H;Z�H;C�H;<�H;3�H;�H;�H;-�H;�H;��H;t�H;w�H;��H;;�H;      P�H;q�H;�H;��H;��H;L�H;��H;��H;��H;��H;�H;K�H;��H;��H;��H;��H;e�H;&�H;��H;�H;P�H;`�H;[�H;.�H;��H;��H;"�H;��H;��H;#�H;a�H;��H;��H;��H;��H;��H;��H;��H;��H;��H;��H;��H;_�H;�H;��H;��H;�H;��H;��H;,�H;^�H;X�H;H�H;�H;��H;(�H;e�H;��H;��H;��H;��H;K�H;�H;��H;��H;��H;�H;H�H;��H;��H;�H;y�H;      ߹H;A�H;˺H;��H;�H;��H;��H;��H;��H;R�H;��H;<�H;��H;�H;t�H;��H;��H;��H;`�H;��H;q�H;��H;��H;��H;��H;2�H;��H;P�H;��H; �H;T�H;��H;��H;��H;��H;��H;��H;��H;��H;��H;��H;��H;Q�H;��H;��H;I�H;��H;4�H;��H;��H;��H;��H;g�H;��H;^�H;��H;��H;��H;o�H;�H;��H;>�H;��H;P�H;��H;��H;��H;��H;�H;��H;ѺH;A�H;      }�H;��H;w�H;��H;T�H;H�H;��H;>�H;��H;��H;�H;��H;��H;��H;��H;U�H;��H;#�H;<�H;%�H;��H;r�H;��H;��H;��H;��H;@�H;��H;u�H;��H;�H;[�H;��H;��H;��H;��H;��H;��H;��H;��H;��H;X�H;�H;��H;l�H;��H;:�H;��H;��H;��H;��H;p�H;��H;!�H;9�H;�H;��H;V�H;��H;��H;��H;��H;��H;��H;��H;@�H;��H;F�H;]�H;��H;�H;°H;      �H;ߢH;ͣH;C�H;L�H;ԩH;��H;��H;��H;N�H;3�H;�H;��H;��H;%�H;t�H;��H;��H;�H;y�H;��H;y�H;/�H;��H;��H;��H;��H;]�H;��H;o�H;��H;�H;Q�H;��H;��H;��H;��H;��H;��H;��H;Q�H;�H;��H;g�H;��H;U�H;��H;��H;��H;��H;5�H;u�H;��H;u�H;�H;��H;��H;t�H;"�H;��H;��H;�H;2�H;L�H;��H;��H;��H;ΩH;R�H;J�H;ڣH;آH;      ��H;�H;7�H;F�H;�H;S�H;4�H;y�H;&�H;��H;��H;�H;ظH;��H;j�H;��H;��H;g�H;��H;��H;��H;��H;��H;��H;B�H;��H;��H;��H;R�H;��H;d�H;��H;�H;X�H;��H;�H;��H;��H;��H;Z�H;�H;��H;`�H;��H;H�H;��H;��H;��H;>�H;��H;��H;��H;��H;��H;��H;f�H;��H;��H;g�H;��H;ظH;�H;��H;��H;(�H;z�H;:�H;F�H;�H;G�H;<�H;�H;      �sH;)tH;�uH;ZxH;�{H;X�H;��H;;�H;s�H;�H;��H;;�H;��H;��H;�H;��H;��H;��H;#�H;��H;e�H;q�H;�H;U�H;a�H;
�H;]�H;��H;��H;N�H;��H;l�H;��H;�H;Z�H;b�H;[�H;c�H;W�H;�H;��H;i�H;��H;I�H;��H;��H;[�H;�H;^�H;O�H;�H;n�H;]�H;��H;%�H;��H;��H;��H;�H;��H;��H;9�H;��H;�H;s�H;B�H;��H;T�H;�{H;exH;�uH;*tH;      nOH;)PH;dRH;�UH;�ZH;�`H;�gH;GoH;�wH;�H;ǈH;��H;3�H;��H;\�H;��H;��H;�H;��H;��H;�H;�H;x�H;n�H;��H;�H;��H;e�H;��H;��H;I�H;��H;e�H;��H;��H;�H;4�H;�H;��H;��H;h�H;��H;H�H;|�H;��H;^�H;��H;�H;��H;h�H;��H;�H;�H;��H;��H;ݾH;��H;��H;Y�H;��H;2�H;��H;ƈH;�H;}wH;EoH;�gH;�`H;�ZH;�UH;wRH; PH;      GH;F H;A#H;�'H;m.H;�6H;�?H;JH;2UH;�`H;`lH;xH;^�H;b�H;טH;��H;h�H;��H; �H;��H;��H;��H;��H;��H;��H;��H;��H;��H;5�H;��H;��H;P�H;��H;s�H;��H;��H;��H;��H;��H;r�H;��H;N�H;��H;��H;-�H;��H;��H;��H;��H;��H;��H;��H;��H;��H; �H;��H;e�H;�H;֘H;`�H;`�H;xH;alH;�`H;4UH;!JH;�?H;�6H;|.H;�'H;@#H;A H;      !�G;��G;��G;��G;��G;��G;0H;�H;�(H;�7H;yGH;WH;$fH;�tH;=�H;�H;��H;w�H;��H;x�H;��H;��H;-�H;�H;�H;x�H;Y�H;��H;��H;a�H;��H;��H;U�H;��H;P�H;��H;��H;��H;O�H;��H;W�H;��H;��H;a�H;��H;��H;X�H;}�H;�H;�H;6�H;��H;��H;v�H;��H;p�H;��H;�H;?�H;�tH;"fH;WH;yGH;�7H;�(H;�H;-H;��G;��G;��G;��G;��G;      OvG;yG;�G;��G;��G;��G;��G;��G;~�G;iH;H;�,H;�@H;�SH;�eH;]vH;��H;��H;�H;�H;s�H;׼H;�H;G�H;j�H;��H;`�H;]�H;��H;��H;]�H;��H;��H;A�H;��H; �H;#�H; �H;��H;B�H;��H;��H;`�H;��H;��H;Y�H;]�H;��H;k�H;A�H;)�H;ּH;p�H;�H;�H;{�H;��H;\vH;�eH;�SH;�@H;�,H;H;hH;}�G;��G;��G;��G;ŝG;��G;
�G;	yG;      B�F;�F;��F;��F;n�F;iG;IGG;�pG;�G;0�G;��G;j�G;�H;*H;�AH;OWH;/kH;}H;�H;E�H;��H;+�H;I�H;(�H;��H;-�H;��H;��H;��H;�H;�H;��H;��H;��H;:�H;��H;��H;��H;7�H;��H;��H;��H;�H;�H;��H;|�H;��H;2�H;��H;%�H;P�H;(�H;��H;D�H;�H;}H;0kH;NWH;�AH;*H;�H;f�G;��G;1�G;�G;�pG;JGG;[G;v�F;��F;��F;�F;      �mD;�~D;M�D;��D;`\E;��E;p0F;ƔF;��F;�8G;�vG;�G;<�G;M�G;4H;s0H;6JH;haH;�uH;�H;��H;;�H;��H;��H;��H;��H;e�H;�H;��H;��H;\�H;A�H;��H;��H;��H;��H;(�H;��H;��H;��H;��H;A�H;b�H;��H;��H;�H;g�H;��H;��H;��H;��H;8�H;��H;��H;�uH;aaH;5JH;p0H;4H;L�G;<�G;�G;�vG;�8G;��F;ǔF;r0F;��E;j\E;��D;O�D;�~D;      (`?;��?;��?;�@;��A;}�B;��C;�D;CiE;�F;'�F;�G;KnG;�G;��G;I H;j!H;?H;hYH;^pH;I�H;x�H;�H;E�H;��H;!�H;?�H;�H;��H;p�H;S�H;��H;��H;��H;��H;7�H;O�H;9�H;��H;��H;��H;��H;W�H;p�H;��H;�H;A�H;&�H;��H;E�H;�H;v�H;F�H;^pH;iYH;?H;j!H;H H;��G;�G;JnG;�G;&�F;�F;>iE;�D;��C;p�B;��A;�@;��?;��?;      1�4;��4;�5;�l7;z_9;P�;;��=;
�?;[�A;ɚC;m�D;~�E;̨F;_)G;��G;�G;��G;DH;�6H;�SH;mH;u�H;��H;
�H;��H;K�H;�H;3�H;��H;z�H;�H;��H;0�H;��H;��H;a�H;��H;_�H;��H;��H;0�H;��H;�H;��H;��H;2�H;"�H;O�H;��H;�H;��H;r�H;mH;�SH;�6H;=H;��G; �G;��G;[)G;̨F;y�E;j�D;ǚC;U�A;�?;��=;P�;;w_9;�l7;�5;��4;      e; ;f";\%;��(;(j-;82;Ƅ6;��:;�0>;�A;FYC;.�D;
F;�F;�XG;��G;I�G;�H;W1H;�PH;�kH;r�H;z�H;6�H;'�H;ӼH;��H;��H;�H;m�H;��H;s�H;n�H;��H;[�H;��H;]�H;��H;k�H;u�H;��H;p�H;�H;��H;��H;ԼH;,�H;1�H;}�H;t�H;�kH;�PH;W1H;�H;F�G;��G;�XG;�F;	F;.�D;AYC;�A;�0>;��:;Ȅ6;02;j-;�(;N%;f";  ;      ��:�B�:��:yx;��
;�;4�;�}$;:|,;b�3;�_9;=>;zA;��C;�E;�F;5G;v�G;U�G;?H;�/H;�PH;mH;H�H;��H;��H;h�H;��H;��H;�H;]�H;��H;��H;��H;j�H;G�H;��H;H�H;i�H;��H;��H;��H;^�H;�H;��H;��H;l�H;��H;��H;H�H;mH;�PH;�/H;?H;W�G;t�G;5G;�F;�E;��C;zA;8>;�_9;c�3;6|,;�}$;9�;�;��
;wx;���:�B�:      �w[:�Bd: �}:��:C�:��:�:�;�;X ;�+;��3;ܡ:;�?;��B;�E;FZF;�G;�G;p�G;DH;X1H;�SH;`pH;݇H;E�H;ߪH;x�H;��H;��H;��H;��H;s�H;#�H;��H;�H;[�H;�H;��H;�H;p�H;��H;��H;��H;��H;v�H;�H;G�H;ׇH;bpH;�SH;U1H;AH;p�G;�G;�G;EZF;�E;��B;�?;١:;��3;�+;W ;�;�;�:ϳ�:M�:��:$�}:^Bd:      <�S���D�Ė�؆�� (7��9��R:/��:O��:��:�>;�";�P.;(m7;��=;YB;ݰD;z9F;G;�G;X�G;�H;�6H;iYH;�uH;�H;�H;��H;��H;��H;�H;��H;�H;6�H;a�H;��H;��H;��H;]�H;5�H;�H;��H;"�H;��H;��H;��H;�H;�H;�uH;lYH;�6H;�H;U�G;�G;G;v9F;۰D;SB;��=;%m7;�P.;�";�>;��:K��:1��:��R:��9 (7؆��ܖ���D�       E^��/X�
rF�/}*����P����D�`ˬ�|i:��:R��::�;��;H�);��4;�<;�A;$�D;v9F;�G;r�G;F�G;AH;?H;^aH;}H;x�H;t�H;��H;�H;��H;`�H;�H;�H;��H;&�H;��H;&�H;��H;�H;�H;_�H;��H;�H;��H;s�H;{�H;}H;XaH;?H;>H;C�G;m�G;�G;t9F;#�D;�A;�<;��4;D�);��;7�;V��:��:ti:�ˬ���D��P����3}*�rF��/X�      ��ﻫ��e�ܻF�ƻd󩻶���FL� ������`��P�-:�:���:�;�>&;��3;U9<;�A;ڰD;EZF;!5G;��G;��G;l!H;2JH;-kH;��H;��H;h�H;��H;��H;��H;��H;��H;��H;c�H;��H;c�H;��H;��H;��H;��H;��H;��H;g�H;��H;��H;*kH;,JH;l!H;��G;��G;5G;FZF;ڰD;�A;T9<;��3;�>&;�;���:�:L�-:����������FL����i�I�ƻj�ܻ���      i�V��5S��6H���6�C� �Q,��?ػ4G���D^������D����9�4�:	�:1�;�%;��3;�<;SB;�E;�F;�XG;�G;F H;l0H;LWH;XvH;�H;~�H;��H;��H;��H;p�H;T�H;��H;��H;8�H;��H;��H;M�H;m�H;��H;��H;��H;|�H;�H;VvH;IWH;g0H;E H;�G;�XG;��F;�E;SB;�<;��3;�%;.�;�:�4�:���9��D�����D^�6G���?ػQ,�E� ���6��6H��5S�      ��
.��JȤ���������:�f�s�=����:�ܻ�*��Lo5�\��� (7|�}:�n�:.�;�>&;��4;��=;��B;�E;�F;��G;��G;/H;�AH;�eH;=�H;טH;Y�H;޷H;g�H; �H;��H;j�H;��H;Q�H;��H;j�H;��H;�H;b�H;۷H;X�H;טH;:�H;�eH;}AH;-H;��G;��G;�F;�E;��B;��=;��4;�>&;*�;�n�:t�}: |(7\���Oo5��*��9�ܻ���s�=�9�f���������JȤ�
.��      �c��8���������Ҽ����������r�FE:�D,�Hߵ�{/X���º�Ƭ���}:�:�;F�);$m7;�?;��C;	F;Y)G;�G;L�G;*H;�SH;�tH;b�H;�H;�H;��H;��H;��H;�H;��H;M�H;��H;�H;��H;��H;��H;�H;��H;b�H;�tH;�SH;�)H;E�G;�G;\)G;F;��C;�?;#m7;F�);�;�:p�}:�Ƭ���º|/X�Jߵ�D,�GE:���r�����������Ҽ�켵����8�      "'K���G��>��0�[y��c����S��� ��U�V�'���ƻ�od�x�º �(7�4�:���:��;�P.;ա:;zA;-�D;̨F;QnG;>�G;�H;�@H;"fH;c�H;/�H;��H;ָH;��H;��H;��H;}�H;6�H;{�H;��H;��H;��H;иH;��H;0�H;c�H;"fH;�@H;�H;8�G;NnG;̨F;-�D;
zA;ڡ:;�P.;��;���:�4�: �(7~�º�od��ƻ(��U�V� ��S�����伔c�\y��0��>���G�      ���1Z��ΐ����}��c���D�1/%��8���Ҽ0c��1�f�����ƻz/X�R������9	�:9�;�";��3;A>;BYC;y�E;�G;�G;e�G;�,H;WH;xH;��H;4�H;�H;�H;��H;0�H;B�H;.�H;D�H;.�H;��H;�H;�H;1�H;��H;xH; WH;�,H;c�G;�G;�G;{�E;BYC;8>;��3;�";:�;�:���9R���}/X��ƻ���2�f�/c����Ҽ�8�1/%���D��c���}�ΐ��1Z��      �Pν�ʽN8���������ΐ��`�f���;�1����AȤ�2�f�(��Jߵ�Oo5���D�4�-:B��:�>;�+;�_9;�A;i�D;!�F;�vG;��G;H;vGH;^lH;ÈH;��H;��H;-�H;��H;��H;�H;$�H;�H;��H;��H;)�H;�H;��H;ňH;`lH;uGH;H;��G;�vG;#�F;j�D;�A;�_9;�+;�>;B��:<�-:��D�Qo5�Lߵ�(��3�f�AȤ����1����;�`�f�ΐ���������N8���ʽ      ���g9�Z[��s�z�ؽ���t����}���G�����/c��U�V�D,��*����������:��:T ;h�3;�0>;ƚC;�F;�8G;*�G;hH;�7H;�`H;
�H;�H;��H;I�H;��H;E�H;��H;�H;��H;E�H;��H;G�H;��H;�H;�H;�`H;�7H;fH;+�G;�8G;�F;ɚC;�0>;^�3;X ;��:��:�������*��E,�V�V�/c��������G���}�t�����{�ؽ�s�Z[�g9�      ��=�׀:���0��Q"�~������Pν�榽?����G�1����Ҽ ��GE:�:�ܻ�D^�����Xi:E��:�;:|,;��:;O�A;?iE;��F;�G;~�G;�(H;2UH;{wH;p�H; �H;��H;�H;��H;��H;�H;��H;��H;�H;��H;!�H;o�H;wH;5UH;�(H;~�G;�G;��F;CiE;N�A;��:;2|,;�;?��:\i:�����D^�;�ܻGE:� ����Ҽ1����G�?���榽�Pν����~��Q"���0�ր:�      0Dx�4�s���f�tS�ր:����Z[��7ս�榽��}���;��8�T�����r����9G�����ͬ�'��:�;�}$;ń6;�?;��D;ȔF;�pG;��G;�H; JH;>oH;:�H;u�H;��H;7�H;��H;��H;%�H;��H;��H;7�H;��H;s�H;:�H;EoH;"JH;�H;��G;�pG;ƔF;�D;�?;Ä6;�}$;�;!��: ͬ���:G�������r�T����8���;���}��榽�7սZ[����׀:�tS���f�4�s�      �*���0��ޥ��;����k��H��#%�Z[��Pνt��`�f�1/%���伅���t�=��?ػ�FL���D�h�R:��:3�;42;��=;��C;e0F;FGG;��G;"H;�?H;�gH;��H;)�H;��H;��H;}�H;��H;r�H;��H;��H;��H;��H;*�H;��H;�gH;�?H;%H;��G;MGG;e0F;��C;��=;22;/�;��:`�R:��D��FL��?ػt�=��������2/%�`�f�t���PνZ[��#%��H��k�;���ޥ���0��      '�þ�������R��{쏾5�s��H�����������ΐ����D��c�����;�f�S,�����P��H�9ѳ�:�;j-;P�;;u�B;��E;YG;��G;��G;�6H;�`H;Z�H;L�H;ҩH;N�H;��H;P�H;��H;R�H;��H;N�H;ҩH;L�H;W�H;�`H;�6H;��G;��G;cG;��E;v�B;M�;;j-;�;ճ�:8�9�P�����S,�;�f������c���D�ΐ�������������H�5�s�|쏾�R��������      @��/�待Yؾ(�þ
Ī�|쏾�k�ր:�~�z�ؽ�����c�\y���Ҽ����B� �h�,�� !(7I�:��
;��(;�_9;��A;h\E;k�F;��G;��G;�.H;�ZH;�{H;�H;G�H;Q�H;�H;��H;v�H;��H;�H;O�H;G�H;�H;�{H;�ZH;�.H;��G;��G;u�F;g\E;��A;}_9;��(;��
;M�: (7(��h�C� �������Ҽ\y��c�����z�ؽ~�׀:��k�|쏾
Ī�(�þ�Yؾ/��      #��O������<I�(�þ�R��;���tS��Q"��s������}��0��켈�����6�F�ƻ8}*������:{x;X%;�l7;ڳ@;��D;��F;��G;��G;�'H;�UH;^xH;K�H;C�H;��H;��H;��H;x�H;��H;��H;��H;D�H;M�H;]xH;�UH;�'H;��G;��G;��F;��D;ڳ@;�l7;X%;zx;��:���4}*�E�ƻ��6��������0���}�����s��Q"�tS�;����R��(�þ<Iᾣ���O��      ���R��8�
������Yؾ���ޥ����f���0�Z[�N8��ϐ���>�����IȤ��6H�`�ܻrF�Ȗ��}:��:b";/�5;��?;T�D;��F;�G;��G;/#H;_RH;�uH;E�H;��H;t�H;��H;�H;��H;�H;ĺH;v�H;��H;E�H;�uH;gRH;2#H;��G;�G;��F;T�D;��?;)�5;`";��:(�}:̖�rF�a�ܻ�6H�IȤ������>�ϐ��N8��Z[���0���f�ޥ������Yؾ����8�
�R��      �� ����R��N��/������0��4�s�ր:�g9��ʽ1Z����G��8�
.���5S�����/X�x�D�nBd:�B�: ;��4;ʈ?;�~D;�F;
yG;��G;M H;)PH;tH;�H;ˢH;ŰH;+�H;n�H;5�H;n�H;,�H;ǰH;ˢH;�H;tH;3PH;P H;��G;yG;�F;�~D;ǈ?;��4; ;�B�:~Bd:��D��/X���껭5S�	.���8���G�1Z���ʽg9�׀:�4�s��0�����/��N��R�����      FEb�`]��N��7����s� ���˾��(�j��!,�o���K��Bm�+��7,˼��x�[���1�����T�:l�:�;�1;9,>;c�C;UwF;�G;m H;�>H;�hH;*�H;A�H;�H;��H;��H;�H;l�H;�H;��H;��H;�H;A�H;)�H;�hH;�>H;p H;��G;_wF;c�C;3,>;
�1;�;n�:`�:����1��[����x�7,˼+��Bm�K��o����!,�(�j�����˾s� �����7��N�`]�      `]�d�W��TI�v3��D�������Ǿv����f�7)�$��r;���Fi��k���Ǽ�[t�M�	�*Ȅ� X��Р:��:��;.J2;TZ>;%	D;=F;7�G;�H;�?H;viH;H;��H;P�H;�H;��H;5�H;��H;1�H;��H;�H;P�H;��H;��H;}iH;�?H;�H;8�G;FF;%	D;OZ>;$J2;��;��:ܠ: X��(Ȅ�M�	��[t���Ǽ�k��Fi�r;��$��7)��f�v�����Ǿ�����D�v3��TI�d�W�      �N��TI���;�/�'�l��쾀���y󐾴Z��K ��s�@����&^���"����g����Ϩu�� ���2<:��:�
;<g3;��>;TBD;u�F;ܔG;iH;BH;ZkH;,�H;��H;�H;��H;?�H;��H;!�H;��H;A�H;��H;�H;��H;)�H;ckH;BH;lH;ߔG;��F;UBD;��>;4g3;�
;��:�2<:� ��Ψu������g��"����&^�@����s潥K ��Z�y󐾀�����l�/�'���;��TI�      �7�v3�/�'����s� ��{Ծ���H���y�F�����ӽ���^�L�Jv��뮼PT����PV���=�Z)i:t��:�z ;�$5;��?;�D;��F;�G;rH;bFH;qnH;a�H;J�H;H�H;��H;�H;/�H;��H;+�H;�H;��H;H�H;J�H;^�H;xnH;fFH;rH;�G;��F;�D;��?;y$5;�z ;t��:j)i:��=��PV���PT��뮼Jv�^�L�����ӽ���y�F�H�������{Ծs� ����/�'�v3�      ����D�l�s� �U�ݾj���U͓��f��>/�����'���섽O�6�~t�w��]�:�&Tʻz.�8۷�@t�:�;��$;�Y7;S�@;�	E;��F;)�G;�H;LH;�rH;��H;��H;��H;��H;�H;"�H;��H;!�H;�H;��H;��H;��H;��H;�rH;	LH;�H;)�G;��F;�	E;L�@;�Y7;��$;�;Jt�:@۷�z.�&Tʻ^�:�w��~t�O�6��섽�'������>/��f�U͓�j���V�ݾs� �l��D�      s� ��������{Ծj���v���Z�x��SC��^��޽?���w�e�'��B�Ѽ$G������R������ݤ8Ç�:�Y;E�);��9;��A;��E;G;�G;>!H;	SH;�wH;H�H;W�H;�H;��H;I�H;V�H;��H;R�H;K�H;��H;�H;Y�H;G�H;�wH;
SH;A!H;	�G;�G;��E;��A;��9;C�);�Y;ˇ�:�ݤ8����R�����#G��B�Ѽ'��w�e�?����޽�^��SC�Z�x�v���j����{Ծ�쾟���      ��˾��Ǿ�������U͓�Z�x���J��K �l���������?����뮼(�[����3|��W����:=�:�';a/;Bg<;�C;FF;�NG;��G;-H;9[H;�}H;��H;��H;��H;�H;��H;��H;��H;��H;��H;�H;��H;��H;��H;�}H;=[H;-H;��G;�NG;DF;�C;=g<;`/;�';E�:|�:�W��3|����(�[��뮼���?������l����K ���J�Y�x�U͓����������Ǿ      ��v���y�H����f��SC��K �nn����Ž���
�Z��k�}ռ,X��`y-�+���n.����P�:�+�:|�;4;�>;�D;�wF;��G;��G;�9H;&dH;S�H;~�H;0�H;H�H;��H;~�H;+�H;E�H;)�H;��H;��H;E�H;/�H;~�H;Z�H;*dH;�9H;��G;�G;�wF;�D;�>;4;y�;�+�:�P�:p��m.�+���_y-�,X��}ռ�k�
�Z������Žmn���K ��SC��f�H���y�v���      (�j��f��Z�y�F��>/��^�l�����ŽF ���Fi��Q+�zt�mT��m�W�����1��,ȺX�9wP�:�Y;��(;��8;�A;�E;��F;9�G;pH;�FH;�mH;h�H;��H;�H;G�H;��H;`�H;��H;��H;��H;a�H;��H;D�H;�H;��H;o�H;�mH;�FH;pH;6�G;��F;�E;�A;��8;~�(;�Y;wP�:X�9$Ⱥ�1�����l�W�mT��zt�Q+��Fi�F ����Žl����^��>/�y�F��Z��f�      �!,�7)��K ��������޽������Fi��0����鷼��x�����.��Q�(� ���*i:x��:%�;��0;8�<;rC;��E;�<G;��G;�$H;8TH;�wH;ŒH;�H;!�H;X�H;�H;c�H;s�H;O�H;q�H;f�H;�H;U�H;�H;�H;ΒH;�wH;;TH;�$H;��G;�<G;�E;tC;8�<;��0;,�;z��:�*i:���P�(��.�������x�鷼����0��Fi�������޽�������K �7)�      n���$��s��ӽ�'��?������
�Z��Q+�����"��G����0���׻ʕb�:W���X�9ԡ�:`;~*';�Y7;�#@;�D;��F;�G;��G;8H;�aH;ˁH;3�H;z�H;G�H;l�H;x�H;W�H;%�H;�H;&�H;Z�H;y�H;i�H;F�H;|�H;<�H;ҁH;�aH;8H;��G;�G;ߖF;�D;�#@;�Y7;�*'; `;ҡ�: Y�96W��ȕb���׻��0�G���"������Q+�
�Z����?����'���ӽ�s�$��      J��r;��@�������섽w�e��?��k�{t�鷼G���e7�����Ǆ�p0���t�u�:�+�:j;l1;B�<;K�B;�E;�G;��G;2H;PJH;2oH;ЋH;��H;�H;m�H;��H;��H;j�H;��H;��H;��H;j�H;��H;��H;k�H;�H;��H;ۋH;4oH;QJH;0H;��G;�G;�E;N�B;D�<;w1;n;�+�:&u�:@�t�l0��Ǆ���껂e7�G��鷼zt��k��?�v�e��섽���@���r;��      Bm��Fi��&^�_�L�N�6�'����}ռmT����x���0����������ط��n`:��:�;�*;�8;��@;�D;D�F;�}G;y�G;k1H;�[H;B|H;��H;��H;Y�H;��H;��H;^�H;h�H;��H;E�H;��H;g�H;^�H;��H;��H;]�H;��H;��H;F|H;�[H;h1H;�G;�}G;G�F;!�D;��@;'�8;�*;�;��:�n`:xط��������껾�0���x�lT��}ռ��'��O�6�_�L��&^��Fi�      )���k��Jv�{t�D�Ѽ�뮼,X��m�W������׻ Ȅ����� 5<:V��:�Y;�t%;�$5;�Z>;�`C;��E;*G;@�G;�H;�GH;ClH;ƈH;ҞH;��H;��H;n�H;��H;��H;K�H;F�H;�H;F�H;J�H;��H;��H;m�H;��H;��H;ܞH;ʈH;FlH;�GH;�H;A�G;*G;��E;�`C;�Z>;�$5;�t%;�Y;Z��:5<:������Ǆ���׻���k�W�+X���뮼B�Ѽ}t�Jv���k�      5,˼��Ǽ�"���뮼w��#G��'�[�]y-�����.��ȕb�x0㺨ط� 5<:�L�:�\;p�!;�J2;�g<;-0B;CE;�F;%�G;��G;\4H;u\H;�{H;}�H;v�H;/�H;��H;�H;i�H;$�H;&�H;��H;��H;��H;%�H;&�H;h�H;�H;��H;5�H;|�H;��H;�{H;r\H;b4H;��G;'�G;�F;CE;70B;�g<;�J2;x�!;�\;�L�:5<:�ط�p0�ĕb��.�����]y-�'�[�"G��w���뮼�"����Ǽ      ��x��[t���g�MT�]�:�������'����1��M�(�4W��@�t��n`:V��:�\;{ ;��0;R;;�<A;��D;�wF;�cG;+�G;�!H;MH;WoH;H�H;Y�H;��H;e�H;9�H;��H;/�H;D�H;��H;m�H;��H;j�H;��H;D�H;,�H;��H;=�H;i�H;��H;]�H;M�H;RoH;�MH;�!H;0�G;�cG;�wF;��D;�<A;M;;��0;{ ;�\;Z��:�n`:��t�0W��L�(��1��&���������_�:�OT���g��[t�      W��J�	������!Tʻ�R��3|�g.� Ⱥ���Y�9u�:��:�Y;v�!;��0;Օ:;��@;�BD;e2F;X8G;��G;�H;?@H;�cH;��H;H�H;�H;�H;!�H;d�H;��H;��H;@�H;��H;��H;W�H;��H;�H;@�H;��H;��H;i�H;$�H;�H;�H;K�H;��H;�cH;B@H;�H;��G;Z8G;j2F;�BD;��@;ؕ:;��0;x�!;�Y;��:$u�: Y�9���Ⱥf.�3|��R��$Tʻ�����H�	�      �1��$Ȅ�Ψu��PV�l.�����W��H��(X�9+i:ء�:�+�:�;�t%;�J2;K;;��@;\D;�F;G;W�G;gH;X5H;UZH;xH;�H;��H;�H;�H;-�H;?�H;��H;�H;��H;�H;0�H;��H;.�H;�H;��H;��H;��H;C�H;3�H;�H;�H;��H;�H;
xH;UZH;U5H;hH;X�G;	G;�F;YD;��@;H;;�J2;�t%;�;�+�:桼:+i:PX�9(��W�����h.��PV�Ĩu�%Ȅ�      ܥ��.X��� ��t�=�8۷��ߤ8��:�P�:P�:���:$`;j;�*;�$5;�g<;�<A;�BD;�F;�G;V�G;@�G;w-H;�RH;+qH;��H;��H;P�H;�H;�H;��H;��H;��H;%�H;��H;r�H;j�H;��H;g�H;p�H;��H;"�H;��H;��H;��H;�H;�H;Q�H;��H;��H;/qH;�RH;z-H;C�G;Z�G;�G;�F;�BD;�<A;�g<;�$5;�*;n;)`;���:�P�:�P�:��:�ޤ8 ۷���=�� ��0X��      D�:Р:�2<:�)i:Bt�:ɇ�:Y�:�+�:�Y;+�;�*';t1;#�8;�Z>;70B;��D;i2F;G;Y�G;��G;W)H;ZNH;IlH;�H;6�H;W�H;p�H;�H;Z�H;��H;�H;��H;�H;/�H;��H;��H;��H;��H;��H;.�H;�H;��H;	�H;��H;X�H;�H;p�H;U�H;<�H; �H;HlH;]NH;Y)H;��G;\�G;	G;i2F;��D;:0B;�Z>;$�8;w1;�*';,�;�Y;�+�:S�:ه�:Ht�:V)i:�2<:��:      ��:���:���:d��:�;�Y;�';w�;~�(;��0;�Y7;>�<;��@;�`C;CE;�wF;X8G;a�G;C�G;U)H;�LH;�iH;�H;.�H;x�H;��H;��H;7�H;��H;��H;��H;,�H;��H;o�H;��H;}�H;��H;v�H;��H;n�H;��H;(�H;��H;��H;��H;7�H;��H;��H;|�H;.�H;�H;�iH;�LH;W)H;C�G;\�G;Z8G;�wF;CE;�`C;��@;A�<;�Y7;��0;~�(;w�;�';�Y;�;d��:��:���:      �;��;;�z ;��$;G�);^/;
4;��8;<�<; $@;I�B;�D;��E;�F;�cG;��G;lH;z-H;]NH;�iH;�H;��H;��H;��H;��H;x�H;v�H;�H;��H;G�H;�H;�H;��H;��H;F�H;��H;@�H;��H;��H;�H;�H;J�H;��H;�H;v�H;t�H;��H;��H;��H;��H;�H;�iH;]NH;{-H;jH;��G;�cG;�F;��E;!�D;L�B;$@;:�<;��8;4;d/;C�);��$;�z ;�
;��;      ,�1;,J2;5g3;�$5;�Y7;��9;Qg<;�>;�A;xC;�D;�E;G�F;*G;'�G;1�G;�H;^5H;�RH;FlH;	�H;��H; �H;��H;^�H;?�H;3�H;	�H;��H;�H;`�H;��H;]�H;��H;��H;�H;I�H;��H;��H;��H;Z�H;��H;b�H;�H;��H;�H;/�H;?�H;a�H;��H;��H;��H;�H;FlH;�RH;X5H;�H;0�G;(�G;*G;G�F;	�E;�D;tC;�A; �>;Mg<;��9;�Y7;�$5;2g3;J2;      9,>;^Z>;��>;��?;H�@;��A;�C;�D;�E;��E;��F;�G;�}G;D�G;��G;�!H;B@H;\ZH;/qH;�H;.�H;��H;��H;��H;��H;��H;�H;��H;��H;��H;:�H;�H;�H;x�H;>�H;��H;��H;��H;;�H;x�H;~�H;�H;<�H;��H;��H;��H;�H;��H;��H;�H;��H;��H;.�H;�H;-qH;XZH;C@H;�!H;��G;@�G;�}G;�G;�F;��E;�E;�D;�C;��A;S�@;��?;��>;VZ>;      ��C;'	D;SBD;��D;�	E;��E;QF;�wF;��F;�<G;�G;��G;}�G;�H;c4H;�MH;dH;xH;��H;C�H;��H;��H;d�H;��H;$�H;��H;��H;P�H;V�H;��H;��H;X�H;x�H;0�H;��H;<�H;>�H;7�H;��H;2�H;t�H;S�H;��H;��H;R�H;M�H;��H;��H;%�H;��H;a�H;��H;��H;?�H;��H;xH;dH;�MH;e4H;�H;��G;��G;��G;�<G;��F;�wF;OF;��E;�	E;�D;QBD;%	D;      LwF;DF;~�F;��F;��F;�G;�NG;	�G;8�G;��G;��G;4H;l1H;�GH;s\H;\oH;��H;�H;��H;U�H;��H;��H;>�H;��H;��H;A�H;�H;�H;��H;y�H;�H;G�H;(�H;��H;e�H;��H;��H;��H;b�H;��H;&�H;C�H;�H;x�H;��H;�H;�H;E�H;��H;��H;;�H;��H;��H;S�H;��H;�H;��H;YoH;u\H;�GH;l1H;6H;��G;��G;;�G;�G;�NG;|G;��F;��F;{�F;FF;      �G;?�G;ڔG;�G; �G;
�G;��G;��G;lH;�$H;8H;MJH;�[H;FlH;�{H;K�H;N�H;�H;U�H;r�H;��H;x�H;6�H;%�H;��H;�H;��H;Z�H;A�H;��H;'�H;�H;��H;}�H;��H;��H;	�H;��H;��H;}�H;��H;�H;'�H;��H;;�H;U�H;��H;�H;��H;�H;4�H;z�H;��H;p�H;S�H;��H;L�H;K�H;�{H;BlH;�[H;PJH;8H;�$H;mH;��G;��G;�G;5�G;�G;۔G;*�G;      q H;�H;gH;zH;�H;A!H;-H;�9H;�FH;ATH;�aH;9oH;C|H;̈H;|�H;]�H;�H;�H;�H;�H;;�H;v�H;�H;��H;L�H;�H;X�H;P�H;��H;��H;��H;��H;o�H;��H;�H;W�H;[�H;S�H;�H;��H;l�H;��H;��H;��H;��H;N�H;T�H;�H;P�H;��H;�H;v�H;9�H;�H;�H;�H;�H;\�H;}�H;ʈH;E|H;9oH;�aH;?TH;�FH;�9H;-H;5!H;�H;wH;gH;�H;      �>H;}?H;BH;vFH;�KH;
SH;@[H;"dH;�mH;�wH;сH;׋H;��H;؞H;y�H;��H;�H;�H;�H;\�H;��H;�H;��H;��H;S�H;��H;:�H;��H;�H;��H;��H;d�H;��H;.�H;h�H;��H;��H;��H;f�H;/�H;��H;^�H;��H;��H;�H;��H;6�H;��H;V�H;��H;��H;�H;��H;X�H;�H;�H;�H;��H;x�H;֞H;��H;֋H;ՁH;�wH;�mH;&dH;>[H;SH;LH;rFH;BH;?H;      �hH;liH;hkH;pnH;�rH;�wH;�}H;S�H;k�H;˒H;9�H;��H;��H;��H;/�H;g�H;%�H;0�H;��H;��H;��H;��H;~�H;��H;��H;r�H;��H;��H;��H;��H;h�H;��H;�H;t�H;��H;��H;��H;��H;��H;t�H;�H;��H;h�H;��H;��H;��H;��H;x�H;��H;��H;�H;��H;��H;��H;��H;/�H;%�H;g�H;0�H;��H;��H;��H;:�H;ΒH;k�H;V�H;�}H;�wH;�rH;rnH;hkH;oiH;      1�H;ԈH;3�H;d�H;��H;K�H;��H;��H;��H;�H;��H;�H;a�H;��H;��H;@�H;n�H;G�H;��H;�H;��H;M�H;b�H;?�H;��H;	�H;)�H;��H;��H;p�H;��H;(�H;�H;��H;��H;��H;��H;��H;��H;��H;��H;&�H;��H;n�H;��H;��H;%�H;�H;��H;<�H;e�H;M�H;��H;�H;��H;F�H;p�H;A�H;��H;��H;c�H;�H;��H;�H;��H;��H;��H;@�H;��H;d�H;5�H;ֈH;      I�H;��H;��H;J�H;��H;P�H;��H;2�H;�H;!�H;K�H;q�H;��H;w�H;�H;��H;��H;��H;��H;�H;4�H;	�H;��H;�H;X�H;C�H;�H;��H;b�H;��H;#�H;v�H;��H;��H;��H;��H;�H;��H;��H;��H;��H;t�H; �H;��H;^�H;��H; �H;G�H;[�H;�H;��H;	�H;/�H;�H;��H;��H;��H;��H;�H;t�H;��H;r�H;O�H;!�H;�H;3�H;��H;P�H;��H;J�H;��H;��H;      �H;]�H;�H;M�H;�H;�H;��H;D�H;A�H;Z�H;o�H;��H;��H;��H;k�H;3�H;��H;�H;,�H;
�H;��H;"�H;^�H;�H;z�H;&�H;��H;u�H;��H;!�H;~�H;��H;��H;��H;�H;�H;��H;�H;�H;��H;��H;��H;{�H;�H;��H;o�H;��H;)�H;|�H;�H;a�H;!�H;��H;�H;,�H;�H;��H;6�H;l�H;��H;��H;��H;r�H;Z�H;D�H;D�H;��H;�H;
�H;F�H;�H;^�H;      �H;�H;��H;��H;��H;��H;��H;��H;��H;�H;��H;��H;h�H;��H;*�H;I�H;G�H;�H;��H;6�H;x�H;��H;��H;r�H;2�H;��H;z�H;��H;/�H;x�H;��H;��H;��H;��H;(�H;/�H;�H;/�H;%�H;��H;��H;��H;��H;t�H;+�H;��H;y�H;��H;4�H;q�H;��H;��H;o�H;/�H;��H;�H;L�H;K�H;+�H;��H;e�H;��H;��H;�H;��H;��H;��H;��H; �H;��H;��H;�H;      ��H;��H;L�H;�H;�H;B�H;��H;��H;d�H;m�H;b�H;t�H;u�H;T�H;-�H;��H;��H;�H;t�H;��H;��H;��H;�H;2�H;��H;^�H;��H;�H;j�H;��H;��H;��H;�H;)�H;�H;'�H;D�H;(�H;	�H;)�H;�H;��H;��H;��H;c�H;	�H;��H;`�H;��H;2�H;��H;��H;��H;��H;q�H;�H;��H;��H;,�H;R�H;s�H;t�H;d�H;n�H;h�H;��H;��H;B�H;�H;�H;M�H;��H;      �H;0�H;��H;.�H;�H;K�H;��H;,�H;��H;z�H;-�H;��H;��H;J�H;��H;m�H;��H;0�H;k�H;��H;��H;D�H;��H;��H;7�H;��H;��H;W�H;��H;��H;��H;��H;�H;3�H;)�H;�H;0�H;�H;(�H;6�H;�H;��H;��H;��H;��H;S�H;��H;��H;5�H;��H;�H;A�H;z�H;��H;j�H;2�H;��H;o�H;��H;L�H;��H;��H;/�H;{�H;��H;/�H;��H;L�H;!�H;+�H;��H;?�H;      q�H;��H;9�H;��H;��H;��H;��H;G�H;��H;R�H;�H;��H;P�H;�H;��H;��H;b�H;��H;��H;��H;��H;��H;I�H;��H;A�H;��H;�H;a�H;��H;��H;��H;�H;�H;�H;F�H;.�H; �H;0�H;C�H;�H;�H;�H;��H;��H;��H;\�H;�H;��H;>�H;��H;N�H;��H;��H;��H;��H;��H;b�H;��H;��H;�H;O�H;��H;�H;T�H;��H;I�H;��H;��H;��H;��H;:�H;��H;      �H;5�H;��H;.�H; �H;P�H;��H;+�H;��H;z�H;,�H;��H;��H;M�H;��H;m�H;��H;0�H;k�H;��H;��H;F�H;��H;��H;7�H;��H;��H;W�H;��H;��H;��H;��H;�H;5�H;,�H;�H;0�H;�H;(�H;5�H;�H;��H;��H;��H;��H;Q�H;��H;��H;5�H;��H;�H;?�H;z�H;��H;g�H;2�H;��H;n�H;��H;J�H;��H;��H;/�H;w�H;��H;0�H;��H;L�H;$�H;/�H;��H;<�H;      ��H;��H;E�H;�H;�H;>�H;��H;��H;d�H;n�H;b�H;t�H;s�H;T�H;.�H;��H;��H;�H;t�H;��H;��H;��H;�H;3�H;��H;]�H;��H;�H;j�H;��H;��H;��H;�H;)�H;�H;(�H;D�H;(�H;�H;)�H;�H;��H;��H;��H;c�H;�H;��H;`�H;��H;0�H;��H;��H;��H;��H;p�H;�H;��H;��H;*�H;R�H;s�H;u�H;a�H;m�H;e�H;��H;��H;;�H;�H;	�H;L�H;��H;      �H;�H;��H;��H;��H;��H;��H;��H;��H;�H;��H;��H;g�H;��H;-�H;I�H;J�H;�H;��H;5�H;x�H;��H;��H;t�H;4�H;��H;|�H;��H;1�H;w�H;��H;��H;��H;��H;(�H;.�H;�H;/�H;%�H;��H;��H;��H;��H;q�H;&�H;��H;w�H;��H;/�H;m�H;��H;��H;k�H;/�H;��H;�H;G�H;K�H;+�H;��H;e�H;��H;��H;�H;��H;��H;��H;��H; �H;��H;��H;�H;      �H;d�H;�H;H�H; �H;�H;��H;H�H;C�H;Z�H;p�H;��H;��H;��H;o�H;4�H;��H;�H;,�H;�H;��H;"�H;[�H;�H;|�H;"�H;��H;u�H;��H;!�H;{�H;��H;��H;��H;�H;�H;��H;�H;�H;��H;��H;��H;z�H;�H;��H;l�H;��H;&�H;x�H;{�H;a�H;�H;��H;�H;(�H;�H;��H;4�H;l�H;��H;��H;��H;p�H;W�H;A�H;E�H;��H;�H;�H;N�H; �H;]�H;      9�H;��H;��H;C�H;��H;`�H;��H;6�H;�H; �H;K�H;r�H;��H;u�H;�H;��H;��H;��H;��H;�H;6�H;�H;��H;�H;[�H;A�H;�H;��H;d�H;��H; �H;v�H;��H;��H;��H;��H;�H;��H;��H;��H;��H;t�H;�H;��H;[�H;��H;��H;D�H;W�H;�H;��H;�H;,�H;��H;��H;��H;��H;��H;�H;t�H;��H;r�H;M�H;!�H;�H;5�H;��H;S�H;��H;F�H;��H;��H;      %�H;ԈH;3�H;^�H;��H;I�H;��H;��H;��H;�H;��H;�H;a�H;��H;��H;A�H;p�H;G�H;��H;�H;��H;N�H;a�H;=�H;��H;�H;%�H;��H;��H;n�H;��H;(�H;��H;��H;��H;��H;��H;��H;��H;��H;��H;'�H;��H;i�H;��H;��H;"�H;	�H;��H;7�H;e�H;K�H;��H;�H;��H;C�H;n�H;@�H;��H;��H;a�H;�H;��H;�H;��H;��H;��H;E�H;��H;k�H;:�H;ԈH;      �hH;siH;akH;znH;�rH;�wH;�}H;[�H;o�H;ΒH;9�H;��H;��H;��H;3�H;h�H;%�H;2�H;��H;��H;��H;��H;{�H;��H;��H;q�H;��H;��H;��H;��H;i�H;��H;�H;t�H;��H;��H;��H;��H;��H;t�H;�H;��H;g�H;��H;��H;��H;��H;t�H;��H;��H;��H;��H;��H;��H;��H;,�H;"�H;g�H;0�H;��H;��H;��H;:�H;ΒH;m�H;Z�H;�}H;�wH;�rH;|nH;rkH;liH;      �>H;z?H;#BH;oFH;�KH;SH;;[H;%dH;�mH;�wH;сH;׋H;��H;؞H;|�H;��H;�H;�H;�H;Z�H;�H;�H;��H;��H;U�H;{�H;7�H;��H;�H;��H;��H;d�H;��H;.�H;h�H;��H;��H;��H;f�H;.�H;��H;a�H;��H;��H;�H;��H;4�H;�H;R�H;��H;��H;�H;��H;Z�H;�H;�H;�H;��H;y�H;֞H;��H;֋H;ҁH;�wH;�mH;'dH;A[H;	SH;LH;mFH;!BH;s?H;      { H;�H;]H;zH;�H;L!H;-H;�9H;�FH;?TH;�aH;7oH;C|H;͈H;~�H;\�H;�H;�H;�H;�H;;�H;w�H;�H;��H;O�H;�H;S�H;L�H;��H;��H;��H;��H;l�H;��H;�H;T�H;\�H;U�H;�H;��H;o�H;��H;��H;��H;��H;H�H;S�H;
�H;L�H;��H;�H;v�H;6�H; �H;�H;�H;�H;Z�H;~�H;ʈH;C|H;7oH;�aH;>TH;�FH;�9H;-H;9!H;�H;wH;hH;�H;      �G;E�G;ܔG;��G;.�G;�G;��G;��G;oH;�$H;8H;RJH;�[H;FlH;�{H;M�H;L�H;�H;S�H;p�H;��H;z�H;0�H;%�H;��H;�H;��H;W�H;@�H;��H;%�H;�H;��H;}�H;��H;��H;	�H;��H;��H;~�H;��H;�H;'�H;��H;:�H;T�H;��H;�H;��H; �H;9�H;z�H;��H;r�H;Q�H;��H;K�H;K�H;�{H;ClH;�[H;NJH;8H;�$H;lH;��G;��G;	�G;4�G;��G;�G;6�G;      AwF;AF;��F;��F;��F;�G;�NG;�G;?�G;��G;��G;9H;o1H;�GH;w\H;\oH;��H;�H;��H;T�H;��H;��H;:�H;��H;��H;>�H;�H;�H;��H;u�H;�H;G�H;&�H;��H;e�H;��H;��H;��H;b�H;��H;(�H;G�H;	�H;u�H;�H;
�H;�H;C�H;��H;��H;?�H;��H;��H;U�H;��H;�H;��H;ZoH;w\H;�GH;l1H;4H;��G;��G;5�G;�G;�NG;}G;��F;��F;m�F;1F;      ��C; 	D;NBD;�D;�	E;��E;QF;�wF;��F;�<G;��G;��G;�G;�H;h4H;�MH;dH;xH;��H;@�H;��H;��H;`�H;��H;%�H;��H;��H;M�H;V�H;��H;��H;X�H;u�H;2�H;��H;:�H;?�H;:�H;��H;3�H;x�H;X�H;��H;��H;P�H;H�H;��H;��H;$�H;��H;e�H;��H;��H;?�H;��H;xH;dH;�MH;h4H;�H;�G;��G;�G;�<G;��F;�wF;OF;��E;�	E;�D;PBD;!	D;      ,>;BZ>;��>;��?;B�@;��A;�C;�D;�E;��E;�F;�G;�}G;D�G;��G;�!H;B@H;]ZH;.qH;�H;/�H;��H;��H;��H;��H;��H;�H;��H;��H;��H;<�H;�H;�H;z�H;=�H;��H;��H;��H;;�H;x�H;��H;�H;?�H;��H;��H;��H;�H;��H;��H;��H;��H;��H;.�H;�H;.qH;XZH;B@H;�!H;��G;B�G;�}G;�G;�F;��E;�E;�D;�C;��A;Z�@;į?;��>;-Z>;      �1;$J2;'g3;�$5;|Y7;��9;Ig<;�>;�A;uC;
�D;	�E;G�F;*G;,�G;4�G;�H;^5H;�RH;HlH;�H;��H;��H;��H;a�H;8�H;/�H;	�H;��H;{�H;a�H;��H;[�H;��H;��H;�H;L�H;�H;��H;��H;^�H;��H;e�H;�H;��H;�H;3�H;<�H;]�H;��H;��H;��H;�H;HlH;�RH;W5H;�H;0�G;+�G;*G;G�F;�E;	�D;tC;�A;�>;Jg<;��9;|Y7;�$5;'g3;J2;      �;��;�
;�z ;��$;K�);d/;4;��8;8�<; $@;O�B;�D;��E;�F;�cG;��G;lH;z-H;]NH;�iH;�H;��H;��H;��H;��H;v�H;v�H;�H;��H;H�H;�H;�H;��H;��H;A�H;��H;D�H;��H;��H;�H;�H;K�H;��H;�H;s�H;x�H;��H;��H;��H;��H;�H;�iH;^NH;y-H;hH;��G;�cG;�F;��E;�D;I�B;�#@;8�<;��8;4;]/;4�);��$;�z ; ;��;      ��:��:��:r��:�;�Y;�';y�;��(;��0;�Y7;A�<;��@;�`C;CE;�wF;Z8G;_�G;A�G;W)H;�LH;�iH;�H;/�H;|�H;��H;��H;6�H;��H;��H;��H;-�H;��H;o�H;��H;x�H;��H;z�H;��H;k�H;��H;,�H;��H;��H;��H;4�H;��H;��H;x�H;/�H;�H;�iH;�LH;W)H;A�G;[�G;W8G;�wF;CE;�`C;��@;=�<;�Y7;��0;��(;|�;�';�Y;�;r��:#��:���:      ��:�:�2<:�)i:@t�:ه�:_�:�+�:�Y;+�;�*';w1;'�8;�Z>;:0B; �D;i2F;G;Y�G;��G;Y)H;^NH;IlH; �H;<�H;T�H;k�H;�H;Z�H;��H;�H;��H;�H;0�H;��H;��H;��H;��H;��H;,�H;�H;��H;�H;��H;Z�H;�H;p�H;U�H;8�H;#�H;IlH;\NH;X)H;��G;Y�G;	G;i2F;��D;80B;�Z>;$�8;s1;�*';)�;�Y;�+�:S�:Ň�:Ht�:j)i:�2<:Ġ:      ڥ��2X��� ����=�X۷�`ߤ8��:�P�:�P�:���:&`;n;�*;�$5;�g<;�<A;�BD;�F;�G;Y�G;C�G;z-H;�RH;-qH;��H;��H;N�H;�H;�H;��H;��H;��H;%�H;��H;r�H;h�H;��H;h�H;p�H;��H;%�H;��H;��H;��H;
�H;�H;P�H;��H;��H;/qH;�RH;w-H;C�G;Z�G;�G;�F;�BD;�<A;�g<;�$5;�*;j;$`;z��:�P�:�P�:��: ߤ8X۷���=�!��,X��      �1�� Ȅ�Ҩu��PV�g.�����W����XX�9+i:ࡼ:�+�:�;�t%;�J2;N;;��@;ZD;�F;G;X�G;hH;Z5H;XZH;xH;�H;��H;�H;�H;,�H;A�H;��H; �H;��H;�H;0�H;��H;2�H;�H;��H; �H;��H;C�H;2�H;�H;�H;��H;�H;xH;VZH;X5H;hH;W�G;	G;�F;YD;��@;H;;�J2;�t%;�;�+�:ࡼ:
+i:@X�9 ��W�����i.��PV�ڨu�"Ȅ�      X��K�	������!Tʻ�R��3|�f.�Ⱥ��� Y�9$u�:��:�Y;z�!;��0;ו:;��@;�BD;h2F;Z8G;��G;�H;C@H;�cH;��H;H�H;�H;�H; �H;g�H;��H;��H;B�H;��H;��H;Z�H;��H;��H;@�H;��H;��H;i�H;"�H;�H;�H;H�H;��H;�cH;@@H;�H;��G;W8G;j2F;�BD;��@;ו:;��0;x�!;�Y;��:u�:Y�9���Ⱥg.�3|��R��&Tʻ�����J�	�      ��x��[t���g�NT�]�:�������%����1��M�(�.W�� �t��n`:Z��:�\;{ ;��0;N;;�<A;��D;�wF;�cG;1�G;�!H;�MH;YoH;H�H;Y�H;��H;e�H;<�H;��H;/�H;G�H;��H;m�H;��H;k�H;��H;B�H;,�H;��H;<�H;e�H;��H;Y�H;G�H;UoH;�MH;�!H;1�G;�cG;�wF;��D;�<A;M;;��0; { ;�\;T��:�n`:��t�4W��O�(��1��&���������`�:�NT���g��[t�      5,˼��Ǽ�"���뮼w��#G��'�[�]y-�����.��ŕb�t0㺐ط�5<:�L�:�\;t�!;�J2;�g<;30B;CE;�F;+�G;��G;b4H;v\H;�{H;��H;{�H;0�H;��H;�H;i�H;'�H;&�H;��H;��H;��H;%�H;&�H;h�H;�H;��H;0�H;|�H;}�H;�{H;s\H;^4H;��G;(�G;�F;CE;40B;�g<;�J2;v�!;�\;�L�: 5<:�ط�x0�ƕb��.�����]y-�(�[�"G��w���뮼�"����Ǽ      )���k��Jv�|t�C�Ѽ�뮼+X��k�W������׻�Ǆ������5<:b��:�Y;�t%;�$5;�Z>;�`C;��E;*G;E�G;�H;�GH;ClH;ɈH;؞H;��H;��H;n�H;��H;��H;J�H;E�H;�H;H�H;H�H;��H;��H;k�H;��H;��H;ٞH;ǈH;AlH;�GH;�H;D�G;*G;��E;�`C;�Z>;�$5;�t%;�Y;T��:5<:�����Ǆ���׻���l�W�+X���뮼B�Ѽ}t�Jv���k�      Bm��Fi��&^�_�L�N�6�'����}ռmT����x���0���������hط��n`:��:�;�*; �8;��@;�D;H�F;�}G;�G;l1H;�[H;C|H;��H;��H;\�H;��H;��H;a�H;h�H;��H;E�H;��H;g�H;^�H;��H;��H;Z�H;��H;��H;B|H;�[H;i1H;y�G;�}G;H�F;�D;��@;$�8;�*;�;��:�n`:xط��������껾�0���x�mT��}ռ��'��P�6�_�L��&^��Fi�      K��r;��@�������섽w�e��?��k�zt�鷼G���e7�����Ǆ�j0� �t�u�:�+�:l;s1;H�<;K�B;�E;�G;��G;3H;NJH;3oH;֋H;��H;�H;k�H;��H;��H;i�H;��H;��H;��H;i�H;��H;��H;j�H;�H;��H;ًH;3oH;KJH;3H;��G;�G;	�E;K�B;@�<;t1;j;�+�: u�:@�t�l0� Ȅ���껃e7�G��鷼zt��k��?�v�e��섽���@���r;��      n���$��s��ӽ�'��?������
�Z��Q+�����"��G����0���׻Ǖb�6W���X�9ҡ�:`;�*';�Y7;�#@;	�D;��F;�G;��G;8H;�aH;ЁH;6�H;}�H;H�H;l�H;{�H;W�H;&�H;�H;&�H;X�H;y�H;i�H;F�H;z�H;9�H;ԁH;�aH;8H;��G;�G;�F;	�D;�#@;�Y7;�*';`;ҡ�:�X�98W��ɕb���׻��0�G���"������Q+�
�Z����?����'���ӽ�s�$��      �!,�7)��K ��������޽������Fi��0����鷼��x�����.��O�(�����*i:x��:(�;��0;8�<;tC;��E;�<G;��G;�$H;8TH;�wH;ʒH;�H; �H;X�H;�H;c�H;q�H;O�H;q�H;d�H;�H;U�H; �H;�H;˒H;�wH;:TH;�$H;��G;�<G;��E;uC;8�<;��0;+�;t��:�*i:���P�(��.�������x�鷼����0��Fi�������޽�������K �7)�      (�j��f��Z�y�F��>/��^�l�����ŽF ���Fi��Q+�zt�mT��m�W�����1��(ȺX�9wP�:�Y;��(;��8;�A;�E;��F;6�G;oH;�FH;�mH;m�H;��H;�H;H�H;��H;^�H;��H;��H;��H;`�H;��H;D�H;�H;��H;m�H;�mH;�FH;mH;9�G;��F;�E;�A;��8;~�(;�Y;uP�:X�9(Ⱥ�1�����m�W�mT��zt�Q+��Fi�F ����Žl����^��>/�y�F��Z��f�      ��v���x�H����f��SC��K �mn����Ž���
�Z��k�}ռ,X��`y-�*���m.����P�:�+�:��;4;�>;�D;�wF;��G;��G;�9H;%dH;S�H;��H;2�H;H�H;��H;~�H;+�H;E�H;)�H;�H;��H;E�H;/�H;��H;X�H;*dH;�9H;��G;�G;�wF;�D;�>;4;y�;�+�:�P�:p��l.�+���`y-�-X��}ռ�k�
�Z������Žmn���K ��SC��f�H���y�v���      ��˾��Ǿ�������U͓�Y�x���J��K �l���������?����뮼(�[����3|��W����:A�:�';a/;@g<;�C;DF;�NG;��G;-H;:[H;�}H;��H;��H;��H;��H;��H;��H;��H;��H;��H;�H;��H;��H;��H;�}H;>[H;-H;��G;�NG;DF;�C;Bg<;`/;�';I�:x�:�W��3|����(�[��뮼���?������l����K ���J�Z�x�U͓����������Ǿ      s� ��������{Ծj���v���Z�x��SC��^��޽?���w�e�'��B�Ѽ#G������R������ݤ8ɇ�:�Y;D�);��9;��A;��E;}G;	�G;>!H;SH;�wH;L�H;Z�H;�H;��H;I�H;V�H;��H;V�H;K�H;��H;�H;Z�H;H�H;�wH;SH;C!H;
�G;�G;��E;��A;��9;D�);�Y;χ�:�ݤ8����R�����#G��B�Ѽ'��w�e�?����޽�^��SC�Z�x�v���j����{Ծ�쾟���      ����D�l�s� �U�ݾj���U͓��f��>/�����'���섽N�6�~t�w��]�:�&Tʻ|.�8۷�Dt�:�;��$;�Y7;R�@;�	E;��F;&�G;�H;LH;�rH;��H;��H;��H;��H;�H;%�H;��H;!�H;�H;�H;��H;��H;��H;�rH;
LH;�H;+�G;��F;�	E;S�@;�Y7;��$;�;Ht�:@۷�x.�&Tʻ]�:�w��~t�O�6��섽�'������>/��f�V͓�j���V�ݾs� �l��D�      �7�v3�/�'����s� ��{Ծ���H���y�F�����ӽ���^�L�Jv��뮼PT����PV���=�^)i:v��:�z ;�$5;��?;�D;��F;�G;pH;bFH;pnH;d�H;J�H;G�H;��H;�H;/�H;��H;-�H;	�H;��H;J�H;M�H;`�H;znH;fFH;sH;�G;��F;�D;��?;{$5;�z ;t��:v)i:��=��PV���PT��뮼Jv�^�L�����ӽ���y�F�H�������{Ծs� ����/�'�v3�      �N��TI���;�/�'�l��쾀���y󐾴Z��K ��s�@����&^���"����g����Шu�� ���2<:��:�
;;g3;��>;WBD;u�F;۔G;iH;BH;ZkH;.�H;��H;�H;��H;>�H;��H;!�H;��H;A�H;��H;�H;��H;)�H;ckH;BH;nH;�G;��F;UBD;��>;4g3;�
;��:�2<:� ��Ψu������g��"����&^�@����s潥K ��Z�y󐾀�����l�/�'���;��TI�      `]�d�W��TI�v3��D�������Ǿv����f�7)�$��r;���Fi��k���Ǽ�[t�M�	�*Ȅ�X��Ԡ:��:��;.J2;TZ>;%	D;;F;7�G;�H;�?H;viH;H;��H;P�H;�H;��H;4�H;��H;1�H;��H;�H;P�H;��H;��H;}iH;�?H;�H;:�G;HF;$	D;PZ>;&J2;��;��:�:"X��)Ȅ�M�	��[t���Ǽ�k��Fi�r;��$��7)��f�v�����Ǿ�����D�v3��TI�d�W�      �?��|h��=v��� ��6�X��O/�0y�@�;ఖ��+X��� �ѽ����^n;�Z�������B(�ښ��X��`�e9�:�;�Y.;S�<;cWC;�ZF;��G;�/H;1jH;8�H;E�H;~�H;%�H;��H;V�H;��H;��H;��H;T�H;��H;%�H;�H;C�H;?�H;4jH;0H;��G;�ZF;eWC;P�<;�Y.;�;�:��e9^��ؚ���B(�����Z��^n;����� �ѽ���+X�ఖ�@�;0y��O/�6�X�� ��=v��|h��      |h��/���a�����y�VvS�pM+��v�9ɾ�����T� ]�\ν����x\8�����x��%�N���v��`�9n-�:g�;��.;�<;�nC;�dF;�G;�1H;�jH;��H;��H;ǵH;f�H;��H;a�H;��H;��H;��H;d�H;��H;d�H;ɵH;��H;��H;�jH;�1H;�G;�dF;�nC;�<;��.;f�;n-�:��9v��L���%��x�����x\8�����\ν ]��T�����9ɾ�v�pM+�VvS���y�a���/���      =v��b���W ��`�h�6E�W��i���{㼾}���nH�ӈ�x�ý�Ȅ��s/��o��#�����$J��*кX	�9Qg�:�l;$0;]=;زC;׀F;n�G;6H;mH;%�H;��H;|�H;��H;>�H;��H;�H;��H; �H;��H;=�H;��H;|�H;��H;,�H;mH;6H;n�G;�F;ٲC;]=;0;�l;Ug�:�	�90к#J������#���o��s/��Ȅ�x�ýӈ��nH�}��{㼾i���W��6E�`�h�W ��a���      � ����y�`�h���N��O/����B�߾B���*|��6�p}�䳽iSt�<�!�nrμ@F{��_��X��̓��D:(��:�Z;�2;�O>;lD;)�F;y�G;=H;�pH;��H;G�H;ȷH;��H;��H;[�H;z�H;\�H;v�H;[�H;��H;��H;ȷH;B�H;��H;�pH;=H;w�G;0�F;lD;�O>;�2;�Z;(��:`:Г���X���_�@F{�nrμ<�!�iSt�䳽p}��6��*|�B��B�߾����O/���N�`�h���y�      6�X�VvS�6E��O/��S�HW����������LS\��� ���9����Y�z��σ����]�����"�b���Y�D�Y:��:d`;9�4;�?;8�D;��F;	�G;FH;DuH;��H;��H;�H;�H;��H;�H;�H;��H;�H;�H;��H;�H;~�H;��H;œH;DuH;FH;�G;��F;9�D;�?;3�4;d`;��:P�Y:��Y�"�b�������]�΃��z���Y�9����彑� �LS\���������HW���S��O/�6E�VvS�      �O/�pM+�W�����HW��9ɾ@���Mw�� :�i��w�ý�L��[n;�\���rv���E<��˻��-�(��jy�:�^;�%;��7;u�@;5E;�"G;
�G;7PH;�zH;��H;W�H;x�H;��H;��H;	�H;��H;��H;��H;
�H;��H;��H;v�H;S�H;��H;�zH;7PH;�G;�"G;5E;q�@;~�7;�%;�^;ny�:0����-��˻�E<�rv��\���[n;��L��w�ýi��� :��Mw�@��9ɾHW�����X��pM+�      0y��v�i���B�߾����@��?����nH���B὜u����d�/O�hrμI"�����	�����Pr89];�:`�;�+;U|:;x7B;��E;�aG;qH;�ZH;c�H;*�H;��H;�H;F�H;B�H;�H;��H;t�H;��H;�H;B�H;C�H;�H;��H;.�H;e�H;�ZH;jH; bG;��E;u7B;Q|:;�+;]�;c;�:Pr89���	�����I"��hrμ/O���d��u��B����nH�?���@������B�߾i����v�      @�;9ɾ{㼾B�������Mw��nH�����Z�䳽ʕ��q\8�m#������^N�L���b��Hx�<5:��:0�;��0;]=;?�C;�[F;՞G;�)H;�eH;r�H;!�H;;�H;��H;�H;��H;'�H;��H;l�H;��H;*�H;��H;�H;~�H;9�H;'�H;r�H;�eH;�)H;֞G;�[F;9�C;]=;��0;,�;��:85:�Hx��b�K��^N�����m#��q\8�ʕ��䳽�Z񽰯��nH��Mw�����B��{㼾9ɾ      ఖ�����}���*|�LS\�� :����Z�k$������ �K�u���Oļ����������>&����C/�:�^;��#;�G6;9�?;��D;G�F;��G;@H;�pH;ޏH;t�H;�H;I�H;.�H;j�H;n�H;��H;x�H;��H;q�H;k�H;*�H;I�H;�H;u�H;ݏH;�pH; @H;��G;G�F;��D;<�?;�G6;��#;�^;C/�:���<&������������Oļu�� �K�����k$���Z���� :�LS\��*|�|������      �+X��T��nH��6��� �i��B�
䳽�����mR����ټ�����E<��?ݻ3d\������ :�d�:��;'�,;x�:;Y7B;��E;nLG;/H;ZSH;�{H;|�H;�H;�H;<�H;R�H;
�H;��H;��H;��H;��H;��H;�H;Q�H;9�H;�H;�H;�H;�{H;VSH;+H;oLG;��E;Z7B;y�:;$�,;��;�d�:� :����2d\��?ݻ�E<�����ټ����mR�����
䳽B�i���� ��6��nH��T�      �� ]�ӈ�p}���w�ý�u��ʕ�� �K�����o�hv���&R���T^��x�� �>����:]B;:";f�4;��>;AD;��F;�G;�)H;fdH;q�H;�H;_�H;&�H;+�H;��H;��H;�H;�H;��H;�H;�H;��H;~�H;*�H;(�H;b�H;
�H;q�H;ddH;�)H;�G;��F;BD;��>;f�4;C";_B;���: �>�z��S^�����&R�hv���o���� �K�ʕ���u��w�ý��p}�ӈ�]�       �ѽ\νx�ý䳽9����L����d�p\8�u��ټhv����Y��_� ���;���[���Y:W��:Im;�r-;
�:;n�A;,oE;�"G;J�G;XGH;�sH;�H;��H;�H;#�H;�H;��H;v�H;~�H;'�H;��H;'�H;~�H;{�H;��H;�H;&�H;�H;��H;�H;�sH;WGH;K�G;�"G;2oE;n�A;�:;�r-;Mm;]��:��Y:�[�8�������_���Y�gv��ټu��p\8���d��L��9���䳽x�ý\ν      ���������Ȅ�iSt��Y�[n;�.O�l#���Oļ�����&R��_������N3�ԅY��3:��:կ;�?&;�G6;~X?;�D;$xF;��G;,!H;�^H;��H;�H;íH;<�H;��H;��H;��H;	�H;��H;P�H;�H;P�H;��H;	�H;��H;��H;�H;E�H;ǭH;�H;��H;�^H;0!H;��G;'xF;�D;X?;�G6;�?&;ӯ;	�: 4:ȅY��N3������_��&R������Oļl#��/O�[n;��Y�iSt��Ȅ�����      \n;�w\8��s/�<�!�y��^���grμ��������E<�������N3�DHx���9��:�^;R ;)2;a�<;�B;��E;$5G;�G;'FH;{qH;��H;>�H;��H;F�H;��H;��H;��H;��H;�H;n�H;�H;n�H;�H;��H;��H;��H;��H;N�H;��H;A�H;��H;uqH;+FH; �G;)5G;��E;�B;i�<;-2;R ;�^;��:��98Hx��N3� ������E<��������hrμ\���z��<�!��s/�w\8�      X������o�nrμ΃��rv��H"��	^N�����?ݻS^��?��܅Y���9��:ڦ�:��;O�.;{|:;�>A;��D;%�F;��G;�)H;aH;�H;u�H;۬H;,�H;�H;/�H;W�H;��H;�H;O�H;��H;��H;��H;N�H;�H;��H;V�H;0�H;�H;0�H;ެH;t�H;�H;aH;�)H;��G;&�F;��D;�>A;|:;K�.;��;ڦ�:��:��9ЅY�;��R^���?ݻ���
^N�H"��pv��σ��nrμ�o����      �����x���#��=F{���]��E<����G�뻨���.d\�v�뺴[��3:��:ަ�:z[;a�,;��8;!@;�0D;p[F;{G;�
H;;PH;vH;ڐH;5�H;�H;�H;]�H;q�H;��H;��H;t�H;o�H;��H;��H;��H;k�H;s�H;��H;��H;s�H;b�H;!�H;�H;6�H;ӐH;vH;;PH;�
H;{G;s[F;�0D;!@;��8;h�,;z[;��:��:�3:�[�p��-d\�����F�뻠���E<���]�>F{��#���x��      �B(� %�����_�����˻ 	����b�7&����� |>���Y:�:�^;��;f�,;`8;a�?;��C;mF;�FG;@�G;�?H;kH;�H;��H;�H;L�H;��H;b�H;k�H;�H;u�H;��H;��H;}�H;��H;x�H;~�H;��H;p�H;�H;n�H;b�H;��H;M�H;�H;��H;��H;kH;�?H;B�G;�FG;uF;��C;[�?;`8;f�,;��;�^;�:��Y: p>�����3&���b�	���˻�����_�����%�      ʚ��F���"J���X���b���-�����Hx����!:���:O��:ί;P ;K�.;��8;U�?;��C;��E;+#G;��G;�1H;�aH;@�H;j�H;m�H;��H;��H;R�H;�H;(�H;0�H;��H;�H;��H;3�H;��H;0�H;~�H;�H;��H;-�H;*�H;�H;S�H;��H;��H;h�H;o�H;>�H;�aH;�1H;��G;0#G;��E;��C;Z�?;��8;M�.;P ;ϯ;U��:��:!:����Hx������-��b��X��J��G���       �����(к������Y���� s89T5:M/�:�d�:eB;Im;�?&;-2;|:;!@;��C;��E;pG;��G;L(H;�ZH;`zH;/�H;ǤH;��H;Z�H;��H;��H;T�H;��H;��H;B�H;$�H;C�H;��H;u�H;��H;@�H;!�H;@�H;��H;��H;X�H;��H;��H;Y�H;��H;ͤH;0�H;]zH;�ZH;O(H;��G;rG;��E;��C;!@;�|:;-2;�?&;Jm;hB;�d�:Q/�:X5:�r89�����Y�Г��(к���      `�e9h�9�	�9�:@�Y:py�:w;�:��:�^;��;C";�r-;�G6;f�<;�>A;�0D;sF;5#G;��G;�$H;RWH;�vH;i�H;4�H;5�H;n�H;�H;��H;o�H;.�H;��H;w�H;��H;!�H;�H;��H;��H;��H;�H; �H;��H;u�H;��H;.�H;n�H;��H;�H;l�H;;�H;5�H;f�H;�vH;VWH;�$H;��G;1#G;sF;�0D;�>A;d�<;�G6;�r-;E";��;�^;��:q;�:|y�:X�Y:\:h	�9�9      U�:X-�:#g�:��:��:�^;^�;*�;��#;&�,;c�4;�:;}X?;�B;��D;u[F;�FG;��G;O(H;PWH;\uH;~�H;�H;�H;�H;��H;��H;��H;��H;��H;��H;��H;��H;��H;��H;Q�H;L�H;J�H;��H;��H;��H;��H;��H;��H;��H;��H;��H;��H;�H;�H;�H;��H;`uH;RWH;Q(H;��G;�FG;s[F;��D;�B;X?;�:;j�4;&�,;��#;)�;d�;�^;��:��:?g�:T-�:      �;u�;�l;[;d`;�%;�+;��0;�G6;|�:;��>;m�A;�D;��E;&�F;{G;D�G;�1H;�ZH;�vH;��H;?�H;��H;øH;|�H;K�H;��H;��H;��H;��H;2�H;2�H;��H;��H;d�H;��H;��H;��H;a�H;��H;��H;.�H;4�H;��H;��H;��H;��H;J�H;�H;¸H;��H;@�H;��H;�vH;�ZH;�1H;G�G;{G;'�F;��E;�D;n�A;��>;z�:;�G6;��0;�+;�%;x`;�Z;�l;k�;      �Y.;��.;0;�2;2�4;��7;c|:;&]=;?�?;]7B;ED;/oE;'xF;25G;��G;�
H;�?H;�aH;azH;g�H;
�H;��H;B�H;��H;[�H;��H;��H;��H;�H;��H;��H;V�H;P�H;?�H;��H;�H;?�H;�H;��H;?�H;L�H;T�H;��H;��H;�H;��H;��H;��H;_�H;��H;<�H;��H;�H;i�H;dzH;�aH;�?H;�
H;��G;.5G;)xF;2oE;HD;Y7B;E�?;)]=;_|:;��7;A�4;�2;0;��.;      V�<;)�<;]=;�O>;�?;{�@;|7B;?�C;�D;��E;��F;�"G;��G;�G;�)H;APH; kH;G�H;0�H;4�H;�H;��H;��H;2�H;)�H;,�H;>�H;��H;�H;4�H;��H;�H;�H;��H;=�H;z�H;��H;s�H;;�H;��H; �H;�H;��H;1�H;�H;��H;:�H;.�H;,�H;-�H;��H;¸H;�H;2�H;0�H;A�H;!kH;?PH;�)H;��G;��G;�"G;��F;��E;��D;D�C;x7B;h�@;�?;�O>;]=; �<;      �WC;�nC;ղC;hD;8�D;$5E;��E;�[F;H�F;rLG;��G;P�G;0!H;2FH;aH;vH;��H;x�H;פH;B�H;�H;��H;c�H;6�H;��H;��H;:�H;��H;��H;��H;��H;��H;��H;.�H;��H;��H;��H;��H;��H;.�H;��H;��H;��H;��H;��H;��H;6�H;��H;��H;2�H;a�H;��H;�H;>�H;֤H;u�H;��H;vH;aH;0FH;1!H;T�G;��G;rLG;L�F;�[F;��E;5E;B�D;lD;ӲC;�nC;      �ZF;�dF;�F;)�F;��F;�"G;bG;ߞG;��G;2H;�)H;[GH;�^H;qH;�H;ݐH;��H;o�H;��H;l�H;��H;G�H;��H;3�H;��H;�H;��H;��H;f�H;��H;��H;��H;�H;q�H;��H;�H;�H;�H;��H;q�H;�H;��H;��H;��H;c�H;��H;��H;!�H;��H;.�H;��H;J�H;��H;l�H;��H;l�H;��H;ސH;�H;|qH;�^H;\GH;�)H;2H;��G;�G;bG;�"G;��F;4�F;ހF;�dF;      �G;�G;k�G;~�G;�G;	�G;zH;�)H;�?H;YSH;fdH;�sH;��H;��H;r�H;8�H;�H;��H;^�H;�H;��H;��H;��H;E�H;9�H;��H;��H;<�H;|�H;��H;]�H;��H;m�H;��H;��H;3�H;N�H;,�H;��H;��H;l�H;��H;[�H;��H;x�H;8�H;�H;��H;;�H;?�H;��H;��H;��H;�H;]�H;��H;�H;8�H;q�H;��H;��H;�sH;gdH;WSH; @H;�)H;tH;�G;�G;v�G;m�G;ݪG;      0H;�1H;6H;=H;�EH;8PH;�ZH;�eH;�pH;�{H;q�H;�H;�H;C�H;جH;��H;L�H;��H;��H;��H;��H;��H;��H;��H;��H;��H;8�H;t�H;Z�H;I�H;��H;a�H;��H;�H;?�H;T�H;?�H;O�H;=�H;�H;��H;[�H;��H;H�H;W�H;q�H;5�H;��H;��H;��H;��H;��H;��H;��H;��H;��H;L�H;��H;جH;A�H;�H;�H;u�H;�{H;�pH;�eH;�ZH;-PH;FH;=H;6H;�1H;      -jH;�jH;mH;�pH;6uH;�zH;j�H;o�H;ԏH;|�H;	�H;��H;ǭH;��H;,�H;#�H;��H;Y�H;��H;r�H;��H;��H;�H;�H;��H;e�H;x�H;\�H;Q�H;��H;L�H;��H;��H;/�H;_�H;f�H;V�H;`�H;[�H;0�H;��H;��H;M�H;��H;M�H;Y�H;q�H;e�H;��H;�H;�H;��H;��H;o�H;��H;V�H;��H;$�H;,�H;��H;ǭH;��H;�H;��H;ُH;r�H;h�H;�zH;DuH;�pH;mH;�jH;      8�H;��H;2�H;��H;œH;��H;-�H;!�H;t�H;�H;a�H;�H;A�H;N�H;�H;_�H;g�H;�H;S�H;.�H;��H;��H;��H;4�H;��H;��H;��H;H�H;��H;B�H;��H;��H;/�H;X�H;c�H;x�H;��H;w�H;`�H;V�H;+�H;��H;��H;?�H;��H;H�H;}�H;��H;��H;0�H;��H;��H;��H;-�H;S�H;�H;d�H;b�H;�H;L�H;B�H;�H;c�H;�H;t�H;&�H;0�H;��H;ƓH;��H;2�H;��H;      L�H;��H;��H;K�H;��H;W�H;��H;=�H;�H;�H;-�H;,�H;�H;��H;3�H;w�H;u�H;0�H;��H;��H;��H;7�H;��H;��H;��H;��H;]�H;��H;Q�H;��H;��H;"�H;Y�H;g�H;��H;�H;z�H;|�H;~�H;i�H;X�H;!�H;��H;��H;L�H;��H;X�H;��H;��H;��H;��H;6�H;��H;��H;��H;/�H;u�H;x�H;5�H;��H;�H;-�H;-�H;�H;�H;A�H;��H;M�H;��H;I�H;��H;��H;      ��H;ѵH;~�H;ȷH;}�H;o�H;�H;��H;O�H;:�H;-�H;�H;��H;��H;W�H;��H;�H;4�H;��H;|�H;��H;5�H;X�H;�H;��H;��H;��H;b�H;��H;��H;�H;:�H;c�H;�H;��H;��H;��H;��H;��H;��H;c�H;9�H;�H;��H;��H;_�H;��H;��H;��H;�H;Y�H;5�H;��H;z�H;��H;6�H;�H;��H;W�H;��H;��H;�H;1�H;<�H;O�H;��H;��H;o�H;��H;ɷH;��H;εH;      .�H;q�H;	�H;��H;�H;��H;F�H;�H;'�H;R�H;��H;��H;��H;��H;��H;��H;y�H;��H;I�H;��H;��H;��H;P�H;�H;��H;�H;p�H;��H;��H;2�H;U�H;d�H;x�H;��H;��H;��H;��H;��H;��H;��H;u�H;d�H;T�H;.�H;��H;��H;l�H;�H;��H;�H;S�H;��H;��H;��H;I�H;��H;|�H;��H;��H;��H;��H;��H;��H;T�H;,�H;�H;F�H;|�H;�H;��H;�H;r�H;      ��H;��H;>�H;��H;��H;��H;H�H;��H;m�H;�H;��H;}�H;�H;��H;�H;w�H;��H;�H;(�H;(�H;��H;��H;>�H;��H;+�H;p�H;��H;�H;/�H;Y�H;b�H;��H;��H;��H;��H;��H;��H;��H;��H;��H;��H;��H;b�H;V�H;+�H;�H;��H;q�H;.�H;��H;C�H;��H;��H;!�H;'�H;�H;��H;x�H;�H;��H;�H;}�H;��H;�H;p�H;��H;L�H;��H;��H;��H;G�H;��H;      P�H;u�H;��H;b�H;+�H;�H;�H;+�H;t�H;��H;#�H;��H;��H;�H;U�H;q�H;��H;��H;C�H;	�H;��H;b�H;��H;4�H;��H;��H;��H;?�H;`�H;f�H;z�H;��H;��H;��H;��H;��H;��H;��H;��H;��H;��H;��H;x�H;`�H;Y�H;:�H;��H;��H;��H;4�H;��H;a�H;��H;�H;C�H;��H;��H;u�H;V�H;�H;��H;��H;&�H;��H;x�H;.�H;�H;�H;+�H;c�H;��H;v�H;      ��H;��H;�H;w�H;�H;��H;��H;��H;��H;��H;�H;*�H;P�H;q�H;��H;��H;}�H;0�H;��H;��H;T�H;��H;�H;l�H;��H;	�H;/�H;T�H;j�H;~�H;|�H;��H;��H;��H;��H;��H;��H;��H;��H;��H;��H;��H;{�H;x�H;d�H;O�H;.�H;�H;��H;m�H;�H;��H;O�H;��H;��H;6�H;��H;��H;��H;r�H;Q�H;)�H;�H;��H;��H;��H;��H;��H;�H;v�H;�H;��H;      ��H;��H;��H;^�H;��H;��H;y�H;l�H;{�H;��H;��H;��H;�H;�H;��H;��H;��H;��H;y�H;��H;V�H;��H;B�H;��H;��H;�H;M�H;G�H;]�H;��H;u�H;��H;��H;��H;��H;��H;��H;��H;��H;��H;��H;��H;u�H;��H;V�H;A�H;K�H;	�H;��H;��H;D�H;��H;O�H;��H;y�H;��H;��H;��H;��H;�H;�H;��H;��H;��H;~�H;p�H;�H;��H;��H;_�H;��H;��H;      ��H;��H;��H;y�H;�H;��H;��H;��H;��H;��H;�H;*�H;S�H;t�H;��H;��H;~�H;2�H;��H;��H;V�H;��H;�H;l�H;��H;�H;/�H;T�H;k�H;|�H;|�H;��H;��H;��H;��H;��H;��H;��H;��H;��H;��H;��H;{�H;w�H;d�H;N�H;,�H;�H;��H;l�H;�H;��H;O�H;��H;��H;6�H;�H;��H;��H;q�H;S�H;)�H;�H;��H;��H;��H;��H;��H;�H;z�H;�H;��H;      F�H;w�H;��H;[�H;)�H;��H;�H;.�H;t�H;��H;#�H;��H;��H;�H;V�H;r�H;��H;��H;C�H;	�H;��H;d�H;��H;4�H;��H;��H;��H;?�H;_�H;d�H;x�H;��H;��H;��H;��H;��H;��H;��H;��H;��H;��H;��H;x�H;_�H;Y�H;7�H;��H;��H;��H;2�H;��H;b�H;��H;�H;C�H;��H;��H;u�H;U�H;�H;��H;��H;#�H;��H;u�H;2�H;�H;��H;/�H;\�H;��H;y�H;      ��H;��H;;�H;��H;��H;��H;E�H;��H;n�H;�H;��H;}�H;�H;��H;�H;x�H;��H;�H;(�H;'�H;��H;��H;>�H;��H;/�H;o�H;��H;�H;/�H;Y�H;b�H;��H;��H;��H;��H;��H;��H;��H;��H;��H;��H;��H;`�H;V�H;(�H;�H;��H;q�H;-�H;��H;C�H;��H;��H;"�H;(�H;�H;��H;{�H;�H;��H;�H;}�H;��H;�H;q�H;��H;N�H;��H;��H;��H;D�H;��H;      .�H;x�H;�H;��H;�H;��H;C�H;�H;)�H;R�H;��H;��H;��H;��H;��H;��H;|�H;��H;H�H;��H;��H;��H;N�H;�H;��H;�H;o�H;��H;��H;2�H;T�H;b�H;w�H;��H;��H;��H;��H;��H;��H;��H;u�H;d�H;T�H;,�H;��H;��H;l�H;�H;��H;��H;U�H;��H;��H;��H;G�H;��H;z�H;��H;��H;��H;��H;��H;��H;Q�H;*�H;�H;L�H;~�H;�H;��H;�H;p�H;      v�H;ҵH;p�H;��H;z�H;}�H;��H;��H;N�H;:�H;.�H;�H;��H;��H;Z�H;��H;�H;6�H;��H;|�H;��H;8�H;U�H;�H;��H;��H;��H;b�H;��H;��H;�H;9�H;d�H;~�H;��H;��H;��H;��H;��H;�H;c�H;9�H;�H;��H;��H;\�H;��H;��H;��H; �H;[�H;5�H;��H;x�H;��H;3�H;�H;��H;X�H;��H;��H;�H;-�H;=�H;P�H;��H;��H;q�H;~�H;ķH;u�H;͵H;      ?�H;��H;��H;D�H;��H;V�H;��H;>�H;�H;�H;,�H;/�H;�H;��H;5�H;x�H;v�H;0�H;��H;��H;��H;9�H;��H;��H;��H;��H;X�H;��H;Q�H;��H;��H;"�H;Y�H;g�H;��H;~�H;z�H;�H;~�H;i�H;[�H;"�H;��H;��H;J�H;��H;W�H;��H;��H;��H;��H;7�H;��H;��H;��H;/�H;v�H;x�H;6�H;��H;�H;-�H;,�H;�H;�H;B�H;��H;S�H;��H;O�H;��H;��H;      H�H;��H;,�H;��H;��H;ƗH;,�H;*�H;w�H;�H;a�H;�H;C�H;M�H;�H;b�H;g�H;�H;T�H;0�H;��H;��H;��H;1�H;��H;��H;��H;I�H;��H;B�H;��H;��H;)�H;X�H;c�H;w�H;��H;x�H;`�H;X�H;,�H;��H;��H;?�H;��H;E�H;}�H;��H;��H;-�H;��H;��H;��H;,�H;T�H;�H;d�H;`�H;�H;L�H;A�H;�H;a�H;�H;t�H;(�H;.�H;��H;ȓH;��H;=�H;��H;      ;jH;�jH;,mH;�pH;.uH; {H;f�H;r�H;ޏH;{�H;�H;��H;ɭH;��H;0�H;$�H;��H;Z�H;��H;q�H;��H;��H;�H;�H;��H;_�H;r�H;Z�H;Q�H;��H;L�H;��H;��H;/�H;]�H;d�H;V�H;c�H;[�H;.�H;��H;��H;M�H;��H;L�H;U�H;r�H;c�H;��H;�H;�H;��H;��H;o�H;��H;V�H;��H;$�H;/�H;��H;ƭH;��H;�H;{�H;ޏH;s�H;i�H;�zH;>uH;�pH;,mH;�jH;      0H;�1H;6H;=H;�EH;EPH;�ZH;�eH;�pH;�{H;t�H;�H;�H;C�H;۬H;��H;M�H;��H;��H;��H;��H;��H;��H;��H;��H;��H;5�H;r�H;\�H;E�H;��H;a�H;��H;�H;=�H;Q�H;@�H;R�H;<�H;�H;��H;^�H;��H;F�H;V�H;n�H;4�H;��H;��H;��H;��H;��H;��H;�H;��H;��H;M�H;��H;ڬH;?�H;�H;�H;t�H;�{H;�pH;�eH;�ZH;1PH;FH;=H;6H;�1H;      �G;��G;m�G;��G;�G;�G;zH;�)H;@H;YSH;gdH;�sH;��H;��H;t�H;;�H;�H;��H;]�H;�H;��H;��H;��H;E�H;:�H;��H;�H;9�H;|�H;��H;Z�H;��H;m�H;��H;��H;/�H;N�H;/�H;��H;��H;o�H;��H;[�H;��H;x�H;6�H;}�H;��H;9�H;?�H;��H;��H;��H;�H;]�H;��H;�H;9�H;t�H;��H;�H;�sH;ddH;VSH;�?H;�)H;|H;
�G;�G;��G;q�G;�G;      �ZF;�dF;�F;%�F;��F;�"G;�aG;�G;��G;5H;�)H;`GH;�^H;}qH;�H;ߐH;��H;q�H;��H;n�H;��H;H�H;��H;1�H;��H;�H;��H;��H;h�H;��H;��H;��H;�H;q�H;��H;�H;�H;�H;��H;q�H;�H;��H;��H;��H;b�H;��H;��H;�H;��H;.�H;��H;G�H;��H;k�H;��H;j�H;��H;ސH;�H;yqH;�^H;XGH;�)H;2H;��G;ܞG;�aG;�"G;��F;'�F;ЀF;�dF;      �WC;�nC;ҲC;iD;4�D;(5E;��E;�[F;O�F;tLG;��G;T�G;1!H;1FH;aH;vH;��H;y�H;פH;?�H;�H;��H;_�H;4�H;��H;��H;6�H;��H;��H;��H;��H;��H;��H;.�H;��H;��H;��H;��H;��H;/�H;��H;��H;��H;��H;��H;��H;9�H;��H;��H;2�H;c�H;��H;�H;?�H;פH;t�H;��H;vH;aH;.FH;0!H;N�G;��G;qLG;I�F;�[F;��E;5E;?�D;hD;ҲC;�nC;      7�<;�<;]=;�O>;݁?;��@;|7B;A�C;��D;��E;��F;�"G;��G;�G;�)H;BPH;!kH;H�H;0�H;2�H;�H;��H;��H;/�H;,�H;'�H;:�H;��H;�H;1�H;��H;
�H;�H;��H;<�H;w�H;��H;x�H;;�H;��H;�H;	�H;��H;3�H;�H;��H;>�H;-�H;*�H;1�H;��H;��H;�H;4�H;2�H;A�H;!kH;?PH;�)H;�G;��G;�"G;��F;��E;��D;9�C;x7B;v�@;�?;�O>;]=;��<;      �Y.;��.;0;�2;.�4;��7;\|:;(]=;E�?;\7B;BD;3oE;)xF;05G;��G;�
H;�?H;�aH;czH;g�H;�H;��H;<�H;��H;_�H;��H;��H;��H;�H;��H;��H;V�H;N�H;?�H;��H;�H;B�H;�H;��H;<�H;O�H;V�H;��H;��H;�H;��H;��H;��H;\�H;��H;A�H;��H;�H;i�H;czH;�aH;�?H;�
H;��G;,5G;'xF;/oE;BD;Z7B;B�?;(]=;[|:;��7;.�4;�2;0;��.;      �;t�;�l;�Z;``;�%;�+;��0;�G6;z�:;��>;s�A;�D;��E;*�F;{G;F�G;�1H;�ZH;�vH;��H;@�H;��H;¸H;��H;F�H;��H;��H;��H;��H;3�H;2�H;��H;��H;a�H;��H;��H;��H;a�H;��H;��H;2�H;6�H;��H;��H;��H;��H;J�H;~�H;ŸH;��H;@�H;��H;�vH;�ZH;�1H;D�G;{G;'�F;��E;�D;l�A;��>;y�:;�G6;��0;�+;�%;x`;�Z;�l;g�;      G�:�-�:Gg�:&��:��:�^;`�;-�;��#;$�,;i�4;�:;X?;�B;��D;v[F;�FG;��G;O(H;PWH;]uH;��H;	�H;�H;�H;��H;��H;��H;��H;��H;��H;��H;��H;��H;��H;M�H;M�H;O�H;��H;��H;��H;��H;��H;��H;��H;��H;��H;��H;�H;�H;
�H;~�H;_uH;SWH;O(H;��G;�FG;r[F;��D;�B;~X?;�:;g�4;$�,;��#;.�;b�;�^;��:,��:[g�:X-�:      �e9��9�	�9�:@�Y:|y�:};�:���:�^;��;G";�r-;�G6;f�<;�>A;�0D;sF;4#G;��G;�$H;VWH;�vH;g�H;4�H;;�H;k�H;��H;��H;n�H;*�H;��H;w�H;��H;"�H;�H;��H;��H;��H;�H;�H;��H;w�H;��H;,�H;o�H;�H;�H;n�H;7�H;8�H;j�H;�vH;UWH;�$H;��G;0#G;pF;�0D;�>A;a�<;�G6;�r-;D";��;�^;��:o;�:jy�:X�Y:`:�	�9X�9       �����(к������Y�����r89X5:U/�:�d�:fB;Jm;�?&;-2;�|:;!@;��C;��E;pG;��G;O(H;�ZH;azH;/�H;ͤH;��H;V�H;��H;��H;S�H;��H;��H;A�H;$�H;D�H;��H;u�H;��H;C�H;#�H;A�H;��H;��H;W�H;��H;��H;Z�H;��H;ɤH;2�H;azH;�ZH;N(H;��G;oG;��E;��C;!@;�|:;)2;�?&;Hm;dB;�d�:O/�:T5:�r89�����Y�����6к���      Қ��B���$J���X���b���-�����Hx�`��!:��:U��:ѯ;P ;O�.;��8;X�?;��C;��E;-#G;��G;�1H;�aH;@�H;o�H;j�H;��H;��H;U�H;�H;)�H;-�H;��H;�H;�H;2�H;��H;3�H;}�H;�H;��H;-�H;*�H;�H;S�H;��H;��H;j�H;j�H;@�H;�aH;�1H;��G;.#G;��E;��C;W�?;��8;O�.;K ;ί;O��:��:� :����Hx������-��b��X��(J��D���      �B(�%�����_�����˻	����b�6&����� t>���Y:	�:�^;��;i�,;`8;^�?;��C;pF;�FG;B�G;�?H;kH;��H;��H;�H;I�H;��H;]�H;l�H;�H;s�H;��H;��H;{�H;��H;{�H;~�H;��H;r�H;�H;n�H;b�H;��H;I�H;�H;��H;�H;kH;�?H;@�G;�FG;tF;��C;[�?;
`8;f�,;��;�^;�:��Y: |>�����3&���b�	���˻�����_���� %�      �����x���#��>F{���]��E<����F�뻦���.d\�p�뺠[��3:��:��:}[;b�,;��8;!@;�0D;u[F;{G;�
H;>PH;vH;ڐH;4�H;�H; �H;\�H;q�H;��H;��H;t�H;o�H;��H;��H;��H;m�H;s�H;��H;��H;s�H;`�H; �H;�H;2�H;אH;vH;;PH;�
H;{G;o[F;�0D;!@;��8;d�,;y[;��:��:�3:�[�t��0d\�����G�뻢���E<���]�>F{��#���x��      X������o�nrμ΃��qv��H"��	^N�����?ݻR^��=��ЅY���9��:��:��;M�.;||:;�>A;��D;%�F;��G;�)H;aH;	�H;p�H;۬H;/�H;�H;2�H;W�H;��H;�H;O�H;��H;��H;��H;O�H;�H;��H;T�H;0�H;�H;2�H;۬H;p�H;�H;aH;�)H;��G;&�F;��D;�>A;{|:;K�.;��;ئ�:��:��9܅Y�>��S^���?ݻ���	^N�H"��qv��σ��orμ�o����      ]n;�w\8��s/�<�!�y��]���hrμ��������E<��� ����N3�<Hx���9��:�^;Q ;*2;b�<;��B;��E;(5G;�G;-FH;{qH;��H;>�H;��H;G�H;��H;��H;��H;��H;�H;m�H;�H;p�H;�H;��H;��H;��H;��H;M�H;��H;A�H;��H;vqH;'FH;�G;,5G;��E;�B;h�<;'2;Q ;�^;��:��9@Hx��N3� ������E<��������hrμ\���z��<�!��s/�w\8�      ���������Ȅ�iSt��Y�[n;�.O�l#���Oļ�����&R��_������N3���Y� 4:�:ү;�?&;�G6;�X?;�D;)xF;��G;0!H;�^H;��H;�H;ƭH;?�H;�H;��H;��H;�H;��H;P�H;�H;P�H;��H;	�H;��H;��H; �H;B�H;ɭH;�H;��H;�^H;,!H;��G;)xF;�D;{X?;�G6;�?&;ѯ;�:�3:ąY��N3������_��&R������Oļl#��/O�[n;��Y�iSt��Ȅ�����       �ѽ\νx�ý䳽9����L����d�p\8�u��ټgv����Y��_� ���8���[���Y:K��:Jm;�r-;�:;m�A;0oE;�"G;M�G;XGH;�sH;�H;��H;�H;(�H;�H;��H;y�H;~�H;&�H;��H;'�H;|�H;x�H;��H;�H;%�H;�H;��H;�H;�sH;XGH;I�G;�"G;2oE;n�A;�:;�r-;Hm;U��:��Y:�[�8������_���Y�hv��ټu��p\8���d��L��:���䳽x�ý\ν      ��]�ӈ�p}���w�ý�u��ʕ�� �K�����o�hv���&R���S^��x�� �>����:[B;>";j�4;��>;ED;��F;�G;�)H;adH;p�H;�H;a�H;)�H;-�H;��H;��H;�H;�H;��H;�H;�H;��H;~�H;*�H;&�H;b�H;�H;q�H;adH;�)H;�G;��F;ED;��>;b�4;>";[B;���: �>�z��T^�����&R�hv���o���� �K�ʕ���u��v�ý��p}�ӈ� ]�      �+X��T��nH��6��� �i��B�
䳽�����mR����ټ�����E<��?ݻ1d\������ :�d�:��;*�,;x�:;]7B;��E;oLG;.H;VSH;�{H;}�H;�H;�H;:�H;R�H;�H;��H;��H;��H;��H;��H;�H;Q�H;:�H;�H;�H;��H;�{H;VSH;/H;mLG;��E;]7B;y�:;"�,;��;�d�:� :����3d\��?ݻ�E<�����ټ����mR�����
䳽B�i���� ��6��nH��T�      ఖ�����|���*|�LS\�� :����Z�k$������ �K�u���Oļ����������=&���A/�:�^;��#;�G6;;�?;��D;I�F;��G;�?H;�pH;ޏH;t�H;�H;H�H;0�H;m�H;p�H;��H;z�H;��H;p�H;k�H;,�H;I�H;�H;u�H;�H;�pH;�?H;��G;H�F;��D;>�?;�G6;��#;�^;?/�:���<&������������Oļu�� �K�����k$���Z���� :�LS\��*|�|������      @�;9ɾ{㼾B�������Mw��nH�����Z�䳽ʕ��q\8�m#������^N�K���b�Ix�<5:��:0�;��0;!]=;@�C;�[F;ӞG;�)H;�eH;p�H;!�H;;�H;��H;�H;��H;(�H;��H;l�H;��H;*�H;��H;�H;��H;;�H;'�H;u�H;�eH;�)H;ٞG;�[F;@�C;]=;��0;,�;��:85:�Hx��b�K��^N�����m#��q\8�ʕ��䳽�Z񽰯��nH��Mw�����B��{㼾9ɾ      0y��v�i���B�߾����@��?����nH���B὜u����d�/O�hrμI"�����	�����Pr89a;�:`�;�+;T|:;y7B;��E;�aG;kH;�ZH;c�H;*�H;��H;�H;F�H;E�H;�H;��H;t�H;��H;�H;D�H;E�H;�H;��H;.�H;f�H;�ZH;nH;bG;��E;y7B;W|:;�+;]�;i;�:0r89���	�����I"��hrμ/O���d��u��B����nH�?���@������B�߾j����v�      �O/�pM+�X�����HW��9ɾ@���Mw�� :�i��w�ý�L��[n;�\���rv���E<��˻��-� ��jy�:�^;�%;��7;v�@;5E;�"G;�G;6PH;�zH;��H;X�H;x�H;��H;��H;	�H;��H;��H;��H;
�H;��H;��H;y�H;V�H;��H;�zH;:PH;�G;�"G;5E;x�@;��7;�%;�^;ry�:8����-��˻�E<�rv��\���[n;��L��w�ýi��� :��Mw�@��9ɾHW�����X��pM+�      6�X�VvS�6E��O/��S�HW����������LS\��� ���9����Y�z��΃����]�����$�b���Y�L�Y:��:b`;9�4;�?;9�D;��F;�G; FH;AuH;��H;��H;~�H;�H;��H;�H;�H;��H;�H;�H;��H;�H;�H;��H;ƓH;GuH;FH;�G;��F;9�D;�?;6�4;f`;��:P�Y:��Y��b�������]�΃��z���Y�9����彑� �LS\���������HW���S��O/�6E�VvS�      � ����y�`�h���N��O/����B�߾B���*|��6�p}�䳽iSt�<�!�nrμ@F{��_��X��̓��P:,��:�Z;�2;�O>;lD;%�F;s�G;=H;�pH;��H;H�H;ȷH;��H;��H;Z�H;y�H;\�H;w�H;[�H;��H;��H;˷H;G�H;��H;�pH;=H;z�G;1�F;mD;�O>;�2;�Z;(��:h:Г���X���_�@F{�nrμ<�!�iSt�䳽p}��6��*|�B��B�߾����O/���N�`�h���y�      =v��b���W ��`�h�6E�W��j���{㼾}���nH�ӈ�x�ý�Ȅ��s/��o��#�����$J��,кX	�9Ug�:�l;"0;]=;ٲC;րF;j�G;6H;mH;%�H;��H;|�H;��H;=�H;��H;�H;��H;�H;��H;>�H;��H;|�H;��H;,�H; mH;6H;q�G;�F;ڲC;]=;0;�l;Ug�:�	�9,к"J������#���o��s/��Ȅ�x�ýӈ��nH�}��{㼾j���W��6E�`�h�W ��b���      |h��/���b�����y�VvS�pM+��v�9ɾ�����T� ]�\ν����x\8�����x��%�N���t��h�9n-�:g�;��.;�<;�nC;�dF;�G;�1H;�jH;��H;��H;ɵH;f�H;��H;b�H;��H;��H;��H;e�H;��H;d�H;ʵH;��H;��H;�jH;�1H;�G;�dF;�nC;�<;��.;f�;n-�:��9z��L���%��x�����x\8�����\ν ]��T�����9ɾ�v�pM+�VvS���y�b���/���      dܿ3�ֿ�aǿ=^��/���Xo���7����iþ�(���-=��` �
A���_�0]�.p����I�R�ѻ��)���R���:.�
;�*;"�:;��B;�HF;$�G;�lH;�H;r�H;<�H;��H;|�H;L�H;{�H;�H;��H;�H;{�H;L�H;{�H;��H;:�H;{�H;��H;�lH;(�G;IF;��B;�:;�*;,�
;��:0�R���)�P�ѻ��I�.p��0]��_�
A���` ��-=��(���iþ����7�Xo�/���=^���aǿ3�ֿ      2�ֿCpѿ�¿������_Xi�ϕ3��
�UD��Fl��A�9�.���R�� \� �dx��0�E��ͻ�$�@ �ۍ�:<�;L�*;4�:;�B;�TF;��G;&nH;��H;��H;j�H;��H;��H;Z�H;}�H;�H;��H;�H;��H;X�H;��H;��H;f�H;ķH;��H;(nH;��G;�TF;�B;1�:;E�*;;�;ۍ�: ��$��ͻ0�E�dx�� � \��R��.��A�9�Fl��UD���
�ϕ3�_Xi��������¿Cpѿ      �aǿ�¿����������"Y��f'�����6o���.}��k/����$ڟ�!<Q�-#�ע��(;�,���9�� g7���:�;s,;��;;�C;�vF;�G;�rH;�H;��H;�H;��H;��H;��H;��H;L�H;��H;D�H;��H;��H;��H;��H;�H;��H;�H;�rH;�G;wF;�C;��;;l,;�;��: c7�=��,����(;�ע�-#�!<Q�$ڟ�����k/��.}�7o�������f'��"Y�����������¿      =^������k���Xo���@�(�#�޾����9ce�0����ڽ���� g@������R���O*�IG������C^9,��:;]d.;��<;��C;�F;��G;�yH;��H;�H;�H;��H;h�H;��H;��H;��H;�H;{�H;��H;��H;g�H;��H;�H;�H;��H;�yH;��G;��F;��C;��<;Vd.; ;*��:�C^9���GG���O*��R������ g@�������ڽ0��9ce�����#�޾(���@�Xo�k�������      /����������Xo��!J�K�#��\��VD������zPH�����b��C��� +���ټ(����뿐����d�:$��:C�;�Y1;>;�0D;|�F;^H;C�H;¨H;
�H;[�H;��H;�H;b�H;H�H;��H;_�H;��H;H�H;_�H;�H;��H;U�H;�H;ĨH;C�H;`H;��F;�0D;>;�Y1;D�;$��:|�:���꿐���(����ټ� +�C���b�����zPH�����VD���\��K�#��!J�Xo��������      Xo�_Xi��"Y���@�K�#��
��о�A���i���(�~��ur��
�_��5��ɺ�o�`��<��d�d�h�\�T�X:�P�:�`;˱4;��?;��D;u8G;j0H;��H;k�H;r�H;�H;��H;��H;��H;��H;�H;��H;�H;��H;��H;��H;��H; �H;u�H;k�H;��H;i0H;{8G;��D;��?;Ǳ4;�`;�P�:X�X:h�\�b�d��<��p�`��ɺ��5�
�_�ur��~����(��i��A���о�
�K�#���@��"Y�_Xi�      ��7�ϕ3��f'�(��\���о�����.}��-=�{
���Ľ[��+:��������� �7�"GĻ$�O�����:�{;�D&;�+8;JA;�E;��G;{LH;�H;u�H;2�H;��H;��H;��H;��H;�H;��H;�H;~�H;�H;��H;��H;��H;��H;5�H;v�H;�H;vLH;��G;�E;JA;�+8;�D&;�{;ǿ�: O��Ã$�"GĻ �7���������+:�[����Ľ{
��-=��.}������о�\��(��f'�ϕ3�      ���
�����#�޾VD���A���.}�(�D�ht���ڽ�!��\����Z�ļ�
v�<��ȿ���IɺS�9���:(;�-;��;;��B;fIF;��G;fH;��H;�H;,�H;��H;c�H;��H;Z�H;��H;��H;g�H;��H;��H;Z�H;��H;b�H;��H;0�H;�H;��H;fH;��G;hIF;��B;��;;�-;(;���:�R�9�Iɺǿ��<���
v�Z�ļ���\��!����ڽht�(�D��.}��A��VD��#�޾�����
�      �iþUD��6o�����������i��-=�ht�����R��gys�y +����w񗼒(;�(�ѻ�s@�ԅ!�4j:�P�:��;�D3;3�>;FD;��F;�	H;:|H;��H;q�H;4�H;��H;��H;��H;�H;.�H;n�H;��H;m�H;/�H;�H;��H;��H;��H;6�H;s�H;��H;8|H;�	H;��F;FD;4�>;�D3;��;�P�:4j:؅!��s@�(�ѻ�(;�w����y +�hys��R�����ht��-=��i���������6o��UD��      �(��Fl���.}�9ce�zPH���(�{
���ڽ�R����{�B�6�� �,p��]�`�̨��,��BIҺPL^9���:ۣ;�~(;-�8;�IA;|E;jG;�=H;B�H;լH;�H;]�H;%�H;i�H;��H;��H;��H;��H;J�H;��H;��H;��H;��H;h�H;%�H;`�H;�H;լH;A�H;�=H;jG;�{E;�IA;0�8;�~(;�;���:pL^98IҺ�,��˨�\�`�,p��� �B�6���{��R����ڽ{
���(�zPH�9ce��.}�Fl��      �-=�A�9��k/�0�����~��Ľ�!��hys�B�6�$#��ɺ��vz����>^��f�$��~�D�r:���:��;�Y1;�H=;)xC;'wF;�G;�eH;H�H;��H;��H;��H;P�H;��H;��H;��H;d�H;w�H;��H;y�H;e�H;��H;��H;��H;P�H;��H;��H;��H;H�H;�eH;�G;$wF;*xC;�H=;�Y1;��;��:H�r:�~�e�$�>^������vz��ɺ�$#�B�6�gys��!����Ľ~���0���k/�A�9�      �` �.�����ڽ�b��ur��[��\�y +�� ��ɺ�>��O*�Bͻ�5R�ǅ�Ȝ:,��:��;�);�t8;d�@;W*E;m8G;>$H;@�H;A�H;�H;�H;��H;m�H;a�H;�H;N�H;��H;��H; �H;��H;��H;Q�H;�H;^�H;n�H;��H;&�H;�H;>�H;<�H;?$H;j8G;^*E;f�@;�t8;�);��;,��:��:ǅ��5R�@ͻ�O*�>��ɺ�� �y +�\�[��ur���b����ڽ���.��      
A���R��$ڟ�����C��
�_�*:�������+p���vz��O*��4ֻk�(���P�09.�:1;O� ;�D3;H�=;��C;�kF;��G;�\H;��H;N�H; �H;9�H;��H;w�H;��H;��H;	�H;��H;W�H;��H;W�H;��H;
�H;��H;��H;z�H;��H;>�H; �H;L�H;��H;�\H;��G;�kF;��C;H�=;�D3;T� ;
1;<�:`�09 ���k��4ֻ�O*��vz�+p����輣��*:�
�_�C������$ڟ��R��      �_�\� <Q� g@� +��5�����Y�ļw�\�`����Cͻk��Hɺ �6�?�:�P�:)�;�d.;F�:;#�A;&|E;xNG;B'H;��H;ǥH;[�H;��H;#�H;J�H;Y�H;4�H;��H;��H;�H;��H;��H;��H;�H;��H;��H;4�H;\�H;O�H;*�H;��H;[�H;��H; �H;B'H;~NG;*|E;#�A;N�:;�d.;)�;�P�:?�: �6��Hɺk�Aͻ���\�`�v�Y�ļ�����5�� +� g@� <Q�\�      /]� �-#�������ټ�ɺ������
v��(;�˨�>^���5R�,��� �6����:���:��;)�*;�+8;�!@;U�D;`�F;��G;�eH;}�H;��H;��H;��H;��H;��H; �H;s�H;��H;e�H;}�H;.�H;Y�H;+�H;z�H;g�H;��H;p�H;!�H;��H;��H;��H;��H;��H;��H;�eH;��G;c�F;X�D;�!@;�+8;#�*;��;���:���: �6�$����5R�;^��˨��(;��
v������ɺ���ټ����-#� �      +p��cx��
ע��R��'��p�`���7�:��*�ѻ�,��b�$�ǅ� �09C�:���:�;�~(;�Z6;��>;̨C;�HF;٠G;�DH;F�H;��H;��H;�H;)�H;�H;��H;��H;��H;��H;�H;��H;��H;��H;��H;��H;�H;��H;��H;��H;��H;�H;*�H;�H;��H;��H;E�H;�DH;ܠG;�HF;ҨC;��>;�Z6;�~(;�;���:?�:@�09ǅ�`�$��,��%�ѻ:����7�m�`�(���R��
ע�ax��      �I�-�E��(;��O*����<��GĻ¿���s@�,IҺ�~�Ԝ:<�:�P�:��;�~(;�5;�>;7C;/�E;wcG;8$H;�{H;8�H;�H;��H;��H;9�H;��H;�H;W�H;��H;P�H;��H;A�H;��H;��H;��H;=�H;��H;J�H;��H;Z�H; �H;��H;;�H;��H;��H;�H;8�H;�{H;:$H;zcG;7�E;8C;�>;�5;�~(;��;�P�::�:��:`~�.IҺ�s@�¿�� GĻ�<�����O*��(;�,�E�      B�ѻ�ͻ*���>G��俐�]�d���$��Iɺԅ!��L^9H�r:"��:1;(�;$�*;�Z6;�>;<�B;��E;�8G;�	H;�mH;�H;I�H;��H;b�H;��H;��H;G�H;��H;��H;v�H;��H;��H;��H;�H;!�H;�H;��H;��H;��H;t�H;��H;�H;H�H;��H;��H;`�H;��H;E�H;�H; nH;�	H;�8G;��E;8�B;�>;�Z6;&�*;(�;1;(��:d�r:�L^9��!��Iɺ��$�[�d�ῐ�AG��$����ͻ      i�)�&�$�8���������(�\��N��@S�94j:���:��:��;T� ;�d.;�+8;��>;7C;��E;�)G;��G;dH;�H;��H;\�H;��H;6�H;��H;��H;��H;��H;��H;I�H;{�H;`�H; �H;7�H;I�H;4�H;��H;]�H;x�H;F�H;��H;��H;��H;��H;��H;/�H;��H;\�H;��H;��H;dH;��G;�)G;��E;:C;��>;�+8;�d.;V� ;��;��:���:(4j:@S�9�N��@�\�������7��(�$�      `�R�@ � Y7�E^9t�:`�X:׿�:���:�P�:�;��;�);�D3;L�:;�!@;ҨC;4�E;�8G;��G;�`H;o�H;�H;�H;x�H;:�H;2�H;L�H;]�H;��H;��H;��H;�H;��H;��H;0�H;n�H;c�H;h�H;,�H;��H;��H;	�H;��H;��H;��H;^�H;H�H;-�H;>�H;x�H;�H;�H;s�H;�`H;��G;�8G;4�E;ϨC;�!@;J�:;�D3;�);��;�;�P�:���:տ�:|�X:��:�C^9 c7�� �      ��:���:��: ��:��:�P�:�{;(;��;�~(;�Y1;�t8;E�=; �A;V�D;�HF;wcG;�	H;dH;l�H;G�H;ӶH;0�H;��H;��H;;�H;H�H;��H;!�H;��H;}�H;��H;U�H;��H;H�H;��H;��H;��H;H�H;��H;R�H;��H;~�H;��H; �H;��H;B�H;7�H;��H;��H;.�H;ֶH;K�H;n�H;dH;�	H;zcG;�HF;X�D;�A;F�=;�t8;�Y1;�~(;��;(;�{;�P�:&��: ��:��:���:      0�
;L�;�;;C�;�`;�D&;�-;�D3;2�8;I=;b�@;��C;+|E;c�F;ߠG;=$H;nH;��H;�H;ٶH;��H;7�H;�H;f�H;��H;��H;s�H;j�H;�H;�H;��H;��H;�H;e�H;��H;��H;��H;a�H;�H;��H;��H; �H;�H;g�H;r�H;��H;��H;i�H;�H;3�H;��H;ڶH;�H;��H;nH;>$H;ޠG;d�F;'|E;��C;f�@;I=;2�8;�D3;�-;�D&;�`;Y�;;��;B�;      �*;L�*;n,;jd.;�Y1;ӱ4;,8;��;;:�>;�IA;0xC;[*E;�kF;�NG;��G;�DH;�{H;�H;��H;�H;/�H;6�H;��H;��H;��H;^�H;
�H;��H;��H;��H;��H;n�H;��H;:�H;��H;��H;��H;��H;��H;:�H;��H;j�H;��H;��H;��H;��H;�H;_�H;��H;��H;��H;7�H;2�H;�H;��H;�H;�{H;�DH;��G;NG;�kF;^*E;3xC;�IA;>�>;��;;�+8;α4;�Y1;ld.;k,;6�*;      "�:;@�:;��;;�<;�>;��?;JA;��B;	FD;|E;%wF;k8G;��G;E'H;�eH;L�H;:�H;N�H;_�H;v�H;��H;�H;��H;��H;�H;��H;��H;4�H;w�H;p�H;�H;��H;�H;\�H;}�H;��H;��H;��H;{�H;\�H;�H;��H;�H;m�H;p�H;3�H;��H;��H;�H;��H;��H;�H;��H;u�H;]�H;G�H;:�H;K�H;�eH;@'H;��G;j8G;(wF;|E;FD;��B;JA;��?;>;��<;��;;5�:;      ңB;�B;�C;��C;�0D;��D;��E;fIF;��F;jG;!�G;E$H;�\H;�H;��H;��H;"�H;��H;��H;F�H;��H;k�H;��H;!�H;��H;q�H;��H;E�H;+�H;��H;��H;��H;,�H;q�H;��H;��H;��H;��H;��H;r�H;(�H;��H;��H;��H;$�H;B�H;��H;s�H;��H;�H;��H;n�H;��H;A�H;��H;��H;%�H;��H;��H;�H;�\H;F$H;&�G;jG;��F;jIF;��E;��D;�0D;��C;�C;�B;      �HF;�TF;wF;��F;u�F;~8G;��G;��G;�	H;�=H;�eH;?�H;��H;˥H;��H;��H;��H;g�H;5�H;/�H;=�H;��H;a�H;��H;p�H;��H;#�H;	�H;��H;D�H;��H;!�H;4�H;o�H;��H;��H;��H;��H;��H;n�H;2�H;�H;��H;A�H;��H;	�H;�H;��H;s�H;��H;[�H;��H;=�H;-�H;3�H;b�H;��H;��H;��H;ȥH;��H;@�H;fH;�=H;�	H;��G;��G;r8G;��F;��F;�vF;�TF;      <�G;��G;�G;��G;YH;k0H;�LH;fH;5|H;B�H;I�H;>�H;G�H;Z�H;��H;�H;��H;��H;��H;M�H;O�H;��H;�H;��H;��H;"�H;��H;��H;Q�H;��H;��H;0�H;O�H;r�H;��H;��H;��H;}�H;��H;t�H;L�H;,�H;��H;��H;J�H;��H;��H;'�H;��H;��H;
�H;��H;N�H;J�H;��H;��H;��H;�H;��H;V�H;H�H;@�H;J�H;A�H;:|H;fH;}LH;f0H;oH;��G;�G;��G;      �lH;*nH;�rH;�yH;>�H;��H;�H;��H;��H;ܬH;��H;��H;��H;��H;��H;*�H;;�H;��H;��H;]�H;��H;s�H;��H;9�H;A�H;�H;��H;5�H;��H;��H;�H;:�H;^�H;c�H;|�H;��H;}�H;��H;{�H;c�H;\�H;4�H;�H;��H;��H;3�H;��H;�H;B�H;4�H;��H;s�H;��H;]�H;��H;��H;;�H;,�H;��H;��H;��H;��H;��H;٬H;��H;��H;�H;��H;I�H;�yH;�rH;!nH;      �H;��H;�H;��H;��H;j�H;|�H;�H;h�H;�H;��H;%�H;=�H;&�H;��H;�H;��H;N�H;��H;��H;+�H;i�H;��H;y�H;'�H;��H;J�H;��H;��H;�H;(�H;K�H;^�H;c�H;a�H;m�H;j�H;h�H;`�H;d�H;`�H;G�H;*�H;�H;��H;��H;D�H;��H;(�H;s�H;��H;g�H;'�H;��H;��H;K�H;��H;�H;��H;&�H;;�H;#�H;��H;�H;o�H;�H;{�H;g�H;ŨH;��H;�H;��H;      u�H;��H;��H;�H;�H;q�H;4�H;,�H;3�H;`�H;��H;��H;��H;R�H;��H;��H;#�H;�H;��H;��H;��H;�H;��H;q�H;��H;=�H;��H;��H;�H;#�H;@�H;B�H;P�H;c�H;K�H;Z�H;o�H;Y�H;H�H;c�H;L�H;@�H;>�H;!�H;
�H;��H;��H;A�H;��H;m�H;��H;�H;��H;��H;��H; �H;#�H;��H;��H;O�H;��H;��H;��H;c�H;4�H;-�H;6�H;n�H;�H;�H;��H;��H;      C�H;��H;�H;%�H;Z�H;�H;��H;��H;��H;)�H;T�H;t�H;~�H;`�H;$�H;��H;`�H;��H;��H;��H;��H;$�H;��H;�H;��H;��H;��H;�H;/�H;E�H;U�H;N�H;@�H;>�H;`�H;N�H;-�H;K�H;\�H;A�H;>�H;N�H;U�H;D�H;)�H;�H;��H;��H;��H;�H;��H;#�H;��H;��H;��H;��H;a�H;��H;$�H;`�H;~�H;u�H;T�H;*�H;��H;��H;��H;��H;h�H;#�H;�H;��H;      ��H;��H;��H;��H;��H;��H;�H;c�H;��H;h�H;��H;e�H;��H;9�H;s�H;��H;��H;{�H;O�H;�H;��H;��H;p�H;��H;��H;�H;/�H;;�H;K�H;D�H;H�H;U�H;=�H;6�H;I�H;*�H;#�H;-�H;G�H;7�H;>�H;U�H;G�H;B�H;E�H;9�H;,�H;"�H;��H;��H;t�H;��H;��H;�H;M�H;|�H;��H;��H;s�H;9�H;��H;e�H;��H;i�H;��H;d�H;�H;��H;��H;��H;��H;��H;      ��H;��H;�H;n�H;�H;��H;��H;��H;��H;��H;��H;�H;��H;��H;��H;��H;T�H;�H;��H;��H;_�H;��H;��H;�H;/�H;3�H;R�H;e�H;g�H;S�H;:�H;>�H;E�H;=�H;�H;�H;K�H;�H;�H;@�H;B�H;A�H;9�H;O�H;`�H;`�H;O�H;4�H;2�H;�H;��H;��H;Y�H;��H;��H;�H;V�H;��H;��H;��H; �H;�H;��H;��H;��H;��H;��H;��H;�H;e�H;�H;��H;      H�H;Z�H;��H;��H;c�H;��H;��H;Z�H;�H;��H;��H;U�H;�H;��H;i�H;�H;��H;��H;c�H;��H;��H;#�H;;�H;Y�H;r�H;n�H;q�H;e�H;e�H;e�H;9�H;9�H;>�H;&�H;�H;�H;%�H;�H;�H;(�H;>�H;9�H;9�H;c�H;`�H;a�H;o�H;o�H;t�H;V�H;>�H;!�H;��H;��H;c�H;�H;��H;�H;h�H;��H;�H;T�H;��H;��H;�H;\�H;��H;��H;l�H;��H;��H;b�H;      u�H;��H;��H;��H;V�H;��H;!�H;��H;2�H;��H;m�H;��H;��H;�H;��H;��H;G�H;��H; �H;3�H;L�H;d�H;��H;u�H;��H;��H;��H;}�H;e�H;O�H;W�H;K�H;�H;�H;"�H;�H;��H;�H;!�H;�H;!�H;N�H;V�H;I�H;^�H;x�H;��H;��H;��H;t�H;��H;`�H;G�H;,�H;��H;��H;G�H;��H;��H;�H;��H;��H;o�H;��H;6�H;��H;$�H;��H;W�H;��H;��H;��H;      �H;�H;J�H;~�H;��H;�H;��H;��H;k�H;��H;}�H;��H;W�H;��H;.�H;��H;��H;�H;7�H;m�H;��H;��H;��H;��H;��H;��H;��H;��H;o�H;^�H;I�H;/�H;"�H;�H;�H;�H;�H;�H;�H;!�H;"�H;2�H;H�H;Z�H;k�H;��H;�H;��H;��H;��H;��H;��H;��H;h�H;7�H;	�H;��H;��H;+�H;��H;U�H;��H;~�H;��H;o�H;��H;��H;�H;��H;~�H;I�H;+�H;      ��H;��H;��H;�H;\�H;��H;�H;h�H;��H;J�H;��H;(�H;��H;�H;`�H;��H;��H;(�H;N�H;k�H;��H;��H;��H;��H;��H;��H;��H;��H;q�H;v�H;*�H;(�H;O�H;#�H;��H;�H;��H;�H;��H;%�H;R�H;*�H;*�H;r�H;j�H;��H;��H;��H;��H;��H;��H;��H;��H;g�H;N�H;)�H;��H;��H;]�H;�H;��H;'�H;��H;J�H;��H;k�H;!�H;��H;_�H;�H;��H;��H;      �H;!�H;D�H;�H;��H;�H;��H;��H;k�H;��H;|�H;��H;X�H;��H;.�H;��H;��H;�H;7�H;m�H;��H;��H;��H;��H;��H;��H;��H;��H;q�H;]�H;I�H;0�H;#�H;�H;�H;�H;�H;�H;�H;�H;"�H;2�H;H�H;Y�H;k�H;��H;�H;��H;��H;��H;��H;��H;��H;h�H;7�H;�H;��H;��H;+�H;��H;W�H;��H;~�H;��H;n�H;��H;��H;�H;��H;��H;L�H;'�H;      m�H;��H;��H;��H;V�H;��H;!�H;��H;2�H;��H;m�H;��H;��H;�H;��H;��H;F�H;��H; �H;2�H;N�H;d�H;��H;r�H;��H;��H;��H;}�H;e�H;L�H;V�H;K�H;�H;�H;#�H;�H;��H;�H;#�H;�H;"�H;K�H;V�H;H�H;^�H;v�H;��H;��H;��H;r�H;��H;a�H;E�H;-�H;��H;��H;G�H;��H;�H;�H;��H;��H;k�H;��H;5�H;��H;(�H;��H;Z�H;��H;��H;��H;      F�H;W�H;��H;��H;e�H;��H;��H;]�H;�H;��H;��H;T�H;�H;��H;k�H;�H;��H;�H;c�H;��H;��H;#�H;:�H;Y�H;u�H;m�H;r�H;e�H;g�H;e�H;9�H;9�H;>�H;&�H;�H;�H;%�H;�H;�H;&�H;@�H;9�H;7�H;a�H;]�H;a�H;n�H;o�H;q�H;S�H;>�H;"�H;��H;��H;d�H;�H;��H;�H;i�H;��H;�H;R�H;��H;��H;�H;]�H;��H;��H;l�H;��H;��H;W�H;      ��H;��H;�H;g�H;�H;��H;��H;��H;��H;��H;��H;�H; �H;��H;��H;��H;T�H;�H;�H;��H;_�H;��H;��H;�H;2�H;/�H;P�H;e�H;g�H;S�H;9�H;;�H;D�H;;�H;�H;�H;K�H;�H;�H;>�H;A�H;@�H;9�H;N�H;]�H;^�H;L�H;3�H;-�H;�H;��H;��H;V�H;��H;��H;�H;S�H;��H;��H;��H;��H;�H;��H;��H;��H;��H;��H;��H;�H;o�H;�H;��H;      |�H;��H;��H;��H;��H;��H;�H;f�H;��H;h�H;��H;e�H;��H;:�H;v�H;��H;��H;|�H;M�H;�H;��H;��H;p�H;��H;��H;�H;,�H;;�H;N�H;B�H;G�H;S�H;=�H;4�H;I�H;)�H;#�H;-�H;G�H;7�H;=�H;U�H;E�H;A�H;E�H;6�H;)�H;�H;��H;��H;t�H;��H;��H;�H;M�H;{�H;��H;��H;r�H;7�H;��H;d�H;��H;h�H;��H;f�H;	�H;��H;��H;��H;��H;��H;      6�H;��H;�H;�H;_�H;�H;��H;��H;��H;)�H;T�H;v�H;}�H;a�H;'�H;��H;a�H;��H;��H;��H;��H;$�H;��H;�H;��H;��H;��H;
�H;/�H;D�H;S�H;N�H;>�H;>�H;`�H;L�H;-�H;L�H;\�H;A�H;>�H;N�H;S�H;A�H;(�H;�H;��H;��H;��H;�H;��H;#�H;��H;��H;��H;��H;a�H;��H;$�H;^�H;{�H;t�H;S�H;(�H;��H;��H;��H;��H;l�H;'�H;�H;�H;      ��H;��H;��H;�H; �H;{�H;4�H;3�H;7�H;b�H;��H;��H;��H;Q�H;��H;��H;#�H;�H;��H;��H;��H;�H;��H;o�H;��H;:�H;��H;��H;�H;!�H;>�H;A�H;L�H;c�H;K�H;Y�H;o�H;Y�H;H�H;a�H;L�H;@�H;=�H;!�H;	�H;��H;��H;A�H;��H;i�H;��H;�H;��H;��H;��H; �H;!�H;��H;��H;N�H;��H;��H;��H;b�H;4�H;1�H;5�H;k�H;�H;"�H;��H;��H;       �H;��H;*�H;��H;��H;p�H;y�H;�H;s�H;�H;��H;&�H;=�H;)�H;��H;�H;��H;O�H;��H;��H;-�H;j�H;��H;y�H;*�H;��H;F�H;��H;��H;
�H;(�H;K�H;^�H;d�H;a�H;k�H;j�H;j�H;`�H;c�H;^�H;I�H;)�H;
�H;��H;��H;D�H;��H;&�H;p�H;��H;i�H;&�H;��H;��H;K�H;��H;�H;��H;&�H;;�H;!�H;��H;�H;p�H;�H;|�H;j�H;��H;��H;*�H;~�H;      �lH;nH;�rH;�yH;7�H;��H;�H;��H;��H;ܬH;��H;��H;��H;��H;��H;,�H;;�H;��H;��H;^�H;��H;u�H;��H;7�H;B�H;�H;��H;3�H;��H;��H;�H;:�H;]�H;a�H;{�H;��H;�H;��H;{�H;d�H;`�H;7�H;�H;��H;��H;0�H;��H;�H;>�H;3�H;��H;r�H;��H;[�H;��H;��H;:�H;*�H;��H;��H;��H;��H;��H;جH;��H;��H;�H;��H;I�H;�yH;�rH;nH;      -�G;��G;�G;��G;gH;r0H;�LH;fH;8|H;A�H;I�H;B�H;H�H;Z�H;��H;�H;��H;��H;��H;J�H;P�H;��H;�H;��H;��H;�H;��H;��H;O�H;��H;��H;0�H;L�H;r�H;��H;��H;��H;��H;��H;u�H;O�H;0�H;��H;��H;H�H;��H;��H;&�H;��H;��H;�H;��H;K�H;M�H;��H;��H;��H;�H;��H;V�H;E�H;=�H;H�H;>�H;7|H;fH;�LH;k0H;lH;��G;�G;��G;      �HF;�TF;	wF;�F;y�F;�8G;��G;��G;�	H;�=H;fH;E�H;��H;ʥH;��H;��H;��H;h�H;5�H;/�H;@�H;��H;Z�H;��H;q�H;��H; �H;�H;��H;@�H;��H;!�H;2�H;o�H;��H;��H;��H;��H;��H;o�H;3�H;!�H;��H;A�H;��H;�H;"�H;��H;p�H;��H;_�H;��H;=�H;/�H;5�H;a�H;��H;��H;��H;ǥH;��H;>�H;fH;�=H;�	H;��G;��G;t8G;��F;�F;�vF;�TF;      ΣB;�B;�C;��C;�0D;��D;��E;iIF;��F;jG;$�G;F$H;�\H;�H;��H;��H;$�H;��H;��H;B�H;��H;n�H;��H; �H;��H;l�H;��H;C�H;*�H;��H;��H;��H;)�H;q�H;��H;��H;��H;��H;��H;t�H;,�H;��H;��H;��H;$�H;?�H;��H;s�H;��H;�H;��H;n�H;��H;B�H;��H;��H;$�H;��H;��H;�H;�\H;B$H;�G;jG;��F;hIF;��E;��D;�0D;��C;�C;�B;      ��:;#�:;}�;;�<;�>;ȧ?;JA;��B;FD;|E;(wF;m8G;��G;C'H;�eH;M�H;:�H;N�H;]�H;u�H;��H;�H;��H;��H;�H;��H;��H;4�H;v�H;l�H;�H;��H;�H;\�H;{�H;��H;��H;��H;{�H;\�H;�H;��H;�H;o�H;r�H;0�H;��H;��H;�H;��H;��H;�H;��H;x�H;]�H;I�H;:�H;K�H;�eH;@'H;��G;g8G;%wF; |E;FD;��B;JA;��?;>;�<;}�;;�:;      �*;A�*;d,;rd.;�Y1;˱4;�+8;��;;?�>;�IA;+xC;^*E;�kF;�NG;��G;�DH;�{H;�H;��H;�H;0�H;7�H;��H;��H;��H;X�H;�H;��H;��H;��H;��H;n�H;��H;:�H;��H;��H;��H;��H;��H;9�H;��H;n�H;��H;��H;��H;��H;�H;_�H;��H;��H;��H;7�H;3�H;�H;��H;�H;�{H;�DH;��G;}NG;�kF;X*E;*xC;�IA;<�>;��;;�+8;˱4;�Y1;sd.;c,;,�*;      ,�
;L�;��;
;C�;�`;�D&;�-;�D3;0�8;I=;g�@;��C;)|E;g�F;�G;=$H;nH;��H;�H;ٶH;��H;3�H;�H;j�H;��H;��H;s�H;i�H;�H;�H;��H;��H;�H;a�H;��H;��H;��H;`�H;�H;��H;��H;#�H;�H;i�H;r�H;��H;��H;g�H;!�H;7�H;��H;ڶH;�H;��H; nH;;$H;ܠG;c�F;'|E;��C;b�@;I=;-�8;�D3;�-;�D&;�`;X�;�;��;?�;      ��:鍨:��:*��:��:�P�:�{;(;��;�~(;�Y1;�t8;F�=; �A;[�D;�HF;ycG;�	H;dH;n�H;G�H;ضH;.�H;��H;��H;4�H;B�H;��H; �H;��H;~�H;��H;R�H;��H;G�H;��H;��H;��H;G�H;��H;V�H;��H;��H;��H; �H;��H;G�H;9�H;��H;��H;0�H;ֶH;I�H;o�H;dH;�	H;ycG;�HF;X�D;�A;E�=;�t8;�Y1;�~(;��;(;�{;�P�:.��:.��:��:Í�:      ��R�� � ^7��D^9p�:|�X:ݿ�:���:�P�:�;��;�);�D3;J�:;�!@;ӨC;4�E;�8G;��G;�`H;q�H;�H;�H;x�H;>�H;,�H;E�H;]�H;��H;��H;��H;�H;��H;��H;/�H;j�H;d�H;k�H;,�H;��H;��H;�H;��H;��H;��H;]�H;L�H;2�H;;�H;|�H;�H;�H;r�H;�`H;��G;�8G;2�E;ШC;�!@;G�:;�D3;�);��;ޣ;�P�:���:Ͽ�:T�X:|�:0D^9 ]7�0 �      i�)�'�$�7�����"���,�\��N��0S�9(4j:���:��:��;U� ;�d.;�+8;��>;7C;��E;�)G;��G;dH;��H;��H;[�H;��H;0�H;��H;��H;��H;��H;��H;H�H;{�H;`�H;��H;6�H;I�H;6�H;��H;]�H;{�H;I�H;��H;��H;��H;��H;��H;3�H;��H;`�H;��H;�H;dH;��G;�)G;��E;6C;��>;�+8;�d.;R� ;��;��:���:4j:0S�9�N��8�\� ������>��#�$�      J�ѻ�ͻ,���BG��࿐�T�d���$��Iɺ��!��L^9`�r:(��:1;&�;)�*;�Z6;�>;9�B;��E;�8G;�	H; nH;�H;I�H;��H;a�H;��H;��H;H�H;��H;��H;u�H;��H;��H;��H;�H;"�H;�H;��H;��H;��H;t�H;��H;�H;H�H;��H;��H;a�H;��H;G�H;�H;�mH;�	H;�8G;��E;8�B;�>;�Z6;&�*;$�;1;"��:d�r:�L^9ą!��Iɺ��$�Y�d�⿐�DG��0����ͻ      �I�.�E��(;��O*����<��GĻÿ���s@�.IҺx~��::�:�P�:��;�~(;�5;�>;6C;2�E;zcG;:$H;�{H;:�H;�H;��H;��H;9�H;��H;�H;X�H;��H;O�H;��H;@�H;��H;��H;��H;?�H;��H;L�H;��H;[�H;�H;��H;9�H;��H;��H;�H;:�H;�{H;:$H;vcG;5�E;4C;�>;�5;�~(;��;�P�::�:Ԝ:�~�4IҺ�s@�ÿ�� GĻ�<�����O*��(;�-�E�      +p��cx��ע��R��(��m�`���7�9��&�ѻ�,��`�$�ǅ�@�09?�:���:�;�~(;�Z6;��>;ΨC;�HF;ܠG;�DH;I�H;��H;��H;�H;(�H;�H;��H;��H;��H;��H;�H;��H;��H;��H;��H;��H;�H;��H;��H;��H;��H;�H;)�H;�H;��H;��H;H�H;�DH;۠G;�HF;ШC;~�>;�Z6;�~(;�;���:=�: �09ǅ�b�$��,��(�ѻ:����7�n�`�)���R��ע�cx��      0]� �-#�������ټ�ɺ������
v��(;�˨�<^���5R�(��� �6����:���:��;$�*;�+8;�!@;Y�D;c�F;��G;�eH;��H;��H;��H;��H;��H;��H; �H;r�H;��H;h�H;}�H;+�H;Y�H;+�H;{�H;g�H;��H;p�H; �H;��H;��H;��H;��H;��H;~�H;�eH;��G;c�F;T�D;�!@;�+8;#�*;��;���:���: �6�,����5R�=^��̨��(;��
v������ɺ���ټ����-#� �      �_�\� <Q� g@� +��5�����Y�ļv�\�`����Bͻk��Hɺ �6�I�:�P�:&�;�d.;I�:;'�A;)|E;~NG;F'H;�H;ȥH;X�H;��H;&�H;K�H;\�H;4�H;��H;��H;�H;��H;��H;��H;�H;��H;��H;3�H;Z�H;O�H;*�H;��H;W�H;ƥH;��H;F'H;�NG;'|E;�A;M�:;�d.;(�;�P�:C�: �6��Hɺk�Bͻ���\�`�w�Y�ļ�����5�� +� g@� <Q�\�      
A���R��$ڟ�����C��
�_�*:�������+p���vz��O*��4ֻ	k����`�096�:	1;Q� ;�D3;L�=;��C;�kF;��G;�\H;��H;H�H;��H;=�H;��H;x�H;��H;��H;�H;��H;W�H;��H;W�H;��H;
�H;��H;��H;x�H;��H;@�H; �H;I�H;��H;�\H;��G;�kF;��C;D�=;�D3;O� ;	1;6�:P�09���k��4ֻ�O*��vz�,p����輣��+:�
�_� C������$ڟ��R��      �` �.�����ڽ�b��ur��[��\�y +�� ��ɺ�>��O*�Bͻ�5R�ǅ�М:"��:��;�);�t8;d�@;^*E;n8G;B$H;?�H;=�H;�H;"�H;��H;o�H;a�H;�H;Q�H;��H;��H;!�H;��H;��H;O�H; �H;`�H;n�H;��H;(�H;�H;=�H;?�H;=$H;n8G;^*E;d�@;�t8;�);��;*��:؜:ǅ��5R�Cͻ�O*�?��ɺ�� �y +�\�[��ur���b����ڽ���.��      �-=�A�9��k/�0�����~��Ľ�!��hys�B�6�$#��ɺ��vz����=^��f�$��~�<�r:���:��;�Y1;�H=;-xC;'wF;�G;�eH;C�H;��H;��H;��H;Q�H;��H;��H;��H;d�H;z�H;��H;y�H;d�H;��H;��H;��H;P�H;��H;��H;��H;E�H;�eH;�G;'wF;+xC;�H=;�Y1;��;���:H�r:�~�g�$�>^������vz��ɺ�$#�B�6�gys��!����Ľ}���0���k/�A�9�      �(��Fl���.}�9ce�zPH���(�{
���ڽ�R����{�B�6�� �,p��]�`�̨��,��<IҺ@L^9���:ޣ;�~(;/�8;�IA;|E;jG;�=H;?�H;ԬH;�H;_�H;&�H;f�H;��H;��H;��H;��H;L�H;��H;��H;��H;��H;h�H;&�H;`�H;!�H;֬H;?�H;�=H;jG;|E;�IA;-�8;�~(;�;���:PL^98IҺ�,��˨�]�`�,p��� �B�6���{��R����ڽ{
���(�zPH�9ce��.}�Fl��      �iþUD��6o�����������i��-=�ht�����R��gys�y +����w񗼒(;�(�ѻ�s@��!�4j:�P�:��;�D3;5�>;FD;��F;�	H;8|H;��H;s�H;4�H;��H;��H;��H;�H;.�H;n�H;��H;m�H;/�H;�H;��H;��H;��H;6�H;v�H;��H;:|H;�	H;��F;FD;7�>;�D3;��;�P�:�3j:ԅ!��s@�(�ѻ�(;�w����y +�gys��R�����ht��-=��i���������6o��UD��      ���
�����#�޾VD���A���.}�(�D�ht���ڽ�!��\����Z�ļ�
v�<��ǿ���IɺS�9���:(;�-;��;;��B;iIF;��G;fH;��H;�H;,�H;��H;c�H;��H;\�H;��H;��H;h�H;��H;��H;Y�H;��H;c�H;��H;1�H;�H;��H;fH;��G;hIF;��B;��;;�-;(;���:�R�9�Iɺƿ��<���
v�Z�ļ���\��!����ڽht�(�D��.}��A��VD��#�޾�����
�      ��7�ϕ3��f'�(��\���о�����.}��-=�{
���Ľ[��+:��������� �7�"GĻŃ$� O��ÿ�:�{;�D&;�+8;JA;�E;��G;vLH;�H;u�H;2�H;��H;��H;��H;��H;�H;��H;�H;��H;�H;��H;��H; �H;��H;6�H;{�H;�H;{LH;��G;�E;JA;�+8;�D&;�{;ɿ�: O����$� GĻ �7���������+:�[����Ľ{
��-=��.}������о�\��(��f'�ϕ3�      Xo�_Xi��"Y���@�K�#��
��о�A���i���(�~��ur��
�_��5��ɺ�p�`��<��e�d�`�\�X�X:�P�:�`;˱4;��?;��D;t8G;i0H;��H;j�H;t�H;�H;��H;��H;��H;��H;�H;��H;�H;��H;��H;��H;��H;�H;w�H;n�H;��H;k0H;~8G;��D;��?;ʱ4;�`;�P�:`�X:p�\�c�d��<��p�`��ɺ��5�
�_�ur��~����(��i��A���о�
�K�#���@��"Y�_Xi�      /����������Xo��!J�K�#��\��VD������zPH�����b��C��� +���ټ(����쿐����p�:&��:C�;�Y1;>;�0D;x�F;]H;B�H;��H;�H;Z�H;��H;�H;c�H;C�H;��H;]�H;��H;F�H;_�H;�H;��H;X�H;�H;ŨH;H�H;dH;��F;�0D;>;�Y1;E�;$��:|�:���꿐���(����ټ� +�C���b�����zPH�����VD���\��K�#��!J�Xo��������      =^������k���Xo���@�(�$�޾����9ce�0����ڽ���� g@������R���O*�HG������C^9,��: ;[d.;��<;��C;�F;��G;�yH;��H;�H;�H;��H;h�H;��H;��H;�H;�H;~�H;��H;��H;i�H;��H;�H; �H;��H;�yH;��G;��F;��C;��<;Wd.; ;,��:D^9���FG���O*��R������ g@�������ڽ0��9ce�����#�޾(���@�Xo�k�������      �aǿ�¿����������"Y��f'�����6o���.}��k/����$ڟ�!<Q�-#�ע��(;�-���9�� e7���:��;r,;��;;�C;�vF;�G;�rH;�H;��H;�H;��H;��H;��H;��H;J�H;��H;F�H;��H;��H;��H;��H;�H;��H;�H;�rH;�G;wF;�C;��;;l,;�;��: a7�9��+����(;�ע�-#�!<Q�$ڟ�����k/��.}�6o�������f'��"Y�����������¿      2�ֿCpѿ�¿������_Xi�ϕ3��
�UD��Fl��A�9�.���R�� \� �dx��0�E��ͻ�$�0 �ۍ�:<�;L�*;5�:;�B;�TF;��G;%nH;��H;��H;j�H;��H;��H;Z�H;�H;�H;��H;�H;��H;Z�H;��H;��H;f�H;ķH;��H;(nH;��G;�TF;�B;2�:;E�*;;�;ۍ�:  � �$��ͻ1�E�dx�� � \��R��.��A�9�Fl��UD���
�ϕ3�_Xi��������¿Cpѿ      �� $������꿯�ſ�ޞ�%3s��2�>����� j���yHͽƸ����'�B<ͼr�n�e���BQ^��-.�n��:nW;aS%;fo8;��A;DF;�H;z�H;��H;��H;�H;�H;"�H;��H;��H;��H;�H;��H;��H;��H;"�H;�H;�H;��H;��H;}�H;�H;DF;��A;bo8;XS%;jW;p��:�-.�CQ^�d���r�n�B<ͼ��'�Ƹ��yHͽ�� j���>����2�%3s��ޞ���ſ������ $�       $�������忇�����cm�V�-�����Ph��Vde�"-�֪ɽ�v��(�$��ɼzmj�8���X�$���ņ:fx;�%;2�8;EB; RF;�H;�H;�H;��H;C�H;�H;�H;v�H;��H;��H;�H;��H;��H;u�H;�H;�H;A�H;��H;�H;�H;�H;*RF;CB;.�8;�%;dx;�ņ:��X�6���zmj��ɼ(�$��v��תɽ"-�Vde�Ph������V�-�cm��������忝����      ����������ԿLw�����:�\�"����k��Y0X�����;����w����������]� ���F�����ɒ:��;�';��9;�oB;�zF;�!H;s�H;��H;�H;o�H;�H;�H;�H;��H;��H;��H;��H;��H;}�H;�H;�H;k�H;�H;��H;t�H;�!H;�zF;�oB;��9;��';��;�ɒ:����F� �黫�]����������w��;�����Y0X�k�����"�:�\����Lw���Կ��𿝏�      ������Կp���ޞ�`F�h�C�-E�"�;�I��D���"��f�c�|��֯���J��ѻТ)��K���:
�
;�M*;m�:;�C;ʸF;�8H;-�H;H�H;Z�H;��H;�H;�H;��H;��H;��H;��H;��H;��H;}�H;�H;�H;��H;^�H;K�H;+�H;�8H;иF;�C;i�:;�M*;�
;��:�K�Ѣ)��ѻ��J��֯�|�f�c�"����D��I��"�;-E�g�C�`F��ޞ�p���Կ��      ��ſ���Lw���ޞ�����?�W�5�%�����hɰ��|x�e{+�ѱ����J��  �ζ��Y�1�*���+�  
9��:��;�-;��<;]�C;�G;�TH;$�H;��H;��H;��H;)�H;�H;d�H;��H;t�H;��H;o�H;��H;c�H;�H;)�H;��H;��H;��H;&�H;�TH;�G;Z�C;��<;ܷ-;��;��:P 
9!+�)���Z�1�ζ���  ��J���ѱ�e{+��|x�hɰ�����5�%�>�W������ޞ�Lw�����      �ޞ�������_F�>�W�W�-���?Kɾ�G����O����ƽǸ��̈́-���ۼㄼ44�ǐ�϶�]:��:};|�1;�c>;D�D;x\G;,sH;v�H;7�H;D�H;��H;J�H;�H;I�H;j�H;]�H;��H;Y�H;h�H;D�H;
�H;K�H;��H;H�H;5�H;w�H;*sH;|\G;B�D;�c>;x�1;|;��:$]:϶�ǐ�44�ㄼ��ۼ̈́-�Ǹ��ƽ�����O��G��?Kɾ��W�-�>�W�_F�������      %3s�cm�:�\�h�C�5�%����TҾj��	 j��C(����]P����[�|������Y�:��eX�l�<���k:2��:�� ;֟5;1R@;5uE;ϲG;�H; �H;��H;��H;!�H;F�H;	�H;A�H;N�H;7�H;m�H;4�H;L�H;@�H;�H;D�H;�H;��H;��H;�H;�H;ҲG;5uE;-R@;ҟ5;�� ;(��:�k:p�<�eX�8����Y����|���[�]P����콪C(�	 j�j���TҾ��5�%�h�C�:�\�cm�      �2�U�-�"�-E�����?Kɾj����s�8�5���u㻽�v��	z0��;��+���*����56�@BS�CM�:M�	;p�(;�9;�/B;HDF; H;��H;]�H;��H;��H;M�H;c�H;��H;�H;�H;�H;9�H;�H;�H;�H;��H;`�H;J�H;��H;��H;\�H;��H; H;HDF;�/B;�9;p�(;H�	;OM�:�BS�26�����*��+���;�	z0��v��u㻽��8�5���s�j��?Kɾ����-E�"�U�-�      >����������"�;hɰ��G��	 j�8�5��	�ΪɽY����J�s���沼��]�����	x�V	��n:���:�v;��/;f-=;��C;�F;�HH;{�H;��H;��H;�H;}�H;f�H;��H;��H;��H;��H;�H;��H;��H;��H;��H;f�H;{�H;�H;��H;��H;x�H;�HH;�F;��C;g-=;��/;�v;���:n:V	���	x������]��沼r���J�Y���Ϊɽ�	�8�5�	 j��G��hɰ�"�;��徶���      ��Ph��k���I���|x���O��C(���Ϊɽ����RDX�G��&<ͼㄼ�X!��s���W��uK���:�y;��#;�H6;R@;�PE;g�G;\�H;��H;�H;��H;}�H;��H;T�H;��H;��H;��H;��H;��H;��H;��H;��H;��H;R�H;��H;��H;��H;�H;��H;X�H;i�G;�PE;
R@;�H6;��#;�y;��:�uK��W��s���X!�ㄼ&<ͼG��RDX�����Ϊɽ���C(���O��|x��I��k��Ph��       j�Vde�Y0X�D�e{+�������t㻽Y���RDX������ۼ˾����;�F>ۻX�l�y��>":���:��;��-;��;;��B;lzF;�H;`�H;X�H;��H;��H;��H;��H;N�H;��H;|�H;r�H;��H;[�H;��H;r�H;|�H;��H;K�H;��H;��H;��H;��H;W�H;[�H;�H;hzF;��B;��;;��-;��;���:�>":T�y�X�D>ۻ��;�ʾ����ۼ���RDX�Y���t㻽��콂��f{+�D�Y0X�Vde�      ��!-������ѱ�ƽ]P���v���J�G����ۼ��c�J������+���rѺ (
9�M�:��;r $;��5;��?;\�D;>\G;�eH;��H;��H;��H;��H;��H;��H;5�H;T�H;<�H;5�H;G�H;�H;F�H;3�H;=�H;R�H;2�H;��H;�H;��H;��H;��H;��H;�eH;=\G;b�D;��?;��5;| $;��;�M�:`(
9�rѺ�+������b�J�����ۼG���J��v��]P��ƽѱ轃����!-�      yHͽ֪ɽ�;��"����Ǹ����[�z0�r��%<ͼʾ��b�J�����j��}*�p�訂::b�:5�;��/;|L<;�C;mF;m�G;ڡH;��H;��H;��H;�H;2�H;��H;�H;�H;��H;��H;��H;��H;��H;��H;��H;�H;�H;��H;8�H;�H;��H;��H;��H;ޡH;l�G;mF;�C;~L<;��/;9�;2b�:���:P�z*��j�����b�J�ʾ��%<ͼr��z0���[�Ǹ����"���;��֪ɽ      Ÿ���v����w�f�c��J�΄-�{��;缄沼ㄼ��;������j���5�`���>Q:2��:Oi;�M*;d�8;d�@;�PE;�uG;iH;��H;��H;��H;��H;��H;U�H;��H;��H;��H;��H;��H;��H;��H;��H;��H;��H;��H;��H;��H;\�H;��H; �H;��H;��H;��H;iH;�uG;�PE;d�@;l�8;�M*;Oi;@��:�>Q:H�깤5��j��������;�ㄼ�沼�;�{�̈́-��J�f�c���w��v��      ��'�'�$����{��  ���ۼ����+����]��X!�D>ۻ�+��~*�`����>:���:��;!�%;Ο5;w�>;�(D;��F;T!H;�H;)�H;��H;��H;��H;��H;M�H;��H;��H;l�H;p�H;L�H;6�H;Q�H;4�H;I�H;p�H;j�H;��H;��H;Q�H;��H;��H;��H;��H;+�H;�H;U!H;��F;�(D;~�>;ҟ5;�%;��;���:��>:P��{*��+��B>ۻ�X!���]��+�������ۼ�  �|����(�$�      ><ͼ~�ɼ�����֯�Ͷ��ㄼ��Y��*�����s��X��rѺ���>Q:���:��
;2�#;O�3;sc=;�#C;DF;��G;�H;��H;��H;�H;��H;5�H;��H;F�H;p�H;I�H;�H;4�H;��H;��H;��H;��H;��H;2�H;�H;F�H;s�H;I�H;�H;8�H;��H;�H;��H;��H;�H;��G;DF;�#C;tc=;K�3;8�#;��
;���:�>Q:���rѺX��s������*���Y�ㄼζ���֯�����|�ɼ      m�n�vmj���]���J�X�1�34�4������	x��W�D�y�P(
9�:>��:��;8�#;:�2;�<;MpB;�E;��G;�eH;��H;�H;��H;��H;��H;��H;�H;*�H;�H;��H;��H;��H;��H;��H;��H;��H;��H;��H;��H;��H;�H;+�H;�H;��H;��H;��H;��H;�H;��H;�eH;��G;�E;MpB;�<;<�2;8�#;��;@��:�:`(
98�y��W��	x����6��34�Y�1���J���]�umj�      V���0������ѻ$���ǐ�XX�+6�P	��PuK��>":�M�:,b�:Ki;�%;I�3;߆<;,0B;��E;T\G;�HH;!�H;w�H;>�H;��H;�H;�H;��H;��H;��H;��H;��H;��H;E�H;8�H;8�H;�H;5�H;4�H;C�H;��H;��H;��H;��H;��H;��H;�H;�H;��H;9�H;s�H;#�H;�HH;Y\G;��E;)0B;�<;H�3; �%;Li;0b�:�M�:?":puK�B	��)6�]X�ǐ� ����ѻ��2���      *Q^�X��F�Ƣ)�$+��ζ�D�<�@@S�(n:��:���:��;9�;�M*;ҟ5;uc=;MpB;��E;�JG;-8H;J�H;d�H;��H;�H;b�H;��H;s�H;��H;��H;��H;u�H;[�H;7�H;��H;��H;��H;��H;��H;��H;��H;5�H;Z�H;v�H;��H;��H;��H;n�H;��H;f�H;�H;��H;e�H;M�H;38H;�JG;��E;QpB;qc=;ҟ5;�M*;;�;��;���:��:4n:�@S�T�<��ζ�+�Ӣ)��F�X�      �-.�$�����@~K�@ 
9,]:4�k:IM�:���:�y;��;z $;��/;j�8;��>;�#C;�E;]\G;28H;��H;��H;��H;m�H;�H;g�H;3�H;��H;��H;��H;d�H;�H;��H;��H;��H;�H;v�H;]�H;q�H;{�H;��H;��H;��H;�H;a�H;��H;��H;��H;-�H;j�H;�H;i�H;��H;��H;��H;38H;Y\G;�E;�#C;��>;h�8;��/;| $;��;�y;���:OM�: �k:@]:� 
9PK����L��      ���:�ņ:�ɒ:��:��:���:*��:I�	;�v;��#;��-;��5;zL<;c�@;�(D;DF;��G;�HH;M�H;��H;��H;(�H;��H;=�H;��H;n�H;��H;��H;B�H;�H;��H;��H;U�H;H�H;�H;�H;�H;�H;�H;G�H;R�H;��H;��H;�H;>�H;��H;��H;i�H;��H;9�H;��H;*�H;��H;��H;K�H;�HH;��G;DF;�(D;`�@;}L<;��5;·-;��#;�v;H�	;6��:��:��:��:�ɒ:�ņ:      nW;tx;��;�
;��;�;�� ;n�(;��/;�H6;��;;��?;�C;�PE;��F;��G;�eH;'�H;h�H; �H;,�H;��H;�H;��H;A�H;e�H;i�H;J�H;��H;��H;��H;/�H;��H;��H;��H;��H;��H;��H;��H;��H;��H;)�H;��H;��H;��H;I�H;d�H;b�H;C�H;��H;
�H;��H;,�H;��H;g�H;$�H;�eH;��G;��F;�PE;�C;��?;��;;�H6;��/;t�(;�� ;};��;�
;��;jx;      {S%;�%;��';�M*;۷-;��1;�5;��9;n-=;R@;��B;b�D;mF;�uG;W!H;��H;��H;{�H;��H;j�H;��H;�H;��H;I�H;`�H;W�H;�H;��H;��H;y�H;	�H;��H;��H;�H;p�H;X�H;9�H;T�H;j�H;�H;��H;��H;	�H;x�H;��H;��H;�H;X�H;b�H;E�H;��H;�H;��H;j�H;��H;w�H;��H;�H;W!H;�uG;mF;d�D;��B;
R@;o-=;��9;��5;��1;�-;�M*;��';��%;      fo8;<�8;��9;p�:;{�<;�c>;2R@;�/B;��C;�PE;hzF;=\G;k�G;iH;�H;��H;�H;B�H;
�H;�H;=�H;��H;H�H;S�H;J�H;,�H;��H;��H;S�H;��H;��H;��H;D�H;�H;�H;�H;��H;�H;�H;�H;A�H;��H;��H;��H;N�H;��H;��H;-�H;L�H;O�H;A�H;��H;=�H;�H;�H;>�H;�H;��H;�H;iH;k�G;>\G;lzF;�PE;��C;�/B;0R@;�c>;��<;l�:;��9;2�8;      ��A;EB;�oB;�C;W�C;T�D;@uE;HDF;�F;l�G;�H;�eH;ޡH;��H;.�H;��H;��H;��H;p�H;r�H;�H;F�H;h�H;T�H;�H;��H;��H;Y�H;��H;��H;_�H;0�H;��H;��H;��H;��H;��H;��H;��H;��H;��H;+�H;`�H;��H;��H;W�H;��H;��H;�H;Q�H;d�H;H�H;�H;n�H;n�H;��H;��H;��H;0�H;��H;�H;�eH;�H;l�G;�F;KDF;@uE;K�D;d�C;�C;�oB;FB;      DF;.RF;�zF;͸F;�G;�\G;ղG;*H;�HH;`�H;^�H;��H;��H;��H;��H;�H;��H;�H;��H;0�H;p�H;b�H;Z�H;1�H;��H;v�H;I�H;��H;��H;R�H;�H;��H;��H;��H;e�H;T�H;a�H;N�H;b�H;��H;��H;��H;�H;Q�H;��H;��H;D�H;y�H;��H;.�H;W�H;d�H;o�H;.�H;��H;�H;��H;�H;��H;��H;��H;��H;d�H;`�H;�HH;-H;ԲG;w\G;�G;ԸF;�zF;,RF;      �H;H;�!H;�8H;�TH;-sH;!�H;��H;z�H;��H;W�H;��H;��H;��H;��H;��H;��H;�H;v�H;��H;��H;i�H;�H;��H;��H;H�H;��H;z�H;?�H;�H;��H;��H;U�H;6�H;!�H;��H;�H;��H;�H;8�H;S�H;��H;��H;�H;6�H;w�H;��H;L�H;��H;��H;�H;k�H;��H;��H;s�H;�H;��H;��H;��H;��H;��H;��H;X�H;��H;|�H;��H;�H;'sH;�TH;�8H;�!H;�H;      ��H;
�H;q�H;8�H;�H;z�H;-�H;\�H;��H;�H;��H;��H;��H;��H;��H;7�H;��H;��H;��H;��H;��H;J�H;��H;��H;U�H;��H;w�H;K�H;��H;��H;f�H;<�H;�H;��H;��H;��H;��H;��H;��H;��H;�H;9�H;f�H;��H;��H;H�H;q�H;��H;W�H;��H;��H;I�H;��H;��H;��H;��H;��H;8�H;��H;��H;��H;��H;�H;�H;��H;_�H;+�H;o�H;*�H;6�H;s�H;��H;      ��H;�H;��H;\�H;��H;4�H;��H;��H;��H;��H;��H;��H;�H;��H;��H;�H;�H;��H;��H;��H;I�H;��H;��H;V�H;��H;��H;6�H;��H;��H;b�H;+�H;��H;��H;��H;��H;��H;u�H;��H;��H;��H;��H;��H;+�H;a�H;��H;��H;0�H;��H;��H;P�H;��H;��H;F�H;��H;��H;��H;�H;�H;��H;��H;�H;��H;��H;��H;��H;��H;��H;0�H;��H;\�H;��H;�H;      ��H;��H;�H;T�H;��H;D�H;��H;��H; �H;��H;��H;�H;4�H;\�H;L�H;F�H;.�H;��H;��H;g�H;�H;��H;y�H;��H;��H;M�H;�H;��H;c�H;$�H;��H;��H;��H;~�H;^�H;C�H;7�H;B�H;Z�H;��H;��H;��H;��H;!�H;^�H;��H;��H;O�H;��H;��H;{�H;��H;�H;d�H;��H;��H;.�H;J�H;L�H;[�H;5�H;�H;��H;��H;�H;��H;��H;A�H;��H;X�H;�H;��H;      '�H;]�H;y�H;��H;��H;��H;'�H;S�H;�H;��H;��H;��H;��H;��H;��H;w�H;!�H;��H;z�H;&�H;��H;��H;�H;��H;b�H;	�H;��H;m�H;1�H;��H;��H;}�H;r�H;8�H;�H; �H;�H;�H;�H;;�H;p�H;|�H;��H;��H;+�H;i�H;��H;�H;d�H;��H;�H;��H;��H;�H;z�H;��H;!�H;w�H;��H;��H;��H;��H;��H;��H;��H;T�H;.�H;��H;��H;��H;y�H;[�H;      �H;�H;�H;�H;"�H;@�H;H�H;c�H;j�H;R�H;N�H;7�H;	�H;��H;��H;I�H;��H;��H;`�H; �H;��H;2�H;��H;��H;2�H;��H;��H;?�H;��H;��H;w�H;[�H;;�H;�H;��H;��H;��H;��H;��H;�H;<�H;Z�H;v�H;��H;��H;<�H;��H;��H;3�H;��H;��H;2�H;��H;��H;^�H;��H;��H;L�H;��H;��H;�H;6�H;Q�H;T�H;i�H;b�H;N�H;C�H;2�H;�H;�H;�H;      /�H;%�H;*�H;�H;�H;�H;�H;��H;��H;��H;��H;U�H;�H;��H;l�H;�H;��H;��H;;�H;��H;a�H;�H;��H;G�H;��H;��H;X�H;�H;��H;��H;l�H;;�H;��H;��H;��H;��H;��H;��H;��H;��H;��H;>�H;k�H;��H;��H;�H;U�H;��H;��H;G�H;��H;�H;Z�H;��H;<�H;��H;��H;�H;l�H;��H;�H;U�H;��H;��H;��H;��H;�H;��H;!�H;�H;2�H;#�H;      |�H;v�H;�H;{�H;d�H;=�H;D�H;�H;��H;��H;��H;@�H;�H;��H;t�H;8�H;��H;H�H;��H;��H;P�H;��H;��H;�H;��H;��H;5�H;��H;��H;��H;3�H;�H;��H;��H;��H;��H;��H;��H;��H;��H;��H;�H;4�H;~�H;��H;��H;4�H;��H;��H;�H;��H;��H;K�H;��H;��H;L�H;��H;8�H;s�H;��H;�H;?�H;��H;��H;��H;�H;I�H;=�H;k�H;{�H;��H;��H;      ��H;��H;��H;��H;��H;c�H;U�H;!�H;��H;��H;{�H;=�H;�H;��H;S�H;��H;��H;8�H;��H;��H;!�H;��H;n�H;�H;��H;_�H;�H;��H;��H;a�H;�H;��H;��H;��H;��H;��H;��H;��H;��H;��H;��H;��H;�H;]�H;��H;��H;�H;b�H;��H;�H;q�H;��H;�H;|�H;��H;;�H;��H;��H;P�H;��H;�H;=�H;|�H;��H;��H;"�H;W�H;c�H;��H;��H;��H;��H;      ��H;��H;��H;��H;j�H;V�H;@�H;�H;��H;��H;��H;H�H;��H;��H;5�H;��H;��H;5�H;��H;u�H;�H;��H;T�H;�H;��H;J�H;��H;��H;��H;H�H;�H;��H;��H;��H;��H;��H;��H;��H;��H;��H;��H;��H;�H;C�H;��H;��H;��H;L�H;��H;�H;X�H;��H;�H;r�H;��H;:�H;��H;��H;5�H;��H;��H;G�H;��H;��H;��H;�H;E�H;W�H;m�H;��H;��H;��H;      �H;�H;
�H;��H;��H;��H;r�H;;�H;�H;��H;c�H;!�H;��H;��H;X�H;��H;��H;�H;��H;d�H;�H;��H;=�H;��H;��H;^�H;�H;��H;|�H;>�H;�H;��H;��H;��H;��H;��H;y�H;��H;��H;��H;��H;��H;�H;:�H;v�H;��H;�H;_�H;��H;��H;?�H;��H;�H;`�H;��H;�H;��H;��H;X�H;��H;��H; �H;f�H;��H;	�H;=�H;y�H;��H;��H;��H;
�H;�H;      ��H;��H;��H;��H;k�H;Y�H;>�H;�H;��H;��H;��H;H�H;��H;��H;5�H;��H;��H;5�H;��H;u�H;�H;��H;T�H;�H;��H;J�H;��H;��H;��H;F�H;�H;��H;��H;��H;��H;��H;��H;��H;��H;��H;��H;��H;�H;B�H;��H;��H;��H;M�H;��H;�H;X�H;��H;�H;r�H;��H;:�H;��H;��H;5�H;��H;��H;G�H;��H;��H;��H;�H;D�H;V�H;q�H;��H;��H;��H;      ��H;��H;��H;��H;��H;^�H;S�H;#�H;��H;��H;z�H;=�H;�H;��H;S�H;��H;��H;:�H;��H;��H;!�H;��H;n�H;�H;��H;^�H;�H;��H;��H;`�H;�H;��H;��H;��H;��H;��H;��H;��H;��H;��H;��H;��H;�H;Z�H;��H;��H;�H;a�H;��H;�H;p�H;��H;�H;|�H;��H;;�H;��H;��H;N�H;��H;�H;?�H;z�H;��H;��H;(�H;\�H;]�H;��H;��H;��H;��H;      |�H;u�H;}�H;|�H;e�H;B�H;B�H;�H;��H;��H;��H;@�H;�H;��H;v�H;6�H;��H;J�H;��H;��H;O�H;��H;��H;�H;��H;��H;6�H;��H;��H;��H;3�H;�H;��H;��H;��H;��H;��H;��H;��H;��H;��H;�H;3�H;~�H;��H;��H;2�H;��H;��H;�H;��H;��H;H�H;��H;��H;J�H;��H;9�H;t�H;��H;�H;?�H;��H;��H;��H;�H;K�H;>�H;m�H;}�H;��H;u�H;      -�H;)�H;*�H;�H;�H;�H;�H;��H;��H;��H;��H;X�H;�H;��H;o�H;�H;��H;��H;>�H;��H;^�H;�H;��H;G�H;��H;��H;T�H;�H;��H;��H;k�H;:�H;��H;��H;��H;��H;��H;��H;��H;��H;��H;>�H;l�H;��H;��H;�H;T�H;��H;��H;C�H;��H;�H;W�H;��H;>�H;��H;��H;�H;l�H;��H;�H;T�H;��H;��H;��H;��H;�H; �H;�H;"�H;3�H;#�H;      �H;�H;�H;�H;"�H;O�H;K�H;d�H;i�H;R�H;O�H;6�H;�H;��H;��H;L�H;��H;��H;`�H;��H;��H;4�H;��H;��H;3�H;��H;�H;?�H;��H;��H;u�H;X�H;;�H;�H;��H;��H;��H;��H;��H;�H;;�H;Z�H;u�H;��H;��H;;�H;~�H;��H;0�H;��H;��H;2�H;��H;��H;`�H;��H;��H;J�H;��H;��H;�H;6�H;N�H;T�H;j�H;c�H;N�H;C�H;(�H;�H;�H;�H;      �H;]�H;v�H;��H;��H;��H;$�H;S�H;��H;��H;��H;��H;��H;��H;��H;x�H;#�H;��H;z�H;"�H;��H;��H;�H;��H;d�H;�H;��H;j�H;1�H;��H;��H;|�H;p�H;8�H;�H;�H;�H; �H;�H;:�H;o�H;|�H;��H;��H;*�H;h�H;��H;�H;_�H;��H;�H;��H;��H;"�H;|�H;��H;#�H;w�H;��H;��H;��H;��H;��H;��H;�H;U�H;*�H;��H;��H;��H;~�H;[�H;      ��H;��H;
�H;^�H;��H;N�H;��H;��H;�H;��H;��H;�H;5�H;\�H;P�H;J�H;/�H;��H;��H;h�H;�H;��H;x�H;��H;��H;H�H;�H;��H;c�H;#�H;��H;��H;��H;~�H;^�H;B�H;5�H;C�H;Z�H;~�H;��H;��H;��H; �H;\�H;��H;��H;O�H;��H;��H;|�H;��H;�H;b�H;��H;��H;-�H;I�H;L�H;[�H;4�H; �H;��H;��H;�H;��H;��H;@�H;��H;c�H;�H;��H;      ��H;�H;	�H;Y�H;��H;8�H;��H;��H;��H;��H;��H;��H;�H;��H;��H;�H;�H;��H;��H;��H;J�H;��H;��H;V�H;��H;��H;3�H;��H;��H;_�H;*�H;��H;��H;��H;��H;��H;s�H;��H;��H;��H;��H;��H;+�H;_�H;��H;��H;2�H;��H;��H;N�H;��H;��H;E�H;��H;��H;��H;�H;�H;��H;��H;�H;��H;��H;��H;��H;��H;��H;3�H;��H;Y�H;	�H;�H;      ��H;��H;f�H;6�H;�H;��H;+�H;d�H;�H;�H;�H;��H;��H;�H;��H;:�H;��H;��H;��H;��H;��H;L�H;��H;��H;W�H;��H;t�H;J�H;��H;��H;h�H;<�H;�H;��H;��H;��H;��H;��H;��H;��H;�H;;�H;h�H;��H;��H;F�H;r�H;��H;S�H;��H;��H;I�H;��H;��H;��H;��H;��H;7�H;��H;��H;��H;��H;�H;�H;��H;]�H;+�H;q�H;*�H;6�H;s�H;��H;      �H;H;�!H;�8H;�TH;4sH;!�H;��H;|�H;��H;X�H;��H;��H;��H;��H;��H;��H; �H;u�H;��H;��H;l�H;�H;��H;��H;E�H;��H;z�H;=�H;�H;��H;��H;S�H;5�H; �H;��H;�H;��H;�H;8�H;T�H;��H;��H;�H;6�H;t�H;��H;L�H;��H;��H;�H;l�H;��H;��H;s�H;�H;��H;��H;��H;��H;��H;��H;W�H;��H;{�H;��H;"�H;.sH;�TH;�8H;�!H;�H;      DF;,RF;�zF;øF;�G;�\G;βG;-H;�HH;`�H;d�H;��H;��H;��H;��H;�H;��H;�H;��H;.�H;s�H;b�H;V�H;1�H;��H;r�H;E�H;��H;��H;O�H;�H;��H;��H;��H;e�H;P�H;b�H;S�H;b�H;��H;��H;��H;	�H;Q�H;��H;��H;G�H;y�H;��H;0�H;Z�H;d�H;p�H;0�H;��H;�H;��H;�H;��H;��H;��H;��H;a�H;_�H;�HH;&H;βG;w\G;�G;ɸF;}zF;RF;      ��A;AB;�oB;�C;V�C;W�D;@uE;JDF; �F;n�G;�H;�eH;ޡH;��H;4�H;��H;��H;��H;p�H;o�H;�H;H�H;d�H;T�H;�H;��H;��H;W�H;��H;��H;_�H;/�H;��H;��H;��H;��H;��H;��H;��H;��H;��H;0�H;d�H;��H;��H;U�H;��H;��H;�H;S�H;h�H;I�H;�H;o�H;p�H;��H;��H;��H;1�H;��H;ޡH;�eH;�H;k�G;�F;JDF;?uE;I�D;`�C;�C;�oB;AB;      Co8;"�8;��9;t�:;x�<;�c>;1R@;�/B;��C;�PE;lzF;A\G;l�G;iH;�H;��H;�H;B�H;�H;�H;>�H;��H;A�H;Q�H;L�H;%�H;��H;��H;R�H;��H;��H;��H;D�H;�H;�H;�H;��H;�H;�H;�H;G�H;��H;��H;��H;P�H;��H;��H;,�H;I�H;S�H;E�H;��H;=�H;�H;
�H;>�H;�H;��H;�H;iH;i�G;<\G;kzF;�PE;��C;�/B;1R@;�c>;��<;��:;��9;�8;      bS%;��%;�';�M*;շ-;~�1;ܟ5;��9;t-=;R@;��B;d�D;mF;�uG;Y!H;�H;��H;{�H;��H;j�H;��H;�H;��H;H�H;b�H;P�H;�H;��H;��H;u�H;	�H;��H;��H;~�H;m�H;X�H;<�H;V�H;k�H;~�H;��H;��H;�H;{�H;��H;��H;�H;X�H;`�H;F�H;��H;�H;��H;l�H;��H;v�H;��H;��H;X!H;�uG;mF;`�D;��B;
R@;n-=;��9;ڟ5;~�1;׷-;�M*;�';��%;      jW;tx;��;�
;��;�;�� ;t�(;��/;�H6;��;;��?;�C;�PE;��F;��G;�eH;'�H;g�H;��H;,�H;��H;�H;��H;E�H;]�H;g�H;J�H;��H;��H;��H;,�H;��H;��H;��H;��H;��H;��H;��H;��H;��H;/�H;��H;��H;��H;I�H;i�H;d�H;A�H;��H;�H;��H;.�H; �H;g�H;$�H;�eH;��G;��F;�PE;�C;��?;��;;�H6;��/;r�(;�� ;n;��;�
;��;jx;      ���:�ņ:�ɒ:��:��: ��:0��:I�	;�v;��#;��-;��5;|L<;a�@;�(D;DF;��G;�HH;K�H;��H;��H;*�H;��H;;�H;��H;g�H;��H;��H;?�H;�H;��H;��H;S�H;I�H;�H;
�H;�H;�H;�H;E�H;U�H;��H;��H;�H;?�H;��H;��H;k�H;��H;=�H;��H;(�H;��H;��H;K�H;�HH;��G;DF;�(D;`�@;zL<;��5;��-;��#;�v;L�	;0��:��:��:!��:�ɒ:�ņ:      �-.�����깐~K�  
9@]:4�k:]M�:���:�y;��;| $;��/;h�8;��>;�#C;�E;[\G;08H;��H;��H;��H;j�H;�H;j�H;,�H;��H;��H;��H;`�H;�H;��H;��H;��H;}�H;r�H;^�H;t�H;|�H;��H;��H;��H; �H;b�H;��H;��H;��H;0�H;g�H;�H;m�H;��H;��H;��H;08H;Y\G;�E;�#C;��>;d�8;��/;x $;��;�y;���:MM�:�k: ]:` 
90K������      )Q^�X��F�ʢ)�&+��ζ�T�<��@S�4n:��:���:��;9�;�M*;ԟ5;uc=;MpB;��E;�JG;/8H;M�H;e�H;��H;�H;f�H;��H;n�H;��H;��H;��H;v�H;[�H;7�H;��H;��H;��H;��H;��H;��H;��H;7�H;[�H;y�H;��H;��H;��H;r�H;��H;b�H;�H;��H;d�H;K�H;28H;�JG;��E;KpB;pc=;ҟ5;�M*;8�;��;���:��:(n: AS�`�<��ζ�&+�ɢ)��F�X�      \���,��� ���ѻ ���ǐ�ZX�&6�F	��puK��>":�M�:,b�:Ki;!�%;K�3;��<;)0B;��E;V\G;�HH;#�H;y�H;>�H;��H;�H;�H;��H;��H;��H;��H;��H;��H;E�H;5�H;5�H;�H;7�H;4�H;C�H;��H;��H;��H;��H;��H;��H;�H;�H;��H;<�H;z�H;!�H;�HH;Y\G;��E;)0B;��<;I�3;!�%;Ii;*b�:�M�:?":�uK�H	��)6�^X�ǐ� ����ѻ$��.���      n�n�wmj���]���J�X�1�34�5������	x��W�@�y�`(
9ꨂ:<��:��;8�#;;�2;�<;KpB;�E;��G;�eH;��H;�H;��H;��H;��H;��H;�H;'�H;�H;��H;��H;��H;��H;��H;��H;��H;��H;��H;��H;��H;�H;*�H;�H;��H;��H;��H;��H;�H;��H;�eH;��G;�E;KpB;�<;;�2;8�#;��;<��:�:0(
9L�y��W��	x����8��34�Z�1���J���]�vmj�      ><ͼ~�ɼ�����֯�ζ��ㄼ��Y��*�����s��X��rѺ���>Q:���:��
;2�#;K�3;qc=;�#C;DF;��G;��H;��H;��H;�H;��H;4�H; �H;D�H;q�H;G�H;�H;6�H;��H;��H;��H;��H;��H;2�H;�H;F�H;s�H;G�H; �H;7�H;��H;�H;��H;��H;�H;��G;DF;�#C;pc=;I�3;4�#;��
;���:�>Q:���rѺX��s������*���Y�ㄼζ���֯�����~�ɼ      ��'�'�$����{��  ���ۼ����+����]��X!�C>ۻ�+��}*�`����>:���:��;�%;Ο5;|�>;�(D;��F;[!H;�H;+�H;��H;��H;��H;��H;M�H;��H;��H;j�H;q�H;J�H;2�H;Q�H;4�H;I�H;p�H;j�H;��H;��H;M�H;��H;��H;��H;��H;)�H;�H;Y!H;��F;(D;~�>;̟5;�%;��;���:��>:h��~*��+��D>ۻ�X!���]��+�������ۼ�  �|����(�$�      Ÿ���v����w�f�c��J�̈́-�{��;缄沼ㄼ��;������j���5�H��?Q:8��:Ki;�M*;f�8;h�@;�PE;�uG;iH;��H;��H;��H;��H;��H;W�H;��H;��H;��H;��H;��H;��H;��H;��H;��H;��H;��H;��H;��H;\�H;��H;��H;��H;��H;��H;iH;�uG;�PE;`�@;j�8;�M*;Li;<��:�>Q:P�깦5��j��������;�ㄼ�沼�;�|�̈́-��J�f�c���w��v��      yHͽ֪ɽ�;��"����Ǹ����[�z0�r��%<ͼʾ��b�J�����j��z*�p�訂:0b�:6�;��/;�L<;�C;mF;o�G;ޡH;��H;��H;��H;�H;4�H;��H;�H;�H;��H;��H;��H;��H;��H;��H;��H;�H;�H;��H;6�H; �H;��H;��H;��H;ۡH;m�G;mF;�C;yL<;��/;5�;0b�:ꨂ:��z*��j�����b�J�ʾ��&<ͼr��z0���[�Ǹ����"���;��֪ɽ      ��!-������ѱ�ƽ]P���v���J�G����ۼ��b�J������+���rѺ (
9�M�:��;x $;��5;��?;b�D;@\G;�eH;��H;��H;��H;��H;��H;��H;2�H;U�H;=�H;3�H;D�H;�H;F�H;2�H;=�H;T�H;2�H;��H;�H;��H;��H;��H;��H;�eH;@\G;f�D;��?;��5;z $;��;�M�:0(
9�rѺ�+������b�J�����ۼG���J��v��]P��ƽұ轃����!-�       j�Vde�Y0X�D�e{+�������t㻽Y���RDX������ۼʾ����;�D>ۻX�h�y��>":���:��;·-;��;;��B;lzF;�H;`�H;S�H;��H;��H;��H;��H;M�H;��H;~�H;q�H;��H;\�H;��H;q�H;~�H;��H;M�H;��H;��H;��H;�H;T�H;^�H;�H;mzF;��B;��;;��-;��;���:�>":\�y�X�E>ۻ��;�˾����ۼ���RDX�Y���t㻽��콂��f{+�D�Y0X�Vde�      ��Ph��k���I���|x���O��C(���Ϊɽ����RDX�G��&<ͼㄼ�X!��s���W��uK���:�y;��#;�H6;R@;�PE;i�G;\�H;��H;�H;��H;��H;��H;R�H;��H;��H;��H;��H;��H;��H;��H;��H;��H;R�H;��H;��H;��H;
�H;��H;\�H;g�G;�PE;R@;�H6;��#;�y;��:�uK��W��s���X!�ㄼ&<ͼG��RDX�����Ϊɽ���C(���O��|x��I��k��Ph��      >����������"�;hɰ��G��	 j�8�5��	�ΪɽY����J�s���沼��]�����	x�\	��n:���:�v;��/;g-=;��C;�F;�HH;x�H;��H;��H;�H;~�H;f�H;��H;��H;��H;��H;�H;��H;��H;��H;��H;g�H;}�H;�H;��H;��H;|�H;�HH;�F;��C;j-=;��/;�v;���:n:T	���	x������]��沼s���J�Y���Ϊɽ�	�8�5�	 j��G��hɰ�"�;��徶���      �2�U�-�"�-E�����?Kɾj����s�8�5���u㻽�v��	z0��;��+���*����86�@BS�GM�:O�	;n�(;�9;�/B;HDF;H;��H;Z�H;��H;��H;M�H;c�H;��H;�H;�H;�H;9�H;�H;�H;�H;��H;b�H;M�H;��H;��H;]�H;��H;#H;HDF;�/B;��9;p�(;I�	;QM�:�BS�16�����*��+���;�	z0��v��u㻽��8�5���s�j��?Kɾ����-E�"�U�-�      %3s�cm�:�\�h�C�5�%����TҾj��	 j��C(����]P����[�|������Y�8��hX�p�<� �k:2��:�� ;ԟ5;0R@;5uE;ͲG;�H;�H;��H;��H;!�H;F�H;�H;B�H;L�H;7�H;m�H;6�H;N�H;A�H;�H;G�H;!�H;��H;��H;"�H;�H;ԲG;5uE;2R@;؟5;�� ;*��:�k:p�<�dX�8����Y����|���[�]P����콪C(�	 j�j���TҾ��5�%�h�C�:�\�cm�      �ޞ�������_F�>�W�W�-���?Kɾ�G����O����ƽǸ��̈́-���ۼㄼ44�ǐ�϶� ]:��:z;|�1;�c>;B�D;w\G;)sH;v�H;4�H;F�H;��H;K�H;
�H;I�H;j�H;\�H;��H;^�H;k�H;H�H;
�H;M�H;��H;H�H;:�H;{�H;.sH;\G;D�D;�c>;~�1;|;��:0]:϶�ǐ�44�ㄼ��ۼ̈́-�Ǹ��ƽ�����O��G��?Kɾ��W�-�>�W�_F�������      ��ſ���Lw���ޞ�����?�W�5�%�����hɰ��|x�e{+�ѱ����J��  �ζ��Y�1�+���!+�@ 
9��:��;߷-;��<;[�C;�G;�TH;!�H;��H;��H;��H;)�H;�H;g�H;��H;u�H;��H;q�H;��H;a�H;�H;)�H;��H;��H;��H;'�H;�TH;�G;[�C;��<;߷-;��;��:` 
9!+�(���Z�1�ζ���  ��J���ѱ�e{+��|x�hɰ�����5�%�>�W������ޞ�Lw�����      ������Կp���ޞ�`F�g�C�-E�"�;�I��D���"��f�c�|��֯���J��ѻТ)��K���:�
;�M*;j�:;�C;ƸF;�8H;+�H;G�H;X�H;��H;�H;�H;��H;��H;��H;��H;��H;��H;|�H;�H;�H;��H;_�H;K�H;-�H;�8H;ѸF;�C;m�:;�M*;�
;��:pK�Ѣ)��ѻ��J��֯�|�f�c�"����D��I��"�;-E�h�C�`F��ޞ�p���Կ��      ����������ԿLw�����:�\�"����k��Y0X�����;����w����������]�!���F�����ɒ:��; �';��9;�oB;�zF;�!H;s�H;��H;�H;p�H;�H;�H;�H;��H;��H;��H;��H;��H;}�H;�H;�H;l�H;�H;��H;u�H;�!H;�zF;�oB;��9;��';��;�ɒ:����F� �黫�]����������w��;�����Y0X�k�����"�:�\����Lw���Կ��𿝏�       $�������忇�����cm�V�-�����Ph��Vde�"-�תɽ�v��'�$��ɼzmj�9���X� ���ņ:dx;�%;2�8;EB;RF;�H;�H;�H;��H;C�H;�H;�H;v�H;��H;��H;�H;��H;��H;v�H;�H;�H;A�H;��H;�H;�H;�H;-RF;BB;0�8;�%;dx;�ņ:��X�6���zmj��ɼ'�$��v��֪ɽ"-�Vde�Ph������V�-�cm��������忝����      �>���8���*�O������˿p��E�b�C\�4m־^��Q�:��J�)��E�B�<��������1/��R���ܑ>:kt�:p ;�J6;�DA;[IF;�NH;��H;�!I;�I;�I;|I;NI;�I;I I;��H;�H;��H;H I;�I;NI;|I;�I;�I;�!I;��H;�NH;hIF;�DA;�J6;
p ;it�:ܑ>:F���1/���������<��E�B�)���J�Q�:�^��4m־C\�E�b�p���˿����O���*���8�      ��8��4��g&�6��<����<ƿ񲗿�>]����O�Ѿ�p���*7����%W��LR?��|�q8�������օ����G:s �:�!;�6;�kA;fYF;�TH;D�H;�!I;�I;�I;eI;(I;�I;; I;��H;��H;��H;> I;�I;)I;gI;�I;�I;�!I;F�H;�TH;rYF;�kA;�6;�!;q �:��G:̅�������q8�� }�LR?�%W�����*7��p��O�Ѿ����>]�񲗿�<ƿ<���6���g&��4�      ��*��g&��#�t�T[�qL�������M�r5��>ľ����,��D�蒐��5�2�ݼ���q
��x�(uk���b:'l�:�#;ė7;V�A;��F;�dH;�I;""I;�I;GI;I;�I;�I;��H;Y�H;��H;R�H;��H;�I;�I;I;AI;�I;#"I;�I;�dH;��F;T�A;��7;�#;%l�:��b:uk��x��q
���2�ݼ�5�蒐��DὫ�,����>ľr5���M����qL��T[�t��#��g&�      O�6��t����˿@1��7�y�Î6��z �����2�l�+��ͽ#�����&���˼?�k�#�����X��� �t��:8�;�&;~9;m�B;��F;�}H;�	I;/"I;I;�I;{I;UI;%I;��H;�H;a�H;��H;��H;"I;RI;{I;�I;I;2"I;�	I;�}H;��F;j�B;y9;�&;6�;p��:� ���X�!���?�k���˼��&�#����ͽ+�2�l������z �Î6�7�y�@1���˿���t�6��      ����<���T[忶˿�T���{�R�����E۾ӗ����M���	������j��3�d����O�<�׻��/�`��=��:� 
;�*;P;;�jC;�'G;ԛH;�I;�!I;�I;wI;�
I;�I;�I;!�H;��H;��H;��H;"�H;�I;�I;�
I;sI;�I;�!I;�I;כH;�'G;�jC;H;;�*;� 
;9��:(����/�:�׻��O�d���3���j������	���M�ӗ���E۾���{�R���T���˿T[�<���      �˿�<ƿqL��@1����>]���)��$��ֳ���{���,�q��'��Q`I��J���,���3/�,��� ��,69�4�:҄;�o.;.=;?aD;��G;Q�H;�I;!I;AI;,I;�	I;�I;� I;��H;��H;C�H;��H;��H;� I;�I;�	I;)I;CI;!I;�I;P�H;��G;=aD;.=;�o.;΄;�4�: -69� � ,���3/��,���J��Q`I�'��q�齥�,���{�ֳ��$����)��>]��@1��qL���<ƿ      p��񲗿���7�y�{�R���)�nv��>ľ^���I�Xl����������&�ӮҼ�}�2B�̮�����p�!:�*�: z;[3;Kj?;s\E;��G;��H;KI;I;mI;�I;XI;�I;��H;��H;C�H;��H;A�H;��H;��H;�I;WI;�I;pI;I;HI;��H;��G;s\E;Dj?;W3; z;�*�:��!:���̮��1B��}�ӮҼ��&��������Xl��I�^���>ľnv���)�{�R�7�y����񲗿      E�b��>]���M�Î6�����$���>ľ#q��y�Z�+�Q9ݽ W����L����"F���G��׻;�@o�zȊ:�i; P$;��7;T�A;�IF;CH;��H;� I;EI;WI;�I;	I;�I;��H;��H;t�H;��H;r�H;��H;��H;I;I;�I;ZI;EI;� I;��H;CH;�IF;M�A;��7; P$;zi;�Ȋ:Ho�;��׻�G�"F�������L� W��Q9ݽ+�y�Z�#q���>ľ�$�����Î6���M��>]�      C\����r5��z ��E۾ֳ�^��y�Z�K?#����A����j�%��Dϼ�����˵���lۺX9�9^4�:>�;A�,;U�;;�C;~G;�H;�I;�!I;�I;%I;I;sI;$I;��H;��H;��H;�H;��H;��H;��H;#I;sI;I;'I;�I;�!I;I;�H;G;�C;W�;;D�,;;�;n4�:X9�9�lۺʵ�������Dϼ%����j��A�����K?#�y�Z�^��ֳ��E۾�z �r5����      4m־O�Ѿ�>ľ����җ����{��I�+����V���{�>�/�%���,��?=�D�һp�@�L� ���k:��:�a;��3;	j?;Q2E;��G;A�H;I;P I;�I;�I; 	I;�I;��H;��H;��H;��H;9�H;��H;��H;��H;��H;�I; 	I;�I;�I;N I;I;>�H;��G;M2E;	j?;��3;�a;��:��k:@� �k�@�B�һ>=��,��$��>�/��{��V�����+��I���{�җ�������>ľO�Ѿ      ^���p����2�l���M���,�Xl�Q9ݽ�A���{���5��J��	;���T[�"?�����bP�� P�9��:��;
*;�9;4kB;��F;TNH;V�H; I;iI;�I; I;�I;!I;F�H;��H;��H;��H;I�H;��H;��H;��H;D�H;!I;�I;I;�I;iI;�I;S�H;YNH;��F;5kB;�9;
*;��;��:P�9VP������"?��T[�;���J����5��{��A��Q9ݽXl���,���M�2�l����p��      Q�:��*7���,�+���	�q�齂��� W����j�>�/��J���I���k�l�.��e��H���Ȋ:)o�:�;@r3;��>;�D;M�G;!�H;�I;!I;�I;cI;b
I;�I;A I;��H;z�H;��H;��H;A�H;��H;��H;|�H;��H;? I;�I;g
I;mI;�I;!I;�I;%�H;L�G;�D; �>;Br3;�;-o�:�Ȋ:��d��.��k��k��I���J��>�/���j� W������q�齂�	�+���,��*7�      �J�����D��ͽ���'�������L�%��$��;���k����kI����/��/��>:��:�B;=�,;��:;
�B;jxF;u<H;��H;�I;tI;�I;I;�I;�I;p�H;Z�H;�H;O�H;�H;N�H;�H;N�H;�H;W�H;n�H;�I;�I;I;�I;pI;�I;��H;t<H;kxF;�B;��:;H�,;�B;��:4�>:�/���/�jI������k�;��$��$����L����'������ͽ�D����      (��$W��璐�"�����j�Q`I���&����Dϼ�,���T[�k�lI��e;��nk�x:�4�:�;�&;��6;�!@;2E;��G;�H;�I;� I;2I;�I;�
I;I;Q I;��H;��H;��H;@�H;v�H;'�H;v�H;@�H;��H;��H;��H;V I;I;�
I;�I;.I;� I;�I;|�H;��G;2E;�!@;��6;�&;�;�4�:t:�nk�a;�kI��k��T[��,��Cϼ�����&�Q`I���j�#���璐�$W��      D�B�LR?��5���&��3��J��ӮҼ!F����>=�"?�.����/��nk�ح�9 ׳:��;!;93;��=;��C;��F;�cH;��H;lI;�I;�I;I;�I;�I;"�H;��H;u�H;`�H;!�H;g�H;�H;e�H; �H;b�H;u�H;��H;%�H;�I;�I;I;�I;�I;nI;��H;�cH;��F;��C;��=;=3;!;��;"׳:ح�9�nk���/�.�� ?�>=� ��!F��ҮҼ�J���3���&��5�LR?�      9���|�0�ݼ��˼d���,���}� �G����B�һ����f���/�t:&׳:��;Pb;��0;m<;�B;�IF;IH;�H;�I;M I;�I;I;9
I;�I; I;�H;8�H;��H;	�H;�H;]�H;�H;\�H;�H;�H;��H;6�H;�H; I;�I;:
I;I;�I;O I;�I;�H;IH;�IF;��B;p<;��0;Sb;��;(׳:t:�/�d������A�һ��� �G��}��,��d����˼0�ݼ�|�      ���o8����>�k���O��3/�/B��׻ǵ��d�@�NP�� ��4�>:�4�:��;Tb;��/;;;�A;g�E;��G;ЭH;�
I;E I;�I;�I;�I;�I;�I;f�H;�H;��H;}�H;��H;��H;Q�H;�H;M�H;��H;��H;x�H;��H;�H;i�H;�I;�I;�I;�I;�I;D I;�
I;ЭH;��G;k�E;�A;;;��/;Tb;��;�4�:0�>:��FP��d�@�ŵ���׻0B��3/���O�@�k���n8��      ������q
����4�׻�+��Ʈ�� ;��lۺ0� � P�9�Ȋ:��:�;!;��0;;;��A;�pE;M�G;��H;��H;�I;I;.I; I;�I;VI;��H;#�H;X�H;��H; �H;��H;��H;G�H;�H;D�H;��H;��H;��H;��H;[�H;(�H;��H;SI;�I;�I;0I;I;�I;��H;��H;S�G;�pE;��A;;;��0;!;�;��:�Ȋ:XP�90� ��lۺ�;�Ȯ���+��1�׻����q
���      $/��"����x���X���/�� ���� o치9�9��k:��:/o�:�B;�&;=3;p<;�A;�pE;BtG;�|H;�H;I;RI;#I;�I;K
I;�I;3 I;-�H;�H;��H;`�H;��H;��H;��H;X�H;E�H;W�H;��H;��H;��H;]�H;��H;�H;*�H;3 I;�I;G
I;�I;#I;JI;I;
�H;�|H;BtG;�pE; �A;m<;?3;�&;�B;/o�:��:��k:�9�9o����� ���/���X��x�"���      F���օ���tk��� �H��@-69��!:�Ȋ:n4�:��:��;�;C�,;��6;��=;��B;n�E;W�G;�|H;u�H;WI;�I;bI;9I;�I;I;hI;'�H;��H;�H;��H;��H;��H;��H;��H;n�H;U�H;j�H;��H;��H;��H;��H;��H;�H;��H;*�H;cI;I;�I;6I;\I;�I;ZI;u�H;�|H;T�G;m�E;��B;��=;��6;C�,;�;��;��:z4�:�Ȋ:��!:�-69(��� �$uk��      l�>:D�G:t�b:n��:%��:�4�:�*�:�i;;�;�a;
*;=r3;��:;�!@;��C;�IF;��G;��H;�H;TI;�I;I;I;�I;�I;<I;��H;m�H;��H;X�H;*�H;��H;}�H;��H;��H;��H;c�H;��H;��H;��H;y�H;��H;-�H;[�H;��H;k�H;��H;7I;�I;�I;I;I;�I;TI;
�H;��H;��G;�IF;��C;�!@;��:;?r3;*;�a;;�;|i;�*�:�4�:=��:h��:��b:D�G:      kt�:� �:Gl�:N�;� 
;Ԅ;"z;�O$;J�,;��3;�9; �>;�B;2E; �F;PH;խH;��H;	I;�I;$I;\I;I;�I;�I;��H;�H;0�H;��H;x�H;��H;��H;t�H;��H;�H;��H;��H;��H;�H;��H;o�H;��H;��H;x�H;��H;0�H;��H;��H;�I;�I;I;]I;$I;�I;I;��H;խH;LH; �F;2E;�B;�>;�9;��3;J�,;P$;&z;҄;� 
;B�;1l�: �:      *p ;�!;�#;�&;�*;�o.;j3;��7;^�;;j?;;kB;	�D;kxF;��G;�cH;�H;�
I;�I;RI;aI;I;I;�I;:I;�H;q�H;p�H;�H;��H;��H;��H;d�H;u�H;��H;9�H;�H;��H;��H;5�H;��H;q�H;c�H;��H;��H;��H;�H;k�H;q�H;�H;6I;�I;I;I;aI;QI;�I;�
I;�H;�cH;��G;kxF;�D;@kB;
j?;a�;;��7;g3;�o.;�*;�&;�#;�!;      �J6;�6;��7;~9;B;;.=;Kj?;Q�A;�C;N2E;��F;M�G;r<H;�H;��H;�I;E I;I;%I;6I;�I;�I;:I;0�H;��H;��H;A�H;�H;�H;��H;h�H;T�H;v�H;�H;��H;T�H;*�H;O�H;��H;	�H;s�H;Q�H;h�H;��H;�H;�H;:�H;��H;��H;,�H;2I;�I;�I;3I;"I;I;D I;�I;��H;|�H;o<H;L�G;��F;N2E;�C;X�A;Ej?;.=;P;;|9;��7;�6;      EA;�kA;O�A;k�B;�jC;PaD;{\E;�IF;�G;��G;]NH;+�H;��H;�I;rI;V I;�I;9I;�I;�I;�I;�I;�H;��H;��H;b�H;�H;/�H;��H;y�H;M�H;e�H;��H;?�H;��H;��H;��H;��H;��H;B�H;��H;_�H;N�H;x�H;��H;/�H;�H;`�H;��H;��H;�H;�I;�I;�I;�I;5I;�I;W I;qI;�I;��H;.�H;aNH;��G;�G;�IF;{\E;CaD;�jC;m�B;M�A;�kA;      [IF;sYF;��F;��F;v'G;��G;��G;CH; �H;F�H;W�H;�I;�I;� I;�I;�I;�I; I;J
I;I;=I;��H;r�H;��H;_�H;8�H;D�H;��H;|�H;\�H;F�H;��H;�H;}�H;6�H;�H;�H;�H;2�H;}�H;�H;��H;F�H;Y�H;x�H;��H;?�H;<�H;`�H;��H;n�H;��H;<I;I;J
I;�I;�I;�I;�I;� I;�I;�I;^�H;H�H;#�H;CH;��G;��G;�'G;��F;��F;pYF;      �NH;�TH;�dH;�}H;ϛH;T�H;��H;��H;�I;I;�I;!I;lI;.I;�I;I;�I;�I;�I;jI;�H;�H;s�H;G�H;�H;C�H;��H;�H;N�H;M�H;��H;��H;U�H;��H;��H;��H;w�H;��H;��H;��H;S�H;��H;��H;J�H;G�H;}�H;��H;F�H;�H;C�H;p�H;�H;�H;hI;�I;�I;�I;I;�I;,I;oI;!I;  I;I;�I;��H;��H;O�H;�H;�}H;�dH;{TH;      ��H;L�H;�I;�	I;�I;�I;VI;� I;�!I;U I;lI;�I;�I;�I;�I;:
I;�I;PI;4 I;(�H;n�H;.�H;	�H;�H;+�H;��H;�H;]�H;D�H;u�H;��H;2�H;��H;q�H;3�H;�H;��H;��H;0�H;r�H;��H;/�H;��H;s�H;?�H;\�H;x�H;��H;/�H;�H;	�H;0�H;m�H;'�H;1 I;PI;�I;:
I;�I;�I;�I;�I;mI;R I;�!I;� I;UI;�I;�I;�	I;�I;@�H;      �!I;�!I;"I;D"I;�!I;!I;�I;GI;�I;�I;�I;lI;I;�
I;�I;�I;�I;��H;3�H;��H;��H;��H;��H;!�H;��H;v�H;G�H;D�H;��H;��H;#�H;��H;A�H;��H;��H;��H;��H;��H;��H;��H;@�H;��H;"�H;��H;��H;C�H;C�H;v�H;��H;�H;��H;��H;��H;��H;1�H;��H;�I;�I;�I;�
I;I;jI;�I;�I;�I;GI;�I;!I;�!I;D"I;!"I;�!I;      �I;I;�I;I;�I;?I;nI;ZI;%I;�I;I;i
I;�I;I;�I; I;l�H;"�H;�H;!�H;b�H;y�H;��H;��H;x�H;V�H;L�H;w�H;��H;�H;��H;<�H;��H;��H;a�H;@�H;/�H;@�H;\�H;��H;��H;:�H;��H;�H;��H;v�H;F�H;X�H;y�H;��H;��H;y�H;[�H;�H;�H;!�H;l�H; I;�I;I;�I;g
I;I;�I;$I;WI;qI;<I;�I;I;�I;I;      �I;�I;LI;�I;vI;,I;�I;�I;
I;	I;�I;�I;�I;X I;(�H;�H;%�H;`�H;��H;��H;6�H;��H;��H;n�H;Q�H;I�H;��H;��H;)�H;��H;�H;��H;m�H;1�H;�H;��H;��H;��H;�H;4�H;m�H;��H;�H;��H;"�H;��H;��H;I�H;Q�H;j�H;��H;��H;0�H;��H;��H;^�H;$�H;�H;%�H;W I;�I;�I;�I;	I;I;�I;�I;"I;�I;�I;NI;�I;      }I;pI;I;vI;�
I;�	I;XI;
I;wI;�I;"I;C I;q�H;��H;��H;9�H;��H;��H;e�H;��H;��H;��H;e�H;U�H;h�H;��H;��H;7�H;��H;?�H;��H;L�H;�H;��H;��H;��H;��H;��H;��H;��H;�H;J�H;��H;=�H;��H;2�H;��H;��H;h�H;N�H;j�H;��H;��H;��H;d�H;��H;��H;<�H;��H;��H;p�H;C I;%I;�I;vI;I;`I;�	I;�
I;yI;I;oI;      YI;6I;�I;XI;�I;�I;�I;|I;I;��H;F�H;��H;Y�H;��H;u�H;��H;�H;�H;��H;��H;��H;x�H;w�H;x�H;��H;�H;W�H;��H;H�H;��H;j�H;�H;��H;��H;��H;g�H;`�H;g�H;��H;��H;��H;�H;i�H;��H;D�H;��H;U�H;�H;��H;v�H;z�H;u�H;��H;��H;��H;�H;��H;��H;v�H;��H;Y�H;��H;H�H;��H;I;{I;�I;�I;�I;RI;�I;6I;      �I;�I;�I;I;�I;� I;��H;��H;��H;��H;��H;��H;�H;��H;d�H;�H;��H;��H;��H;��H;��H;��H;��H;�H;?�H;{�H;��H;w�H;��H;��H;.�H;��H;��H;g�H;Q�H;B�H;4�H;C�H;P�H;g�H;��H;��H;/�H;��H;��H;r�H;��H;{�H;A�H;�H;��H;��H;��H;��H;��H;��H;��H;�H;d�H;��H;�H;~�H;��H;��H;��H;��H;  I;� I;�I; I;�I;�I;      B I;P I; I;��H;0�H;{�H;��H;��H;��H;��H;��H;��H;W�H;H�H;*�H;�H;��H;��H;��H;��H; �H;�H;8�H;��H;��H;/�H;��H;5�H;��H;b�H;��H;��H;��H;P�H;.�H;�H;#�H; �H;*�H;P�H;��H;��H;��H;_�H;��H;/�H;��H;0�H;��H;��H;9�H;�H;��H;��H;��H;��H;��H;
�H;(�H;H�H;W�H;��H;��H;��H;��H;��H;��H;z�H;0�H;��H;  I;Q I;      ��H;��H;X�H;�H;��H;��H;J�H;x�H;��H;��H;��H;��H;��H;w�H;h�H;Z�H;R�H;C�H;Z�H;n�H;��H;��H; �H;H�H;��H;�H;��H;�H;��H;F�H;��H;��H;l�H;B�H;#�H;�H;�H;�H; �H;H�H;k�H;��H;��H;B�H;��H;��H;��H;�H;��H;F�H;�H;��H;��H;j�H;X�H;G�H;T�H;^�H;g�H;z�H;��H;��H;��H;��H;��H;v�H;Q�H;��H;��H;�H;T�H;��H;      �H;��H;��H;f�H;��H;>�H;��H;��H;�H;6�H;S�H;I�H;T�H;.�H;�H;�H;�H;�H;I�H;\�H;m�H;��H;��H;%�H;��H;��H;u�H;��H;��H;6�H;��H;��H;d�H;3�H;%�H;�H;�H;�H;"�H;4�H;e�H;��H;��H;1�H;��H;��H;u�H;�H;��H;#�H;��H;��H;g�H;W�H;I�H;!�H;�H;"�H;�H;1�H;T�H;E�H;T�H;9�H;�H;��H;��H;<�H;��H;j�H;��H;��H;      ��H;��H;R�H;�H;��H;��H;I�H;u�H;��H;��H;��H;��H;��H;z�H;h�H;Z�H;R�H;C�H;Z�H;n�H;��H;��H;��H;E�H;��H;�H;��H;�H;��H;F�H;��H;��H;n�H;C�H;#�H;�H;�H;�H; �H;F�H;k�H;��H;��H;?�H;��H;��H;��H;�H;��H;F�H;�H;��H;��H;j�H;X�H;I�H;R�H;`�H;g�H;w�H;�H;��H;��H;��H;��H;x�H;Q�H;��H;��H;�H;Y�H;��H;      7 I;P I;��H;��H;/�H;u�H;��H;��H;��H;��H;��H;��H;Y�H;H�H;+�H;�H;��H;��H;��H;��H; �H;�H;5�H;��H;��H;,�H;��H;5�H;��H;a�H;��H;��H;��H;P�H;-�H;�H;#�H;"�H;,�H;Q�H;��H;��H;��H;\�H;��H;,�H;��H;0�H;��H;��H;9�H;�H;��H;��H;��H;��H;��H;
�H;'�H;G�H;V�H;��H;��H;��H;��H;��H;��H;t�H;4�H;��H; I;V I;      �I;�I;�I; I;I;� I;��H;��H;��H;��H;��H;�H;�H;��H;f�H;�H;��H;��H;��H;��H;��H;��H;��H;�H;?�H;y�H;��H;w�H;��H;��H;-�H;��H;��H;e�H;Q�H;A�H;4�H;B�H;P�H;e�H;��H;��H;-�H;��H;��H;p�H;��H;|�H;A�H;�H;��H;��H;��H;��H;��H;��H;��H;�H;f�H;��H;�H;|�H;��H;��H;��H;��H; I;� I;�I;"I;�I;�I;      VI;;I;�I;RI;�I;�I;�I;�I;I;��H;F�H;��H;Z�H;��H;w�H;��H;�H;�H;��H;��H;��H;v�H;t�H;v�H;��H;�H;U�H;��H;H�H;��H;f�H;�H;��H;��H;��H;g�H;`�H;g�H;��H;��H;��H;�H;h�H;��H;?�H;��H;S�H;�H;��H;s�H;{�H;u�H;~�H;��H;��H;�H;��H;��H;v�H;��H;Y�H;��H;F�H;��H;I;I;�I;�I;�I;]I;�I;6I;      rI;pI;I;rI;�
I;�	I;]I;	I;tI;�I;%I;E I;q�H;��H;��H;;�H;��H;��H;d�H;��H;��H;��H;g�H;R�H;h�H;��H;��H;4�H;��H;<�H;��H;I�H;�H;��H;��H;��H;��H;��H;��H;��H;�H;J�H;��H;:�H;��H;/�H;��H;��H;e�H;K�H;k�H;��H;��H;��H;d�H;��H;��H;=�H;��H;��H;q�H;C I;$I;�I;vI;	I;^I;�	I;�
I;xI;I;lI;      �I;�I;KI;�I;{I;)I;�I;�I;
I;	I;�I;�I;�I;Z I;)�H;�H;'�H;`�H;��H;��H;7�H;��H;��H;k�H;R�H;C�H;��H;��H;(�H;��H;�H;��H;l�H;2�H;�H;��H;��H;��H;�H;4�H;m�H;��H;�H;��H;"�H;��H;��H;J�H;N�H;h�H;��H;��H;/�H;��H;��H;^�H;%�H;�H;'�H;W I;�I;�I;�I;	I;I; I;�I;'I;�I;�I;PI;�I;      �I;�I;�I;I;�I;JI;nI;`I;)I;�I;I;i
I;�I;I;�I; I;l�H;#�H;�H;�H;a�H;{�H;��H;��H;{�H;R�H;I�H;w�H;��H;�H;��H;9�H;��H;��H;_�H;?�H;/�H;B�H;\�H;��H;��H;:�H;��H;�H;��H;s�H;F�H;Y�H;v�H;��H;��H;y�H;\�H;�H;�H;!�H;l�H; I;�I;I;�I;d
I; I;�I;%I;]I;nI;<I;�I;'I; I;�I;      �!I;�!I;2"I;@"I;�!I;!I;�I;GI;�I;�I;�I;lI;I;�
I;�I;�I;�I;��H;0�H;��H;��H;��H;��H; �H;��H;q�H;D�H;F�H;��H;��H;!�H;��H;@�H;��H;��H;��H;��H;��H;��H;��H;A�H;��H;"�H;��H;��H;@�H;C�H;x�H;��H;�H;��H;��H;��H;��H;1�H;��H;�I;�I;�I;�
I;I;iI;�I;�I;�I;HI;�I;!I;�!I;C"I;2"I;�!I;      ��H;B�H;|I;�	I;�I;�I;UI;� I;�!I;U I;lI;�I;�I;�I;I;<
I;�I;SI;3 I;'�H;p�H;0�H;�H;�H;/�H;��H;{�H;]�H;D�H;r�H;��H;0�H;��H;q�H;0�H;�H;��H;�H;0�H;r�H;��H;0�H;��H;r�H;@�H;Y�H;y�H;��H;+�H;�H;�H;0�H;k�H;&�H;3 I;OI;�I;9
I;�I;�I;�I;�I;kI;R I;�!I;� I;VI;�I;�I;�	I;�I;B�H;      �NH;�TH;�dH;�}H;ݛH;X�H;��H;��H;�I;I;  I;!I;oI;0I;�I;I;�I;�I;�I;hI;�H;�H;n�H;H�H;�H;@�H;��H;�H;M�H;I�H;��H;��H;S�H;��H;��H;��H;w�H;��H;��H;��H;U�H;��H;��H;J�H;H�H;|�H;��H;G�H;�H;D�H;u�H;�H;�H;iI;�I;�I;�I;I;�I;,I;lI;!I;�I;I;�I;��H;��H;T�H;�H;�}H;�dH;�TH;      OIF;sYF;��F;��F;z'G;ňG;��G;CH;)�H;F�H;[�H;�I;�I;� I;�I;�I;�I;I;J
I;I;?I;��H;m�H;��H;_�H;5�H;A�H;��H;}�H;Y�H;F�H;��H;�H;{�H;6�H;�H;�H;�H;3�H;}�H;�H;��H;I�H;[�H;v�H;��H;A�H;>�H;\�H;��H;q�H;��H;<I;I;K
I;�I;�I;�I;�I;� I;�I;�I;[�H;E�H;�H;CH;��G;��G;�'G;��F;��F;dYF;      �DA;�kA;J�A;d�B;�jC;PaD;}\E;�IF;�G;��G;^NH;.�H;��H;�I;uI;X I;�I;9I;�I;�I;�I;�I;�H;��H;��H;X�H;�H;/�H;��H;v�H;M�H;c�H;��H;?�H;��H;��H;��H;��H;��H;A�H;��H;c�H;R�H;x�H;��H;,�H;�H;b�H;��H;��H;�H;�I;�I;�I;�I;5I;�I;X I;uI;�I;��H;)�H;[NH;��G;�G;�IF;{\E;CaD;�jC;j�B;J�A;�kA;      �J6;�6;��7;�9;>;;.=;Ej?;T�A;�C;M2E;��F;O�G;q<H;~�H;��H;�I;G I;I;#I;3I;�I;�I;3I;-�H;��H;��H;=�H;�H;�H;��H;h�H;R�H;t�H;�H;��H;P�H;,�H;Q�H;��H;	�H;x�H;T�H;m�H;��H;�H;�H;@�H;��H;��H;0�H;7I;�I;�I;6I;#I;I;G I;�I;��H;|�H;o<H;J�G;��F;K2E;�C;L�A;Fj?;.=;V;;�9;��7;�6;      p ;�!;�#;�&;�*;�o.;_3;��7;b�;;j?;8kB;	�D;kxF;��G;�cH;�H;�
I;�I;OI;_I;I;I;�I;7I;�H;h�H;l�H;�H;��H;��H;��H;e�H;r�H;��H;8�H;�H;��H; �H;4�H;��H;t�H;d�H;��H;��H;��H;	�H;o�H;q�H;�H;:I;�I;I;I;bI;RI;�I;�
I;�H;�cH;��G;kxF;�D;8kB;j?;a�;;��7;_3;�o.;�*;�&;�#;�!;      ct�:� �:1l�:>�;� 
;܄;(z;P$;K�,;��3;	�9;�>;�B;2E;�F;RH;խH;��H;I;�I;"I;ZI;I;�I;�I;��H;��H;0�H;��H;v�H;��H;��H;o�H;��H;�H;��H;��H;��H;�H;��H;r�H;��H;��H;{�H;��H;.�H;�H;��H;�I;�I;I;]I;$I;�I;	I;��H;ԭH;OH; �F;2E;�B; �>;�9;��3;K�,;P$;z;;� 
;4�;1l�:� �:      8�>:��G:��b:t��:%��:�4�:�*�:~i;@�;�a;*;@r3;��:;�!@;��C;�IF;��G;��H;�H;SI;�I;I;I;�I;�I;3I;��H;j�H;��H;W�H;,�H;��H;z�H;��H;��H;��H;d�H;��H;��H;��H;|�H;��H;-�H;[�H;��H;j�H;��H;:I;�I;�I;I;I;�I;VI;
�H;��H;��G;�IF;��C;�!@;��:;<r3;*;�a;;�;~i;�*�:�4�:G��:z��:��b:`�G:      ���̅��uk��� �`���-69��!:�Ȋ:z4�:��:��;�;G�,;��6;��=;��B;m�E;V�G;�|H;t�H;WI;�I;^I;6I;�I;�I;bI;'�H;��H;�H;��H;��H;��H;��H;��H;j�H;V�H;m�H;��H;��H;��H;��H;��H;�H;��H;'�H;fI;I;�I;=I;cI;�I;XI;u�H;�|H;T�G;k�E;��B;��=;��6;D�,;�;��;��:p4�:�Ȋ:��!: -69@��ؙ �uk�Ѕ��      $/��"����x���X���/�� ����o치9�9��k:��:-o�:�B;�&;C3;q<;�A;�pE;BtG;�|H;�H;I;OI;"I;�I;G
I;�I;1 I;,�H;�H;��H;^�H;��H;��H;��H;W�H;E�H;W�H;��H;��H;��H;^�H;��H;�H;*�H;1 I;�I;H
I;�I;(I;QI;I;
�H;�|H;@tG;�pE;�A;m<;@3;�&;�B;)o�:��:��k:�9�9o����� ���/���X��x� ���      ������q
����2�׻�+��Ʈ���;��lۺ,� �(P�9�Ȋ:��:�; !;��0;;;��A;�pE;P�G;��H;��H;�I;I;3I;�I;�I;SI;��H;"�H;[�H;��H;��H;��H;��H;F�H;�H;G�H;��H;��H;��H;��H;]�H;#�H;��H;UI;�I;�I;.I;I;�I;��H;��H;S�G;�pE;��A;;;��0;!;�;��:�Ȋ:@P�9<� ��lۺ�;�Ȯ���+��4�׻����q
���      ����p8����>�k���O��3/�0B�	�׻Ƶ��d�@�HP����(�>:�4�:��;Vb;��/;;;�A;h�E;��G;ЭH;�
I;E I;�I;�I;�I;�I;�I;e�H;�H;��H;z�H;��H;��H;O�H;�H;O�H;��H;��H;x�H;��H;�H;h�H;�I;�I;�I;�I;�I;E I;�
I;ѭH;��G;k�E;�A;;;�/;Vb;��;�4�:0�>:(��NP��f�@�ŵ���׻0B��3/���O�?�k���o8��      9���|�0�ݼ��˼d���,���}� �G����B�һ����d���/�p:*׳:�;Ob;��0;m<;��B;�IF;KH;�H;�I;Q I;�I;I;6
I;�I; I;�H;6�H;��H;�H;�H;\�H;�H;\�H;�H;�H;��H;4�H;�H; I;�I;:
I;I;�I;L I;�I;�H;LH;�IF;��B;k<;��0;Rb;��;(׳:t:�/�h������B�һ����G��}��,��d����˼2�ݼ�|�      D�B�LR?��5���&��3��J��ӮҼ!F����>=�!?�.����/��nk���9&׳:��;!;<3;��=;��C;��F;�cH;��H;oI;�I;�I;I;�I;�I;%�H;��H;s�H;c�H;#�H;d�H;�H;e�H;!�H;b�H;s�H;��H;$�H;�I;�I;I;�I;�I;kI;��H;�cH; �F;��C;��=;93;!;��; ׳:��9�nk���/�.��!?�?=� ��!F��ӮҼ�J���3���&��5�LR?�      (��$W��蒐�"�����j�Q`I���&����Dϼ�,���T[�k�kI��a;��nk��:�4�:�;�&;��6;�!@;2E;��G;��H;�I;� I;.I;�I;�
I;I;V I;��H;��H;��H;A�H;t�H;'�H;w�H;?�H;��H;��H;��H;S I;I;�
I;�I;.I;� I;�I;��H;��G;2E;�!@;��6;�&;�;�4�:t:�nk�c;�lI��k��T[��,��Dϼ�����&�Q`I���j�"���璐�$W��      �J�����D��ͽ���'�������L�%��$��;���k����jI����/��/��>:��:�B;C�,;��:;�B;mxF;v<H;��H;�I;mI;�I; I;�I;�I;n�H;Y�H;�H;P�H;�H;N�H;�H;O�H;�H;V�H;m�H;�I;�I;!I;�I;oI;�I;��H;t<H;pxF;�B;��:;F�,;�B;��:$�>:�/���/�kI������k�;��$��$����L����'������ͽ�D����      Q�:��*7���,�+���	�q�齂��� W����j�>�/��J���I���k�l�.��e��H���Ȋ:)o�:�;Fr3;��>;�D;O�G;'�H;�I;!I;�I;iI;b
I;�I;? I;��H;|�H;��H;��H;B�H;��H;��H;{�H;��H;> I;�I;d
I;mI;�I;!I;�I;!�H;M�G;�D; �>;=r3;�;#o�:�Ȋ:(��h��.��l��k��I���J��>�/���j� W������q�齂�	�+���,��*7�      ^���p����2�l���M���,�Xl�Q9ݽ�A���{���5��J��;���T[�"?�����\P���O�9��:��;*;�9;7kB;��F;YNH;W�H;�I;iI;�I; I;�I;"I;D�H;��H;��H;��H;J�H;��H;��H;��H;D�H; I;�I;I;�I;kI;�I;V�H;TNH;��F;;kB;�9;*;��;��: P�9ZP������"?��T[�	;���J����5��{��A��Q9ݽXl���,���M�2�l����p��      4m־O�Ѿ�>ľ����җ����{��I�+����V���{�>�/�$���,��>=�B�һm�@�T� ���k:��:�a;��3;
j?;Q2E;��G;A�H;I;M I;�I;�I;	I;�I;��H;��H;��H;��H;9�H;��H;��H;��H;��H;�I; 	I;�I;�I;Q I;I;B�H;��G;P2E;j?;��3;�a;��:��k:H� �j�@�C�һ>=��,��$��>�/��{��V�����+��I���{�җ�������>ľO�Ѿ      C\����r5��z ��E۾ֳ�^��y�Z�K?#����A����j�%��Eϼ�����ʵ���lۺX9�9h4�:B�;C�,;U�;;�C;�G;�H;I;�!I;�I;%I;	I;sI;$I;��H;��H;��H;�H;��H;��H;��H;#I;sI;I;$I;�I;�!I;�I;"�H;~G;�C;Y�;;G�,;:�;l4�:P9�9�lۺʵ�������Dϼ%����j��A�����K?#�y�Z�^��ֳ��E۾�z �r5����      E�b��>]���M�Î6�����$���>ľ#q��y�Z�+�Q9ݽ W����L����"F���G��׻;�Ho칀Ȋ:�i;�O$;��7;T�A;�IF;CH;��H;� I;BI;VI;�I;
I;�I;��H;��H;t�H;��H;r�H;��H;��H;I;I;�I;ZI;EI;� I;��H;CH;�IF;S�A;��7;P$;zi;�Ȋ:Ho�;��׻�G�"F�������L� W��Q9ݽ+�y�Z�#q���>ľ�$�����Î6���M��>]�      p��񲗿���7�y�{�R���)�nv��>ľ^���I�Xl����������&�ԮҼ�}�1B�ͮ��"���|�!:�*�: z;X3;Fj?;r\E;��G;��H;GI;I;mI;�I;WI;�I;��H;��H;C�H;��H;C�H;��H;��H;�I;XI;�I;pI;�I;LI;��H;��G;r\E;Ij?;_3; z;�*�:��!:"���̮��0B��}�ԮҼ��&��������Xl��I�^���>ľnv���)�{�R�7�y����񲗿      �˿�<ƿqL��@1����>]���)��$��ֳ���{���,�q��'��Q`I��J���,���3/�,��� � -69�4�:Є;�o.;.=;=aD;��G;O�H;�I;!I;BI;,I;�	I;�I;� I;��H;��H;E�H;��H;��H;� I;�I;�	I;*I;BI;!I;�I;T�H;��G;=aD;.=;�o.;Є;�4�: -69� � ,���3/��,���J��Q`I�'��q�齥�,���{�ֳ��$����)��>]��@1��qL���<ƿ      ����<���T[忶˿�T���{�R�����E۾ӗ����M���	������j��3�d����O�<�׻��/�@��?��:� 
;�*;K;;�jC;}'G;ћH;�I;�!I;�I;wI;�
I;�I;�I;�H;��H;��H;��H;"�H;�I;�I;�
I;vI;�I;�!I;�I;ۛH;�'G;�jC;O;;�*;� 
;7��:0����/�:�׻��O�d���3���j������	���M�ӗ���E۾���{�R���T���˿T[�<���      O�6��t����˿@1��7�y�Î6��z �����2�l�+��ͽ#�����&���˼?�k�#�����X�� �z��:6�;�&;z9;j�B;��F;�}H;�	I;."I;I;�I;yI;TI;%I;��H;�H;c�H;�H;��H;"I;TI;|I;�I;I;3"I;�	I;�}H;��F;j�B;}9;�&;8�;p��:� ���X� ���>�k���˼��&�#����ͽ+�2�l������z �Î6�7�y�@1���˿���t�6��      ��*��g&��#�t�T[�qL�������M�r5��>ľ����,��D�蒐��5�1�ݼ���q
��x�$uk���b:%l�:�#;×7;T�A;��F;�dH;�I;!"I;�I;EI;I;�I;�I;��H;Y�H;��H;T�H;��H;�I;�I;I;BI;�I;%"I;�I;�dH;��F;Q�A;7;�#;%l�:��b:uk��x��q
���1�ݼ�5�蒐��DὫ�,����>ľr5���M����qL��T[�t��#��g&�      ��8��4��g&�6��<����<ƿ񲗿�>]����O�Ѿ�p���*7����%W��LR?��|�q8�������҅����G:s �:�!;�6;�kA;eYF;�TH;C�H;�!I;�I;�I;eI;(I;�I;> I;��H;��H;��H;> I;�I;)I;hI;�I;�I;�!I;F�H;�TH;sYF;�kA;�6;�!;q �:��G:ʅ�������q8�� }�LR?�%W�����*7��p��O�Ѿ����>]�񲗿�<ƿ<���6���g&��4�      �Aq���i���U�F:�@�����<���u���{A�d5�� ��~^Z�����A���]�����d��K",��5����Ѻ(��9���:�;[Y4;H�@;LVF;~�H;�GI;�bI;OI;:I;�)I;I;~I;�I;�I;�I;}I;�I;~I;I;�)I;:I;OI;�bI;�GI;��H;XVF;E�@;ZY4;�;���: ��9��Ѻ�5��K",��d������]��A�����~^Z�� ��d5�{A�u���<�������@�F:���U���i�      ��i���b�Z�O�.5�1i�������������q<�����e��`
V�GE	�!���IY�j9�D�����(��R���Ⱥ`�:P��:�;?�4;>�@;hF;��H;
II;vbI;�NI;�9I;�)I;�I;[I;�I;`I;]I;ZI;�I;ZI;�I;�)I;�9I;�NI;ybI;II;��H;(hF;<�@;<�4;ݔ;J��:T�: �Ⱥ�R����(�D���j9��IY�!��GE	�`
V��e������q<������������1i�.5�Z�O���b�      ��U�Z�O�H-?�.�'���M�ῴ欿a�{�ea/���뾝���I����c���ZN�\5������=H�d ��n�����":��:z�;��5;�`A;��F;K�H;MI;�aI;�MI;�8I;�(I;BI;�I;:I;I;I;�I;9I;�I;BI;�(I;�8I;�MI;�aI;MI;L�H;��F;�`A;��5;v�;��:|�":h���f ��=H�����\5���ZN�c������I�������ea/�a�{��欿M����.�'�H-?�Z�O�      F:�.5�.�'��������jȿ���l$_���W�Ҿە���6�����*���`=�<�漮)��IG�(6�����$�Q:��:�/";	�7;_&B;��F;��H;�RI;�`I;xKI;7I;�'I;>I;I;�I;qI;p
I;kI;�I;I;<I;�'I;7I;zKI;�`I;�RI;��H;��F;[&B;�7;�/";��:�Q:���(6��HG��)��<���`=��*������6�ܕ��W�Ҿ��l$_����jȿ�������.�'�.5�      @�1i�������I�ѿk��� ���q<��:��a����q����Wн罅���'�Tb̼�zl��.��N�X�`����:��;Ύ&;ū9;$C;;MG;��H;8YI;�^I;�HI;�4I;�%I;�I;I;�I;�
I;�	I;�
I;�I;I;�I;�%I;�4I;�HI;�^I;8YI;��H;@MG;!C;��9;ˎ&;��;��:T��P�X��.���zl�Ub̼��'�罅��Wн����q��a���:��q<� ��k���I�ѿ������1i�      �������L��jȿk���������O���{]׾z����I�����A��>�d�n�}֮�RH��jλQ�$��(�n��:EN;��+;�<;�3D;��G;�I;�^I;l[I;�DI;"2I;�#I;CI;�I;]I;�	I;�I;�	I;]I;�I;CI;�#I; 2I;�DI;j[I;�^I;�I;��G;�3D;�<;��+;BN;d��:�(�Q�$��jλRH�}֮�n�>�d��A������I�z���{]׾����O�����k���jȿL�Ῡ��      <��������欿��� ����O��x����� ���l���"��ܽ���`=����u���k"�/R��Dۺ���9�?�:ZL;~�0;��>;�ME;H#H;�%I;�aI;�VI;�@I;�.I;=!I;>I;I;
I;MI;�I;JI;
I;I;@I;=!I;�.I;�@I;�VI;�aI;�%I;M#H;�ME;��>;}�0;XL;|?�:Г�9Dۺ/R���k"�u������`=����ܽ��"��l�� ����뾁x���O� ������欿����      u�������a�{�l$_��q<�������}��w��	�6�����!���h����ⷾ�� d��.���^e�I[���Z:^��:�, ;��5;�A;�VF;��H;�@I;obI;�QI;�;I;=+I;mI;I;7I;}	I;�I;,I;�I;	I;7I;I;kI;;+I;�;I;�QI;rbI;�@I;��H;�VF;�A;��5;�, ;T��:��Z:I[��^e�~.��� d�ⷾ�����h�!������	�6�w���}��������q<�l$_�a�{�����      {A��q<�ea/����:�{]׾� ��w��>�DE	�����ڽ����3�^�꼙���",��W��a�� Q�t��:�M
;�f);��:;$@C;�?G;O�H;ETI;�_I;$KI;�6I;N'I;eI;�I;;I;�I;oI;�I;lI;�I;;I;�I;gI;O'I;�6I;)KI;�_I;DTI;M�H;�?G;!@C;��:;�f);�M
;���: Q�c���W��",�����^�꼘�3�ڽ������DE	�>�w��� ��{]׾�:���ea/��q<�      d5�������W�Ҿ�a��z����l�	�6�DE	���Ƚk���aG����d֮��W����p�k�2���c,:���:��;��1;<�>;=E;�G;I;#_I;AZI;3DI;�1I;0#I;EI; I;
I;I;�I;I;�I;I;
I;�I;AI;0#I;�1I;7DI;DZI;#_I;I;"�G;9E;>�>;��1;��;���:�c,:0��l�k�����W�d֮�����aG�k����ȽDE	�	�6��l�z����a��W�Ҿ������      � ���e�����ە����q��I���"���������k���ZN�[�!¼P�y��$��Q���� � pX���:0;$�&;�w8;j B;��F;АH;T@I;�aI;jRI;=I;,I;�I;�I;\I;�I;4I;I;eI;I;5I;�I;[I;�I;�I;,I;=I;mRI;�aI;R@I;ԐH;��F;l B;�w8;#�&;0;��: dX��� ��Q���$�N�y� ¼Z��ZN�k������������"��I���q�ە������e��      ~^Z�`
V��I��6�������ܽ!��ڽ���aG�Z�
�ȼ�)��}�(�h��LG5������Z:�:S;
'1;��=;��D;,�G;��H;�XI;^I;~II;�5I;�&I;�I;�I;�
I;�I;MI;a I;��H;a I;MI;�I;�
I;�I;�I;�&I;�5I;II;^I;�XI;��H;+�G;��D;��=;'1;S;�:��Z:���JG5�f��|�(��)��
�ȼZ��aG�ڽ��!���ܽ������6��I�`
V�      ���GE	��������Wн�A�����h���3���� ¼�)��1x/��һu�X�x#����9N��:�>;,f);c`9;Z&B;��F;d}H;�6I;NaI;�UI;`@I;�.I;� I;GI;(I;�I;NI;Q I;��H;��H;��H;P I;NI;�I;(I;KI;!I;�.I;a@I;�UI;KaI;�6I;b}H;��F;^&B;b`9;7f);�>;H��:��9r#��r�X��һ0x/��)�� ¼�����3��h��󑽠A���Wн��콺��FE	�      �A��!��c���*��潅�>�d��`=����]��c֮�N�y�|�(��һ�]e����f9���:6�;A1";�4;�m?;�E;��G;e�H;�WI;}^I;KI;q7I;�'I;�I;$I;�
I;$I;I;m�H;��H;;�H;��H;k�H;I;!I;�
I;(I;�I;�'I;t7I;KI;y^I;�WI;d�H;��G;�E;�m?;�4;G1";4�;���:p�f9ꄮ��]e��һ|�(�M�y�c֮�]�꼗���`=�>�d�潅��*��c��!��      �]��IY��ZN��`=���'�m����᷾������W��$�h��u�X�����09x��:Y��:o�;��0;��<;N�C;G;��H;�?I;#aI;�TI;>@I;/I;U!I;�I;I;yI;�I;��H;}�H;�H;��H;�H;|�H;��H;�I;vI;I;�I;Z!I;/I;;@I;�TI;&aI;�?I;��H;G;P�C;��<;��0;l�;e��:t��: 9ꄮ�r�X�f���$��W�����᷾����m���'��`=��ZN��IY�      ���i9�Z5��:��Tb̼}֮�t��� d�",�����Q��KG5�z#����f9|��:��:�;��-;��:;�KB;8VF;KH;�I;�\I;\I;�HI;6I;'I;I;�I;
I;BI;��H;��H;��H;Z�H;��H;X�H;��H;��H;��H;AI;
I;�I;I;'I;6I;�HI;\I;�\I;�I;KH;:VF;�KB;��:;��-;�;��:|��:p�f9|#��HG5��Q�����",�� d�u��|֮�Ub̼:��Z5��h9�      �d��B��������)���zl�RH��k"�{.���W��e�k��� ������9���:e��:�;�-;̫9;BaA;��E;%�G;u�H;�RI;`I;�OI;�<I;�,I;�I;.I;I;zI;TI;��H;��H;��H;��H;a�H;��H;��H;��H;��H;TI;~I;I;.I;�I;�,I;�<I;�OI;`I;�RI;t�H;%�G;��E;DaA;ƫ9;�-;�;g��:���:��9����� �e�k��W��z.���k"�RH��zl��)������A���      D",���(�<H�EG��.���jλ(R���^e�_��"�� XX���Z:F��:2�;m�;��-;ū9;wA;�cE;�G;��H;OGI;�`I;�UI;8BI;�1I;�#I;�I;�I;�I;�I;��H;H�H;��H;�H;�H;��H;�H;	�H;��H;E�H;��H;�I;�I;�I;�I;�#I;�1I;;BI;�UI;�`I;NGI;��H; �G;�cE;tA;ȫ9;��-;m�;2�;B��:��Z: DX�"��Y���^e�*R���jλ�.��FG�:H���(�      �5���R��d ��$6��R�X�B�$�.ۺ�H[� 
Q��c,:��:�:�>;G1";��0;��:;BaA;�cE;��G;r�H;�=I;+`I;qYI;�FI;�5I;�'I;�I;�I;�
I;�I;��H;�H;�H;��H;�H;��H;<�H;��H;}�H;��H;�H;�H;��H;�I;�
I;�I;�I;�'I;�5I;�FI;gYI;+`I;�=I;u�H;��G;�cE;GaA;��:;��0;E1";�>;�:��:�c,: 
Q��H[�6ۺH�$�P�X�)6��d ���R��      ��Ѻ�ȺZ������d���(���9��Z:���:���:%0;S;3f);�4;��<;�KB;��E;%�G;v�H;]:I;O_I;[I;#JI;9I;�*I;�I;�I; I;]I;I;��H;��H;�H;/�H;��H;7�H;��H;2�H;��H;.�H;�H;��H;��H;I;YI; I;�I;�I;�*I;9I;JI;~[I;Q_I;\:I;v�H;�G;��E;�KB;��<;�4;2f);S;%0;���:���:��Z:�9@(�H�����p���"�Ⱥ      X��9�:�":�Q:��:r��:�?�:Z��:�M
;��;#�&;'1;b`9;�m?;P�C;<VF;&�G;��H;�=I;N_I;\I;�KI;;I;�,I;� I;�I;�I;�I;HI;��H;5�H;x�H;5�H;��H;��H;��H;��H;��H;��H;��H;2�H;r�H;7�H;��H;DI;�I;�I;�I;� I;�,I;;I;�KI;\I;L_I;�=I;��H;&�G;<VF;P�C;�m?;c`9;'1;(�&;��;�M
;X��:�?�:f��:��:�Q:H�":�:      ���:p��:��:��:��;FN;ZL;�, ;�f);��1;�w8;��=;_&B;�E;#G;KH;x�H;SGI;1`I;�[I;�KI;�;I;�-I;0"I;-I;I;	I;aI;��H;��H;��H;j�H;y�H;�H;F�H;��H;e�H;��H;C�H;�H;x�H;f�H;��H;��H;��H;cI;	I;I;0I;,"I;�-I;�;I;�KI;[I;.`I;OGI;x�H;KH;#G;�E;^&B;��=;�w8;��1;�f);�, ;_L;BN;��;��:��:T��:      7�;�;t�;�/";Î&;��+;��0;��5;��:;D�>;v B;��D;��F;��G;��H;�I;SI;�`I;qYI;!JI;;I;�-I;�"I;I;�I;�	I;,I;G�H;o�H;W�H;��H;��H;��H;��H;��H;��H;a�H;��H;��H;��H;��H;��H;��H;V�H;j�H;K�H;%I;�	I;�I;�I;�"I;�-I;;I;JI;nYI;�`I;�RI;�I;��H;��G;��F;��D;y B;?�>;��:;��5;��0;��+;Վ&;�/";q�;ɔ;      XY4;H�4;��5;�7;��9;�<;��>;�A;@C;=E;��F;.�G;b}H;e�H;�?I;�\I;`I;�UI;�FI;�8I;�,I;+"I; I;#I;[
I;�I;��H;��H;��H;��H;��H;��H;��H;��H;��H;��H;f�H;��H;��H;��H;��H;��H;��H;��H;��H;��H;��H;�I;\
I; I;�I;+"I;�,I;�8I;�FI;�UI;`I;�\I;�?I;a�H;b}H;,�G;��F;<E; @C;�A;��>;�<;ū9;�7;��5;?�4;      h�@;>�@;�`A;]&B;C;4D;�ME;�VF;�?G;%�G;ڐH;��H;�6I;�WI;*aI;&\I;�OI;CBI;�5I;�*I;� I;3I;�I;d
I;�I; I;0�H;��H;$�H;��H;��H;��H;K�H;z�H;��H;��H;e�H;��H;��H;z�H;G�H;��H;��H;��H;�H;��H;*�H; I;�I;`
I;�I;4I;� I;�*I;�5I;?BI;�OI;*\I;'aI;�WI;�6I;��H;ڐH;%�G;�?G;�VF;�ME;�3D;'C;[&B;�`A;?�@;      NVF;.hF;��F;��F;1MG;��G;N#H;��H;R�H;I;W@I;�XI;PaI;�^I;�TI;�HI;�<I;�1I;�'I;�I;�I;I;�	I;�I; I;?�H;�H;X�H;��H;��H;w�H;H�H;=�H;x�H;�H;��H;|�H;��H;�H;x�H;<�H;D�H;w�H;��H;��H;V�H;�H;A�H; I;�I;�	I;I;�I;�I;�'I;�1I;�<I;�HI;�TI;~^I;PaI;�XI;]@I;I;R�H;��H;P#H;��G;GMG;��F;��F;(hF;      ��H;��H;E�H;��H;��H;�I;�%I;�@I;HTI;$_I;�aI;^I;�UI;	KI;;@I;6I;�,I;�#I;�I;�I;�I;	I;-I;��H;-�H;�H;J�H;�H;.�H;n�H;&�H;�H;8�H;��H;7�H;��H;��H;��H;4�H;��H;6�H;�H;&�H;l�H;'�H;�H;@�H;�H;.�H;��H;,I;	I;�I;�I;�I;�#I;�,I;6I;:@I;KI;�UI;^I;�aI;#_I;GTI;�@I;�%I;�I;��H;��H;E�H;��H;      �GI;II;MI;�RI;.YI;�^I;�aI;pbI;�_I;GZI;oRI;�II;]@I;t7I;/I;'I;�I;�I;�I;�I;�I;aI;G�H;��H;��H;T�H;�H;�H;|�H;&�H;��H;�H;e�H;��H;t�H;>�H;3�H;=�H;r�H;��H;d�H;�H;��H;#�H;w�H;�H;�H;V�H;��H;��H;E�H;aI;�I;�I;�I;�I;�I;!'I;/I;r7I;[@I;�II;qRI;GZI;�_I;nbI;�aI;w^I;:YI;�RI;MI;II;      �bI;ubI;�aI;�`I;�^I;k[I;WI;�QI;KI;6DI;=I;�5I;�.I;�'I;Z!I;I;4I;�I;�
I;`I;NI;��H;n�H;��H;�H;��H;%�H;z�H;!�H;��H;��H;8�H;��H;)�H;��H;��H;��H;��H;��H;*�H;��H;5�H;��H;��H;�H;y�H; �H;��H;�H;��H;n�H;��H;JI;\I;�
I;�I;2I;I;W!I;�'I;�.I;�5I;=I;9DI;&KI;�QI;WI;d[I;�^I;�`I;�aI;sbI;      OI;�NI;�MI;sKI;�HI;�DI;�@I;�;I;�6I;�1I;,I;�&I; !I;�I;�I;�I;I;�I;�I;I;��H;��H;X�H;��H;��H;��H;n�H;*�H;�H;��H;#�H;|�H;��H;��H;D�H;�H;�H;�H;@�H;��H;��H;{�H;#�H;��H;��H;%�H;g�H;��H;��H;��H;X�H;��H;��H;I;�I;�I;I;�I;�I;�I; !I;�&I;,I;�1I;�6I;�;I;�@I;�DI;�HI;yKI;�MI;�NI;       :I;�9I;�8I;&7I;�4I;!2I;�.I;H+I;P'I;6#I;�I;�I;NI;,I;I; 
I;�I;�I;��H;��H;@�H;��H;��H;��H;��H;v�H;)�H;�H;��H;*�H;��H;��H;\�H;	�H;��H;��H;��H;��H;��H;�H;\�H;��H;��H;&�H;��H;�H;#�H;w�H;��H;��H;��H;��H;9�H;��H;��H;�I;�I;!
I;I;+I;OI;�I;�I;7#I;S'I;G+I;�.I;2I;�4I;(7I;�8I;�9I;      �)I;�)I;�(I;�'I;�%I;�#I;=!I;mI;jI;EI;�I;�I;+I;�
I;{I;EI;ZI;��H;�H;��H;��H;l�H;��H;��H;��H;B�H;�H;�H;;�H;�H;��H;t�H;��H;��H;t�H;L�H;6�H;N�H;p�H;��H;��H;t�H;��H;|�H;5�H;	�H;	�H;B�H;��H;��H;��H;l�H;x�H;��H;�H;��H;[I;HI;{I;�
I;(I;�I;�I;EI;hI;jI;F!I;�#I;�%I;�'I;�(I;�)I;      %I;�I;MI;AI;�I;9I;;I;I;�I;�I;\I;�
I;�I;&I;�I;��H;��H;K�H;#�H;�H;B�H;}�H;��H;��H;N�H;<�H;9�H;l�H;��H;��H;V�H;��H;��H;S�H;�H; �H;�H;�H;	�H;U�H;��H;��H;X�H;��H;��H;g�H;5�H;9�H;N�H;��H;��H;{�H;9�H;�H;#�H;K�H;��H; I;�I;&I;�I;�
I;_I;�I;�I;	I;=I;4I;�I;;I;WI;�I;      vI;\I;�I;I;I;�I;I;:I;;I;	
I;�I;�I;SI;!I;��H;��H;��H;��H;��H;5�H;��H;�H;��H;��H;u�H;t�H;��H;��H;-�H;��H;�H;��H;U�H;�H;��H;��H;��H;��H;��H;�H;W�H;��H;�H;��H;(�H;��H;��H;t�H;x�H;��H;��H;�H;��H;.�H;��H;��H;��H;��H;��H;!I;RI;�I;�I;
I;>I;7I;
I;�I;	I;I;�I;eI;      �I;�I;@I;�I;�I;WI;I;�	I;�I;I;>I;XI;Z I;u�H;��H;��H;��H;�H;��H;��H;��H;D�H;��H;��H;��H;��H;1�H;u�H;��H;F�H;��H;s�H;�H;��H;��H;��H;��H;��H;��H;��H;�H;w�H;��H;@�H;��H;q�H;1�H;��H;��H;��H;��H;B�H;��H;��H;��H;�H;��H;��H;��H;u�H;[ I;VI;?I;I;�I;�	I;I;WI;�I;�I;@I;�I;      ~I;dI;I;nI;�
I;	I;SI;�I;lI;�I;"I;e I;��H;��H;�H;W�H;��H;�H;��H;6�H;��H;��H;��H;x�H;��H;��H;��H;A�H;��H;$�H;��H;M�H;�H;��H;��H;z�H;y�H;}�H;��H;��H;�H;P�H;��H;�H;��H;=�H;��H;��H;��H;z�H;��H;��H;��H;3�H;��H;�H;��H;[�H;�H;��H;��H;d I;%I;�I;oI;�I;ZI;�	I;�
I;oI; I;rI;      �I;WI;I;q
I;�	I;�I;�I;2I;�I;I;mI;��H;��H;B�H;��H;��H;j�H;��H;A�H;��H;��H;h�H;`�H;]�H;b�H;u�H;��H;:�H;��H;!�H;��H;8�H;�H;��H;��H;u�H;~�H;w�H;��H;��H;�H;;�H;��H;�H;��H;3�H;��H;w�H;f�H;]�H;d�H;h�H;��H;��H;A�H;��H;j�H;��H;��H;E�H;��H;��H;mI;I;�I;2I;�I;�I;�	I;u
I;I;dI;      ~I;eI; I;nI;�
I;�	I;QI;�I;lI;�I;!I;g I;��H;��H;�H;W�H;��H;�H;��H;6�H;��H;��H;��H;w�H;��H;��H;��H;A�H;��H;!�H;��H;M�H;�H;��H;��H;z�H;y�H;}�H;��H;��H;�H;P�H;��H;�H;��H;:�H;��H;��H;��H;x�H;��H;��H;��H;3�H;��H;�H;��H;\�H;�H;��H;��H;b I;"I;�I;mI;�I;XI;�	I;�
I;uI;I;lI;      �I;�I;;I;�I;�I;SI;I;�	I;�I;I;?I;XI;Z I;u�H;��H;��H;��H;�H;��H;��H;��H;D�H;��H;��H;��H;��H;0�H;t�H;��H;D�H;��H;s�H;�H;��H;��H;��H;��H;��H;��H;��H;�H;v�H;��H;=�H;��H;n�H;1�H;�H;��H;��H;��H;C�H;��H;��H;�H;�H;��H;��H;��H;t�H;Z I;VI;>I;I;�I;�	I;I;SI;�I;�I;AI;�I;      vI;[I;�I;I;I;�I;I;=I;>I;
I;�I;�I;RI;!I;��H;��H;��H;��H;��H;4�H;��H;�H;��H;��H;w�H;t�H;��H;��H;-�H;��H;�H;��H;U�H;�H;��H;��H;��H;��H;��H;�H;W�H;��H;�H;��H;&�H;��H;��H;w�H;w�H;��H;��H;�H;��H;/�H;��H;��H;��H;��H;��H; I;PI;�I;�I;
I;<I;<I;I;�I;	I;I;�I;\I;      "I;�I;PI;:I;�I;<I;:I;I;�I;�I;^I;�
I;�I;&I;�I;��H;��H;I�H;!�H;�H;?�H;|�H;��H;��H;N�H;6�H;5�H;k�H;��H;��H;U�H;��H;��H;S�H;�H;�H;�H; �H;�H;T�H;��H;��H;V�H;��H;��H;e�H;4�H;:�H;K�H;��H;��H;|�H;8�H;�H; �H;K�H;��H; I;�I;$I;�I;�
I;\I;�I;�I;I;AI;8I;�I;EI;XI;�I;      �)I;�)I;�(I;�'I;�%I;�#I;B!I;kI;gI;EI;�I;�I;(I;�
I;}I;EI;ZI;��H;
�H;��H;�H;l�H;��H;��H;��H;A�H;	�H;�H;<�H;|�H;��H;q�H;��H;��H;t�H;G�H;6�H;L�H;p�H;��H;��H;t�H;��H;{�H;5�H;�H;�H;D�H;��H;��H;��H;l�H;y�H;��H;
�H;��H;[I;HI;yI;�
I;)I;�I;�I;EI;gI;kI;C!I;�#I;�%I;�'I;�(I;�)I;      :I;�9I;�8I;7I;�4I;!2I;�.I;G+I;R'I;4#I;�I;�I;NI;.I;I; 
I;�I;�I;��H;��H;@�H;��H;��H;��H;��H;s�H;%�H;�H;��H;'�H;��H;��H;[�H;�H;��H;��H;��H;��H;��H;�H;\�H;��H;��H;%�H;��H;��H;#�H;y�H;��H;��H;��H;��H;9�H;��H;��H;�I;�I;!
I;I;+I;MI;�I;�I;4#I;R'I;G+I;�.I;2I;�4I;*7I;�8I;�9I;      'OI;�NI;�MI;}KI;yHI;�DI;�@I;�;I;�6I;�1I;,I;�&I;� I;�I;�I;�I;I;�I;�I;I;��H;��H;V�H;��H;��H;��H;k�H;(�H;�H;��H;#�H;{�H;��H;��H;C�H;�H;�H;�H;@�H;��H;��H;|�H;#�H;��H;��H;%�H;h�H;��H;��H;��H;Z�H;��H;��H;I;�I;�I;I;�I;�I;�I;� I;�&I;,I;�1I;�6I;�;I;�@I;�DI;�HI;�KI;�MI;�NI;      �bI;sbI;�aI;�`I;{^I;n[I; WI;�QI;)KI;2DI;=I;�5I;�.I;�'I;\!I;I;2I;�I;�
I;]I;OI;��H;m�H;��H;�H;��H;$�H;z�H;!�H;��H;��H;7�H;��H;)�H;��H;��H;��H;��H;��H;)�H;��H;7�H;��H;��H;�H;w�H;!�H;��H;�H;��H;o�H;��H;KI;\I;�
I;�I;2I;I;X!I;�'I;�.I;�5I;=I;3DI;#KI;�QI;WI;j[I;�^I;�`I;�aI;obI;      �GI;II;MI;�RI;'YI;�^I;�aI;ubI;�_I;EZI;lRI;�II;[@I;u7I;/I;"'I;�I;�I;�I;�I;�I;dI;E�H;��H;��H;O�H;�H;�H;|�H;#�H;��H;	�H;b�H;��H;r�H;;�H;4�H;>�H;q�H;��H;e�H;�H;�H;%�H;w�H;�H;
�H;U�H;��H;��H;H�H;cI;�I;�I;�I;�I;�I;'I;/I;r7I;]@I;�II;mRI;DZI;�_I;nbI;�aI;}^I;9YI;�RI;MI;II;      ��H;ȗH;D�H;��H;��H;�I;�%I;�@I;HTI;$_I;�aI;^I;�UI;KI;>@I;6I;�,I;�#I;�I;�I;�I;	I;)I;��H;-�H;�H;D�H;�H;,�H;i�H;%�H;�H;5�H;��H;5�H;��H;��H;��H;4�H;��H;6�H;�H;(�H;k�H;(�H;�H;D�H;�H;,�H;��H;.I;	I;�I;�I;�I;�#I;�,I;6I;<@I;KI;�UI;^I;�aI;#_I;ETI;�@I;�%I;�I;��H;��H;J�H;��H;      @VF;+hF;��F;��F;4MG;��G;F#H;��H;V�H;I;Y@I;�XI;PaI;�^I;�TI;�HI;�<I;�1I;�'I;�I;�I;I;�	I;�I; I;:�H;�H;[�H;��H;��H;v�H;E�H;:�H;x�H;�H;��H;}�H;��H;�H;x�H;=�H;G�H;z�H;��H;��H;X�H;�H;B�H; I;�I;�	I;I;�I;�I;�'I;�1I;�<I;�HI;�TI;�^I;PaI;�XI;Z@I;I;L�H;��H;J#H;��G;CMG;��F;��F;hF;      d�@;<�@;�`A;U&B;C;4D;�ME;�VF;�?G;%�G;ڐH;��H;�6I;�WI;-aI;)\I;�OI;BBI;�5I;�*I;� I;4I;�I;b
I;�I; I;,�H;��H;!�H;��H;��H;��H;G�H;x�H;��H;��H;c�H;��H;��H;{�H;I�H;��H;�H;��H;�H;��H;-�H; I;�I;`
I;�I;5I;� I;�*I;�5I;?BI;�OI;*\I;-aI;�WI;�6I;��H;֐H;%�G;�?G;�VF;�ME;�3D;#C;[&B;�`A;;�@;      7Y4;2�4;��5;	�7;��9;�<;��>;�A;#@C;:E;��F;.�G;b}H;c�H;�?I;�\I;`I;�UI;�FI;�8I;�,I;'"I;�I; I;\
I;�I;��H;��H;��H;��H;��H;��H;��H;��H;��H;��H;g�H;��H;��H;��H;��H;��H;��H;��H;��H;��H;��H;�I;Y
I;$I;�I;+"I;�,I;�8I;�FI;�UI;`I;�\I;�?I;c�H;b}H;+�G;��F;9E;@C;�A;��>;�<;ʫ9;(�7;��5;�4;      "�;��;l�;�/";��&;��+;��0;��5;��:;D�>;r B;��D;��F;��G;��H;�I;�RI;�`I;nYI;JI;;I;�-I;�"I;�I;�I;�	I;&I;I�H;o�H;S�H;��H;��H;��H;��H;��H;��H;d�H;��H;��H;��H;��H;��H;��H;X�H;k�H;H�H;)I;�	I;�I; I;�"I;�-I;;I; JI;pYI;�`I;SI;�I;��H;��G;��F;��D;r B;B�>;��:;��5;��0;��+;��&;�/";i�;Ŕ;      ���:l��:��:��:��;LN;^L;�, ;�f);��1;�w8;��=;^&B;�E;&G;KH;v�H;RGI;.`I;[I;�KI;�;I;�-I;,"I;0I;I;	I;cI;��H;��H;��H;i�H;x�H;�H;B�H;��H;g�H;��H;B�H;�H;x�H;h�H;��H;��H;��H;aI;	I;I;.I;3"I;�-I;�;I;�KI;�[I;/`I;RGI;x�H;KH;"G;�E;^&B;��=;�w8;��1;�f);�, ;WL;5N;��;��:��:Z��:      ���9p�:d�":�Q:��:x��:�?�:T��:�M
;��;'�&;
'1;e`9;�m?;T�C;>VF;%�G;��H;�=I;L_I;\I;�KI;;I;�,I;� I;�I;�I;�I;FI;��H;5�H;v�H;4�H;��H;��H;��H;��H;��H;��H;��H;5�H;u�H;6�H;��H;DI;�I;�I;�I;� I;�,I;;I;�KI;\I;O_I;�=I;��H;&�G;>VF;T�C;�m?;b`9;'1;%�&;��;�M
;^��:�?�:l��:��:�Q:��":8�:      ��Ѻ��Ⱥb������`��0(���9��Z:���:���:#0;S;5f);�4;��<;�KB;��E;"�G;u�H;\:I;R_I;[I;JI;9I;�*I;�I;�I;�I;\I;	I;��H;��H;�H;1�H;��H;3�H;��H;6�H;��H;-�H;�H;��H;��H;I;[I;�I;�I;�I;�*I;9I; JI;[I;Q_I;]:I;v�H;!�G;��E;�KB;��<;�4;2f);S;%0;���:���:��Z:�9�(�T�����d��� �Ⱥ      �5���R��d ��$6��T�X�B�$�8ۺ�H[�@	Q��c,:��:�:�>;D1";��0;��:;DaA;�cE;��G;s�H;�=I;+`I;nYI;�FI;�5I;�'I;�I;�I;�
I;�I;��H;�H;�H;��H;~�H;��H;<�H;��H;{�H;��H;�H;�H;��H;�I;�
I;�I;�I;�'I;�5I;�FI;nYI;+`I;�=I;v�H;��G;�cE;DaA;��:;��0;C1";�>;�:��:�c,: 
Q��H[�8ۺE�$�T�X�$6��g ���R��      G",���(�=H�FG��.���jλ*R���^e�Z��$�� PX���Z:B��:2�;o�;��-;ū9;sA;�cE; �G;��H;OGI;�`I;�UI;<BI;�1I;�#I;�I;�I;�I;�I;��H;G�H;��H;
�H;�H;��H;�H;�H;��H;H�H;�H;�I;�I;�I;�I;�#I;�1I;7BI;�UI;�`I;QGI;��H;!�G;�cE;sA;ë9;��-;m�;2�;B��:��Z: HX�*��\���^e�*R���jλ�.��FG�?H���(�      �d��B��������)���zl�RH��k"�z.���W��f�k��� ������9���:g��:�;�-;ȫ9;?aA;��E;)�G;u�H;�RI;`I;�OI;�<I;�,I;�I;1I;I;|I;TI;��H;��H;��H;��H;c�H;��H;��H;��H;��H;QI;~I;I;/I;�I;�,I;�<I;�OI;`I;SI;u�H;"�G;��E;BaA;ȫ9;�-;�;g��:���:��9����� �f�k��W��z.���k"�RH��zl��)������A���      ���i9�Z5��:��Tb̼|֮�t��� d�",�����Q��HG5�|#��p�f9|��:��:�;��-;��:;�KB;<VF;KH;�I;�\I; \I;�HI;6I;'I;I;�I;
I;BI;��H;��H;��H;X�H;��H;X�H;��H;��H;��H;?I;
I;�I;I;'I;6I;�HI;\I;�\I;�I;KH;6VF;�KB;��:;��-;�;��:x��:��f9z#��LG5��Q�����",�� d�u��|֮�Ub̼:��\5��i9�      �]��IY��ZN��`=���'�m����᷾������W��$�h��s�X��`9|��:]��:k�;��0;��<;T�C; G;��H;�?I;&aI;�TI;:@I;/I;[!I;�I;I;yI;�I;��H;}�H;�H;��H;�H;z�H;��H;�I;uI;I;�I;[!I;/I;:@I;�TI;#aI;�?I;��H;"G;M�C;��<;��0;h�;_��:t��: 9�u�X�h���$��W�����᷾����m���'��`=��ZN��IY�      �A��!��c���*��潅�>�d��`=����]��c֮�N�y�|�(��һ�]e�脮���f9���:2�;C1";�4;�m?;�E;��G;e�H;�WI;~^I;KI;q7I;�'I;�I;(I;�
I;!I;I;m�H;��H;;�H;��H;j�H;I;!I;�
I;%I;�I;�'I;r7I;KI;z^I;�WI;g�H;��G;�E;�m?;�4;@1";2�;���:��f9ꄮ��]e��һ}�(�N�y�d֮�]�꼗���`=�>�d�潅��*��c��!��      ���FE	��������Wн�A�����h���3���� ¼�)��1x/��һp�X�t#����9F��:�>;/f);g`9;]&B;��F;f}H;�6I;NaI;�UI;^@I;�.I;� I;JI;(I;�I;PI;Q I;��H;��H;��H;P I;NI;�I;%I;HI; !I;�.I;`@I;�UI;KaI;�6I;d}H;��F;]&B;``9;5f);�>;@��:��9x#��p�X��һ2x/��)�� ¼�����3��h��󑽠A���Wн��콺��FE	�      ~^Z�`
V��I��6�������ܽ!��ڽ���aG�Z�
�ȼ�)��}�(�h��KG5������Z:�:S;'1;��=;��D;.�G;��H;�XI;^I;{II;�5I;�&I;�I;�I;�
I;�I;MI;` I;��H;a I;KI;�I;�
I;�I;�I;�&I;�5I;~II;^I;�XI;��H;.�G;��D;��=;'1;S;�:��Z:���NG5�f��~�(��)��
�ȼZ��aG�ڽ��!���ܽ������6��I�`
V�      � ���e�����ە����q��I���"���������k���ZN�[�!¼O�y��$��Q���� � pX���:0;*�&;�w8;o B;��F;ԐH;T@I;�aI;lRI;=I;,I;�I;�I;\I;�I;4I;I;eI;I;4I;�I;\I;�I;�I;,I;=I;oRI;�aI;S@I;АH;��F;s B;�w8;�&;0;��: pX��� ��Q���$�O�y�!¼[��ZN�k������������"��I���q�ە������e��      d5�������W�Ҿ�a��z����l�	�6�DE	���Ƚk���aG����d֮��W����l�k�6���c,:���:��;��1;>�>;=E;"�G;I;#_I;@ZI;6DI;�1I;2#I;BI; I;
I;	I;�I;I;�I;	I;
I;�I;BI;2#I;�1I;:DI;EZI;"_I;I;�G;=E;D�>;��1;�;���:�c,:2��j�k�����W�d֮�����aG�k����ȽDE	�	�6��l�z����a��W�Ҿ������      {A��q<�ea/����:�{]׾� ��w��>�DE	�����ڽ����3�^�꼙���",��W��f���Q�z��:�M
;�f);��:;#@C;�?G;M�H;ETI;�_I;'KI;�6I;P'I;eI;�I;>I;�I;oI;�I;mI;�I;<I;�I;gI;O'I;�6I;*KI;�_I;GTI;P�H;�?G;'@C;��:;�f);�M
;���: Q�c���W��",�����^�꼘�3�ڽ������DE	�>�w��� ��{]׾�:���ea/��q<�      u�������a�{�l$_��q<�������}��w��	�6�����!���h����ⷾ�� d��.���^e�I[���Z:`��:�, ;��5;�A;�VF;��H;�@I;nbI;�QI;�;I;>+I;kI;I;9I;~	I;�I;.I;�I;	I;7I;I;kI;>+I;�;I;�QI;rbI;�@I;��H;�VF;�A;��5;�, ;T��:��Z:I[��^e�~.��� d�ⷾ�����h�!������	�6�w���}��������q<�l$_�a�{�����      <��������欿��� ����O��x����� ���l���"��ܽ���`=����u���k"�0R��Fۺ���9�?�:ZL;}�0;��>;�ME;H#H;�%I;�aI;�VI;�@I;�.I;<!I;@I;I;
I;MI;�I;LI;I;I;@I;=!I;�.I;�@I; WI;�aI;�%I;N#H;�ME;��>;��0;ZL;|?�:Г�9Fۺ.R���k"�u������`=����ܽ��"��l�� ����뾁x���O� ������欿����      �������L��jȿk���������O���{]׾z����I�����A��>�d�n�}֮�RH��jλQ�$��(�r��:@N;��+;�<;�3D;��G;�I;~^I;j[I;�DI;%2I;�#I;BI;�I;^I;�	I;�I;�	I;^I;�I;CI;�#I;!2I;�DI;l[I;�^I;�I;��G;�3D;�<;��+;CN;j��:�(�S�$��jλRH�}֮�n�>�d��A������I�z���{]׾����O�����k���jȿL�Ῡ��      @�1i�������I�ѿk��� ���q<��:��a����q����Wн罅���'�Tb̼�zl��.��P�X�\����:��;͎&;«9;!C;5MG;��H;5YI;�^I;�HI;�4I;�%I;�I;
I;�I;�
I;�	I;�
I;�I;I;�I;�%I;�4I;�HI;�^I;:YI;��H;@MG;!C;ƫ9;Ύ&;��;��:T��P�X��.���zl�Tb̼��'�罅��Wн����q��a���:��q<� ��k���I�ѿ������1i�      F:�.5�.�'��������jȿ���l$_���W�Ҿܕ���6�����*���`=�<�漮)��IG�(6�����,�Q:��:�/";�7;]&B;��F;��H;�RI;�`I;sKI;7I;�'I;;I;I;�I;oI;q
I;mI;�I;I;>I;�'I;7I;|KI;�`I;�RI;��H;��F;[&B;	�7;�/";��:�Q:���(6��HG��)��<���`=��*������6�ە��W�Ҿ��l$_����jȿ�������.�'�.5�      ��U�Z�O�H-?�.�'���M�ῴ欿a�{�ea/���뾝���I����d���ZN�\5������<H�f ��j�����":��:x�;��5;�`A;��F;H�H;MI;�aI;�MI;�8I;�(I;@I;�I;7I;I;	I;I;9I;�I;BI;�(I;�8I;�MI;�aI;MI;N�H;��F;�`A;��5;v�;��:|�":d���f ��<H�����[5���ZN�d������I�������ea/�a�{��欿M����.�'�H-?�Z�O�      ��i���b�Z�O�.5�1i�������������q<�����e��`
V�GE	�!���IY�j9�D�����(��R�� �Ⱥ`�:P��:�;?�4;>�@;hF;��H;II;ubI;�NI;�9I;�)I;�I;[I;�I;^I;^I;]I;�I;[I;�I;�)I;�9I;�NI;ybI;II;��H;*hF;;�@;?�4;ݔ;J��:T�:��Ⱥ�R����(�D���j9��IY�!��GE	�`
V��e������q<������������1i�.5�Z�O���b�      ඕ�S���Ѭ��.�_���7�{�}߿����,b��V�-l¾Hx�c.���Ž��t�)��f����?�N��(����x9���:N�;��2;3@@;_fF;6�H;}�I;O�I;|I;�[I;�CI;2I;�%I;[I;�I;2I;�I;ZI;�%I;2I;�CI;�[I;|I;O�I;��I;<�H;mfF;/@@;��2;J�;���: �x9%��N����?�f��)����t���Žc.�Hx�-l¾�V��,b����}߿{���7�.�_�Ѭ��S���      S���D���#}��+Y��3�����$ڿ%��Ľ\����(���s��3�5����p�c�S���<<�<������h��9I��:ϻ;N%3;Ep@;�yF;��H;��I;��I;�{I;H[I;LCI;�1I;P%I;I;WI;I;QI;I;N%I;�1I;NCI;E[I;�{I;�I;��I;��H;�yF;Dp@;L%3;˻;A��:H��9����<���<<�T��c��p�5����3��s�(�����Ľ\�$���$ڿ����3��+Y�#}�D���      Ѭ��#}�>tf��lG�ע%��p�.�ʿZ����>M����T�����d�Ȥ�̷�.�d��
��I���1�f���d�ຠ��9���:;�U4;��@;ұF;1�H;َI;��I;�yI;�YI;6BI;�0I;�$I;�I;�I;I;�I;�I;�$I;�0I;7BI;�YI;�yI;��I;܎I;4�H;߱F;��@;�U4;;���:���9Z��j����1��I���
�.�d�̷�Ȥ���d�T�������>M�Z���.�ʿ�p�ע%��lG�>tf�#}�      .�_��+Y��lG�f.�{���꿲���M䂿��5���󾍰��N�N�V��Q��!�Q����|���i!��g��p�h	:W
�:��;\16;��A;9G;�I;5�I;u�I;jvI;HWI;h@I;k/I;�#I;�I;
I;�I;I;�I;�#I;k/I;k@I;EWI;lvI;w�I;5�I; I;BG;��A;X16;��;O
�:T	:h񳺊g��i!�|������!�Q�Q��V��N�N���������5�M䂿�������{�f.��lG��+Y�      ��7��3�ע%�{��<����ſ	���½\�<����Ͼ����`�3��轻z��}�9�^�Ἓ���z��7}��dt��^:]+�:��#;��8;��B;sG;n%I;��I;�I;rI;TI;�=I;p-I;"I;HI;�I;zI;�I;JI;"I;p-I;�=I;TI;	rI;�I;��I;q%I;sG;��B;��8;��#;Y+�:��^:�dt��7}��z����^��}�9��z����`�3�������Ͼ<��½\�	�����ſ�<��{�ע%��3�      {�����p������ſ$���Ps���1�1r���d���d�|I�ΈŽ��}�_*�JC���^��B�~�D�G์ �:��;l);7;;'D;1�G;SHI;��I;��I;�lI;�OI;�:I;+I; I;�I;yI;,I;uI;�I; I;+I;�:I;�OI;�lI;��I;��I;SHI;7�G;&D;7;;j);��;~ �:G�~�D��B��^�JC��_*���}�ΈŽ|I��d��d��1r����1��Ps�$����ſ��꿃p����      }߿�$ڿ.�ʿ����	����Ps�QX:����%l¾�ǆ���7����85���Q�����t���75�m����� �8�ɼ:��;��.;��=;�EE;�YH;�hI;!�I;��I;%fI;KI;#7I;E(I;�I;�I;�I;wI;�I;�I;�I;E(I;#7I;KI;(fI;��I;#�I;�hI;�YH;�EE;��=;��.;��;�ɼ:��8���n���75��t������Q�85�������7��ǆ�%l¾���QX:��Ps�	�������.�ʿ�$ڿ      ���$��Z���M䂿½\���1�����J˾青�D�N�x��H������V�'�d�Ҽ��|��z��n��Rx����&:�P�:��;�W4;̠@;!gF;^�H;�I;�I;0�I;_I;�EI;3I; %I;BI;�I;�I;�I;�I;�I;BI;!%I;3I;�EI;_I;0�I;�I;�I;`�H;#gF;Ƞ@;�W4;��;�P�:��&:Px���n���z���|�d�ҼV�'����H���x��D�N�青��J˾�����1�½\�M䂿Z���$��      �,b�ý\��>M���5�<��1r��%l¾青�"&W��3�8Sؽ�z��ZG����}I����?���̻��-��
��
��:��;��&;|9;�C;�dG;HI;=�I;M�I;MvI;{WI;)@I;�.I;�!I;�I;UI;�I;�I;�I;VI;�I;�!I;�.I;)@I;|WI;OvI;Q�I;=�I;HI;�dG;�C;|9;��&;��;��:�
����-���̻��?�|I�����ZG��z��8Sؽ�3�"&W�青�%l¾1r��<����5��>M�ý\�      �V������������Ͼ�d���ǆ�D�N��3��c�[����\�3��)C���o���	� 숻\�x��9��:�h;K�/;2�=;EE;�2H;�WI;��I;�I;�kI;�OI;!:I;�)I;"I;�I;�I;�I;xI;�I;�I;�I;!I;�)I;!:I;�OI;�kI;��I;��I;�WI;�2H;BE;5�=;O�/;~h;��:���9`��눻��	��o�)C��3����\�[���c཰3�D�N��ǆ��d����Ͼ���������      ,l¾(��T������������d���7�x��8Sؽ[���d�C*�ckּ-\����'�-���R�p~��j�:�Z;ͣ#;5=7;$�A;�F;Q�H;l�I;�I;��I;�`I;�GI;�3I;'%I;rI;�I;SI;K
I;J	I;M
I;TI;�I;qI;$%I;�3I;�GI;�`I;��I;�I;h�I;V�H;�F;&�A;6=7;̣#;�Z;p�:`~���R�-����'�,\��ckּC*��d�[��8Sؽx����7��d���������T���(��      Gx��s���d�N�N�`�3�|I����H����z����\�C*��ݼI���0<<�
�ڻ�V�Tdt��&:z��:7C;�</;ID=;ψD;��G;�8I;ĘI;��I;tI;$VI;Z?I;�-I;d I;�I;ZI;�
I;�I;I;�I;�
I;]I;�I;b I;�-I;]?I;+VI;tI;��I;��I;�8I;��G;ԈD;LD=;�</;AC;���:�&:<dt��V�
�ڻ/<<�I����ݼC*���\��z��H������|I�`�3�N�N���d��s�      c.��3�Ȥ�V����ΈŽ75�����ZG�2��ckּI���yC��>�l6}������x9^��:	;(�&;�;8;��A;��F;��H;.yI;��I;�I;0fI;�KI;K7I;|'I;�I;�I;XI;I;�I;�I;�I;I;XI;�I;�I;�'I;O7I;�KI;1fI;�I;��I;2yI;��H;��F;��A;�;8;2�&;
	;\��:��x9���j6}��>� yC�H���ckּ3��YG����75��ΈŽ��V��Ȥ��3�      ��Ž5���̷�Q���z����}��Q�U�'����(C��,\��0<<��>n��H�຀�(��:*��:�;�'3;��>;�E;bH;]<I;ȗI;��I;�vI;�XI;�AI;u/I;�!I;�I;�I;S	I;cI;%I;tI;#I;bI;T	I;�I;�I;�!I;{/I;�AI;�XI;�vI;��I;͗I;[<I;dH;�E;��>;�'3;�;(��:6��:��D�ຆn���>�.<<�,\��(C�����U�'��Q���}��z��Q��̷�4���      ��t��p�.�d� �Q�}�9�_*����b�Ҽ|I���o���'�
�ڻl6}�H�ຠ9���:Pm�:��;��.;<;�oC;87G;��H;сI;ќI;хI;fI;<LI;�7I;�'I;�I;uI;OI;HI;�I;� I;Q I;� I;�I;JI;OI;rI;�I;�'I;�7I;BLI;fI;ͅI;ӜI;ρI;��H;<7G;�oC;<;��.;��;Zm�:��:�9�F��l6}��ڻ��'��o�{I��c�Ҽ���^*�}�9� �Q�.�d��p�      (��b��
����^��JC���t����|���?���	�,���V��������:��:�h;�+;��9;��A;wfF;S�H;r_I;��I;��I;sI;�VI;s@I;�.I;� I;TI;I;�I;jI;O I;�H;�H;~�H;L I;jI;�I;I;YI;� I;�.I;v@I;�VI;�rI;��I;��I;p_I;V�H;xfF;��A;��9;�+;�h;��:��:�� ����V�*����	���?���|��t��IC��_������
�b�      c��R���I��|�������^��75��z���̻�눻�R�<dt���x96��:^m�:�h;Y�*;ۍ8;��@;ۼE;5(H;b8I;��I;�I;G~I;�`I;�HI;�5I;[&I;tI;2I;�	I;�I;� I;��H;W�H;��H;S�H;��H;� I;�I;�	I;6I;uI;\&I;�5I;�HI;�`I;K~I;�I;��I;d8I;6(H;�E;��@;ԍ8;[�*;�h;Zm�:4��:��x9<dt��R��눻��̻�z��75��^����}����I��Q��      ��?��<<��1��h!��z��B�h���n����-�N�8~���&:V��:*��:��;�+;ҍ8;=�@;�]E;c�G;BI;�I;O�I;5�I;jiI;8PI;<I;�+I;�I;nI;PI;+I;sI;��H;��H;R�H;��H;O�H;��H;��H;pI;)I;TI;rI;�I;�+I; <I;1PI;liI;1�I;G�I;�I;CI;g�G;�]E;9�@;Ս8;�+;��;"��:R��:�&:(~��N𳺈�-��n��j���B黶z��h!��1��<<�      N��@��f����g���7}�n�D����<x��x
�����9��:���:	;�;��.;��9;��@;�]E;i�G;9I;�I;�I;K�I;�pI;�VI;�AI;|0I;�"I;�I;�I;�I;�I;��H;^�H;w�H;a�H;��H;^�H;t�H;\�H;��H;�I;�I;�I;�I;�"I;w0I;�AI;�VI;�pI;C�I;�I;�I;<I;g�G;�]E;��@;��9;��.;�;	;���:��:���9�
��>x�����u�D��7}��g��f���@��      &������P��N񳺨dt��F�`�8��&:��:��:�Z;?C;/�&;�'3;<;��A;�E;k�G;<I;U|I;��I;��I;~uI;o[I;FI;�4I;)&I;�I;II;�	I;�I;9�H;��H;6�H;u�H;�H;�H;z�H;q�H;5�H;��H;7�H;�I;�	I;FI;�I;%&I;~4I;FI;m[I;vuI;��I;ÜI;U|I;<I;f�G;߼E;��A;<;�'3;.�&;BC;�Z;��:��:��&: �8�F๐dt�h�h��ʎ��      ��x9�9��9X	:��^:� �:�ɼ:�P�:��;�h;Σ#;�</;�;8;��>;�oC;|fF;7(H;JI;�I;��I;��I;�wI;n^I;8II;�7I;)I;I;�I;�I;GI;L I;I�H;S�H;:�H;��H;��H;��H;��H;��H;9�H;Q�H;C�H;O I;II;�I;�I;I;)I;�7I;2II;f^I;�wI;��I;��I;�I;CI;6(H;zfF;�oC;��>;�;8;�</;ӣ#;�h;��;�P�:�ɼ:~ �:�^:L	:@��9�9      ���:c��:���:w
�:O+�:��;��;��;��&;R�/;==7;OD=;��A;�E;?7G;Z�H;h8I;�I;�I;��I;�wI;�_I;�JI;�9I;�*I;�I;4I;9I;I;9I;��H;��H;�H;=�H;��H;�H;��H;�H;��H;<�H;�H;��H;�H;8I;|I;;I;.I;�I;�*I;�9I;�JI;�_I;�wI;��I;�I;�I;g8I;V�H;=7G;�E;��A;PD=;?=7;M�/;��&;��;��;��;+�:_
�:���:G��:      f�;ϻ;;��;��#;t);��.;�W4;"|9;:�=;.�A;ۈD;��F;nH;��H;w_I;��I;R�I;J�I;}uI;m^I;�JI;':I; ,I;5 I;I;NI;�I;!I;��H;��H;4�H;�H;k�H;d�H;��H;T�H;��H;`�H;m�H;�H;0�H;�H;��H;I;�I;JI;I;: I;,I;:I;�JI;m^I;zuI;J�I;K�I;��I;t_I;��H;iH;��F;ڈD;2�A;6�=;"|9;�W4;��.;n);��#;��;;��;      ��2;Y%3;�U4;V16;��8;!7;;��=;ɠ@;�C;EE;�F;��G;��H;^<I;ρI;��I;�I;6�I;�pI;k[I;6II;�9I;,I;� I;I;I;SI;�I;H�H;c�H;Z�H;(�H;:�H;��H;��H;^�H;��H;Z�H;��H;��H;7�H;'�H;]�H;`�H;D�H;�I;LI;I;I;� I;,I;�9I;2II;g[I;�pI;/�I;�I;��I;΁I;X<I;��H;��G;�F;CE;�C;Ϡ@;��=;7;;��8;S16;�U4;Q%3;      R@@;Dp@;��@;��A;��B;4D;�EE;#gF;�dG;�2H;Z�H;�8I;0yI;ԗI;ٜI;��I;Q~I;siI;�VI;FI;�7I;�*I;> I;"I;]I;�I;=I;��H;��H;��H;�H;!�H;��H;n�H;��H;#�H;��H;�H;��H;o�H;��H;�H;�H;��H;��H;��H;6I;�I;^I;I;8 I;�*I;�7I;	FI;�VI;niI;Q~I;��I;֜I;ϗI;0yI;�8I;[�H;�2H;�dG;!gF;�EE;)D;��B;��A;��@;Ep@;      bfF;�yF;ӱF;=G;sG;>�G;�YH;n�H;NI;�WI;q�I;˘I;��I;��I;хI;sI;�`I;7PI;�AI;�4I;)I;�I;~I;I;�I;RI;��H;��H;��H;T�H;-�H;c�H;�H;*�H;r�H;�H;�H;�H;n�H;*�H;�H;a�H;-�H;Q�H;��H;��H;��H;UI;�I;I;{I;�I;)I;~4I;�AI;3PI;�`I;sI;΅I;��I;��I;ʘI;u�I;�WI;PI;l�H;�YH;1�G;sG;DG;ѱF;�yF;      M�H;��H;,�H;I;f%I;SHI;�hI;�I;A�I;��I;�I;��I;��I;�vI;fI;�VI;�HI;<I;~0I;+&I;I;2I;QI;VI;;I;��H;�H;��H;i�H;2�H;l�H;��H;��H;�H;i�H;�H;�H;�H;f�H;�H;��H;��H;l�H;/�H;c�H;��H;��H;��H;=I;QI;NI;4I;I;'&I;|0I;�;I;�HI;�VI;fI;�vI;�I;��I;�I;��I;?�I;�I;�hI;PHI;|%I;�I;+�H;��H;      ��I;�I;َI;?�I;��I;��I;-�I;�I;P�I;��I;��I;tI;-fI;�XI;;LI;u@I;�5I;�+I;�"I;�I;�I;8I;�I;�I;��H;��H;��H;^�H;G�H;\�H;��H;��H;��H;��H;��H;?�H;%�H;<�H;��H;��H;��H;��H;��H;[�H;B�H;\�H;��H;��H;��H;�I;�I;8I;�I;�I;�"I;�+I;�5I;v@I;:LI;�XI;+fI;tI;��I;��I;P�I;�I;+�I;��I;��I;@�I;َI;��I;      R�I;ޛI;��I;��I;ܔI;��I;��I;4�I;HvI;�kI;�`I;,VI;�KI;�AI;�7I;�.I;`&I;�I;�I;LI;�I;{I; I;G�H;��H;��H;c�H;E�H;a�H;��H;��H;��H;��H;#�H;��H;��H;O�H;}�H;��H;&�H;��H;��H;��H;��H;\�H;E�H;\�H;��H;��H;C�H; I;{I;�I;FI;�I;�I;`&I;�.I;�7I;�AI;�KI;(VI;�`I;�kI;LvI;4�I;��I;��I;�I;��I;��I;ۛI;      "|I;�{I;�yI;hvI;rI;�lI;'fI;!_I;{WI;�OI;�GI;d?I;O7I;}/I;�'I;� I;zI;kI;�I;�	I;NI;6I;��H;b�H;��H;M�H;0�H;a�H;��H;��H;��H;��H;��H;��H;�H;��H;��H;��H;	�H;��H;��H;��H;��H;��H;��H;^�H;)�H;P�H;��H;_�H;��H;8I;II;�	I;�I;iI;xI;� I;�'I;{/I;L7I;`?I;�GI;�OI;|WI;_I;,fI;�lI;rI;ovI;�yI;�{I;      �[I;e[I;�YI;UWI;TI;�OI;KI;�EI;-@I;':I;�3I;�-I;�'I;�!I;�I;YI;;I;VI;�I;�I;V I;�H;�H;]�H;�H;,�H;m�H;��H;��H;��H;~�H;��H;V�H;��H;w�H;Y�H;R�H;X�H;r�H;��H;W�H;��H;~�H;��H;��H;��H;i�H;-�H; �H;\�H;�H; �H;P I;�I;�I;SI;;I;[I;�I;�!I;�'I;�-I;�3I;(:I;-@I;�EI;%KI;�OI;TI;SWI;�YI;c[I;      �CI;WCI;6BI;b@I;�=I;�:I;#7I;3I;�.I;�)I;'%I;h I;�I;�I;uI;I;
I;.I;�I;>�H;P�H;��H;4�H;'�H;!�H;^�H;��H;��H;��H;��H;��H;A�H;��H;M�H;�H;��H;��H;��H;�H;O�H;��H;@�H;��H;��H;��H;��H;��H;_�H;#�H;!�H;7�H;��H;J�H;:�H;�I;.I;
I;I;uI;�I;�I;e I;(%I;�)I;�.I;3I;)7I;�:I;�=I;i@I;=BI;ZCI;      2I;�1I;�0I;n/I;p-I;
+I;?(I;%I;�!I;I;tI;�I;�I;�I;PI;�I;�I;tI;��H;��H;^�H;�H;�H;7�H;��H;�H;��H;��H;��H; �H;S�H;��H;2�H;��H;��H;~�H;m�H;~�H;��H;��H;0�H;��H;R�H;��H;��H;��H;��H;�H;��H;7�H;�H;�H;W�H;��H;��H;tI;�I;�I;PI;�I;�I;�I;wI; I;�!I;%I;B(I;+I;v-I;h/I;�0I;�1I;      �%I;S%I;�$I;�#I;"I; I;�I;HI;�I;�I;�I;cI;`I;Z	I;NI;nI;� I;��H;a�H;;�H;A�H;?�H;j�H;��H;i�H;%�H;�H;�H;'�H;��H;��H;N�H;��H;��H;[�H;8�H;$�H;8�H;[�H;��H;��H;O�H;��H;}�H;"�H;��H;�H;%�H;n�H;��H;n�H;<�H;;�H;5�H;^�H;��H;� I;oI;MI;Z	I;]I;`I;�I;�I;�I;EI;�I; I;"I;�#I;�$I;\%I;      NI;4I;�I;�I;TI;�I;�I;�I;[I;�I;^I;�
I;I;jI;�I;Q I;��H;��H;x�H;v�H;��H;��H;`�H;��H;��H;g�H;b�H;��H;��H;�H;n�H;�H;��H;Z�H;�H;�H;�H;�H;�H;\�H;��H;�H;n�H;�H;��H;��H;b�H;i�H;��H;��H;c�H;��H;��H;r�H;v�H;��H;��H;V I;�I;lI;I;�
I;aI;�I;\I;�I;�I;�I;QI;�I;�I;5I;      �I;]I;�I;I;�I;sI;�I;�I;�I;�I;R
I; I;�I;(I;� I;|�H;W�H;N�H;b�H;|�H;��H;�H;��H;O�H;�H;�H;�H;A�H;��H;��H;V�H;��H;��H;6�H;�H;��H;��H;��H;�H;<�H;��H;��H;V�H;��H;��H;>�H;�H;�H;�H;Q�H;��H;�H;��H;z�H;`�H;R�H;Z�H;��H;� I;)I;�I;�I;T
I;�I;�I;�I;�I;sI;�I;
I;�I;kI;      7I;�I;�I;�I;sI;%I;zI;�I;�I;xI;U	I;I;�I;|I;X I;�H;��H;��H;��H; �H;��H;��H;S�H;��H;��H;�H;�H;,�H;V�H;��H;M�H;��H;p�H; �H;�H;��H;��H;��H;�H;!�H;q�H;��H;N�H;��H;P�H;&�H;�H;	�H;��H;��H;W�H;��H;��H;�H;��H;��H;��H;�H;X I;|I;�I;I;U	I;yI;�I;�I;�I;%I;sI;�I;�I;I;      �I;^I;�I;I;�I;vI;�I;�I;�I;�I;Q
I; I;�I;)I;� I;|�H;W�H;N�H;b�H;|�H;��H;�H;��H;O�H;�H;�H;�H;A�H;��H;��H;V�H;��H;��H;8�H;�H;��H;��H;��H;�H;;�H;��H;��H;V�H;��H;��H;<�H;�H;�H;�H;P�H;��H;�H;��H;z�H;`�H;R�H;X�H;��H;� I;&I;�I;�I;R
I;�I;�I;�I;�I;uI;�I;I;�I;eI;      DI;4I;�I;�I;TI;�I;�I;�I;[I;�I;_I;�
I;I;lI;�I;Q I;��H;��H;w�H;v�H;��H;��H;_�H;��H;��H;f�H;b�H;��H;��H;�H;m�H;�H;��H;Z�H;�H;�H;�H;�H;�H;\�H;��H;�H;n�H;�H;��H;��H;b�H;j�H;��H;��H;c�H;��H;��H;r�H;w�H;��H;��H;V I;�I;jI;I;�
I;^I;�I;\I;�I;�I;�I;UI;�I;�I;;I;      �%I;P%I;�$I;�#I;	"I; I;�I;KI;�I;�I;�I;aI;]I;Z	I;OI;nI;� I;��H;`�H;9�H;A�H;?�H;j�H;��H;l�H;%�H;�H;�H;)�H;��H;��H;N�H;��H;��H;\�H;6�H;$�H;8�H;Z�H;��H;��H;O�H;��H;}�H;"�H;��H;�H;(�H;o�H;��H;n�H;=�H;;�H;6�H;a�H;��H;� I;qI;NI;X	I;[I;^I;�I;�I;�I;HI;�I; I;"I;�#I;�$I;T%I;      2I;�1I;�0I;e/I;m-I;+I;?(I;#%I;�!I;I;tI;�I;�I;�I;SI;�I;�I;tI;��H;��H;\�H;�H;�H;7�H;��H;�H;��H;��H;��H;��H;R�H;��H;0�H;��H;��H;~�H;m�H;~�H;��H;��H;/�H;��H;R�H;��H;��H;��H;��H;�H;��H;4�H;�H;�H;U�H;��H;��H;tI;�I;�I;PI;�I;�I;�I;rI;I;�!I; %I;F(I;
+I;t-I;r/I;�0I;�1I;      �CI;YCI;)BI;`@I;�=I;�:I;(7I;3I;�.I;�)I;+%I;h I;�I;�I;xI;I;
I;.I;�I;;�H;Q�H;��H;4�H;&�H;#�H;^�H;��H;��H;��H;��H;��H;>�H;��H;K�H;�H;��H;��H;��H;�H;M�H;��H;@�H;��H;��H;��H;��H;��H;a�H;!�H;�H;9�H;��H;I�H;:�H;�I;.I;
I;I;tI;�I;�I;g I;'%I;�)I;�.I;3I;(7I;�:I;�=I;i@I;/BI;VCI;      �[I;e[I;�YI;LWI;TI;�OI;KI;�EI;-@I;':I;�3I;�-I;�'I;�!I;�I;[I;<I;SI;�I;�I;W I;�H;�H;]�H; �H;)�H;j�H;��H;��H;��H;|�H;��H;V�H;��H;w�H;X�H;Q�H;Y�H;r�H;��H;W�H;��H;}�H;��H;��H;��H;h�H;/�H;�H;Y�H;�H;�H;P I;�I;�I;SI;=I;\I;�I;�!I;�'I;�-I;�3I;%:I;.@I;�EI;"KI;�OI;TI;YWI;�YI;d[I;      +|I;�{I;�yI;qvI;�qI;�lI;'fI;#_I;}WI;�OI;�GI;d?I;N7I;{/I;�'I;� I;zI;lI;�I;�	I;PI;9I;��H;`�H;��H;L�H;-�H;_�H;��H;��H;��H;��H;��H;�H;�H;��H;��H;��H;	�H;�H;��H;��H;��H;��H;��H;\�H;,�H;Q�H;��H;\�H;��H;9I;JI;�	I;�I;kI;xI;� I;�'I;{/I;L7I;^?I;�GI;�OI;yWI;!_I;(fI;�lI;rI;yvI;�yI;�{I;      Y�I;ޛI;��I;��I;˔I;��I;��I;2�I;RvI;�kI;�`I;+VI;�KI;�AI;�7I;�.I;`&I;�I;�I;GI;�I;|I;I;H�H;��H;��H;_�H;G�H;a�H;��H;��H;��H;��H;#�H;��H;�H;N�H;�H;��H;#�H;��H;��H;��H;��H;[�H;A�H;^�H;��H;��H;@�H;!I;|I;�I;GI;�I;�I;_&I;�.I;�7I;�AI;�KI;'VI;�`I;�kI;KvI;4�I;��I;��I;ݔI;��I;��I;؛I;      ��I;��I;̎I;<�I;��I;��I;-�I;"�I;P�I;��I;��I;tI;+fI;�XI;<LI;v@I;�5I;�+I;�"I;�I;�I;9I;�I;�I;��H;��H;��H;^�H;H�H;Z�H;��H;��H;��H;��H;��H;<�H;&�H;>�H;��H;��H;��H;��H;��H;[�H;B�H;Z�H;��H;��H;��H;�I;�I;8I;�I;�I;�"I;�+I;�5I;v@I;;LI;�XI;-fI;tI;��I;��I;N�I;�I;-�I;��I;��I;=�I;ڎI;��I;      ;�H;��H;*�H;I;t%I;ZHI;�hI;�I;@�I;��I;�I;��I;�I;�vI;fI;�VI;�HI;<I;}0I;(&I;I;4I;KI;WI;;I;��H; �H;��H;h�H;-�H;i�H;��H;��H;�H;h�H;�H;�H;�H;e�H;�H;��H;��H;l�H;/�H;e�H;��H;��H;��H;:I;QI;QI;4I;I;)&I;~0I;<I;�HI;�VI;fI;�vI;�I;��I;�I;��I;=�I;�I;�hI;THI;y%I;I;,�H;��H;      XfF;�yF;ݱF;4G;sG;D�G;�YH;n�H;QI;�WI;q�I;̘I;��I;��I;҅I;sI;�`I;7PI;�AI;}4I;	)I;�I;{I;I;�I;NI;��H; �H;��H;P�H;,�H;b�H;�H;*�H;q�H;�H;�H;�H;n�H;*�H;�H;c�H;0�H;Q�H;��H;��H;��H;VI;�I;I;~I;�I;)I;�4I;�AI;4PI;�`I;sI;ԅI;��I;��I;ȘI;t�I;�WI;GI;e�H;�YH;3�G;sG;9G;űF;�yF;      P@@;Dp@;��@;��A;��B;4D;�EE;"gF;�dG;�2H;[�H;�8I;/yI;їI;ۜI;��I;Q~I;riI;�VI;	FI;�7I;�*I;8 I;!I;]I;�I;9I;��H;��H;��H;�H;�H;��H;n�H;��H;�H;��H;�H;��H;o�H;��H;�H;�H;��H;��H;��H;:I;�I;ZI;I;; I;�*I;�7I;FI;�VI;oiI;R~I;��I;ۜI;їI;2yI;�8I;W�H;�2H;�dG;"gF;�EE;)D;��B;��A;��@;Cp@;      ��2;D%3;�U4;Z16;��8;$7;;��=;ˠ@;�C;CE;�F;��G;��H;Z<I;сI;��I;�I;5�I;�pI;h[I;5II;�9I;,I;� I;I;I;OI;�I;G�H;_�H;\�H;(�H;9�H;��H;��H;[�H; �H;]�H;��H;��H;;�H;(�H;`�H;b�H;F�H;�I;PI;I;I;� I;,I;�9I;5II;j[I;�pI;3�I;�I;��I;ρI;Z<I;��H;��G;�F;BE;�C;Š@;��=;7;;��8;x16;�U4;-%3;      V�;λ;
;��;��#;r);��.;�W4;%|9;9�=;(�A;ۈD;��F;jH;��H;x_I;��I;Q�I;H�I;zuI;k^I;�JI; :I;,I;7 I;wI;KI;�I;"I;��H;��H;3�H;�H;k�H;c�H;��H;U�H;��H;`�H;h�H;�H;3�H;�H;��H;I;�I;NI;I;5 I;,I;":I;�JI;n^I;}uI;M�I;L�I;��I;x_I;��H;gH;��F;وD;*�A;9�=;$|9;�W4;��.;p);��#;�;;��;      ���:_��:���:W
�:I+�:��;��;��;��&;M�/;<=7;QD=;��A;�E;@7G;Z�H;g8I;�I;�I;��I;�wI;�_I;�JI;�9I;�*I;�I;1I;;I;~I;6I;��H;��H;�H;<�H;��H;�H;��H;�H;��H;;�H;�H;��H;�H;;I;|I;9I;4I;�I;�*I;�9I;�JI;�_I;�wI;��I;�I;�I;g8I;Z�H;<7G;�E;��A;MD=;==7;M�/;��&;��;��;x�;{+�:G
�:���:O��:      ��x9���9`��9L	:��^:� �:�ɼ:�P�:��;~h;У#;�</;�;8;��>;�oC;{fF;5(H;FI;�I;��I;��I;�wI;i^I;5II;�7I;�(I;I;�I;�I;DI;J I;H�H;Q�H;=�H;��H;��H;��H;��H;��H;9�H;S�H;F�H;O I;II;�I;�I;I;)I;�7I;9II;j^I;�wI;��I;��I;�I;FI;6(H;zfF;�oC;��>;�;8;�</;ѣ#;�h;��;�P�:�ɼ:� �:�^:X	:���9��9      ������V��N񳺨dt��F� �8��&:��:��:�Z;AC;/�&;�'3;<;��A;޼E;g�G;9I;T|I;ÜI;��I;zuI;m[I;FI;|4I;$&I;�I;II;�	I;�I;9�H;��H;6�H;t�H;z�H;�H;{�H;q�H;2�H;��H;7�H;�I;�	I;GI;�I;(&I;�4I;FI;r[I;}uI;��I;ÜI;W|I;=I;f�G;߼E;��A;<;�'3;.�&;>C;�Z;��:��:��&:��8G๤dt�b�Z�຦���      N��@��f����g���7}�p�D����Bx���
�����9~�:���:	;�;��.;��9;��@;�]E;f�G;9I;�I;�I;H�I;�pI;�VI;�AI;w0I;�"I;�I;�I;�I;�I;��H;]�H;w�H;`�H;��H;`�H;t�H;\�H;��H;�I;�I;�I;�I;�"I;z0I;�AI;VI;�pI;J�I;�I;�I;=I;g�G;�]E;��@;��9;��.;�;	;���:~�:���9�
��Bx�����r�D��7}��g��i���=��      ��?��<<��1��h!��z��B�h���n����-�R�8~���&:R��:&��:��;�+;ҍ8;9�@;�]E;d�G;BI;�I;O�I;3�I;liI;1PI;�;I;�+I;�I;kI;SI;+I;qI;��H;��H;O�H;��H;Q�H;��H;��H;sI;(I;TI;nI;�I;�+I;<I;4PI;hiI;3�I;N�I;�I;BI;h�G;�]E;:�@;ҍ8;�+;��;"��:R��:�&:(~��T𳺋�-��n��h���B黶z��h!��1��<<�      c��R���I��|�������^��75��z���̻�눻�R�<dt���x94��:^m�:�h;[�*;Ս8;��@;ܼE;6(H;b8I;��I;�I;L~I;�`I;�HI;�5I;_&I;qI;5I;�	I;�I;� I;��H;V�H;��H;V�H;��H;� I;�I;�	I;6I;tI;]&I;�5I;�HI;�`I;H~I;�I;��I;e8I;3(H;߼E;��@;ԍ8;Y�*;�h;Zm�:4��:��x9Ddt��R��눻��̻�z��75��^����}����I��Q��      (��b��
����^��IC���t����|���?���	�+���V� ���@���:��:�h;�+;��9;��A;zfF;W�H;u_I;��I;��I; sI;�VI;r@I;�.I;� I;XI;I;�I;mI;Q I;~�H;�H;~�H;L I;hI;�I;	I;VI;� I;�.I;u@I;�VI;�rI;��I;��I;u_I;W�H;tfF;��A;��9;�+;�h;��:��:������V�,����	���?���|��t��JC��_������
�b�      ��t��p�.�d� �Q�}�9�^*����c�Ҽ|I���o���'�
�ڻl6}�H�ຠ9���:Xm�:��;��.;<;�oC;:7G;��H;сI;՜I;хI;fI;<LI;�7I;�'I;�I;tI;NI;KI;�I;� I;P I;� I;�I;JI;NI;qI;�I;�'I;�7I;<LI;fI;΅I;ќI;ҁI;��H;=7G;�oC;<;��.;��;Xm�:��:�9�F��m6}�
�ڻ��'��o�|I��c�Ҽ���^*�}�9�!�Q�.�d��p�      ��Ž4���̷�Q���z����}��Q�U�'����)C��,\��/<<��>n��D�຀�.��:&��:�;�'3;��>;�E;fH;^<I;ϗI;��I;�vI;�XI;�AI;v/I;�!I;�I;�I;T	I;cI;"I;tI;%I;aI;T	I;�I;�I;�!I;y/I;�AI;�XI;�vI;��I;ȗI;^<I;jH;�E;��>;�'3;
�;&��:0��:��H�ຆn���>�0<<�,\��)C�����U�'��Q���}��z��Q��̷�4���      c.��3�Ȥ�V����ΈŽ75�����ZG�3��ckּI��� yC��>�i6}������x9\��:	;,�&;�;8;��A;��F;��H;0yI;��I;�I;-fI;�KI;L7I;'I;�I;�I;[I;I;�I;�I;�I;I;XI;�I;�I;}'I;N7I;�KI;.fI;�I;��I;.yI;��H;��F;��A;�;8;/�&;	;V��:��x9���j6}��>�yC�H���ckּ3��ZG����85��ΈŽ��V��Ȥ��3�      Hx��s���d�N�N�`�3�|I����H����z����\�C*��ݼI���0<<�
�ڻ�V�Pdt��&:|��:;C;�</;LD=;ֈD;��G;�8I;ØI;��I;tI;(VI;Y?I;�-I;b I;�I;]I;�
I;�I;I;�I;�
I;\I;�I;a I;�-I;\?I;+VI;tI;��I;��I;�8I;��G;وD;MD=;�</;>C;z��:�&:Hdt��V�	�ڻ0<<�I����ݼC*���\��z��H������|I�`�3�N�N���d��s�      ,l¾(��T������������d���7�x��8Sؽ[���d�C*�ckּ-\����'�.���R�p~��n�:�Z;ѣ#;8=7;*�A;�F;T�H;k�I;�I;��I;�`I;�GI;�3I;'%I;qI;�I;TI;M
I;L	I;M
I;TI;�I;rI;$%I;�3I;�GI;�`I;��I;�I;k�I;S�H;�F;+�A;8=7;ǣ#;�Z;h�:p~���R�.����'�-\��dkּC*��d�[��8Sؽx����7��d���������T���(��      �V������������Ͼ�d���ǆ�D�N��3��c�[����\�3��)C���o���	� 숻b𳺀��9��:�h;L�/;6�=;FE;�2H;�WI;��I;�I;�kI;�OI;":I;�)I;"I;�I;�I;�I;xI;�I;�I;�I;"I;�)I;":I;�OI;�kI;��I;��I;�WI;�2H;FE;9�=;M�/;zh;��:h��9b��눻��	��o�)C��3����\�[���cཱ3�D�N��ǆ��d����Ͼ���������      �,b�ý\��>M���5�<��1r��%l¾青�"&W��3�8Sؽ�z��ZG����|I����?���̻��-��
����:��;��&;|9;�C;�dG;HI;<�I;N�I;PvI;{WI;,@I;�.I;�!I;�I;UI;�I;�I;�I;VI;�I;�!I;�.I;)@I;yWI;RvI;P�I;=�I;JI;�dG;�C;|9;��&;��;��:�
����-���̻��?�|I�����ZG��z��8Sؽ�3�"&W�青�%l¾1r��<����5��>M�ý\�      ���$��Z���M䂿½\���1�����J˾青�D�N�x��H������V�'�d�Ҽ��|��z��n��Px����&:�P�:��;�W4;͠@;"gF;]�H;�I;�I;0�I;_I;�EI;3I;!%I;DI;�I;�I;�I;�I;�I;DI; %I;3I;�EI;_I;1�I;�I;�I;`�H;!gF;̠@;�W4;��;�P�:��&:Rx���n���z���|�d�ҼV�'����H���x��D�N�青��J˾�����1�½\�M䂿Z���$��      }߿�$ڿ.�ʿ����	����Ps�QX:����%l¾�ǆ���7����85���Q�����t���75�o�����`�8�ɼ:��;��.;��=;�EE;�YH;�hI; �I;��I;%fI;KI;#7I;E(I;�I;�I;�I;wI;�I;�I;�I;E(I;%7I;KI;(fI;��I;#�I;�hI;�YH;�EE;��=;��.;��;�ɼ:��8���n���75��t������Q�85�������7��ǆ�%l¾���QX:��Ps�	�������.�ʿ�$ڿ      {�����p������ſ$���Ps���1�1r���d���d�|I�ΈŽ��}�_*�JC���^��B�}�D�G๊ �:��;l);7;;&D;0�G;QHI;��I;��I;�lI;�OI;�:I;+I; I;�I;yI;-I;yI;�I; I;+I;�:I;�OI;�lI;��I;��I;THI;8�G;'D;7;;n);��;� �:�Fเ�D��B��^�JC��_*���}�ΈŽ|I��d��d��1r����1��Ps�$����ſ��꿃p����      ��7��3�ע%�{��<����ſ	���½\�<����Ͼ����`�3��轻z��}�9�^�Ἒ���z��7}��dt��^:Y+�:��#;��8;��B;sG;m%I;��I;�I;rI;TI;�=I;p-I;"I;GI;�I;zI;�I;JI;"I;p-I;�=I;TI;	rI;�I;��I;t%I;sG;��B;��8;��#;]+�:��^:�dt��7}��z����^��}�9��z����`�3�������Ͼ<��½\�	�����ſ�<��{�ע%��3�      .�_��+Y��lG�f.�{���꿲���M䂿��5���󾍰��N�N�V��R��!�Q����|���i!��g��h�h	:Q
�:��;V16;��A;6G;�I;3�I;u�I;hvI;IWI;i@I;j/I;�#I;�I;	I;�I;I;�I;�#I;m/I;k@I;HWI;nvI;w�I;6�I;I;BG;��A;Z16;��;Q
�:T	:h񳺌g�� i!�|������!�Q�Q��V��N�N���������5�M䂿�������{�f.��lG��+Y�      Ѭ��#}�>tf��lG�ע%��p�.�ʿZ����>M����T�����d�Ȥ�̷�.�d��
��I���1�h���`�ຠ��9���:;�U4;��@;ѱF;/�H;َI;��I;�yI;�YI;6BI;�0I;�$I;�I;�I;�I;�I;�I;�$I;�0I;7BI;�YI;�yI;��I;ݎI;5�H;߱F;��@;�U4;;���:���9X��h����1��I���
�.�d�̷�Ȥ���d�T�������>M�Z���.�ʿ�p�ע%��lG�>tf�#}�      S���D���#}��+Y��3�����$ڿ%��Ľ\����(���s��3�5����p�c�S���<<�;������x��9I��:λ;L%3;Ep@;�yF;��H;��I;��I;�{I;I[I;LCI;�1I;Q%I;I;TI;I;QI;I;P%I;�1I;OCI;E[I;�{I;�I;��I;��H;�yF;Cp@;N%3;˻;C��:@��9����=���<<�T��c��p�5����3��s�(�����Ľ\�%���$ڿ����3��+Y�#}�D���      ����,������T���J�Q�ř$�4�����<�}�H(�@�׾�T���L+���սj����L���iO���ͻ���� m8jo�:[�;R�1;��?;�uF;d I;f�I;��I;��I;VvI;�WI;�AI;�1I;�'I;�!I;�I;�!I;�'I;�1I;�AI;�WI;VvI;��I;��I;h�I;g I;�uF;��?;Q�1;W�;do�:�m8�����ͻ�iO�L����j����ս�L+��T��@�׾H(�<�}���4���ƙ$�J�Q�T��������,��      �,��a��#P���{���K��x �����p�����w��$���Ҿf���  (���ѽҷ��'�����K�Fɻ,��`��8x��:z�;��1;�@;k�F;I;ݿI;�I;��I;�uI;#WI;fAI;�1I;�'I;�!I;�I;�!I;�'I;�1I;hAI;%WI;�uI;��I;�I;޿I;I;w�F;�@;��1;v�;p��:���8)��Fɻ�K����'�ҷ����ѽ  (�f�����Ҿ�$���w�p��������x ���K��{�#P��a��      ����#P�������d���;�#���㿲���#f�d��ž��z���<�ƽ%0v�T5�1����o@�����i��`u9AK�:];�73;"�@;��F;FI;��I;M�I;S�I;�sI;�UI;A@I;�0I;�&I;!I;0I;!I;�&I;�0I;A@I;�UI;�sI;V�I;L�I;��I;GI;��F;�@;�73;];7K�:``u9zi������o@�2���T5�%0v�<�ƽ����z�žd��#f�������#����;���d����#P��      T����{���d��F�ř$�:����ɿ.蒿��K�P���j���Yb�F�1���s�a����?�����.��d��r�غ���9�Y�:.X;�25;#�A;Y!G;I7I;s�I;B�I;R�I;�pI;�SI;>I;y/I;�%I;" I;/I; I;�%I;v/I;>I;�SI;�pI;R�I;@�I;q�I;H7I;b!G;�A;�25;*X;�Y�:���9p�غ�d����.�@������s�a�1���F��Yb��j��P����K�.蒿��ɿ:��ř$��F���d��{�      J�Q���K���;�ř$��;
��޿�����w�r,���澝���'�D������I��$�G�����N��������X�����9:Z��:�n!;��7;��B;J�G;�YI;*�I;W�I;��I;�lI;sPI;<I;�-I;$I;�I;�I;�I;$I;�-I;<I;uPI;�lI;��I;W�I;,�I;�YI;Q�G;��B;��7;�n!;V��:t�9:V����������N�����$�G��I������'�D��������r,���w�����޿�;
�ř$���;���K�      ř$��x �#��:���޿o���ʅ���F�}�
��~����z��$���ս���A2+���ϼPp�����P�]� �*���:�;�8';��:;��C;�H;�}I;�I;o�I;׋I;kgI;�LI;9I;7+I;!"I;�I;)I;�I; "I;4+I;9I;�LI;ggI;ًI;p�I;�I;�}I;H;��C;��:;�8';�;��:�*�Q�]�����Pp���ϼA2+������ս�$���z��~��}�
��F�ʅ��o����޿:��"���x �      4��������㿊�ɿ���ʅ����P�d��;�׾�`��S�H����@��R�a���͡���D��ɻ� ��ح��W�:�;`I-;7|=;CE;��H;�I;��I;s�I;��I;haI;"HI;�5I;p(I;�I;�I;QI;�I;�I;p(I;�5I; HI;eaI;��I;s�I;��I;�I;��H; CE;5|=;`I-;�;�W�:@ح�� ��ɻ�D�͡����R�a��@����S�H��`��;�׾d����P�ʅ�������ɿ�㿳���      ��p�������.蒿��w��F�d��ʰ� ����Yb�)����ѽ�%��D4�؟�X�����H���潺���9Br�:��;�93;%Q@;zvF;�H;�I;��I;��I;�zI;�ZI;CI;�1I;b%I;?I;�I;"I;�I;BI;c%I;�1I;CI;�ZI;�zI;��I;��I;�I;�H;}vF;!Q@;�93;��;:r�:Ȓ�9�潺H�����X��؟�D4��%����ѽ)���Yb� ���ʰ�d���F���w�.蒿����p���      <�}���w�#f���K�r,�}�
�;�׾ �����k���'�ez꽝I���;V�<M�	����iO�mG�soE�̱�2��:B� ;��$;��8;[�B;��G;,KI;�I;�I;@�I;qI;�SI;�=I;�-I;"I;jI;I;�I;I;mI;"I;�-I;�=I;�SI;	qI;A�I;�I;�I;+KI;��G;Y�B;��8;��$;>� ;>��:ȱ�soE�jG໫iO�	���<M��;V��I��ez���'���k� ���;�׾}�
�r,���K�#f���w�      H(��$�d��P������~���`���Yb���'��U�G$��D�m�&����ϼ�/��>��������غ08�94��:�F;�G.;|=;GE;�\H;�I;s�I;y�I;��I;gI; LI;�7I;)I;pI;rI;rI;'I;qI;rI;pI;)I;�7I; LI;gI;��I;|�I;q�I;�I;�\H;DE;|=;�G.;�F;B��:88�9��غ����>���/����ϼ&��D�m�G$���U���'��Yb��`���~�����P��d���$�      ?�׾��Ҿž�j��������z�S�H�)��ez�G$���/v�2+�ސ�����5��ɻ<4�P(��~��:T��:5o!;P6;lA;��F;p�H;��I;��I;ߦI;F}I;�\I;[DI;	2I;r$I;�I;HI;�I;�I;�I;II;�I;p$I;2I;]DI;�\I;J}I;�I;��I;��I;s�H;��F;lA;P6;5o!;h��:���:P(��64��ɻ��5���ސ�2+��/v�G$��ez�)��S�H���z������j��ž��Ҿ      �T��f�����z��Yb�&�D��$�����ѽ�I��D�m�2+�������L�K�ﻘ�p�P������9!T�:�/;o�-;d�<;BzD;ZH;�mI;��I;|�I;��I;�oI;�RI;�<I;,I;�I;I;/I;�I;�I;�I;.I;I;�I; ,I;�<I;�RI;�oI;��I;z�I;��I;�mI;WH;FzD;j�<;o�-;�/;'T�:���9D�����p��K�K�������2+�D�m��I����ѽ���$�'�D��Yb���z�f���      �L+�  (���F�������ս�@���%���;V�%��ސ������MS�M��&��xD���n8q�:�;a�$;�^7;(�A;d�F;��H;_�I;b�I;��I;��I;QbI;�HI;5I;(&I;/I;>I;�I;�
I;
I;�
I;�I;>I;/I;$&I;5I;�HI;VbI;�I;��I;]�I;c�I;��H;e�F;.�A;�^7;k�$;�;�p�:��n8tD�&��L���MS�����ސ�%���;V��%���@����ս����F���  (�      ��ս��ѽ;�ƽ1����I�����R�a�D4�<M���ϼ��K�K�O��NG��af���o���:�B�:�Y;��1;Ol>;�E;�/H;qI;��I;��I;ژI;�rI;�UI;�>I;�-I;b I;�I;�I;�
I;I;0I;I;�
I;�I;�I;^ I;�-I;�>I;�UI;sI;טI;��I;��I;qI;�/H;�E;Ol>;��1;�Y;�B�:��:��o�^f�LG��N��K�K�����ϼ<M�D4�Q�a�����I��1���;�ƽ��ѽ      j��ѷ��%0v�r�a�$�G�@2+���ן�	����/����5��'��_f��ج��g:3�:�;I-;g;;�NC;SG;�I;ɶI;�I;��I;	�I;
cI;~II;�5I;n&I;�I;7I;�I;�I;PI;XI;NI;�I;�I;9I;�I;r&I;�5I;�II;cI;�I;��I;�I;ȶI;�I;
SG;�NC;g;;I-;�;;�:�g:�ج�]f�&�����5��/�����ן���@2+�$�G�r�a�%0v�ѷ��      
��&�T5���������ϼ̡��X���iO�>���ɻ��p��D���o��g:�_�:CG;n*;o9;��A;�uF;�H;��I;��I;��I;H�I;�pI;3TI;M>I;-I;�I;}I;�I;VI;�I;�I;�I;�I;�I;VI;�I;xI;�I;-I;Q>I;7TI;�pI;?�I;��I;��I;��I;�H;�uF;��A;p9;j*;CG;�_�:�g:��o��D⺙�p��ɻ>���iO�X��͡����ϼ������T5�&�      L�����2���?����N��Pp��D����gG�����34�>�����n8��:?�:JG;�(;��7;Y�@;��E;KQH;mI;��I;��I;��I;#}I;�^I;�FI;�3I;�$I;\I;�I;�	I;I;�I;��H;P�H;��H;�I;I;�	I;�I;_I;�$I;�3I;�FI;�^I;}I;��I;��I;�I;mI;NQH;��E;Z�@;��7;�(;EG;?�:��:��n8B���04�����hG໇���D�Pp��N��@���3������      �iO���K��o@���.���������ɻ H��loE���غ((�����9�p�:�B�:�;l*;��7;�P@;�\E;�H;�II;~�I;h�I;�I;V�I;<hI;�NI;b:I;9*I;xI;�I;�I;I;I;2�H;b�H;��H;^�H;/�H;I;I;�I;�I;zI;7*I;c:I;�NI;7hI;\�I;�I;a�I;�I;�II;�H;�\E;�P@;��7;h*;�;�B�:�p�:���9 (����غioE� H���ɻ���������.��o@���K�      ��ͻLɻ�����d�����?�]�� ��潺���p8�9���:/T�:�;�Y;I-;v9;Z�@;�\E;��G;/5I;��I;C�I;ڵI;R�I;bpI;�UI;T@I;3/I;{!I;�I;@I;�I;�I;"�H;��H;�H;��H;�H;��H;!�H;�I;�I;AI;�I;z!I;6/I;O@I;�UI;hpI;S�I;ҵI;D�I;��I;25I;��G;�\E;\�@;o9;I-;�Y;�;-T�:���:h8�9����潺� �I�]�����d������Lɻ      ���,��ui�V�غb����*� ׭����9@��:H��:l��:�/;i�$;��1;g;;��A;��E;�H;25I;9�I;��I;L�I;��I;�vI;L[I;^EI;�3I;5%I;�I;�I;P	I;�I;}�H;a�H;'�H;��H;n�H;��H;"�H;^�H;|�H;�I;P	I;�I;�I;6%I;�3I;ZEI;R[I;�vI;��I;J�I;��I;8�I;35I;�H;��E;��A;g;;��1;e�$;�/;n��:B��:@��:���9�׭��*�T���p�غ�i�:��       *m8@��80_u9���9\�9:��:�W�:Jr�:@� ;�F;6o!;q�-;�^7;Pl>;�NC;�uF;PQH;�II;��I;��I;��I;��I;|zI;_I;<II;K7I;a(I;`I;�I;I;�I;, I;u�H;��H;�H;��H;t�H;��H; �H;��H;o�H;% I;�I;I;�I;aI;](I;G7I;@II;|_I;uzI;��I;��I;��I;��I;�II;NQH;�uF;�NC;Kl>;�^7;o�-;;o!;�F;;� ;<r�:�W�:��:��9:x��9�_u9 ��8      \o�:���:WK�:�Y�:F��:�;�;��;��$;�G.;P6;i�<;*�A;�E;SG;!�H;mI;��I;H�I;P�I;��I;�{I;vaI;�KI;�9I;�*I;�I;�I;�I;%I;� I;��H;��H;k�H;��H;�H;��H;�H;��H;h�H;��H;��H;� I;%I;�I;�I;�I;�*I;�9I;�KI;maI;�{I;��I;L�I;G�I;�I;mI;�H;SG;�E;+�A;j�<;P6;�G.;��$;��;�;�;x��:�Y�:CK�:v��:      p�;z�;];<X;�n!;�8';nI-;�93;��8;|=;lA;MzD;f�F;�/H;�I;ȔI;��I;k�I;ڵI;��I;|zI;saI;vLI;;I;^,I;0 I;I;�I;;I;�I;v�H;��H;g�H;o�H;
�H;S�H;!�H;N�H;�H;o�H;d�H;��H;w�H;�I;6I;�I;I;. I;b,I;;I;nLI;saI;|zI;��I;ٵI;d�I;��I;ĔI;�I;�/H;f�F;MzD;lA;|=;��8;�93;jI-;�8';�n!;<X;];\�;      R�1;��1;�73;�25;�7;��:;4|=;$Q@;R�B;HE;��F;ZH;��H; qI;ȶI;��I;��I;�I;R�I;�vI;|_I;�KI;;I;�,I;� I;I;�I;I;tI;��H;q�H;m�H;#�H;��H;p�H;��H;��H;��H;m�H;��H; �H;j�H;t�H;��H;nI;I;�I;I;� I;�,I;;I;�KI;{_I;�vI;N�I;�I;��I;��I;ƶI;qI;��H;ZH;��F;EE;V�B;(Q@;1|=;��:;��7;�25;�73;��1;      ��?;�@;�@;�A;��B;�C;&CE;}vF;��G;�\H;x�H;�mI;b�I;�I;�I;��I;��I;a�I;opI;W[I;GII;�9I;e,I;� I;oI;^I;�I;�I;g�H;��H;��H;-�H;V�H;��H;��H;]�H;1�H;W�H;��H;��H;R�H;&�H;��H;��H;d�H;�I;�I;^I;rI;� I;a,I;�9I;FII;R[I;lpI;\�I;��I;��I;�I; �I;b�I;�mI;x�H;�\H;��G;zvF;'CE;��C;��B;�A;�@;�@;      �uF;y�F;��F;\!G;@�G;
H;��H;�H;0KI;'�I;��I;��I;b�I;��I;��I;I�I;'}I;<hI;�UI;[EI;L7I;�*I;- I;I;\I;�I;GI;��H;��H;��H;&�H;>�H;��H;]�H;��H;�H;��H;�H;��H;]�H;��H;:�H;&�H;��H;��H;��H;@I;�I;^I;I;, I;�*I;I7I;WEI;�UI;8hI;$}I;I�I;��I;��I;b�I;��I;��I;$�I;0KI;�H;��H;�H;W�G;g!G;��F;x�F;      v I;*I;@I;M7I;�YI;�}I;�I;�I;�I;v�I;��I;}�I;��I;ܘI;�I;�pI;�^I;�NI;W@I;�3I;i(I;�I;"I;�I;�I;EI;��H;#�H;��H;1�H;"�H;i�H;�H;�H;��H;�H;��H;�H;|�H;�H;�H;e�H;"�H;/�H;��H;"�H;��H;GI;�I;�I; I;�I;g(I;�3I;S@I;�NI;�^I;�pI;�I;՘I;��I;|�I;��I;r�I;�I;	�I;�I;�}I;�YI;B7I;?I;I;      c�I;�I;��I;z�I;�I;�I;��I;��I;�I;}�I;�I;��I;݃I;sI;	cI;3TI;�FI;_:I;4/I;4%I;dI;�I;�I;I;�I;��H;#�H;��H;D�H;!�H;W�H;��H;��H;�H;Z�H;�H;��H;��H;X�H;�H;��H;��H;W�H;�H;?�H;��H;�H;��H;�I;I;�I;�I;aI;/%I;0/I;Y:I;�FI;4TI;cI; sI;݃I;��I;�I;}�I;�I;��I;��I;�I;'�I;{�I;��I;ڿI;      ��I;��I;F�I;S�I;O�I;p�I;v�I;��I;:�I;��I;L}I;�oI;TbI;�UI;�II;Q>I;�3I;=*I;�!I;�I;�I;�I;7I;pI;c�H;��H;��H;C�H;2�H;U�H;��H;��H;��H;��H;z�H;4�H;-�H;0�H;y�H;��H;��H;��H;��H;S�H;,�H;B�H;��H;��H;f�H;mI;9I;�I;�I;�I;~!I;7*I;�3I;Q>I;II;�UI;QbI;�oI;N}I;��I;=�I;��I;w�I;j�I;Y�I;U�I;K�I;��I;      ��I;��I;a�I;O�I;��I;׋I;��I;�zI;	qI;
gI;�\I;�RI;�HI;�>I;�5I;-I;�$I;vI;�I;�I;#I;"I;�I;��H;��H;��H;1�H;#�H;[�H;��H;��H;��H;��H;�H;��H;{�H;\�H;y�H;��H;�H;��H;��H;��H;��H;W�H;#�H;+�H;��H;��H;��H;�I;$I;I;�I;�I;qI;�$I;-I;�5I;�>I;�HI;�RI;�\I;
gI;qI;�zI;��I;׋I;��I;W�I;_�I;��I;      XvI;�uI;�sI;�pI;�lI;kgI;haI;�ZI;�SI;LI;aDI;�<I;5I;�-I;t&I;�I;eI;�I;FI;W	I;�I;� I;v�H;r�H;��H;$�H;#�H;^�H;��H;��H;��H;��H;��H;Z�H;�H;��H;��H;��H;	�H;]�H;��H;��H;��H;��H;��H;Z�H;�H;$�H;��H;q�H;z�H;� I;�I;S	I;FI;�I;bI;�I;r&I;�-I;5I;�<I;^DI;LI;�SI;�ZI;oaI;cgI;�lI;�pI;�sI;�uI;      �WI;-WI;�UI;�SI;ePI;�LI;"HI;CI;�=I;�7I;	2I;,I;(&I;e I;�I;}I;�I;�I;�I;�I;3 I;��H;��H;j�H;-�H;7�H;f�H;��H;��H;��H;��H;��H;D�H;��H;{�H;@�H;H�H;A�H;x�H;��H;G�H;��H;��H;��H;��H;��H;b�H;6�H;.�H;d�H;�H;��H;, I;�I;�I;�I;�I;~I;�I;e I;'&I;,I;2I;�7I;�=I;CI;&HI;�LI;oPI;�SI;�UI;0WI;      �AI;tAI;C@I;�>I;<I;9I;�5I;�1I;�-I;)I;p$I;�I;-I;�I;:I;�I;�	I;I;�I;��H;}�H;��H;d�H;�H;V�H;��H;�H;��H;��H;��H;��H;B�H;��H;\�H;�H;��H;��H;��H;	�H;_�H;��H;E�H;��H;��H;��H;��H;�H;��H;Y�H;�H;h�H;��H;w�H;�H;�I;I;�	I;�I;:I;�I;/I;�I;u$I;)I;�-I;�1I;�5I;9I;<I;~>I;P@I;tAI;      �1I;�1I;�0I;q/I;�-I;*+I;r(I;i%I;"I;wI;�I;I;DI;�I;�I;XI;I;I;%�H;e�H;��H;j�H;l�H;��H;��H;T�H;�H;�H; �H;�H;W�H;��H;]�H;��H;��H;��H;{�H;��H;��H;��H;_�H;��H;V�H;�H;��H;�H;�H;V�H;��H;��H;q�H;h�H;��H;^�H;#�H;I;I;ZI;�I;�I;BI;I;�I;xI;	"I;e%I;v(I;*+I;�-I;t/I;�0I;�1I;      �'I;�'I;�&I;�%I;$I;"I;�I;JI;pI;}I;QI;<I;�I;�
I;�I;�I;�I;0�H;��H;(�H;�H;��H;�H;b�H;��H;��H;z�H;^�H;~�H;��H;�H;{�H;�H;��H;~�H;Z�H;U�H;^�H;{�H;��H;�H;|�H;�H;��H;w�H;X�H;x�H;��H;��H;c�H;
�H;��H;�H;"�H;��H;3�H;�I;�I;�I;�
I;�I;<I;TI;�I;qI;JI;�I;"I;$I;�%I;�&I;�'I;      �!I;�!I;	!I; I;�I;�I;�I;�I;I;yI;�I;�I;�
I;I;QI;�I;��H;\�H;�H;��H;��H;�H;N�H;��H;T�H;�H;�H;�H;;�H;�H;��H;C�H;��H;��H;^�H;(�H;+�H;-�H;\�H;��H;��H;D�H;��H;x�H;5�H; �H;�H;�H;W�H;��H;R�H;�H;��H;��H;�H;b�H;��H;�I;TI;I;�
I;�I;�I;yI;I;�I;�I;�I;�I;" I;!I;�!I;      �I;�I;@I;+I;�I;!I;TI;(I;�I;(I;�I;�I;
I;9I;`I;�I;Y�H;��H;��H;s�H;��H;��H;�H;��H;-�H;��H;��H;��H;1�H;`�H;��H;J�H;��H;x�H;T�H;&�H;�H;*�H;Q�H;{�H;��H;K�H;��H;Y�H;,�H;��H;��H;��H;.�H;��H;"�H;��H;x�H;o�H;��H;��H;W�H;�I;aI;;I;	
I;�I;�I;)I;�I;(I;ZI;"I;�I;0I;=I;�I;      �!I;�!I;!I; I;�I;�I;�I;�I;I;xI;�I;�I;�
I;I;QI;�I;��H;\�H;�H;��H;��H;�H;N�H;��H;T�H;�H;�H;�H;<�H;}�H;��H;D�H;��H;��H;_�H;(�H;+�H;+�H;\�H;��H;��H;D�H;��H;v�H;5�H;��H;�H;�H;W�H;��H;R�H;�H;��H;��H;�H;b�H;��H;�I;SI;I;�
I;�I;�I;vI;I;�I;�I;�I;�I;& I;	!I;�!I;      �'I;�'I;�&I;�%I;$I;"I;�I;MI;pI;}I;SI;<I;�I;�
I;�I;�I;�I;2�H;��H;(�H;�H;��H;�H;`�H;��H;��H;x�H;\�H;~�H;��H;�H;z�H;�H;��H;~�H;[�H;U�H;^�H;}�H;��H;�H;{�H;�H;��H;w�H;W�H;x�H;��H;��H;b�H;
�H;��H;�H;"�H;��H;3�H;�I;�I;�I;�
I;�I;=I;TI;I;qI;NI;�I;"I;$I;�%I;�&I;�'I;      �1I;�1I;�0I;r/I;�-I;0+I;n(I;i%I;"I;uI;�I;I;AI;�I;�I;WI;I;I;%�H;d�H;��H;k�H;l�H;��H;��H;V�H;�H;�H; �H;�H;U�H;��H;]�H;��H;��H;��H;{�H;��H;��H;��H;]�H;��H;U�H;�H;��H;��H;�H;W�H;��H;��H;q�H;k�H;��H;`�H;&�H;I;I;[I;�I;�I;BI;I;�I;wI;	"I;f%I;y(I;-+I;�-I;v/I;�0I;�1I;      �AI;zAI;H@I;{>I;<I;9I;�5I;�1I;�-I;)I;r$I;�I;-I;�I;:I;�I;�	I;I;�I;��H;}�H;��H;c�H;�H;V�H;��H;�H;��H;��H;��H;��H;A�H;��H;[�H;�H;��H;��H;��H;	�H;\�H;��H;D�H;��H;��H;��H;��H;�H;��H;V�H;�H;j�H;��H;v�H;��H;�I;I;�	I;�I;:I;�I;0I;�I;s$I;)I;�-I;�1I;�5I;9I;<I;�>I;T@I;vAI;      �WI;/WI;�UI;�SI;ePI;�LI;%HI;CI;�=I;�7I;2I;,I;'&I;d I;�I;}I;�I;�I;�I;�I;4 I;��H;��H;g�H;.�H;6�H;c�H;��H;��H;��H;��H;��H;B�H;��H;|�H;@�H;H�H;A�H;x�H;��H;D�H;��H;��H;��H;��H;��H;a�H;7�H;+�H;a�H;�H;��H;, I;�I;�I;�I;�I;I;�I;g I;)&I;,I;2I;�7I;�=I;CI;'HI;�LI;gPI;�SI;�UI;,WI;      MvI;�uI;�sI;�pI;�lI;jgI;iaI;�ZI;�SI;LI;`DI;�<I;5I;�-I;u&I;�I;eI;�I;DI;S	I;�I;� I;w�H;r�H;��H; �H;�H;\�H;��H;��H;��H;��H;��H;Y�H;�H;��H;��H;��H;	�H;\�H;��H;��H;��H;��H;��H;X�H;�H;&�H;��H;n�H;{�H;� I;�I;T	I;GI;�I;eI;�I;u&I;�-I;5I;�<I;aDI;LI;�SI;�ZI;oaI;ggI;�lI;�pI;�sI;�uI;      ��I;��I;Y�I;V�I;��I;�I;��I;�zI;qI;gI;�\I;�RI;�HI;�>I;�5I;-I;�$I;tI;�I;�I;"I;%I;�I;��H;��H;��H;/�H;%�H;[�H;��H;��H;��H;��H;�H;��H;y�H;\�H;{�H;��H;�H;��H;��H;��H;��H;U�H;�H;-�H;��H;��H;��H;�I;%I;I;�I;�I;sI;�$I;-I;�5I;�>I;�HI;�RI;�\I;gI;qI;�zI;��I;ԋI;��I;`�I;c�I;��I;      ��I;��I;W�I;K�I;=�I;v�I;s�I;��I;B�I;�I;J}I;�oI;QbI;�UI;�II;Q>I;�3I;<*I;{!I;�I;�I;�I;6I;qI;f�H;��H;��H;C�H;0�H;Q�H;��H;��H;��H;��H;y�H;3�H;,�H;3�H;y�H;��H;��H;��H;��H;S�H;)�H;=�H;��H;��H;c�H;iI;:I;�I;�I;�I;�!I;9*I;�3I;T>I;�II;�UI;TbI;�oI;L}I;��I;>�I;��I;y�I;p�I;N�I;N�I;Y�I;��I;      p�I;ڿI;��I;y�I;�I;)�I;��I;��I;�I;}�I;ߦI;��I;܃I;sI;
cI;4TI;�FI;]:I;2/I;1%I;bI;�I;�I;I;�I;��H;�H;��H;D�H;�H;U�H;��H;��H;��H;[�H;��H;��H;��H;X�H;�H;��H;��H;W�H;�H;?�H;��H;�H;��H;�I;I;�I;�I;aI;2%I;4/I;\:I;�FI;5TI;	cI;sI;݃I;��I;�I;�I;�I;��I;��I;�I;$�I;{�I;��I;ڿI;      d I;3I;?I;T7I;�YI;�}I;�I;�I;�I;u�I;��I;~�I;��I;٘I;�I;�pI;�^I;�NI;S@I;�3I;h(I;�I;I;�I;�I;@I;��H;#�H;��H;.�H;!�H;h�H;�H;�H;�H;�H;��H;�H;|�H;�H;�H;f�H;"�H;.�H;��H;�H;��H;II;�I;�I;"I;�I;g(I;�3I;V@I;�NI;�^I;�pI;�I;טI;��I;y�I;��I;r�I;�I;�I;�I;�}I;�YI;W7I;@I;I;      �uF;y�F;��F;U!G;F�G;H;��H; �H;5KI;"�I;��I;��I;`�I;��I;��I;K�I;$}I;>hI;�UI;XEI;N7I;�*I;* I;I;\I;�I;DI;��H;��H;��H;$�H;=�H;��H;[�H;��H;�H;��H;�H;��H;[�H;��H;;�H;&�H;��H;��H;��H;DI;�I;\I;I;- I;�*I;L7I;[EI;�UI;:hI;(}I;K�I;��I;��I;`�I;��I;��I;%�I;+KI;�H;��H;�H;Q�G;[!G;��F;k�F;      ��?;�@;�@;�A;��B;�C;$CE;|vF;��G;�\H;x�H;�mI;_�I;�I; �I;��I;��I;`�I;npI;S[I;FII;�9I;a,I;� I;qI;VI;�I;�I;g�H;��H;��H;*�H;S�H;��H;��H;Z�H;1�H;Z�H;��H;��H;V�H;+�H;��H;��H;c�H;�I;�I;`I;oI;� I;e,I;�9I;GII;V[I;rpI;_�I;��I;��I; �I;�I;b�I;�mI;t�H;�\H;��G;zvF;&CE;��C;��B;�A;�@;�@;      3�1;��1;�73;�25;z�7;��:;.|=;!Q@;Y�B;BE;��F;ZH;��H;qI;ɶI;��I;��I;�I;O�I;�vI;}_I;�KI;;I;�,I;� I;I;�I;I;rI;��H;q�H;m�H; �H;��H;k�H;��H;��H;��H;m�H;��H;$�H;n�H;u�H;��H;qI;I;�I;I;� I;�,I;;I;�KI;_I;�vI;S�I;�I;��I;��I;ƶI;qI;��H;YH;��F;DE;U�B;Q@;1|=;��:;��7;�25;�73;��1;      g�;z�;];@X;�n!;�8';dI-;�93;��8;|=;
lA;LzD;d�F;�/H;�I;ǔI;��I;k�I;ٵI;��I;|zI;saI;pLI;;I;a,I;& I;I;�I;;I;�I;v�H;��H;d�H;l�H;�H;S�H;#�H;S�H;�H;l�H;e�H;��H;{�H;�I;7I;�I; I;. I;`,I;;I;sLI;taI;zI;��I;ݵI;g�I;��I;ǔI;�I;�/H;f�F;IzD;lA;|=;��8;�93;dI-;�8';�n!;FX; ];d�;      `o�:���:IK�:�Y�:F��:�;�;��;��$;�G.;P6;m�<;(�A;�E;SG; �H;mI;��I;E�I;O�I;��I;�{I;paI;�KI;�9I;�*I;�I;�I;�I;"I;� I;��H;��H;j�H;��H;�H;��H;�H;��H;h�H;��H;��H;� I;(I;�I;�I;�I;�*I;�9I;�KI;saI;�{I;��I;P�I;H�I;�I;mI; �H;
SG;�E;*�A;i�<;P6;�G.;��$;��;�;�;p��:�Y�:CK�:~��:       &m8���80`u9���9H�9:��:�W�:@r�:A� ;�F;9o!;q�-;�^7;Ll>;�NC;�uF;MQH;�II;��I;��I;��I;��I;xzI;}_I;?II;D7I;](I;`I;�I;I;�I;) I;r�H;��H; �H;��H;t�H;��H; �H;��H;s�H;) I;�I;I;�I;`I;`(I;I7I;=II;�_I;zzI;��I;��I;��I;��I;�II;NQH;�uF;�NC;Ol>;�^7;n�-;;o!;�F;=� ;Dr�:�W�:��:��9:���9�`u9���8      {��%��yi�V�غh����*��׭���9J��:>��:n��:�/;h�$;��1;g;;��A;��E;�H;05I;8�I;��I;M�I;��I;�vI;P[I;WEI;�3I;2%I;�I;�I;P	I;�I;|�H;a�H;%�H;��H;l�H;��H;"�H;]�H;|�H;�I;T	I;�I;�I;4%I;�3I;[EI;N[I;�vI;��I;M�I;��I;9�I;35I;�H;��E;��A;g;;��1;g�$;�/;n��:<��:F��:���9�׭� �*�\���l�غzi�)��      ��ͻLɻ�����d�����B�]�� ��潺���h8�9���:-T�:�;�Y;I-;s9;Y�@;�\E;��G;05I;��I;D�I;ٵI;Q�I;hpI;�UI;O@I;3/I;}!I;�I;@I;�I;�I;�H;��H;�H;��H;�H;��H;�H;�I;�I;DI;�I;{!I;3/I;Q@I;�UI;dpI;V�I;ٵI;G�I;��I;25I;��G;�\E;Z�@;p9;I-;�Y;�;-T�:���:X8�9����潺� �C�]�����d������Hɻ      �iO�ߔK��o@���.���������ɻ�G��joE���غ(�����9�p�:�B�:�;l*;��7;�P@;�\E;�H;�II;�I;h�I;�I;Z�I;8hI;�NI;b:I;<*I;vI;�I;�I;I;I;/�H;^�H;��H;_�H;-�H;I;I;�I;�I;xI;:*I;b:I;�NI;:hI;V�I;�I;g�I;��I;�II;�H;�\E;�P@;��7;l*;�;�B�:�p�:���9(����غjoE��G���ɻ���������.��o@�ߔK�      L�����2���?����N��Pp��D����hG�����34�>��� �n8��:A�:GG;�(;��7;X�@;��E;NQH;mI;��I;��I;��I; }I;�^I;�FI;�3I;�$I;^I;�I;�	I;I;�I;��H;P�H;��H;�I;I;�	I;�I;aI;�$I;�3I;�FI;�^I; }I;��I;��I;��I;mI;JQH;��E;Y�@;��7;�(;GG;A�:��: �n8D���24�����hG໇���D�Pp��N��@���3������      
��'�T5���������ϼ̡��X���iO�>���ɻ��p��D���o��g:�_�:@G;l*;o9;��A;�uF;�H;ĔI;��I;��I;D�I;�pI;3TI;R>I;-I;�I;{I;�I;ZI;�I;�I;�I;�I;�I;TI;�I;xI;�I;-I;Q>I;4TI;�pI;B�I;��I;��I;ǔI; �H;�uF;��A;o9;j*;CG;�_�:�g:��o��D⺙�p��ɻ>���iO�X��͡����ϼ������T5�&�      j��ѷ��%0v�r�a�$�G�@2+���ן�	����/����5��&��^f��ج��g:9�:�;I-;g;;�NC;SG;�I;ȶI;�I;��I;�I;
cI;�II;�5I;q&I;�I;6I;�I;�I;MI;XI;NI;�I;�I;6I;�I;q&I;�5I;�II;
cI;�I;��I;�I;̶I;�I;SG;�NC;g;;I-;�;;�:��g:�ج�_f�(�����5��/�����ן���@2+�$�G�s�a�%0v�ѷ��      ��ս��ѽ;�ƽ1����I�����Q�a�D4�<M���ϼ��K�K�N��MG��]f���o���:�B�:�Y;��1;Rl>;�E;�/H;qI;��I;��I;֘I; sI;�UI;�>I;�-I;a I;�I;�I;�
I;I;/I;I;�
I;�I;�I;^ I;�-I;�>I;�UI; sI;טI;��I;��I;"qI;�/H;�E;Il>;��1;�Y;�B�:��:��o�bf�LG��N��K�K�����ϼ<M�D4�R�a�����I��1���;�ƽ��ѽ      �L+�  (���F�������ս�@���%���;V�%��ސ������MS�M��&��xD���n8�p�:�;g�$;�^7;*�A;h�F;��H;b�I;_�I;��I;߃I;XbI;�HI;5I;%&I;-I;AI;�I;�
I;
I;�
I;�I;>I;/I;"&I;5I;�HI;YbI;��I;��I;\�I;^�I;��H;k�F;-�A;�^7;i�$;�;�p�: �n8|D�&��M���MS�����ސ�%���;V��%���@����ս����F���  (�      �T��f�����z��Yb�&�D��$�����ѽ�I��D�m�2+�������K�K�ﻘ�p�L������9'T�:�/;u�-;d�<;FzD;ZH;�mI;��I;v�I;��I;�oI;�RI;�<I;,I;�I;I;/I;�I;�I;�I;/I;I;�I; ,I;�<I;�RI;�oI;��I;w�I;��I;�mI;ZH;KzD;f�<;k�-;�/;#T�:���9H�����p��L�K�������2+�D�m��I����ѽ���$�'�D��Yb���z�f���      ?�׾��Ҿž�j��������z�S�H�)��ez�G$���/v�2+�ސ�����5��ɻ:4�`(�����:^��:<o!;P6;lA;��F;q�H;��I;��I;ߦI;J}I;�\I;^DI;2I;p$I;�I;HI;�I;�I;�I;HI;�I;r$I;2I;]DI;�\I;M}I;ߦI;��I;��I;p�H;��F;lA;P6;1o!;`��:~��:P(��94��ɻ��5���ސ�2+��/v�G$��ez�)��S�H���z������j��ž��Ҿ      H(��$�d��P������~���`���Yb���'��U�G$��D�m�&����ϼ�/��>��������غ88�9<��:�F;�G.;|=;GE;�\H;�I;q�I;v�I;��I;gI;LI;�7I;	)I;pI;rI;rI;'I;qI;rI;pI;)I;�7I;LI;gI;��I;z�I;s�I;�I;�\H;HE;|=;�G.;�F;>��:88�9��غ����>���/����ϼ&��D�m�G$���U���'��Yb��`���~�����P��d���$�      <�}���w�#f���K�r,�}�
�;�׾ �����k���'�ez꽝I���;V�<M�	����iO�mG�toE����<��:D� ;��$;��8;X�B;��G;+KI;�I;�I;B�I;qI;�SI;�=I;�-I;"I;kI;I;�I;I;kI;"I;�-I;�=I;�SI;qI;B�I;�I;�I;,KI;��G;_�B;��8;��$;;� ;@��:ȱ�soE�lG໫iO�	���<M��;V��I��ez���'���k� ���;�׾}�
�r,���K�#f���w�      ��p�������.蒿��w��F�d��ʰ� ����Yb�)����ѽ�%��D4�؟�X�����H���潺���9Hr�:��;�93;%Q@;|vF;�H;�I;��I;��I;�zI;�ZI;CI;�1I;c%I;?I;�I;"I;�I;BI;b%I;�1I;CI;�ZI;�zI;��I;��I;�I;�H;|vF;'Q@;�93;��;6r�:В�9�潺H�����X��؟�D4��%����ѽ)���Yb� ���ʰ�d���F���w�.蒿����p���      4��������㿊�ɿ���ʅ����P�d��;�׾�`��S�H����@��R�a���͡���D��ɻ� �@ح��W�:�;`I-;5|=;CE;��H;�I;��I;u�I;��I;haI; HI;�5I;r(I;�I;�I;SI;�I;�I;p(I;�5I;"HI;haI;��I;v�I;��I;�I;��H;CE;8|=;fI-;�;�W�:�׭�� ��ɻ�D�͡����R�a��@����S�H��`��;�׾d����P�ʅ�������ɿ�㿳���      ř$��x �"��:���޿o���ʅ���F�}�
��~����z��$���ս���A2+���ϼPp�����P�]��*���:�;�8';��:;��C;�H;�}I;�I;q�I;ًI;mgI;�LI;9I;9+I;!"I;�I;*I;�I;""I;7+I;9I;�LI;jgI;ًI;s�I;"�I;�}I;H;��C;��:;�8';�;��:�*�Q�]�����Pp���ϼA2+������ս�$���z��~��}�
��F�ʅ��o����޿:��"���x �      J�Q���K���;�ř$��;
��޿�����w�r,���澝���'�D������I��$�G�����N��������V�����9:V��:�n!;��7;��B;F�G;�YI;(�I;W�I;��I;�lI;sPI;<I;�-I;
$I;�I;�I;�I;$I;�-I;<I;sPI;�lI;��I;Z�I;.�I;�YI;Q�G;��B;��7;�n!;V��:x�9:T����������N�����$�G��I������'�D��������r,���w�����޿�;
�ř$���;���K�      T����{���d��F�ř$�:����ɿ.蒿��K�P���j���Yb�F�1���s�a����?�����.��d��p�غȰ�9�Y�:,X;�25; �A;U!G;E7I;p�I;@�I;O�I;�pI;�SI;~>I;y/I;�%I;" I;0I; I;�%I;v/I;�>I;�SI;�pI;T�I;B�I;v�I;I7I;c!G;�A;�25;.X;�Y�:���9f�غ�d����.�?������s�a�1���F��Yb��j��P����K�.蒿��ɿ:��ř$��F���d��{�      ����#P�������d���;�#���㿲���#f�d��ž��z���<�ƽ%0v�T5�2����o@�����|i��`u9;K�:];�73;"�@;��F;CI;��I;M�I;S�I;�sI;�UI;?@I;�0I;�&I;!I;0I;!I;�&I;�0I;A@I;�UI;�sI;X�I;M�I;��I;II;��F;�@;�73;];;K�:p`u9yi������o@�2���T5�%0v�<�ƽ����z�žd��#f�������#����;���d����#P��      �,��a��#P���{���K��x �����p�����w��$���Ҿf���  (���ѽҷ��'�����K�Fɻ)�����8x��:x�;��1;�@;i�F;I;ۿI;�I;��I;�uI;%WI;fAI;�1I;�'I;�!I;�I;�!I;�'I;�1I;hAI;&WI;�uI;��I;�I;޿I;!I;x�F;�@;��1;v�;r��:���8'��Hɻ�K����'�ҷ����ѽ  (�f�����Ҿ�$���w�p��������x ���K��{�#P��a��      D(��q'���o��N�d��X1�~x�	Ŀ����3�w���x����4�k��Y+���'���ü:yY��kٻp&���p�H��:8;��0;��?;��F;g I;��I;��I;)�I;g�I;LdI;�KI;�9I;m.I;�'I;�%I;�'I;k.I;�9I;�KI;MdI;d�I;.�I;��I;��I;g I;̀F;��?;��0;4;<��:��p�p&��kٻ:yY���ü�'�Y+��k�ཽ�4��x��w���3����	Ŀ~x��X1�d�N��o��q'��      q'���X��f^�������]]���,�P9�6g��T�����/����o��g1��hܽ���-$�_l���|U�f�Ի�!� �,�u�:�;�51;��?;4�F;?'I;_�I;
�I;=�I;��I;�cI;>KI;x9I;.I;{'I;�%I;v'I; .I;w9I;@KI;�cI;��I;?�I;
�I;b�I;?'I;?�F;��?;51;�;m�: �,��!�f�Ի�|U�_l���-$����hܽg1��o���ྚ�/�T���6g��P9���,��]]�����f^���X��      �o��f^���ē��4z�5K�h��R��&ﱿT�v��X#���Ѿń��&�p�нc̀�_��v���L�I��ǻ�4��"9��:4�; �2;��@;��F;�:I;��I;��I;��I;u�I;KbI;�II;�8I;Z-I;�&I;�$I;�&I;[-I;�8I;�II;KbI;o�I;��I;��I;��I;�:I;��F;��@;�2;2�;��:"9�4��ǻM�I�v���_��c̀�p�н�&�ń���Ѿ�X#�T�v�&ﱿR��h��5K��4z��ē�f^��      N������4z���V��X1��<�tؿ����RZ��	�(���IUo����^y��.l�Y��R��B�7�������ų9��:��;X�4;jtA;\2G;�XI;��I;J�I;�I;�I;�_I;�GI;"7I;�+I;�%I;�#I;�%I;�+I;!7I;�GI;�_I;��I;�I;J�I;��I;�XI;f2G;gtA;W�4;��;���:�ų9�����B�7��R��Y�.l�^y�����IUo�(����	��RZ����tؿ�<��X1���V��4z�����      d��]]�5K��X1�Zf��nQ��S���[58��A���נ���O���_什�Q����@ߓ��� ��V���氺��":Ը�: ;�07;�B;0�G;�{I;��I;��I;��I;:|I;7\I;LEI;5I;3*I;1$I;)"I;-$I;5*I;5I;JEI;5\I;4|I;��I;��I;��I;�{I;7�G;�B;�07; ;и�:��":�氺�V���� �@ߓ�����Q�_什����O��נ��A��[58�S���nQ���Zf��X1�5K��]]�      �X1���,�h���<��5g��e_���U�͂�֌Ⱦń�*�-�i��P ��&�2�?ټb�{�"��n�(�O���u:�P ;�&;+#:;=�C;�%H;�I;!�I;��I;�I;]vI;�WI;�AI;z2I;(I;D"I;^ I;@"I;(I;w2I;�AI;�WI;YvI;�I;��I;$�I;�I;�%H;=�C;&#:;�&;�P ;��u: �O��n�"�b�{�?ټ&�2�P ��i��*�-�ń�֌Ⱦ͂��U�e_��5g��<�h����,�      ~x�P9�R��sؿnQ��e_��6�_��X#�p���f��9�S�{�����l�B�	w�� �M���Ի��+�0=T���:�e;�\,;�/=;�BE;Q�H;z�I;��I;��I;��I;�oI;�RI;>I;]/I;}%I;�I;FI;�I;~%I;\/I;>I;�RI;�oI;��I;��I;��I;v�I;W�H;�BE;�/=;�\,;�e;��: =T���+���Ի�M�	w��B�l�����{�9�S��f��p���X#�6�_�e_��nQ��sؿR��P9�      	Ŀ6g��&ﱿ���S����U��X#�t��d���IUo��#��hܽ����n<����<����� ��᝻F�Ժxt�9`��:�V;̇2;� @;T�F;�I;��I;C�I;)�I;i�I; hI;MI;�9I;�+I;�"I;jI;�I;iI;�"I;�+I;�9I;MI;�gI;l�I;)�I;D�I;��I;�I;W�F;� @;͇2;�V;T��:�t�9J�Ժ�᝻�� �;�������n<�����hܽ�#�IUo�d���t���X#��U�S������&ﱿ6g��      ���T���T�v��RZ�[58�͂�p��d���foy�]1�_O��[什�`�M�����pyY�$�컘�T��1�x�u:���:F#;98;	�B;f�G;�lI;�I;�I;-�I;v�I;�_I;GI;�4I;%(I;�I;�I;I;�I;�I;#(I;�4I;GI;�_I;w�I;-�I;�I;�I;�lI;j�G;�B;98;H#;���:��u:�1���T�$��pyY����M���`�[什_O��]1�foy�d���p��͂�[58��RZ�T�v�T���      �3���/��X#��	��A��֌Ⱦ�f��HUo�]1�˰��|n��Ѽx��'��>ټ�@���k�м��"����39�#�:.R;	e-;�/=;�	E;\xH;��I;�I;p�I;��I;vI;aWI;�@I;�/I;#$I;;I;�I;6I;�I;<I;"$I;�/I;�@I;cWI;vI;�I;s�I;
�I;|�I;_xH;�	E;�/=;e-;*R;�#�:��39"��μ���k��@���>ټ�'�Ѽx�|n��˰��]1�HUo��f��֌Ⱦ�A���	��X#���/�      v���ྃ�Ѿ(����נ�ń�9�S��#�_O��|n��J̀���2���𛼃�>� �Ի��B��#�4m:�G�:^ ;��5;�FA;��F;�I;N�I;Q�I;��I;j�I;njI;�NI;:I;�*I;�I;�I;�I;KI;�I;�I;�I;�*I;:I;�NI;pjI;m�I;��I;P�I;I�I;�I;��F;�FA;��5;[ ;�G�:8m:�#���B� �Ի��>�������2�J̀�|n��_O���#�9�S�ń��נ�(�����Ѿ��      �x���o��ń�IUo���O�*�-�{��hܽ\什Ѽx���2�tb��UR��W|U�Z2��:��$갺�u�9��:D;��,;�h<;crD;N%H;��I;g�I;��I;�I;�I;�^I;FI;V3I;�%I;�I;^I;hI;4I;hI;^I;�I;�%I;R3I;	FI;�^I;
�I;�I;��I;b�I;ďI;M%H;drD;�h<;��,;D;��:�u�9갺:��Z2��V|U�UR��tb����2�Ҽx�[什�hܽ{�*�-���O�IUo�ń��o��      ��4�f1��&������i�ང�������`��'���UR��E�]���"V���X�� Io����:h�;$#;�6;QtA;R�F;�	I;r�I;��I;p�I;�I;�pI;�SI;�=I;�,I;w I;�I;�I;GI;9I;FI;�I;�I;y I;�,I;�=I;�SI;�pI;�I;m�I;��I;v�I;�	I;Q�F;StA;�6;.#;l�;���:�Go��X��"V��~��D�]�TR����'��`��������h��������&�f1�      j�ྲྀhܽo�н]y��^什P ��l��n<�M���>ټ��V|U���������1�������u:Wl�:�;b71;S)>;S	E;
JH;T�I;��I;��I;�I;׃I;YbI;�HI;&5I;c&I;gI;qI;<I;%I;
I;%I;:I;rI;eI;`&I;*5I;�HI;_bI;݃I;�I;��I;��I;Q�I;
JH;W	E;P)>;k71;�;Ol�:��u:�����1��������V|U����>ټM���n<�l�P ��_什^y��o�н�hܽ      Y+����c̀�-l��Q�&�2�B��������@����>�Y2��#V���1�����#R:���:�;t\,;1;;�;C;�eG;U9I;��I;/�I;��I;C�I;�qI;�TI;b>I;8-I;3 I;zI;rI;�
I;I;I;I;�
I;tI;{I;- I;9-I;c>I;�TI;�qI;@�I;��I;1�I;��I;T9I;�eG;�;C;:;;w\,;�;���:�#R:���1�"V��X2����>��@��������B�%�2��Q�-l�c̀���      �'��-$�_��X����?ټw��;���pyY��k���Ի:��Y�������#R:���:�R;�);܍8;��A;��F;3�H;)�I;��I;��I;��I;�I;�`I;�GI;�4I;�%I;JI;�I;�I;qI;I;FI;I;mI;�I;�I;FI;�%I;�4I;�GI;�`I;�I;��I;��I;��I;'�I;6�H;��F;��A;ݍ8;�);�R;���:�#R:����
Y��:����Ի�k�oyY�;���	w��	?ټ���Y�^���-$�      ��ü^l��w����R��?ߓ�a�{��M��� � ��ʼ����B�갺@Ho���u:���:�R;/�';17;��@;��E;�lH;.�I;h�I;��I;�I;x�I;�lI;�QI;&<I;�+I;�I;�I;eI;�I;CI;0I;�I;,I;AI;�I;eI;�I;�I;�+I;'<I;�QI;�lI;p�I;	�I;��I;e�I;/�I;�lH;��E;��@;17;0�';�R;���:��u:�Ho�갺��B�˼�� �컌� ��M�a�{�@ߓ��R��x���\l��      3yY��|U�L�I�?�7��� �"���Ի�᝻��T���#��u�9���:Ql�:�;�);17;/ @;:]E;�$H;dkI;
�I;U�I;��I;'�I;�wI;�ZI;�CI;w1I;N#I;%I;�I;-	I;rI;9I;m�H;��H;j�H;6I;oI;+	I;�I;)I;P#I;w1I;�CI;�ZI;�wI;+�I;��I;O�I;�I;ekI;�$H;;]E;+ @;17;�);�;Ol�:���:�u�9�#����T��᝻��Ի"��� �A�7�K�I��|U�      �kٻl�Ի�ǻ����V���n���+�6�Ժ��1�0�39Tm:��:l�;�;z\,;��8;��@;A]E;�
H;LVI;q�I;��I;��I;c�I;��I;�bI;bJI;%7I;�'I;�I;.I;�
I;8I;;I;i�H;��H;y�H;��H;f�H;8I;6I;�
I;0I;�I;�'I;(7I;]JI;�bI; �I;e�I;��I;��I;t�I;MVI;�
H;:]E;��@;ڍ8;y\,;	�;j�;��:`m: �39�1�8�Ժ��+��n��V������ǻl�Ի      p&��!��4����氺�O��<T�ht�9��u:�#�:�G�:D;*#;i71;;;;��A;��E;�$H;MVI;�I;��I;�I;��I;��I;iI;'PI;<I;�+I;I;�I;�I;�I;�I;5�H;��H;��H;�H;��H;��H;0�H;�I;�I;�I;�I;I;�+I;<I;#PI;iI;��I;}�I;�I;��I;�I;MVI;�$H;��E;��A;:;;d71;&#;D;�G�:�#�:��u:�t�9�<T��O��氺���4��!�      @�p� �,�!9�ų9Ќ":��u:��:`��:���:.R;\ ;��,;�6;S)>;�;C;��F;�lH;lkI;t�I;��I;��I;�I;r�I;�mI;wTI;%@I;�/I;""I;WI;�I;�I;�I;u�H;u�H;��H;V�H;��H;O�H;��H;r�H;r�H;�I;�I;�I;UI;$"I;�/I;"@I;|TI;�mI;k�I;�I;��I;��I;t�I;fkI;�lH;��F;�;C;N)>;�6;��,;` ;.R;���:Z��:��:|�u:�":�ų9p!9 �,�      :��:��:�:��:¸�:�P ;�e;�V;J#;e-;��5;�h<;RtA;X	E;�eG;8�H;2�I;�I;��I;�I;�I;�I;pI;LWI;�BI;@2I;�$I;sI;oI;B	I;tI;��H;��H;�H;Y�H;3�H;��H;.�H;V�H;�H;��H;��H;vI;B	I;lI;tI;�$I;?2I;�BI;HWI;�oI;�I;�I;�I;��I;�I;1�I;6�H;�eG;S	E;QtA;�h<;��5;e-;L#;�V;�e;�P ;��:���:��:y�:      J;�;0�;��;� ;�&;�\,;ۇ2;98;�/=;�FA;orD;U�F;JH;[9I;.�I;n�I;Z�I;��I;��I;p�I;pI;IXI;�DI;�3I;]&I;I;�I;�
I;oI;��H;��H;��H;��H;9�H;H�H;�H;B�H;6�H;��H;��H;��H;��H;lI;{
I;�I;I;\&I;�3I;�DI;BXI;pI;p�I;��I;��I;R�I;k�I;,�I;X9I;JH;R�F;lrD;�FA;�/=;98;ׇ2;�\,;�&; ;��;*�;�;      ��0;�51;�2;T�4;�07;0#:;�/=;� @;�B;�	E;��F;P%H;�	I;U�I;��I;��I;��I;��I;c�I;��I;�mI;DWI;�DI;�4I;='I;-I;�I;{I;;I;. I;,�H;��H;z�H;��H;c�H;��H;i�H;��H;`�H;��H;z�H;��H;.�H;, I;5I;|I;�I;.I;@'I;�4I;~DI;EWI;�mI;��I;`�I;��I;��I;��I;��I;P�I;�	I;N%H;��F;�	E;�B;� @;�/=;#:;�07;P�4;�2;�51;      ��?;��?;��@;atA;��B;I�C;�BE;W�F;j�G;`xH;�I;ˏI;u�I;��I;7�I;��I;�I;1�I;�I;iI;�TI;�BI;�3I;G'I;�I;|I;I;�I;� I;~�H;�H;k�H;a�H;��H;��H;-�H;��H;'�H;��H;��H;^�H;f�H;�H;}�H;� I;�I;I;}I;�I;A'I;�3I;�BI;�TI;iI;�I;+�I;�I;��I;3�I;��I;u�I;ʏI;�I;`xH;h�G;T�F;�BE;:�C;�B;`tA;��@;��?;      ��F;C�F;��F;_2G;'�G;&H;Y�H;�I;�lI;��I;T�I;p�I;��I;��I;��I;��I;x�I;�wI;�bI;&PI;'@I;:2I;\&I;0I;yI;:I;I; I;��H;F�H;x�H;V�H;|�H;'�H;[�H;��H;��H;��H;X�H;&�H;{�H;P�H;w�H;C�H;��H;� I;I;:I;I;-I;X&I;=2I;%@I;"PI;�bI;�wI;x�I;��I;��I;��I;��I;m�I;X�I;��I;�lI;�I;Z�H;�%H;<�G;m2G;��F;C�F;      v I;K'I;�:I;�XI;�{I;�I;}�I;�I;�I;�I;U�I;��I;m�I;�I;@�I;�I;�lI;�ZI;cJI; <I;�/I;�$I;"I;I;I;I;I;��H;v�H;��H;L�H;T�H;��H;��H;�H;��H;n�H;��H;�H;��H;��H;O�H;M�H;��H;p�H;��H;I;I;I;�I;I;�$I;�/I;<I;`JI;�ZI;�lI;�I;=�I;�I;j�I;��I;U�I;�I;�I;��I;v�I;�I;�{I;�XI;�:I;5'I;      ��I;g�I;��I;��I;��I;"�I;��I;C�I;�I;v�I;��I;�I;�I;ۃI;�qI;�`I;�QI;�CI;%7I;�+I;'"I;oI;�I;}I;�I;� I;��H;l�H;��H;V�H;T�H;��H;��H;��H;��H;��H;o�H;��H;��H;��H;��H;��H;T�H;T�H;��H;j�H;��H;� I;�I;yI;�I;oI;""I;�+I;!7I;�CI;~QI;�`I;�qI;ڃI;�I;�I;��I;t�I;��I;@�I;��I;�I;��I;��I;��I;]�I;      ��I;�I;��I;[�I;��I;��I;��I;-�I;'�I;�I;n�I;
�I;�pI;_bI;�TI;�GI;*<I;{1I;�'I;I;^I;iI;~
I;6I;� I;��H;m�H;��H;P�H;O�H;��H;P�H;@�H;��H;��H;��H;��H;��H;��H;��H;A�H;L�H;��H;M�H;L�H;��H;i�H;��H;� I;1I;{
I;gI;WI;I;�'I;v1I;'<I;�GI;�TI;\bI;�pI;
�I;q�I;�I;(�I;,�I;��I;��I;��I;\�I;��I;��I;      /�I;<�I;��I;
�I;��I;�I;��I;r�I;w�I;vI;rjI;�^I;�SI;�HI;b>I;�4I;�+I;N#I;�I;�I;�I;?	I;lI;, I;��H;?�H;��H;X�H;U�H;��H;*�H;�H;8�H;��H;�H;��H;��H;��H;�H;��H;6�H;�H;*�H;��H;O�H;X�H;��H;@�H;��H;) I;oI;@	I;�I;�I;�I;I#I;�+I;�4I;`>I;�HI;�SI;�^I;rjI;vI;v�I;k�I;��I;�I;��I;�I;��I;9�I;      d�I;��I;w�I;��I;4|I;]vI;�oI;hI;�_I;gWI;�NI;FI;�=I;+5I;=-I;�%I;�I;)I;2I;�I;�I;vI;��H;-�H;�H;w�H;M�H;Y�H;��H;-�H;	�H;�H;T�H;��H;u�H;-�H;��H;,�H;t�H;��H;W�H;�H;�H;*�H;��H;V�H;J�H;w�H;�H;,�H;��H;vI;�I;�I;2I;&I;�I;�%I;<-I;*5I;�=I;FI;�NI;jWI;�_I;hI;�oI;VvI;<|I;��I;v�I;��I;      JdI;�cI;DbI;�_I;)\I;�WI;�RI;MI;GI;�@I;:I;Z3I;�,I;f&I;3 I;JI;�I;�I;�
I;�I;�I;��H;��H;��H;k�H;O�H;Q�H;��H;U�H;�H;�H;M�H;��H;%�H;��H;��H;��H;��H;��H;&�H;��H;M�H;�H;�H;O�H;��H;O�H;O�H;n�H;��H;��H;��H;�I;�I;�
I;�I;�I;MI;3 I;g&I;�,I;Y3I;:I;�@I;GI;MI;�RI;�WI;1\I;�_I;NbI;�cI;      �KI;LKI;�II;�GI;IEI;�AI;>I;�9I;�4I;�/I;�*I;�%I;w I;jI;{I;�I;iI;.	I;=I;�I;~�H;��H;��H;u�H;a�H;w�H;��H;��H;H�H;;�H;Q�H;��H;�H;��H;J�H;�H;.�H;�H;F�H;��H;�H;��H;P�H;4�H;C�H;��H;��H;u�H;d�H;u�H;��H;��H;x�H;�I;<I;-	I;iI;�I;|I;hI;y I;�%I;�*I;�/I;�4I;�9I;>I;�AI;LEI;�GI;JI;LKI;      �9I;x9I;�8I;7I;5I;k2I;Z/I;�+I;%(I;*$I; I;�I;�I;uI;xI;�I;�I;pI;?I;7�H;|�H;�H;��H;��H;��H;�H;��H;��H;��H;��H;��H;%�H;��H;5�H;��H;��H;��H;��H;��H;6�H;��H;%�H;��H;��H;�H;��H;��H;�H;��H;��H;��H;�H;u�H;/�H;=I;sI;�I;�I;yI;xI;�I;�I; I;-$I;'(I;�+I;c/I;k2I;5I;7I;�8I;�9I;      ].I;9.I;_-I;�+I;?*I;
(I;%I;�"I;�I;HI;�I;lI;�I;CI;�
I;rI;II;8I;k�H;��H;��H;U�H;5�H;U�H;��H;P�H;�H;��H;��H;�H;o�H;��H;J�H;��H;��H;��H;z�H;��H;��H;��H;J�H;��H;m�H;�H;��H;��H;�H;P�H;��H;V�H;8�H;U�H;��H;��H;j�H;9I;II;tI;�
I;FI;�I;jI;�I;JI;�I;�"I;�%I;(I;9*I;,I;\-I;:.I;      �'I;�'I;�&I;�%I;#$I;="I;�I;pI;�I;�I;�I;pI;HI;&I;I;I;0I;h�H;��H;��H;^�H;.�H;B�H;��H;&�H;��H;��H;��H;��H;��H;,�H;��H;�H;��H;��H;a�H;o�H;c�H;��H;��H;�H;��H;)�H;��H;��H;��H;��H;��H;'�H;��H;F�H;/�H;W�H;��H;��H;m�H;3I;I;I;*I;HI;mI;�I;�I;�I;mI;  I;="I;&$I;�%I;�&I;�'I;      �%I;�%I;�$I;�#I;!"I;W I;GI;�I;I;7I;SI;<I;?I;$
I;I;HI;�I;��H;}�H;	�H;��H;��H;�H;[�H;��H;��H;i�H;s�H;��H;��H;��H;��H;/�H;��H;z�H;j�H;s�H;l�H;w�H;��H;0�H;��H;��H;��H;~�H;p�H;j�H;��H;��H;\�H;�H;��H;��H;�H;}�H;��H;�I;LI;I;'
I;@I;:I;YI;:I;I;�I;NI;W I;"I;�#I;�$I;�%I;      �'I;�'I;�&I;�%I;%$I;?"I;�I;mI;�I;�I;�I;pI;HI;)I;I;I;0I;g�H;��H;��H;`�H;/�H;B�H;��H;&�H;��H;��H;��H;��H;��H;,�H;��H; �H;��H;��H;a�H;o�H;c�H;��H;��H;�H;��H;)�H;��H;��H;��H;��H;��H;'�H;��H;F�H;.�H;W�H;��H;��H;m�H;2I;I;I;(I;HI;mI;�I;�I;�I;oI;�I;@"I;&$I;�%I;�&I;�'I;      T.I;:.I;Z-I;�+I;=*I;(I;~%I;�"I;�I;HI;�I;lI;�I;CI;�
I;qI;HI;8I;k�H;��H;��H;W�H;5�H;S�H;��H;O�H;�H;��H;��H;�H;n�H;��H;H�H;��H;��H;��H;z�H;��H;��H;��H;K�H;��H;m�H;�H;��H;��H;�H;Q�H;��H;S�H;9�H;V�H;��H;��H;j�H;9I;LI;uI;�
I;FI;�I;lI;�I;II;�I;�"I;�%I;
(I;<*I;,I;\-I;?.I;      �9I;x9I;�8I;7I;5I;r2I;Z/I;�+I;&(I;*$I; I;�I;�I;uI;yI;�I;�I;rI;<I;5�H;|�H;�H;��H;��H;��H;�H;��H;��H;��H;��H;��H;#�H;��H;5�H;��H;��H;��H;��H;��H;3�H;��H;#�H;��H;��H;~�H;��H;��H;!�H;��H;��H;��H;�H;q�H;3�H;?I;uI;�I;�I;yI;xI;�I;�I; I;-$I;)(I;�+I;e/I;n2I;5I;7I;�8I;}9I;      �KI;RKI;�II;�GI;FEI;�AI;>I;�9I;�4I;�/I;�*I;�%I;w I;gI;|I;�I;fI;-	I;<I;�I;~�H;��H;��H;u�H;d�H;r�H;��H;��H;H�H;9�H;O�H;��H;�H;��H;J�H;�H;.�H;�H;G�H;��H;�H;��H;O�H;2�H;A�H;��H;��H;u�H;a�H;r�H;��H;��H;w�H;�I;=I;-	I;hI;�I;|I;hI;z I;�%I;�*I;�/I;�4I;�9I;>I;�AI;JEI;HI;JI;OKI;      CdI;�cI;9bI;�_I;)\I;�WI;�RI;MI;GI;�@I;:I;Z3I;�,I;f&I;4 I;JI;�I;�I;�
I;�I;�I;��H;��H;��H;n�H;O�H;Q�H;��H;V�H;�H;�H;L�H;��H;"�H;��H;��H;��H;��H;��H;%�H;��H;L�H;�H;�H;N�H;��H;N�H;P�H;k�H;��H;��H;��H;�I;�I;�
I;�I;�I;MI;5 I;g&I;�,I;\3I;:I;�@I;GI;MI;�RI;�WI;)\I;�_I;?bI;�cI;      Z�I;��I;y�I;��I;8|I;]vI;�oI;
hI;�_I;gWI;�NI;FI;�=I;-5I;=-I;�%I;�I;&I;0I;�I;�I;vI;��H;,�H;�H;r�H;J�H;X�H;��H;,�H;�H;�H;T�H;��H;v�H;,�H;��H;-�H;r�H;��H;T�H;�H;�H;)�H;��H;R�H;I�H;x�H;�H;)�H;��H;xI;�I;�I;3I;&I;�I;�%I;<-I;-5I;�=I;FI;�NI;hWI;�_I;hI;�oI;[vI;B|I;�I;}�I;��I;      5�I;@�I;��I;�I;��I;�I;��I;s�I;w�I;vI;mjI;�^I;�SI;�HI;d>I;�4I;�+I;L#I;�I;�I;�I;?	I;iI;* I;��H;;�H;��H;Z�H;U�H;��H;)�H;�H;4�H;��H;�H;��H;��H;��H;�H;��H;6�H;�H;)�H;��H;N�H;V�H;��H;@�H;��H;& I;pI;@	I;�I;�I;�I;I#I;�+I;�4I;b>I;�HI;�SI;�^I;pjI;vI;t�I;o�I;��I;ޟI;��I;�I;��I;9�I;      ��I;�I;��I;R�I;��I;��I;��I;,�I;/�I;��I;k�I;
�I;�pI;]bI;�TI;�GI;'<I;z1I;�'I;I;]I;hI;z
I;5I;� I;��H;j�H;��H;P�H;J�H;��H;P�H;?�H;��H;��H;��H;��H;��H;��H;�H;@�H;N�H;��H;K�H;J�H;��H;i�H;��H;� I;/I;
I;kI;ZI;I;�'I;v1I;'<I;�GI;�TI;]bI;�pI;�I;n�I;��I;*�I;-�I;��I;��I;��I;V�I;��I;��I;      �I;\�I;��I;��I;��I;.�I;��I;G�I;�I;s�I;��I;	�I;�I;ۃI;�qI;�`I;QI;�CI;!7I;�+I;%"I;oI;�I;|I;�I;� I;��H;j�H;��H;Q�H;U�H;��H;��H;��H;��H;��H;q�H;��H;��H;��H;��H;��H;T�H;Q�H;��H;f�H;��H;� I;�I;xI;�I;oI;""I;�+I;#7I;�CI;�QI;�`I;�qI;ڃI;�I;	�I;��I;v�I; �I;@�I;��I;�I;��I;��I;��I;\�I;      d I;R'I;�:I;�XI;�{I;�I;z�I;�I;�I;�I;S�I;��I;g�I;�I;@�I;�I;�lI;�ZI;`JI;<I;�/I;�$I;I;I;I;I;I;��H;t�H;��H;I�H;T�H;��H;��H;�H;��H;n�H;��H;�H;��H;��H;T�H;L�H;��H;p�H;��H;I;I;I;�I;"I;�$I;�/I;<I;cJI;�ZI;�lI;�I;@�I;�I;i�I;��I;U�I;�I;�I;��I;~�I;�I;�{I;�XI;�:I;='I;      ��F;B�F;��F;Y2G;*�G;&H;T�H;�I;�lI;��I;R�I;p�I;��I;��I;��I;��I;v�I;�wI;�bI;#PI;)@I;:2I;X&I;0I;|I;4I;I; I;��H;@�H;w�H;T�H;{�H;'�H;]�H;��H;��H;��H;Z�H;'�H;|�H;V�H;{�H;B�H;��H;� I;I;;I;{I;.I;[&I;=2I;'@I;&PI;�bI;�wI;x�I;��I;��I;��I;��I;m�I;X�I;��I;�lI;�I;Y�H;�%H;4�G;`2G;��F;5�F;      ��?;��?;��@;]tA;��B;I�C;�BE;U�F;l�G;_xH;�I;͏I;t�I;��I;7�I;��I;�I;0�I;�I;iI;�TI;�BI;�3I;E'I;�I;vI;I;�I;� I;z�H;�H;k�H;]�H;��H;��H;'�H;��H;(�H;��H;��H;a�H;k�H;�H;~�H;� I;�I;I;I;�I;D'I;�3I;�BI;�TI;iI;�I;+�I;�I;��I;7�I;��I;v�I;ʏI;�I;axH;h�G;R�F;�BE;<�C;�B;atA;��@;��?;      ��0;z51;�2;W�4;�07;3#:;�/=;� @;�B;�	E;��F;N%H;	I;Q�I;��I;��I;��I;��I;`�I;��I;�mI;DWI;�DI;�4I;@'I;'I;�I;|I;8I;* I;,�H;��H;z�H;��H;a�H;��H;j�H;��H;`�H;��H;~�H;��H;1�H;0 I;6I;{I;�I;.I;>'I;�4I;�DI;EWI;�mI;��I;e�I;��I;��I;��I;��I;N�I;�	I;M%H;��F;�	E;�B;� @;�/=;*#:;�07;s�4;�2;c51;      C;�;"�;��;� ;�&;�\,;և2;98;�/=;�FA;lrD;P�F;JH;[9I;-�I;i�I;W�I;��I;��I;p�I;pI;CXI;�DI;�3I;U&I;I;�I;�
I;iI;��H;��H;��H;��H;9�H;H�H;�H;H�H;8�H;��H;��H;��H;��H;oI;|
I;�I;I;\&I;�3I;�DI;EXI;pI;s�I;��I;��I;S�I;l�I;,�I;[9I;JH;T�F;krD;�FA;�/=;98;Ӈ2;�\,;�&;� ;��; �;�;      <��:��:��:���:���:�P ;�e;�V;I#;e-;��5;�h<;OtA;T	E;�eG;7�H;.�I;
�I;��I;�I;�I;�I;pI;HWI;�BI;:2I;�$I;sI;nI;?	I;uI;��H;��H;�H;V�H;/�H;��H;3�H;U�H;�H;��H;��H;{I;D	I;lI;qI;�$I;A2I;�BI;NWI;pI;��I;�I;�I;��I;�I;/�I;6�H;�eG;V	E;RtA;�h<;��5;e-;L#;�V;�e;�P ;��:��:��:y�:      ��p� �,��!9�ų9��":��u:��:Z��:���:(R;\ ;��,;�6;P)>;�;C;��F;�lH;hkI;q�I;��I;��I;�I;l�I;�mI;|TI;@I;�/I;""I;VI;�I;�I;�I;r�H;r�H;��H;Q�H;��H;S�H;��H;o�H;u�H;�I;�I;�I;VI;""I;�/I;#@I;yTI;�mI;n�I;�I;��I;��I;t�I;fkI;�lH;��F;�;C;R)>;�6;��,;` ;.R;���:`��:��:��u:�":�ų9�"9 �,�      p&�~!��4����氺�O��<T��t�9��u:�#�:�G�:D;)#;g71;=;;��A;��E;�$H;HVI;�I;��I;�I;��I;��I;iI;"PI;<I;�+I;I;�I;�I;�I;�I;3�H;��H;��H;�H;��H;��H;0�H;�I;�I;�I;�I;I;�+I;<I;&PI;	iI; �I;��I;�I;��I;�I;MVI;�$H;��E;��A;;;;g71;)#;D;�G�:�#�:��u:�t�9�<T�(�O��氺���4��!�      �kٻl�Ի�ǻ����V���n���+�8�Ժ��1��39Pm:��:l�;�;{\,;��8;��@;<]E;�
H;IVI;r�I;��I;��I;`�I;��I;�bI;[JI;#7I;�'I;�I;.I;�
I;6I;9I;i�H;��H;w�H;��H;d�H;8I;8I;�
I;2I;�I;�'I;%7I;`JI;�bI;��I;i�I;��I;��I;t�I;OVI;�
H;;]E;��@;ߍ8;{\,;
�;l�;��:Tm:�39 �1�8�Ժ��+��n��V������ǻh�Ի      6yY��|U�N�I�@�7��� ��!���Ի�᝻��T���#��u�9���:Ol�:�;�);17;, @;:]E;�$H;dkI;
�I;U�I;��I;+�I;�wI;�ZI;�CI;z1I;K#I;&I;�I;+	I;rI;6I;k�H;��H;m�H;5I;pI;-	I;�I;)I;P#I;x1I;�CI;�ZI;�wI;&�I;��I;U�I;�I;dkI;�$H;:]E;, @;17;�);�;Ql�:���:�u�9�#����T��᝻��Ի "��� �@�7�P�I��|U�      ��ü^l��w����R��?ߓ�a�{��M��� �!��˼����B�갺�Ho���u:���:�R;0�';17;��@;��E;�lH;/�I;h�I;��I;	�I;s�I;�lI;QI;*<I;�+I;�I;�I;cI;�I;CI;/I;�I;/I;AI;�I;bI;�I;�I;�+I;)<I;QI;�lI;s�I;�I;��I;k�I;1�I;�lH;��E;��@;17;0�';�R;���:��u:@Ho�갺��B�̼�� �컋� ��M�`�{�@ߓ��R��x���]l��      �'��-$�_��X����
?ټw��:���pyY��k� �Ի:��Y������ $R:���:�R;�);ٍ8;��A;��F;6�H;*�I;��I;��I;��I; �I;�`I;�GI;�4I;�%I;HI;�I;�I;qI;I;EI;I;nI;�I;�I;FI;�%I;�4I;�GI;�`I;�I;��I;��I;��I;-�I;7�H;��F;��A;ڍ8;�);�R;���:�#R:����Y��:����Ի�k�pyY�;���	w��
?ټ���Y�_���-$�      Y+����c̀�-l��Q�%�2�B��������@����>�Z2��#V���1���� $R:���:�;t\,;4;;�;C;�eG;[9I;��I;1�I;��I;=�I;�qI;�TI;`>I;9-I;0 I;xI;tI;�
I;I;I;I;�
I;rI;zI;- I;9-I;`>I;�TI;�qI;@�I;��I;-�I;��I;[9I;�eG;�;C;7;;s\,;�;���:�#R:���1�$V��Z2����>��@��������B�%�2��Q�.l�c̀���      j�ྲྀhܽp�н]y��^什P ��l��n<�M���>ټ��V|U���������1�������u:Ol�:�;d71;U)>;T	E;JH;R�I;��I;��I;�I;փI;]bI;�HI;*5I;b&I;dI;qI;<I;"I;
I;&I;9I;qI;gI;_&I;(5I;�HI;]bI;ڃI;�I;��I;��I;X�I;JH;V	E;L)>;h71;�;Ol�:��u:�����1��������W|U����>ټM���n<�l�P ��_什^y��o�н�hܽ      ��4�f1��&������i�ང�������`��'���UR��E�]���!V���X���Ho����:h�;'#;�6;RtA;T�F;�	I;v�I;��I;j�I;�I;�pI;�SI;�=I;�,I;v I;�I;�I;FI;9I;FI;�I;�I;y I;�,I;�=I;�SI;�pI;�I;n�I;��I;q�I;�	I;U�F;QtA;�6;,#;h�;���: Ho��X��"V��~��F�]�UR����'��`��������h��������&�f1�      �x���o��ń�IUo���O�*�-�{��hܽ[什Ҽx���2�tb��UR��W|U�Z2��:��"갺pu�9��:D;��,;�h<;grD;P%H;ƏI;e�I;��I;�I;�I;�^I;	FI;S3I;�%I;�I;^I;hI;5I;iI;\I;�I;�%I;R3I;FI;�^I;
�I;�I;��I;c�I;��I;P%H;jrD;�h<;��,;D;��:xu�9"갺:��Z2��W|U�UR��tb����2�Ҽx�[什�hܽ{�*�-���O�IUo�ń��o��      v���ྃ�Ѿ(����נ�ń�9�S��#�_O��|n��J̀���2���𛼃�>� �Ի��B��#�4m:�G�:` ;��5;�FA;��F;�I;M�I;M�I;��I;k�I;mjI;�NI;:I;�*I;�I;�I;�I;LI;�I;�I;�I;�*I;:I;�NI;mjI;m�I;��I;N�I;J�I;�I;��F;�FA;��5;U ;�G�:,m:�#���B� �Ի��>�������2�J̀�|n��_O���#�9�S�ń��נ�(�����Ѿ��      �3���/��X#��	��A��֌Ⱦ�f��HUo�]1�˰��|n��Ѽx��'��>ټ�@���k�μ��$����39�#�:.R;e-;�/=;�	E;]xH;�I;
�I;m�I;�I;vI;dWI;�@I;�/I;%$I;:I;�I;6I;�I;<I;#$I;�/I;�@I;aWI;vI;�I;p�I;�I;�I;\xH;�	E;�/=;	e-;$R;�#�:��39"��μ���k��@���>ټ�'�Ҽx�|n��˰��^1�HUo��f��֌Ⱦ�A���	��X#���/�      ���T���T�v��RZ�[58�͂�p��d���foy�]1�_O��[什�`�M�����pyY�$�컚�T��1���u:���:H#;98;�B;j�G;�lI;�I;��I;/�I;v�I;�_I; GI;�4I;%(I;�I;�I;I;�I;�I;%(I;�4I; GI;�_I;q�I;-�I;�I;�I;�lI;h�G;�B;98;C#;���:��u:$�1���T�$��pyY����M���`�\什_O��]1�foy�d���p��͂�[58��RZ�T�v�T���      	Ŀ6g��&ﱿ���S����U��X#�t��d���IUo��#��hܽ����n<����<����� ��᝻F�Ժ�t�9h��:�V;̇2;� @;U�F;�I;��I;A�I;)�I;h�I;�gI;MI;�9I;�+I;�"I;hI;�I;iI;�"I;�+I;�9I;MI;�gI;i�I;(�I;C�I;��I;�I;T�F;� @;Ї2;�V;R��:�t�9F�Ժ�᝻�� �<�������n<�����hܽ�#�IUo�d���t���X#��U�S������&ﱿ6g��      ~x�P9�R��sؿnQ��e_��6�_��X#�p���f��9�S�{�����l�B�	w���M���Ի��+� =T���:�e;�\,;�/=;�BE;Q�H;v�I;��I;��I;��I;�oI;�RI;>I;\/I;{%I;�I;FI;�I;%I;]/I;>I;�RI;�oI;��I;��I;��I;x�I;V�H;�BE;�/=;�\,;�e;��:�<T���+���Ի�M�	w��B�l�����{�9�S��f��p���X#�6�_�e_��nQ��sؿR��P9�      �X1���,�h���<��5g��e_���U�͂�֌Ⱦń�*�-�i��P ��&�2�?ټb�{�"��n� �O���u:�P ;�&;*#:;<�C;�%H;�I;!�I;��I;�I;_vI;�WI;�AI;x2I;(I;C"I;` I;C"I;(I;x2I;�AI;�WI;[vI;�I;��I;'�I;�I;�%H;<�C;-#:;�&;�P ;��u:�O��n�"�b�{�?ټ&�2�P ��i��*�-�ń�֌Ⱦ͂��U�e_��5g��<�h����,�      d��]]�5K��X1�Zf��nQ��S���[58��A���נ���O���_什�Q����@ߓ��� ��V���氺��":Ҹ�: ;�07;�B;,�G;�{I;��I;��I;��I;8|I;4\I;IEI;5I;0*I;1$I;+"I;-$I;5*I;5I;LEI;5\I;5|I;��I;��I;��I;�{I;5�G;�B;�07; ;и�:�":�氺�V���� �@ߓ�����Q�_什����O��נ��A��[58�S���nQ���Zf��X1�5K��]]�      N������4z���V��X1��<�sؿ����RZ��	�(���IUo����^y��.l�Y��R��C�7�������ų9���:��;W�4;itA;Y2G;�XI;��I;K�I;�I;�I;�_I;�GI;"7I;�+I;�%I;�#I;�%I;�+I;7I;�GI;�_I;�I;�I;J�I;��I;�XI;e2G;gtA;X�4;��;���:�ų9
�����B�7��R��Y�.l�^y�����IUo�(����	��RZ����tؿ�<��X1���V��4z�����      �o��f^���ē��4z�5K�h��R��&ﱿT�v��X#���Ѿń��&�p�нc̀�_��v���M�I��ǻ�4��"9��:4�;�2;��@;��F;�:I;��I;��I;��I;v�I;KbI;�II;�8I;X-I;�&I;�$I;�&I;[-I;�8I;�II;KbI;r�I;��I;��I;��I;�:I;��F;��@;�2;2�;��: "9�4��ǻL�I�v���_��c̀�p�н�&�ń���Ѿ�X#�T�v�&ﱿR��h��5K��4z��ē�f^��      q'���X��f^�������]]���,�P9�6g��T�����/����o��g1��hܽ���-$�_l���|U�f�Ի�!� �,�u�:�;�51;��?;2�F;?'I;_�I;
�I;<�I;��I;�cI;>KI;x9I; .I;y'I;�%I;v'I; .I;x9I;@KI;�cI;��I;?�I;
�I;b�I;@'I;@�F;��?;�51;�;o�: �,�~!�g�Ի�|U�_l���-$����hܽg1��o���ྚ�/�T���6g��P9���,��]]�����f^���X��      l����������Т��/�j��5���	� �ȿ&8����7�D�꾂S���7�
3�~L���)���Ƽ��\��ݻ�+��Uɸ��:x;��0;��?;F�F;�+I;��I;��I;ѽI;�I;�hI;�NI;�<I;�0I;�)I;�'I;�)I;�0I;�<I;�NI;�hI;�I;սI;��I;��I;�+I;T�F;��?;�0;x;��:�Vɸ�+��ݻ��\���Ƽ�)�~L��
3��7��S��D�꾨�7�&8�� �ȿ��	��5�/�j�Т����������      ��������B��^�����c�621�%X��ÿiڇ�r�3��s��7��|74�a�>ى���&�Nü(�X���ػ��%� �J�ă�:�b;y�0;r�?;�F;�2I;��I;6�I;�I;E�I;PhI;�NI;0<I;w0I;a)I;�'I;\)I;z0I;.<I;�NI;PhI;A�I;�I;6�I;��I;�2I;�F;r�?;v�0;�b;���:��J���%���ػ(�X�Nü��&�>ى�a�|74��7���s�r�3�iڇ��ÿ%X�621���c�^����B�����      �����B����F��x�P���#�M�������x|��'�YD־�X��o�)�Խ�Ă�J<�9_��}-M���ʻ[��`&�8�:�;K2;v@;L�F;�FI;g�I;��I;'�I;��I;�fI;=MI;B;I;�/I;�(I;�&I;�(I;�/I;A;I;<MI;�fI;��I;*�I; �I;j�I;�FI;X�F;v@;K2;�;���:�%�8[����ʻ~-M�9_��J<��Ă�Խo�)��X��YD־�'��x|����M�����#�x�P�F�����B��      Т��^���F���/]��5�N���,ݿ+8��qm_��K��t��W�s�#>����9�o��3��۩���:�nT�����(�9�f�:�<;�_4;hA;8G;xdI;�I;'�I;Z�I;\�I;&dI;KI;�9I;H.I;�'I;�%I;�'I;K.I;�9I;KI;&dI;X�I;[�I;)�I;�I;wdI;8G;hA;�_4;�<;�f�:�'�9���qT����:��۩��3�9�o����#>�W�s��t���K�qm_�+8���,ݿN���5��/]�F��^���      /�j���c�x�P��5���s��I���hڇ�Fv<�(���p���_S��������
+T��� �+$���G#�ђ��p1���:���:3�;/7;n�B;z�G;��I;�I;c�I;ȮI;��I;�`I;IHI;�7I;a,I;&I; $I;&I;b,I;�7I;IHI;�`I;��I;̮I;a�I;�I;��I;��G;o�B;,7;0�;���:�:n1��Ғ���G#�+$���� �
+T���������_S�p��(���Fv<�hڇ�I���s�����5�x�P���c�      �5�621���#�N��r���ÿ�ҕ�Z������̾�X���0�3�.W����5��zܼA��Z��c�s��U\�h�n:���:ج%;��9;��C;�.H;�I;�I;�I;��I;u{I;\I;�DI;�4I;(*I;$I;"I;$I;(*I;�4I;�DI;\I;r{I;��I; �I;�I;�I;�.H;��C;��9;ج%;���:H�n:�U\�d�s�Z��A���zܼ��5�.W��3��0��X����̾���Z��ҕ��ÿs��N����#�621�      ��	�%X�M����,ݿI����ҕ��d��'�@��#���x�W����k���2�o��G��*���Q���ػ�0���~���:z�;0,;b=;7BE;��H;�I;��I;B�I;�I;`tI;�VI;�@I;�1I;�'I;�!I;�I;�!I;�'I;�1I;�@I;�VI;]tI;�I;D�I;��I;|�I;��H;8BE;`=;.,;x�;��:`�~��0���ػ�Q��*���G�2�o�k������x�W�#���@�꾌'��d��ҕ�I����,ݿM���%X�       �ȿ�ÿ���+8��hڇ�Z��'�����l8��W�s�,�&�X�/i??��V�琼WG#�c7��~Tܺh�9W�:��;L2;P@;ބF;�I;��I;u�I;M�I;A�I;�lI;�PI;[<I;�-I;�$I;%I;DI;"I;�$I;�-I;Z<I;�PI;�lI;F�I;O�I;u�I;��I;�I;�F;L@;L2;��;W�:��9~Tܺd7��WG#�琼�V�i??�/X�,�&�W�s�l8�������'�Z�hڇ�+8������ÿ      &8��iڇ��x|�qm_�Fv<����?��l8��$6~�o74��l��{���7nc�4���^����\��9�JZ���=���n:F��:�#;�8;��B;q�G;�xI;m�I;��I;��I;چI;5dI;xJI;�7I;*I;5!I;PI;�I;LI;5!I;*I;�7I;wJI;5dI;݆I;��I;��I;m�I;�xI;t�G;��B;�8;�#;>��:��n:��=�MZ��9���\��^��4��7nc�{����l��o74�$6~�l8��?�꾎��Fv<�qm_��x|�iڇ�      ��7�r�3��'��K�'�����̾#���W�s�o74����!N��·|���)�9zܼ�Y��@ ����D����S9Љ�:!�; -;=;�E;��H;J�I;/�I;��I;��I;{I;^[I;�CI;X2I;&I;�I;-I;�I;+I;�I;&I;V2I;�CI;`[I;{I;��I;��I;,�I;E�I;�H;�E;=; -;�;ډ�:�S9F������@ ��Y��8zܼ��)�·|�!N�����o74�W�s�#�����̾'����K��'�r�3�      D���s�YD־�t��p���X��x�W�,�&��l��!N���Ă�j�5�����|Q����A�E�ػ��G�"/�f:�a�:��;`�5;�9A;E�F;�*I;��I;��I;
�I;Z�I;/oI;gRI;�<I;-I;�!I;AI;I;�I;I;CI;�!I;-I;�<I;iRI;2oI;^�I;�I;��I;��I;�*I;C�F;�9A;b�5;��;b�:$f: "/���G�F�ػ��A�|Q������i�5��Ă�!N���l��,�&�x�W��X��p���t��YD־�s�      �S���7���X��W�s��_S��0����W�{���·|�i�5�j���ک�5�X� c �z��3����9
��:�;��,;�L<;SoD;.H;I;��I;��I;S�I;N�I;7cI;[II;�5I;�'I;GI;�I;�I;�I;�I;�I;JI;�'I;�5I;\II;:cI;W�I;W�I;��I;��I;ěI;.H;VoD;�L<;��,;�;��:��9�3��z�!c �4�X��ک�i��i�5�·|�{���Wར��~�0��_S�W�s��X���7��      �7�|74�o�)�#>����3�k���/7nc���)������ک�va��Q�T���N���ȸ ��:��;�#;r�6;hA;��F;�I;4�I;]�I;�I;v�I;�uI;mWI;r@I;
/I;c"I;I;�I;gI;[I;gI;�I;I;c"I;/I;v@I;qWI;�uI;z�I;�I;W�I;8�I;�I;��F;hA;o�6;�#;��;��:@�ȸN�T����Q�va��ک�������)�7nc�/k���3����#>�o�)�|74�      	3�`�Խ�������/W��1�o�h??�4��8zܼ|Q��4�X��Q��6�������Ϲx�n:�m�:>;��0;�>;.E;MSH;J�I;��I;^�I;?�I;U�I;�fI;"LI;�7I;e(I;I;�I;^I;I;>I;I;]I;�I;I;`(I;�7I;'LI;�fI;Z�I;=�I;W�I;��I;G�I;NSH;0E;�>;��0;>;�m�:��n:��Ϲ����6���Q�4�X�|Q��8zܼ4��h??�1�o�.W���������Խ`�      }L��>ى��Ă�8�o�
+T���5��G��V��^���Y����A� c �V���������4�J:Yl�:�e;,;��:;5C;lG;�DI; �I;��I;��I;��I;�vI;�XI;BAI;�/I;"I;�I;�I;�I;�I;HI;�I;�I;�I;�I;"I;�/I;FAI;�XI;�vI;��I;��I;��I;��I;�DI;lG;5C;��:; ,;�e;al�:,�J:������V��� c ���A��Y���^���V��G���5�+T�8�o��Ă�>ى�      �)���&�I<��3��� ��zܼ�*��琼��\�@ �E�ػ{�!N���Ϲ0�J:pj�:f�;t�(;�e8;��A;�F;��H;�I;j�I;��I;��I;]�I;\eI;�KI;7I;�'I;�I;I;�I;aI;�I;'I;�I;^I;�I;I;�I;�'I;7I;�KI;aeI;\�I;�I;�I;g�I;�I;��H;�F;��A;�e8;n�(;i�;nj�:0�J:��Ϲ"N�z�D�ػ? ���\�琼�*���zܼ�� ��3�I<���&�      ��ƼNü9_���۩�*$��A���Q�TG#��9�����G��3����ȸ��n:al�:m�;�';�7;qv@;�E;vH;�I;��I;��I;8�I;��I;�qI;qUI;*?I;�-I;y I;I;kI;�I;CI;�I;I;�I;@I;�I;jI;I;} I;�-I;,?I;tUI;�qI;z�I;;�I;��I;��I;�I;vH;!�E;qv@;�7;�';l�;al�:��n:��ȸ�3����G�����9�TG#��Q�@��+$���۩�:_��Nü      ��\�%�X�~-M���:��G#�X����ػ`7��JZ�6���"/���9��:�m�:�e;q�(;7;�@;!]E;}-H;1wI;t�I;��I;��I;��I;�|I;�^I;�FI;�3I;J%I;�I;�I;D
I;?I;"I;- I;r�H;* I;I;<I;C
I;�I;�I;M%I;�3I;�FI;�^I;�|I;��I;��I;��I;t�I;0wI;�-H;!]E;�@;�7;n�(;�e;�m�:��:��9"/�:���EZ�`7����ػX���G#���:�|-M�%�X�      �ݻ��ػ��ʻnT��Ғ��S�s���0�jTܺ��=�@T9@f:��:��;>;",;�e8;qv@;(]E;/H;�aI;�I;��I;=�I;��I;Q�I;�fI;�MI;�9I;�)I;iI;mI;�I;2I;I;G�H;~�H;��H;z�H;B�H;I;0I;�I;oI;iI;�)I;�9I;�MI;�fI;U�I;��I;4�I;��I;�I; bI;,H;!]E;sv@;�e8; ,;>;��;��:@f: T9��=�pTܺ��0�Z�s�ђ��rT����ʻ��ػ      �+���%�T�� ����1���U\���~�P�9��n:ډ�:
b�:�;�#;��0;��:;��A;!�E;�-H; bI;��I;d�I;y�I;�I;��I;�mI;�SI;?I;2.I;� I;VI;�I;^I;uI;��H;o�H;�H;r�H;	�H;l�H;��H;wI;ZI;�I;TI;� I;6.I;?I;�SI;�mI;��I;�I;w�I;e�I;��I;bI;-H; �E;��A;��:;��0;�#;�;
b�:؉�:��n:h�90�~��U\�t1�����b����%�      @Qɸ��J��#�8�'�9Ч:X�n:��:W�:@��: �;��;��,;p�6;�>;
5C;�F;vH;9wI;�I;d�I;3�I;��I;U�I;�rI;�XI;2CI;�1I;'$I;�I;�I;�I;EI;;�H;.�H;��H;��H;r�H;��H;��H;,�H;;�H;>I;�I;�I;�I;'$I;�1I;/CI;�XI;�rI;M�I;¸I;4�I;c�I;�I;4wI;vH;�F;	5C;�>;o�6;��,;��;�;4��:	W�:��:H�n:��:�'�9�$�8 �J�      ��:܃�:ޓ�:�f�:���:���:x�;��;�#;-;f�5;�L<;hA;3E;lG;��H;��I;w�I;��I;}�I;øI;�I;�tI;u[I;FFI;�4I;�&I;2I;�I;O
I;hI;��H;
�H;s�H;��H;��H;d�H;��H;��H;s�H;�H;��H;kI;N
I;�I;2I;�&I;�4I;HFI;r[I;�tI;�I;øI;z�I;��I;t�I;��I;��H;lG;.E;�gA;�L<;f�5;�-;�#;��;��;���:ͱ�:�f�:ȓ�:ă�:      .x;�b;�;�<;%�;�%;;,;+L2;�8;=;�9A;`oD;��F;\SH;�DI;$�I;��I;��I;=�I;�I;T�I;�tI;]\I;�GI;|6I;�(I;�I;=I;�I;MI;B I;r�H;J�H;�H;��H;��H;��H;��H;��H;�H;J�H;o�H;E I;JI;�I;@I;�I;�(I;�6I;�GI;V\I;�tI;T�I;�I;=�I;��I;��I;!�I;�DI;USH;��F;\oD;�9A;=;�8;'L2;8,;۬%;6�;�<;�;�b;      ��0;��0;	K2;�_4;"7;��9;[=;O@;��B;�E;A�F;.H;�I;K�I;��I;i�I;��I;��I;��I;��I;rI;m[I;�GI;7I;m)I;�I;PI;�I;0I;� I;��H;��H;��H;��H;��H;�H;��H;�H;��H;��H;��H;��H;��H;� I;,I;�I;LI;�I;q)I;7I;�GI;n[I;~rI;��I;��I;��I;��I;g�I;��I;D�I;�I;.H;D�F;�E;��B;S@;Y=;��9;*7;�_4;K2;��0;      Ǥ?;s�?;v@;hA;c�B;��C;<BE;�F;u�G;�H;�*I;̛I;4�I;��I;��I;�I;B�I;��I;\�I;�mI;�XI;GFI;�6I;x)I;YI;�I;4I;�I;vI;2�H;��H;��H;��H;(�H;�H;l�H;/�H;f�H;�H;)�H;��H;��H;��H;2�H;oI;�I;.I;�I;[I;s)I;6I;JFI;�XI;�mI;\�I;��I;B�I;�I;��I;��I;5�I;˛I;�*I;�H;t�G;ބF;>BE;��C;n�B;hA;v@;s�?;      H�F;�F;H�F;
8G;p�G;�.H;��H;I;�xI;S�I;��I;��I;`�I;e�I;��I;��I;��I;�|I;�fI;�SI;4CI;�4I;�(I;�I;�I;qI;-I;�I;o�H;��H;��H;��H;��H;��H;��H;��H;��H;��H;��H;��H;��H;��H;��H;��H;j�H;�I;(I;tI;�I;�I;�(I;�4I;2CI;�SI;�fI;�|I;��I;��I;��I;_�I;^�I;��I;��I;R�I;�xI; I;��H;�.H;��G;8G;G�F;�F;      ,I;�2I;�FI;|dI;��I;�I;��I;��I;p�I;1�I;��I;��I;�I;?�I;��I;\�I;�qI;�^I;�MI;?I;�1I;�&I;�I;TI;1I;,I;�I;��H;�H;��H;��H;��H;5�H;�H;)�H;��H;��H;��H;(�H;�H;6�H;��H;��H;��H;�H;��H;�I;-I;5I;OI;�I;�&I;�1I;?I;�MI;�^I;�qI;_�I;��I;;�I;�I;��I;��I;,�I;l�I;��I;~�I;�I;ʇI;pdI;�FI;�2I;      ��I;��I;d�I;�I;�I;�I;��I;u�I;��I;��I;�I;X�I;s�I;[�I;�vI;[eI;pUI;�FI;�9I;3.I;,$I;-I;=I;�I;�I;�I;��H;0�H;�H;��H;~�H;��H;��H;��H; �H;��H;��H;��H; �H;��H;��H;��H;~�H;��H;�H;.�H;��H;�I;�I;~I;;I;,I;'$I;..I;�9I;�FI;oUI;^eI;�vI;Z�I;u�I;X�I;�I;��I;��I;p�I;��I;�I;�I;
�I;d�I;��I;      ��I;+�I;��I;8�I;W�I;�I;H�I;V�I;��I;��I;\�I;W�I;�uI;�fI;�XI;�KI;/?I;�3I;�)I;� I;�I;�I;�I;.I;oI;h�H;�H;�H;��H;|�H;��H;��H;N�H;��H;8�H;��H;��H;��H;6�H;��H;N�H;��H;��H;x�H;��H;�H;	�H;c�H;oI;'I;�I;�I;�I;� I;�)I;�3I;-?I;�KI;�XI;�fI;�uI;U�I;a�I;��I;��I;U�I;I�I;��I;a�I;;�I;��I;'�I;      սI;�I;4�I;Y�I;ŮI;��I;�I;K�I;݆I;{I;4oI;DcI;qWI;*LI;FAI;7I;�-I;G%I;fI;VI;�I;K
I;JI;� I;5�H;��H;��H;��H;��H;��H;��H;F�H;\�H;��H;"�H;��H;��H;��H;�H;��H;Z�H;C�H;��H;��H;|�H;��H;��H;��H;5�H;� I;II;J
I;�I;QI;cI;C%I;�-I;7I;DAI;&LI;nWI;>cI;3oI;!{I;݆I;D�I;�I;��I;ŮI;a�I;2�I;�I;      �I;]�I;�I;f�I;��I;v{I;`tI;�lI;:dI;g[I;nRI;hII;y@I;�7I;�/I;�'I;� I;�I;qI;I;�I;iI;B I;��H;��H;��H;��H;��H;��H;��H;7�H;5�H;��H;��H;k�H;D�H;0�H;B�H;j�H;��H;��H;5�H;9�H;��H;��H;�H;��H;��H;��H;��H;C I;hI;�I;�I;oI;�I;� I;�'I;�/I;�7I;w@I;cII;nRI;h[I;:dI;�lI;htI;o{I;��I;g�I;��I;]�I;      �hI;ZhI;�fI;dI;|`I;�[I;�VI;�PI;|JI;�CI;�<I;�5I;/I;i(I;"I;�I;I;�I;�I;cI;NI;��H;p�H;��H;��H;��H;��H;�H;��H;H�H;2�H;��H;��H;0�H;��H;��H;��H;��H;��H;3�H;��H;~�H;1�H;D�H;��H;��H;��H;��H;��H;��H;s�H;��H;DI;\I;�I;�I;I;�I;"I;g(I;	/I;�5I;�<I;�CI;zJI;�PI;�VI; \I;�`I;%dI;�fI;[hI;      �NI;�NI;<MI;KI;FHI;�DI;�@I;W<I;|7I;R2I;-I;�'I;d"I;I;�I;I;pI;D
I;7I;{I;H�H;�H;I�H;��H;��H;��H;6�H;��H;V�H;_�H;��H;��H;�H;��H;w�H;3�H;.�H;3�H;u�H;��H;�H;��H;��H;W�H;Q�H;��H;5�H;��H;��H;��H;L�H;�H;@�H;tI;6I;C
I;qI;I;�I;I;b"I;�'I;-I;T2I;}7I;T<I;�@I;�DI;IHI;KI;IMI;�NI;      �<I;.<I;;;I;�9I;�7I;�4I;�1I;.I;*I;&I;�!I;SI;I;�I;�I;�I;�I;<I;	I; �H;7�H;t�H;��H;��H;%�H;��H;�H;��H;��H;��H;��H;2�H;��H;O�H;�H;��H;��H;��H;�H;O�H;��H;2�H;��H;��H;��H;��H;�H;��H;(�H;��H;�H;s�H;0�H;��H;I;=I;�I;�I;�I;�I;I;NI;�!I;&I;*I;�-I;�1I;�4I;�7I;�9I;E;I;;<I;      �0I;�0I;�/I;M.I;k,I;!*I;�'I;�$I;9!I;�I;KI;�I;I;gI;�I;dI;GI; I;H�H;s�H;��H;��H;��H;��H;�H;}�H;%�H;!�H;?�H;%�H;e�H;��H;w�H;�H;��H;��H;��H;��H;��H;�H;w�H;��H;c�H;�H;6�H;�H;%�H;|�H;�H;��H;��H;��H;��H;n�H;E�H;!I;GI;eI;�I;gI;I;�I;NI;�I;9!I;�$I;�'I;%*I;e,I;U.I;�/I;�0I;      �)I;i)I;�(I;�'I;�%I;$I;�!I;)I;LI;4I;I;�I;hI;"I; 	I;�I;�I;' I;�H;�H;��H;��H;��H;��H;f�H;��H;��H;��H;��H;��H;B�H;��H;7�H;��H;��H;f�H;f�H;j�H;��H;��H;7�H;��H;@�H;��H;��H;��H;��H;��H;f�H;��H;��H;��H;��H;	�H;~�H;* I;�I;�I; 	I;%I;hI;�I;I;4I;MI;%I;�!I;$I;�%I;�'I;�(I;v)I;      �'I;�'I;�&I;�%I;�#I;"I;�I;LI;�I;�I;�I;�I;_I;GI;QI;*I;%I;t�H;��H;{�H;~�H;g�H;��H;��H;.�H;��H;��H;��H;��H;��H;*�H;��H;.�H;��H;��H;c�H;I�H;e�H;��H;��H;/�H;��H;)�H;��H;��H;��H;��H;��H;.�H;��H;��H;f�H;v�H;w�H;��H;t�H;$I;-I;QI;HI;_I;�I;�I;�I;�I;JI;�I;"I;�#I;�%I;�&I;�'I;      �)I;j)I;�(I;�'I;�%I;$I;�!I;(I;LI;4I;I;�I;jI;%I;�I;�I;�I;' I;�H;�H;��H;��H;��H;��H;f�H;��H;��H;��H;��H;��H;B�H;��H;9�H;��H;��H;f�H;f�H;j�H;��H;��H;7�H;��H;@�H;��H;��H;��H;��H;��H;f�H;��H;��H;��H;��H;
�H;~�H;* I;�I;�I; 	I;#I;hI;�I;I;1I;MI;(I;�!I;$I;�%I;�'I;�(I;q)I;      �0I;�0I;�/I;H.I;k,I;!*I;�'I;�$I;9!I;�I;KI;�I;I;eI;�I;bI;FI;!I;H�H;r�H;��H;��H;��H;��H;�H;|�H;%�H;!�H;=�H;"�H;d�H;��H;x�H;�H;��H;��H;��H;��H;��H;�H;w�H;��H;c�H;�H;8�H;�H;#�H;}�H;�H;��H;��H;��H;��H;n�H;H�H;!I;II;eI;�I;gI;I;�I;NI;�I;9!I;�$I;�'I;"*I;i,I;R.I;�/I;�0I;      �<I;0<I;:;I;�9I;�7I;�4I;�1I;.I;*I;&I;�!I;PI;I;�I;�I;�I;�I;?I;	I;��H;7�H;t�H;��H;��H;(�H;��H;�H;��H;��H;��H;��H;0�H;��H;N�H;�H;��H;��H;��H;�H;N�H;��H;2�H;��H;��H;��H;��H;�H;��H;&�H;��H;�H;t�H;-�H;��H;I;=I;�I;�I;�I;�I;I;NI;�!I;&I;*I;�-I;�1I;�4I;�7I;�9I;B;I;3<I;      �NI;�NI;?MI;KI;CHI;�DI;�@I;]<I;7I;R2I;-I;�'I;b"I;I;�I;I;pI;C
I;5I;xI;G�H;�H;G�H;��H;��H;��H;4�H;��H;V�H;^�H;��H;��H;�H;��H;x�H;3�H;.�H;3�H;w�H;��H;�H;��H;��H;W�H;N�H;��H;4�H;��H;��H;��H;M�H;�H;>�H;xI;5I;A
I;nI;I;�I;I;d"I;�'I;-I;R2I;7I;X<I;�@I;�DI;HHI;#KI;PMI;�NI;      �hI;]hI;�fI;dI;}`I;\I;�VI;�PI;zJI;�CI;�<I;�5I;	/I;g(I;"I;�I;I;�I;�I;^I;LI;��H;o�H;��H;��H;��H;��H;�H;��H;F�H;/�H;}�H;��H;/�H;��H;��H;��H;��H;��H;0�H;��H;~�H;.�H;C�H;��H;��H;��H;��H;��H;��H;u�H;��H;DI;\I;�I;�I;I;�I;"I;h(I;/I;�5I;�<I;�CI;{JI;�PI;�VI;�[I;}`I;)dI;�fI;XhI;      �I;^�I;�I;_�I;��I;v{I;`tI;�lI;8dI;d[I;jRI;fII;v@I;�7I;�/I;�'I;� I;�I;oI;�I;�I;hI;? I;��H;��H;��H;��H;��H;��H;��H;6�H;5�H;��H;��H;n�H;B�H;0�H;E�H;h�H;��H;��H;5�H;5�H;��H;��H;~�H;��H;��H;��H;��H;E I;iI;�I;�I;qI;�I;� I;�'I;�/I;�7I;w@I;cII;mRI;e[I;<dI;�lI;htI;t{I;��I;j�I;�I;`�I;      ۽I;�I;.�I;a�I;��I;��I;�I;K�I;݆I;!{I;/oI;AcI;nWI;'LI;GAI;7I;�-I;F%I;cI;TI;�I;K
I;FI;� I;5�H;��H;��H;��H;��H;��H;��H;F�H;X�H;��H; �H;��H;��H;��H;�H;��H;[�H;F�H;��H;��H;{�H;��H;��H;��H;4�H;� I;MI;K
I;�I;QI;fI;C%I;�-I;7I;GAI;'LI;nWI;>cI;0oI;"{I;܆I;J�I;�I;�I;îI;i�I;6�I;�I;      ��I;,�I;�I;.�I;H�I;�I;E�I;S�I;��I;��I;^�I;W�I;�uI;�fI;�XI;�KI;-?I;�3I;�)I;� I;�I;�I;�I;+I;oI;a�H;�H;�H;��H;w�H;��H;��H;N�H;��H;9�H;��H;��H;��H;6�H;��H;N�H;��H;��H;x�H;��H;�H;�H;f�H;mI;%I;�I;�I;�I;� I;�)I;�3I;-?I;�KI;�XI;�fI;�uI;T�I;_�I;��I;��I;U�I;L�I;�I;W�I;1�I;�I;'�I;      ��I;��I;Y�I;�I;�I;�I;��I;u�I;��I;��I;
�I;Z�I;u�I;Z�I;�vI;\eI;oUI;�FI;�9I;..I;*$I;-I;:I;�I;�I;�I;��H;.�H;�H;��H;|�H;��H;��H;��H; �H;��H;��H;��H;�H;��H;��H;��H;~�H;��H;�H;,�H;��H;�I;�I;~I;@I;-I;'$I;..I;�9I;�FI;qUI;^eI;�vI;X�I;u�I;W�I;�I;��I;��I;p�I;��I;�I;�I;
�I;c�I;��I;      �+I;�2I;�FI;�dI;��I;�I;��I;��I;m�I;/�I;��I;��I;�I;=�I;��I;]�I;�qI;�^I;�MI;?I;�1I;�&I;�I;TI;4I;(I;�I;��H;�H;��H;��H;��H;4�H;�H;*�H;��H;��H;��H;(�H;�H;5�H;��H;��H;��H;�H;��H;�I;/I;2I;PI;�I;�&I;�1I;?I;�MI;�^I;�qI;`�I;��I;=�I;�I;��I;��I;/�I;l�I;��I;��I;�I;ȇI;�dI;�FI;�2I;      ?�F;�F;S�F;8G;v�G;�.H;��H;I;�xI;O�I;��I;��I;`�I;b�I;��I;��I;��I;�|I;�fI;�SI;6CI;�4I;�(I;�I;�I;mI;*I;�I;p�H;��H;��H;��H;��H;��H;��H;��H;��H;��H;��H;��H;��H;��H;��H;��H;i�H;�I;,I;tI;�I;�I;�(I;�4I;3CI;�SI;�fI;�|I;��I;��I;��I;a�I;^�I;��I;��I;R�I;�xI;�I;��H;�.H;~�G;8G;9�F;�F;      Ĥ?;q�?;	v@;hA;a�B;��C;<BE;߄F;u�G;�H;�*I;̛I;4�I;��I;��I;�I;A�I;��I;\�I;�mI;�XI;HFI;6I;w)I;[I;�I;/I;�I;tI;/�H;��H;��H;��H;(�H;�H;i�H;/�H;i�H;�H;)�H;��H;��H;��H;2�H;mI;�I;2I;�I;YI;t)I;�6I;JFI;�XI;�mI;_�I;��I;B�I;�I;��I;��I;5�I;țI;�*I;�H;r�G;ބF;?BE;��C;l�B;hA;
v@;q�?;      f�0;o�0;K2;�_4;7;��9;X=;M@;��B;�E;A�F;.H;�I;F�I; �I;g�I;��I;��I;��I;��I;~rI;k[I;�GI;7I;q)I;�I;MI;�I;/I;� I;��H;��H;��H;��H;��H;�H;��H;�H;��H;��H;��H;��H;��H;� I;/I;�I;PI;�I;p)I;7I;�GI;n[I;�rI;��I;��I;��I;��I;j�I;��I;D�I;�I;.H;C�F;�E;��B;J@;\=;��9;/7;�_4;K2;Z�0;      &x;�b;~;�<;#�;ެ%;1,;$L2;�8;=;�9A;\oD;��F;WSH;�DI;"�I;��I;��I;:�I;�I;R�I;�tI;V\I;�GI;6I;�(I;�I;>I;�I;GI;B I;s�H;I�H;�H;��H;��H;��H;��H;��H;��H;L�H;s�H;H I;NI;�I;=I;�I;�(I;~6I;�GI;Z\I;�tI;U�I;�I;>�I;��I;��I;"�I;�DI;TSH;��F;[oD;�9A;=;�8;$L2;4,;߬%;"�;�<;};�b;      ��:؃�:̓�:�f�:���:���:}�;��;�#;�-;c�5;�L<;�gA;.E;lG;��H;�I;s�I;��I;z�I;øI;�I;�tI;q[I;HFI;�4I;�&I;0I;�I;M
I;hI;��H;
�H;s�H;��H;��H;f�H;��H;��H;q�H;�H;��H;nI;Q
I;�I;2I;�&I;�4I;GFI;v[I;�tI;�I;øI;|�I;��I;s�I;��I;��H;lG;/E;hA;�L<;f�5; -;�#;��;z�;���:Ǳ�:�f�:Ɠ�:���:       Sɸ��J�`%�8�'�9��:l�n:��:	W�:@��:�;��;��,;o�6;�>;5C;�F;vH;2wI;
�I;a�I;2�I;��I;O�I;�rI;�XI;*CI;�1I;%$I;�I;�I;�I;EI;;�H;0�H;��H;��H;s�H;��H;��H;*�H;=�H;BI;�I;�I;�I;'$I;�1I;0CI;�XI;�rI;Q�I;��I;6�I;e�I;�I;1wI;vH;�F;	5C;�>;o�6;��,;��; �;:��:W�:��:\�n:�:�'�9�&�8��J�      {+���%�X������1���U\�P�~���9��n:؉�:
b�:�;�#;��0;��:;��A;�E;�-H;�aI;��I;e�I;y�I;�I;��I;�mI;�SI;�>I;2.I;� I;QI;�I;]I;wI;��H;p�H;
�H;t�H;�H;l�H;��H;uI;]I;�I;TI;� I;2.I;?I;�SI;�mI;��I;�I;z�I;e�I;��I;�aI;-H;!�E;��A;��:;��0;�#;�;b�:҉�:��n:��9 �~��U\�v1�����[����%�      �ݻ��ػ��ʻnT��Ԓ��U�s���0�pTܺ��=� T94f:��:��;>;%,;�e8;qv@;"]E;*H;�aI;�I;��I;:�I;��I;U�I;�fI;�MI;�9I;�)I;fI;mI;�I;0I;I;G�H;{�H;��H;}�H;D�H;I;2I;�I;qI;iI;�)I;�9I;�MI;�fI;R�I;��I;;�I;��I;�I; bI;,H;!]E;rv@;�e8;#,;>;��;��:@f:0T9��=�lTܺ��0�U�s�Ԓ��lT����ʻ��ػ      ��\�$�X�-M���:��G#�V����ػ^7��FZ�:���"/���9��:�m�:�e;r�(;�7;�@;]E;}-H;.wI;t�I;��I;��I;��I;�|I;�^I;�FI;�3I;G%I;�I;�I;C
I;?I; I;* I;q�H;, I;I;<I;F
I;�I;�I;L%I;�3I;�FI;�^I;�|I;��I;��I;��I;s�I;.wI;�-H;!]E;�@;�7;q�(;�e;�m�:��:��9"/�:���FZ�^7����ػX���G#���:��-M�$�X�      ��ƼNü9_���۩�+$��@���Q�UG#��9�����G��3����ȸ��n:el�:n�;�';�7;nv@;�E;vH;�I;��I;��I;=�I;}�I;�qI;mUI;-?I;�-I;z I;I;kI;�I;BI;�I;I;�I;?I;�I;jI;I;} I;�-I;-?I;pUI;�qI;�I;:�I;��I;��I;�I;vH;!�E;ov@;�7;�';m�;el�:��n:��ȸ�3����G�����9�TG#��Q�@��,$���۩�:_��Nü      �)���&�I<��3��� ��zܼ�*��琼��\�@ �D�ػz� N���Ϲ4�J:tj�:f�;o�(;�e8;��A;�F;��H; �I;g�I;�I;��I;X�I;ZeI;�KI;7I;�'I;�I;I;�I;aI;�I;'I;�I;^I;�I;I;�I;�'I;7I;�KI;\eI;[�I;��I;��I;i�I; �I;��H;�F;��A;�e8;n�(;g�;nj�:0�J:��Ϲ!N�{�E�ػ@ ���\�琼�*���zܼ�� ��3�J<���&�      }L��>ى��Ă�8�o�
+T���5��G��V��^���Y����A� c �V���������<�J:_l�:�e;,;��:;	5C;lG;�DI;��I;��I;��I;��I;�vI;�XI;CAI;�/I;"I;�I;�I;�I;�I;HI;�I;�I;�I;�I;"I;�/I;BAI;�XI;�vI;��I;��I;��I;�I;�DI;lG; 5C;��:;,;�e;_l�:0�J:������V��� c ���A��Y���^���V��G���5�+T�9�o��Ă�>ى�      	3�`�Խ�������.W��1�o�h??�4��8zܼ|Q��4�X��Q��6�������Ϲ��n:�m�:>;��0;�>;/E;NSH;H�I;��I;]�I;;�I;T�I;�fI;#LI;�7I;b(I;	I;�I;]I;I;>I; I;\I;�I;I;a(I;�7I;%LI;�fI;U�I;;�I;Z�I;��I;K�I;USH;/E;�>;��0;>;�m�:��n:��Ϲ����6���Q�4�X�|Q��8zܼ4��h??�2�o�.W���������Խ`�      �7�|74�o�)�#>����3�k���/7nc���)������ک�va��Q�T���N���ȸ��:��;�#;t�6;hA;��F;�I;8�I;Z�I;�I;s�I;�uI;nWI;s@I;	/I;b"I;I;�I;gI;[I;gI;�I;I;d"I;/I;s@I;nWI;�uI;u�I;�I;Y�I;2�I;�I;��F;hA;i�6;�#;��;��:`�ȸN�T����Q�wa��ک�������)�7nc�/k���3����#>�o�)�|74�      �S���7���X��W�s��_S��0����W�{���·|�i�5�i���ک�4�X� c �z��3����9��:�;�,;�L<;VoD;.H;śI;��I;��I;P�I;Q�I;6cI;^II;�5I;�'I;JI;�I;�I;�I;�I;�I;II;�'I;�5I;[II;6cI;T�I;Q�I;��I;��I;��I;.H;[oD;�L<;��,;�;��:��9�3��{� c �5�X��ک�i��i�5�·|�{���Wར��~�0��_S�W�s��X���7��      D���s�YD־�t��p���X��x�W�,�&��l��!N���Ă�i�5�����|Q����A�E�ػ��G�$"/�f:�a�:��;b�5;�9A;D�F;�*I;��I;��I;�I;\�I;/oI;iRI;�<I;-I;�!I;@I;I;�I;I;@I;�!I;-I;�<I;fRI;-oI;^�I;	�I;��I;��I;�*I;G�F;�9A;_�5;��;�a�:f:("/���G�E�ػ��A�|Q������i�5��Ă�!N���l��,�&�y�W��X��p���t��YD־�s�      ��7�r�3��'��K�'�����̾#���W�s�o74����!N��·|���)�8zܼ�Y��? ����H����S9։�:"�; -;=;�E;�H;H�I;,�I;��I;��I;{I;a[I;�CI;V2I;&I;�I;*I;�I;*I;�I;&I;V2I;�CI;`[I;{I;��I;��I;,�I;H�I;��H;�E;=;�-;�;؉�:�S9L������@ ��Y��8zܼ��)�·|�!N�����o74�W�s�#�����̾'����K��'�r�3�      &8��iڇ��x|�qm_�Fv<����?��l8��$6~�o74��l��{���7nc�4���^����\��9�NZ���=���n:H��:�#;�8;��B;u�G;�xI;l�I;��I;��I;܆I;:dI;uJI;�7I;*I;2!I;MI;�I;LI;4!I;*I;�7I;uJI;4dI;نI;��I;��I;l�I;�xI;t�G;��B;�8;�#;4��:��n:��=�MZ��9���\��^��4��7nc�{����l��o74�$6~�l8��@�꾎��Fv<�qm_��x|�iڇ�       �ȿ�ÿ���+8��hڇ�Z��'�����l8��W�s�,�&�X�/i??��V�琼WG#�f7��~Tܺh�9W�:��;L2;P@;߄F;�I;��I;o�I;P�I;A�I;�lI;�PI;Z<I;�-I;�$I;!I;DI;!I;�$I;�-I;Z<I;�PI;�lI;C�I;P�I;r�I;��I;�I;ބF;P@;L2;��;W�:��9�Tܺd7��VG#�琼�V�i??�/X�,�&�W�s�l8�������'�Z�hڇ�+8������ÿ      ��	�%X�M����,ݿI����ҕ��d��'�@��#���x�W����k���2�o��G��*���Q���ػ�0�p�~���:{�;-,;`=;7BE;��H;{�I;��I;F�I;�I;atI;�VI;�@I;�1I;�'I;�!I;�I;�!I;�'I;�1I;�@I;�VI;^tI;�I;E�I;��I;~�I;��H;7BE;c=;3,;w�;��:P�~��0���ػ�Q��*���G�2�o�k������x�W�#���@�꾌'��d��ҕ�I����,ݿM���%X�      �5�621���#�N��r���ÿ�ҕ�Z������̾�X���0�3�.W����5��zܼ@��Z��a�s��U\�h�n:���:ج%;��9;��C;�.H;�I;�I;�I;��I;x{I;
\I;�DI;�4I;'*I;$I;"I;$I;(*I;�4I;�DI;\I;t{I;��I;�I;�I;�I;�.H;��C;��9;۬%;���:L�n:�U\�d�s�Z��A���zܼ��5�.W��3��0��X����̾���Z��ҕ��ÿr��N����#�621�      /�j���c�x�P��5���s��I���hڇ�Fv<�(���p���_S��������+T��� �+$���G#�ђ��n1���:���:1�;-7;q�B;v�G;��I;�I;c�I;ȮI;��I;�`I;FHI;�7I;],I;&I;�#I;&I;a,I;�7I;IHI;�`I;��I;ʮI;c�I;�I;I;��G;o�B;07;1�;���:�:l1��Ғ���G#�,$���� �+T���������_S�p��(���Fv<�hڇ�I���s�����5�x�P���c�      Т��^���F���/]��5�N���,ݿ+8��qm_��K��t��W�s�#>����9�o��3��۩���:�nT����� (�9�f�:�<;�_4;hA;8G;udI;�I;)�I;W�I;_�I;#dI;KI;�9I;G.I;�'I;�%I;�'I;H.I;�9I;KI;&dI;[�I;[�I;'�I;�I;wdI;8G;	hA;�_4;�<;�f�:�'�9���pT����:��۩��3�9�o����#>�W�s��t���K�qm_�+8���,ݿN���5��/]�F��^���      �����B����F��x�P���#�M�������x|��'�YD־�X��o�)�Խ�Ă�J<�8_��~-M���ʻ[��`&�8�:�;K2;v@;K�F;�FI;g�I; �I;'�I;��I;�fI;;MI;@;I;�/I;�(I;�&I;�(I;�/I;@;I;<MI;�fI;��I;(�I;��I;k�I;�FI;X�F;v@;K2;�;���:�%�8X����ʻ~-M�8_��J<��Ă�Խo�)��X��YD־�'��x|����M�����#�x�P�F�����B��      ��������B��^�����c�621�%X��ÿiڇ�r�3��s��7��|74�a�>ى���&�Nü(�X���ػ��%���J�ă�:�b;y�0;r�?;�F;�2I;��I;6�I;�I;E�I;OhI;�NI;0<I;y0I;_)I;�'I;\)I;y0I;0<I;�NI;QhI;A�I;�I;6�I;��I;�2I;�F;q�?;w�0;�b;���:��J���%���ػ(�X�Nü��&�>ى�a�|74��7���s�r�3�iڇ��ÿ%X�621���c�^����B�����      D(��r'���o��N�d��X1�~x�	Ŀ����3�x���x����4�l��Z+���'���ü;yY��kٻp&���p�H��:8;��0;��?;��F;g I;��I;��I;+�I;h�I;LdI;�KI;�9I;k.I;�'I;�%I;�'I;k.I;�9I;�KI;LdI;d�I;.�I;��I;��I;f I;ɀF;��?;��0;2;@��:@�p�p&��kٻ;yY���ü�'�Z+��l�ཽ�4��x��x���3����	Ŀ~x��X1�d�N��o��r'��      q'���X��e^�������]]���,�P9�6g��U�����/����o��g1��hܽ���-$�`l���|U�h�Ի�!� �,�u�:�;�51;��?;2�F;?'I;`�I;
�I;<�I;��I;�cI;>KI;x9I;.I;{'I;�%I;v'I; .I;w9I;>KI;�cI;��I;?�I;
�I;b�I;='I;?�F;��?;~51;�;k�: �,��!�j�Ի�|U�_l���-$����hܽg1��o���ྙ�/�U���6g��P9���,��]]�����e^���X��      �o��e^���ē��4z�5K�h��R��'ﱿU�v��X#���Ѿń��&�o�нc̀�_��v���K�I��ǻ�4�P"9��:4�;�2;��@;��F;�:I;��I;��I;��I;v�I;KbI;�II;�8I;Z-I;�&I;�$I;�&I;Z-I;�8I;�II;JbI;o�I;��I;��I;��I;�:I;��F;��@;�2;.�;��:�!9�4��ǻL�I�v���_��c̀�o�н�&�ń���Ѿ�X#�U�v�'ﱿR��h��5K��4z��ē�e^��      N������4z���V��X1��<�uؿ����RZ��	�(���HUo����^y��-l�Z��R��D�7�������ų9���:��;X�4;itA;\2G;�XI;��I;J�I;�I;�I;�_I;�GI;"7I;�+I;�%I;�#I;�%I;�+I;7I;�GI;�_I;�I;�I;J�I;��I;�XI;e2G;gtA;U�4;��;���:�ų9�����D�7��R��Z�-l�^y�����HUo�(����	��RZ����uؿ�<��X1���V��4z�����      d��]]�5K��X1�Zf��nQ��T���[58��A���נ���O���`什�Q����@ߓ��� ��V���氺��":Ҹ�: ;�07;�B;.�G;�{I;��I;��I;��I;8|I;7\I;JEI;5I;3*I;1$I;)"I;.$I;5*I;5I;LEI;5\I;3|I;��I;��I;��I;�{I;5�G;�B;�07;� ;̸�:܌":�氺�V���� �@ߓ�����Q�`什����O��נ��A��[58�T���nQ���Zf��X1�5K��]]�      �X1���,�h���<��5g��e_���U�͂�֌Ⱦ	ń�*�-�j��P ��&�2�?ټb�{�"��n�,�O���u:�P ;�&;)#:;<�C;�%H;�I;!�I;��I;�I;\vI;�WI;�AI;z2I;(I;D"I;^ I;@"I;(I;u2I;�AI;�WI;YvI;�I;��I;$�I;�I;�%H;<�C;$#:;�&;�P ;t�u:,�O��n�"�b�{�?ټ&�2�P ��j��*�-�	ń�֌Ⱦ͂��U�e_��5g��<�h����,�      ~x�P9�R��uؿnQ��e_��6�_��X#�r���f��9�S�{�����l�B�	w�� �M���Ի��+�`=T���:�e;�\,;�/=;�BE;P�H;z�I;��I;��I;��I;�oI;�RI;>I;\/I;~%I;�I;DI;�I;~%I;\/I;>I;�RI;�oI;��I;��I;��I;v�I;W�H;�BE;�/=;�\,;�e;��:0=T���+���Ի �M�	w��B�l�����{�9�S��f��r���X#�6�_�e_��nQ��uؿR��P9�      	Ŀ6g��'ﱿ���T����U��X#�t��d���HUo��#��hܽ����n<����=����� ��᝻J�Ժht�9`��:�V;ˇ2;� @;R�F;�I;��I;A�I;(�I;i�I;�gI;MI;�9I;�+I;�"I;jI;�I;hI;�"I;�+I;�9I;MI;�gI;k�I;(�I;D�I;��I;�I;U�F;� @;̇2;�V;R��:�t�9L�Ժ�᝻�� �=�������n<�����hܽ�#�HUo�d���t���X#��U�T������'ﱿ6g��      ���U���U�v��RZ�[58�͂�q��d���foy�]1�_O��]什�`�M�����pyY�%�컘�T��1�l�u:���:F#;98;�B;f�G;�lI;�I; �I;-�I;t�I;�_I;GI;�4I;#(I;�I;�I;I;�I;�I;#(I;�4I;GI;�_I;v�I;.�I;�I;�I;�lI;j�G;�B;98;E#;���:��u:�1���T�$��pyY����M���`�\什_O��]1�foy�d���q��͂�[58��RZ�U�v�U���      �3���/��X#��	��A��֌Ⱦ�f��GUo�^1�˰��|n��Լx��'��>ټ�@���k�м�� ���39�#�:.R;	e-;�/=;�	E;ZxH;��I;�I;o�I;��I;vI;aWI;�@I;�/I;#$I;<I;�I;7I;�I;<I;#$I;�/I;�@I;cWI;vI;�I;q�I;�I;}�I;]xH;�	E;�/=;e-;*R;�#�:��39(��μ���k��@���>ټ�'�Լx�|n��˰��^1�GUo��f��֌Ⱦ�A���	��X#���/�      w���ྃ�Ѿ(����נ�ń�9�S��#�`O��|n��J̀���2���𛼄�>��Ի��B��#�,m:�G�:\ ;��5;�FA;��F;�I;P�I;S�I;��I;h�I;kjI;�NI;:I;�*I;�I;�I;�I;II;�I;�I;�I;�*I;:I;�NI;pjI;m�I;��I;S�I;K�I;�I;��F;�FA;��5;[ ;�G�:4m:�#���B��Ի��>�������2�J̀�|n��_O���#�9�S�ń��נ�(�����Ѿ��      �x���o��ń�HUo���O�*�-�{��hܽ]什Լx���2�tb��VR��X|U�]2��:��*갺�u�9��:D;��,;�h<;`rD;N%H;��I;g�I;��I;�I;�I;�^I;FI;W3I;�%I;�I;_I;iI;4I;hI;\I;�I;�%I;R3I;FI;�^I;
�I;�I;��I;c�I;ďI;M%H;erD;�h<;��,;D;��:xu�9갺:��^2��W|U�UR��tb����2�Լx�\什�hܽ{�*�-���O�HUo�ń��o��      ��4�g1��&������j�ཅ�������`��'���UR��F�]�~��!V���X�� Io����:h�;$#;�6;QtA;P�F;�	I;t�I;��I;p�I;�I;�pI;�SI;�=I;�,I;w I;�I;�I;GI;;I;GI;�I;�I;w I;�,I;�=I;�SI;�pI;�I;n�I;��I;x�I;�	I;Q�F;UtA;�6;.#;j�;���:@Ho��X��!V��~��F�]�UR����'��`��������j��������&�g1�      k�ྲྀhܽn�н^y��`什P ��l��n<�M���>ټ��X|U���������1�������u:Sl�:�;a71;R)>;S	E;JH;U�I;��I;��I;�I;փI;XbI;�HI;$5I;c&I;gI;qI;<I;#I;
I;#I;:I;qI;eI;_&I;*5I;�HI;_bI;ڃI;�I;��I;��I;R�I;
JH;V	E;R)>;i71;�;Kl�:��u:�����1��������W|U����>ټM���n<�l�P ��`什^y��n�н�hܽ      Y+����c̀�,l��Q�%�2�B��������@����>�^2��"V���1�����#R:���:�;v\,;3;;�;C;�eG;W9I;��I;-�I;��I;C�I;�qI;�TI;`>I;5-I;1 I;zI;qI;�
I;I;I;I;�
I;qI;zI;. I;9-I;d>I;�TI;�qI;B�I;��I;1�I;��I;T9I;�eG;�;C;;;;y\,;�;���:�#R:ȑ�1�!V��\2����>��@��������B�$�2��Q�-l�c̀���      �'��-$�_��Y����?ټw��<���pyY��k� �Ի<��Y�������#R:���:�R;�);܍8;��A;��F;3�H;'�I;��I;��I;��I;�I;�`I;�GI;�4I;�%I;JI;�I;�I;oI;I;EI;I;mI;�I;�I;FI;�%I;�4I;�GI;�`I;�I;��I;��I;��I;&�I;6�H;��F;��A;ݍ8;�);�R;���:�#R:����Y��:�� �Ի�k�pyY�<���	w��
?ټ���Y�_���-$�      ��ü^l��w����R��?ߓ�b�{��M��� � ��˼����B�갺�Ho���u:���:�R;/�';17;��@;��E;�lH;.�I;h�I;��I;�I;v�I;�lI;�QI;&<I;�+I;�I;�I;eI;�I;EI;0I;�I;,I;AI;�I;bI;�I;�I;�+I;%<I;�QI;�lI;p�I;�I;��I;d�I;/�I;�lH;��E;��@;17;/�';�R;���:��u: Io�갺��B�̼��"�컋� ��M�b�{�@ߓ��R��x���]l��      4yY��|U�K�I�@�7��� �"���Ի�᝻��T����#��u�9���:Ql�:�;�);17;/ @;:]E;�$H;ekI;
�I;U�I;��I;'�I;�wI;�ZI;�CI;w1I;N#I;%I;�I;-	I;rI;8I;m�H;��H;j�H;4I;pI;*	I;�I;)I;P#I;v1I;�CI;�ZI;�wI;-�I;��I;N�I;
�I;ekI;�$H;;]E;+ @;17;�);�;Ol�:���:�u�9�#����T��᝻��Ի"��� �B�7�J�I��|U�      �kٻm�Ի�ǻ����V���n���+�8�Ժ��1��39Tm:��:j�;
�;z\,;�8;��@;?]E;�
H;JVI;q�I;��I;��I;c�I;��I;�bI;`JI;%7I;�'I;�I;,I;�
I;8I;;I;i�H;��H;z�H;��H;d�H;6I;6I;�
I;/I;�I;�'I;&7I;_JI;�bI; �I;e�I;��I;��I;r�I;LVI;�
H;8]E;��@;ݍ8;y\,;	�;j�;��:\m:�39�1�6�Ժ��+��n��V������ǻl�Ի      !p&��!��4���氺�O��<T�Xt�9��u:�#�:�G�:D;)#;h71;;;;��A;��E;�$H;JVI;�I;��I;�I;��I;��I;iI;)PI;<I;�+I;I;�I;�I;�I;�I;2�H;��H;��H;�H;��H;��H;0�H;�I;�I;�I;�I;I;�+I;<I;%PI;iI;��I;}�I;�I;��I;�I;MVI;�$H;��E;��A;:;;d71;&#;D;�G�:�#�:��u:�t�9�<T��O��氺���4��!�      @�p� �,�� 9�ų9��":��u:��:b��:���:.R;\ ;��,;�6;S)>;�;C;��F;�lH;kkI;r�I;��I;��I;�I;r�I;�mI;wTI;&@I;�/I;!"I;WI;�I;�I;�I;r�H;r�H;��H;V�H;��H;O�H;��H;q�H;r�H;�I;�I;�I;SI;$"I;�/I;"@I;|TI;�mI;i�I;�I;��I;��I;r�I;ekI;�lH;��F;�;C;O)>;�6;��,;^ ;,R;���:T��:��:p�u:�":�ų9`!9 �,�      8��:��:�:��:���:�P ;�e;�V;J#;e-;��5;�h<;StA;X	E;�eG;7�H;1�I;�I;��I;�I;�I;�I;pI;LWI;�BI;@2I;�$I;qI;lI;@	I;rI;��H;��H;�H;Y�H;3�H;��H;.�H;V�H;�H;��H;��H;vI;@	I;kI;sI;�$I;A2I;�BI;IWI;�oI;�I;�I;�I;��I;�I;1�I;4�H;�eG;S	E;QtA;�h<;��5;e-;J#;�V;�e;�P ;��:���:��:{�:      I;�;.�;��;� ;�&;�\,;ه2;98;�/=;�FA;nrD;T�F;JH;Y9I;-�I;k�I;W�I;��I;��I;p�I;pI;HXI;�DI;�3I;\&I;I;�I;
I;nI;��H;��H;��H;��H;9�H;H�H;
�H;B�H;6�H;��H;��H;��H;��H;lI;z
I;�I;I;\&I;�3I;�DI;AXI;pI;p�I;~�I;��I;P�I;k�I;*�I;W9I;JH;Q�F;krD;�FA;�/=;98;և2;�\,;�&; ;��;(�;�;      ��0;�51;�2;R�4;�07;-#:;�/=;� @;�B;�	E;��F;M%H;�	I;U�I;��I;��I;��I;��I;c�I;��I;�mI;BWI;�DI;�4I;;'I;-I;�I;|I;8I;- I;*�H;��H;z�H;��H;c�H;��H;g�H;��H;`�H;��H;z�H;��H;.�H;, I;4I;{I;�I;.I;@'I;�4I;~DI;EWI;�mI;��I;`�I;��I;��I;��I;��I;N�I;�	I;N%H;��F;�	E;�B;� @;�/=;#:;�07;P�4;�2;�51;      ��?;��?;��@;_tA;��B;F�C;�BE;W�F;j�G;`xH;�I;ˏI;u�I;��I;4�I;��I;�I;1�I;�I;iI;�TI;�BI;�3I;G'I;�I;}I;I;�I;� I;}�H;�H;j�H;`�H;��H;��H;+�H;��H;&�H;��H;��H;^�H;d�H;�H;}�H;� I;�I;I;}I;�I;A'I;�3I;�BI;�TI;iI;�I;+�I;�I;��I;3�I;��I;u�I;͏I;�I;_xH;h�G;R�F;�BE;<�C;�B;`tA;��@;��?;      ��F;@�F;��F;Y2G;%�G;�%H;Y�H;�I;�lI;��I;T�I;p�I;��I;��I;��I;��I;x�I;�wI;�bI;&PI;'@I;:2I;[&I;1I;{I;8I;I;� I;��H;C�H;w�H;T�H;z�H;&�H;Z�H;��H;��H;��H;X�H;$�H;|�H;P�H;w�H;B�H;��H;� I;I;;I;}I;-I;X&I;=2I;&@I;#PI;�bI;�wI;z�I;��I;��I;��I;��I;m�I;X�I;��I;�lI;�I;Z�H;�%H;:�G;m2G;��F;B�F;      r I;K'I;�:I;�XI;�{I;�I;~�I;�I;�I;�I;U�I;��I;j�I;�I;@�I;�I;�lI;�ZI;cJI;<I;�/I;�$I;!I;I;I;I;I;��H;s�H;��H;J�H;T�H;��H;��H;�H;��H;n�H;��H;�H;��H;��H;O�H;J�H;��H;m�H;��H;I;I;I;�I;I;�$I;�/I;<I;`JI;�ZI;�lI;�I;?�I;�I;j�I;��I;U�I;�I;�I;��I;w�I;�I;�{I;�XI;�:I;3'I;      ��I;f�I;��I;��I;��I;"�I;��I;C�I;�I;t�I;��I;�I;�I;݃I;�qI;�`I;�QI;�CI;#7I;�+I;'"I;mI;�I;|I;�I;� I;��H;l�H;��H;T�H;R�H;��H;��H;��H;��H;��H;m�H;��H;��H;��H;��H;��H;R�H;S�H;��H;h�H;��H;� I;�I;yI;�I;oI;$"I;�+I;"7I;�CI;QI;�`I;�qI;ڃI;�I;�I;��I;t�I; �I;A�I;��I;�I;��I;��I;��I;\�I;      ��I;��I;��I;[�I;��I;��I;��I;-�I;'�I;�I;n�I;�I;�pI;`bI;�TI;�GI;*<I;z1I;�'I;I;^I;gI;{
I;5I;� I;��H;m�H;��H;P�H;N�H;��H;O�H;=�H;�H;��H;��H;~�H;��H;��H;��H;@�H;K�H;��H;K�H;L�H;��H;i�H;��H;� I;1I;z
I;gI;YI;I;�'I;v1I;)<I;�GI;�TI;]bI;�pI;�I;r�I;�I;*�I;,�I;��I;��I;��I;]�I;��I;��I;      .�I;<�I;��I;�I;��I;ߟI;��I;p�I;w�I;vI;rjI;�^I;�SI;�HI;b>I;�4I;�+I;K#I;�I;�I;�I;<	I;lI;, I;~�H;=�H;��H;W�H;T�H;��H;)�H;�H;6�H;��H;�H;��H;��H;��H;�H;��H;5�H;�H;)�H;��H;Q�H;V�H;��H;?�H;��H;) I;kI;=	I;�I;�I;�I;H#I;�+I;�4I;b>I;�HI;�SI;�^I;tjI;vI;v�I;l�I;��I;�I;��I;�I;��I;<�I;      d�I;��I;w�I;��I;4|I;\vI;�oI;hI;�_I;jWI;�NI;FI;�=I;.5I;<-I;�%I;�I;'I;0I;�I;�I;tI;��H;-�H;�H;u�H;M�H;Y�H;��H;/�H;	�H;�H;S�H;��H;t�H;,�H;��H;)�H;r�H;��H;T�H;�H;�H;)�H;��H;V�H;I�H;u�H;�H;*�H;��H;uI;�I;�I;/I;&I;�I;�%I;<-I;+5I;�=I;FI;�NI;kWI;�_I;hI;�oI;VvI;<|I;��I;v�I;��I;      MdI;�cI;CbI;�_I;'\I;�WI;�RI;MI;GI;�@I;:I;\3I;�,I;g&I;1 I;JI;�I;�I;�
I;�I;�I;��H;��H;��H;k�H;M�H;Q�H;��H;S�H;�H;�H;M�H;��H;"�H;��H;��H;��H;��H;��H;#�H;��H;L�H;�H;�H;L�H;��H;O�H;M�H;m�H;��H;��H;��H;�I;�I;�
I;�I;�I;MI;3 I;g&I;�,I;Y3I;:I;�@I;GI;MI;�RI;�WI;1\I;�_I;NbI;�cI;      �KI;LKI;�II;�GI;GEI;�AI;>I;�9I;�4I;�/I;�*I;�%I;y I;jI;|I;�I;iI;+	I;<I;�I;�H;��H;��H;w�H;a�H;t�H;��H;��H;H�H;;�H;Q�H;��H;�H;��H;G�H;�H;,�H;�H;F�H;��H;�H;��H;O�H;2�H;C�H;��H;��H;t�H;b�H;t�H;��H;��H;w�H;�I;<I;-	I;jI;�I;~I;jI;w I;�%I;�*I;�/I;�4I;�9I;>I;�AI;LEI;�GI;JI;LKI;      �9I;w9I;�8I;7I;5I;j2I;Z/I;�+I;%(I;,$I; I;�I;�I;xI;xI;�I;�I;pI;<I;6�H;|�H;�H;��H;��H;��H; �H;��H;��H;��H;��H;��H;&�H;��H;5�H;��H;��H;��H;��H;��H;6�H;��H;%�H;��H;��H;~�H;��H;��H;�H;��H;��H;��H; �H;t�H;/�H;<I;sI;�I;�I;xI;vI;�I;�I; I;,$I;&(I;�+I;d/I;j2I;5I;7I;�8I;�9I;      ].I;9.I;^-I;�+I;<*I;(I;%I;�"I;�I;HI;�I;jI;�I;DI;�
I;tI;II;6I;j�H;��H;��H;V�H;5�H;V�H;��H;P�H;�H;��H;��H;�H;o�H;��H;G�H;��H;��H;��H;z�H;��H;��H;��H;H�H;��H;m�H;�H;��H;��H;�H;P�H;��H;U�H;6�H;S�H;��H;��H;i�H;8I;JI;uI;�
I;DI;�I;jI;�I;II;�I;�"I;�%I;(I;9*I;,I;\-I;:.I;      �'I;�'I;�&I;�%I;#$I;="I;�I;pI;�I;�I;�I;oI;JI;(I;I;I;0I;g�H;��H;��H;]�H;.�H;A�H;��H;'�H;��H;��H;��H;��H;��H;,�H;��H;�H;��H;��H;a�H;o�H;c�H;��H;��H;�H;��H;)�H;��H;��H;��H;��H;��H;&�H;��H;E�H;.�H;V�H;��H;��H;j�H;2I;I;I;*I;JI;oI;�I;�I;�I;lI; I;?"I;%$I;�%I;�&I;�'I;      �%I;�%I;�$I;�#I;"I;V I;GI;�I;I;6I;UI;>I;=I;"
I;I;FI;�I;��H;}�H;	�H;��H;��H;�H;\�H;��H;��H;j�H;s�H;��H;��H;��H;��H;.�H;��H;z�H;i�H;s�H;l�H;w�H;��H;0�H;��H;��H;��H;}�H;m�H;k�H;��H;��H;[�H;
�H;��H;��H;�H;}�H;��H;�I;JI;I;'
I;?I;<I;YI;7I;I;�I;MI;W I;"I;�#I;�$I;�%I;      �'I;�'I;�&I;�%I;#$I;@"I;�I;oI;�I;�I;�I;oI;JI;(I;I;I;/I;e�H;��H;��H;^�H;/�H;?�H;��H;'�H;��H;��H;��H;��H;��H;*�H;��H;�H;��H;��H;a�H;o�H;c�H;��H;��H;�H;��H;)�H;��H;��H;��H;��H;��H;&�H;��H;E�H;,�H;T�H;��H;��H;j�H;0I;I;I;)I;HI;oI;�I;�I;�I;mI;�I;@"I;%$I;�%I;�&I;�'I;      U.I;:.I;Z-I;�+I;<*I;(I;%I;�"I;�I;HI;�I;jI;�I;AI;�
I;tI;HI;6I;j�H;��H;��H;U�H;2�H;S�H;��H;O�H;�H;��H;��H;�H;m�H;��H;G�H;��H;��H;��H;z�H;��H;��H;��H;J�H;��H;m�H;�H;��H;��H;�H;S�H;��H;U�H;6�H;U�H;��H;��H;i�H;8I;JI;uI;�
I;DI;�I;mI;�I;HI;�I;�"I;�%I;
(I;<*I;,I;^-I;=.I;      �9I;x9I;�8I;7I;5I;p2I;Z/I;�+I;&(I;*$I; I;�I;�I;uI;xI;�I;�I;sI;<I;5�H;{�H;�H;��H;��H;��H;�H;��H;��H;��H;��H;��H;%�H;��H;5�H;��H;��H;��H;��H;��H;5�H;��H;%�H;��H;��H;~�H;��H;��H; �H;��H;��H;��H;�H;o�H;0�H;=I;rI;�I;�I;yI;xI;�I;�I; I;,$I;&(I;�+I;e/I;p2I;5I;7I;�8I;{9I;      �KI;RKI;�II;�GI;FEI;�AI;>I;�9I;�4I;�/I;�*I;�%I;v I;hI;I;�I;hI;+	I;9I;�I;�H;��H;��H;t�H;b�H;q�H;��H;��H;J�H;9�H;O�H;��H;�H;��H;H�H;�H;,�H;�H;F�H;��H;�H;��H;O�H;4�H;@�H;��H;��H;u�H;a�H;r�H;��H;��H;t�H;�I;<I;+	I;iI;�I;~I;jI;z I;�%I;�*I;�/I;�4I;�9I;>I;�AI;JEI;HI;JI;OKI;      BdI;�cI;7bI;�_I;)\I;�WI;�RI;MI;GI;�@I;:I;Z3I;�,I;d&I;3 I;JI;�I;�I;�
I;�I;�I;��H;��H;��H;m�H;L�H;O�H;��H;U�H;�H;�H;M�H;��H;!�H;��H;��H;��H;��H;��H;#�H;��H;L�H;�H;�H;O�H;��H;O�H;O�H;j�H;��H;��H;��H;�I;�I;�
I;�I;�I;NI;3 I;g&I;�,I;\3I;:I;�@I;GI;MI;�RI;�WI;)\I;�_I;?bI;�cI;      Z�I;��I;w�I;��I;8|I;\vI;�oI;hI;�_I;eWI;�NI;FI;�=I;+5I;;-I;�%I;�I;'I;/I;�I;�I;uI;��H;*�H;�H;q�H;J�H;V�H;��H;,�H;�H;�H;T�H;��H;v�H;*�H;��H;-�H;r�H;��H;T�H;�H;�H;)�H;��H;T�H;I�H;u�H;�H;'�H;��H;vI;�I;�I;2I;'I;�I;�%I;=-I;.5I;�=I;FI;�NI;gWI;�_I;
hI;�oI;YvI;B|I;�I;|�I;��I;      3�I;A�I;��I;�I;��I;�I;��I;p�I;w�I;vI;kjI;�^I;�SI;�HI;c>I;�4I;�+I;L#I;�I;�I;�I;=	I;hI;) I;��H;;�H;��H;W�H;T�H;��H;)�H;�H;5�H;��H;�H;��H;��H;��H;�H;��H;6�H;�H;)�H;��H;O�H;T�H;��H;?�H;}�H;& I;pI;=	I;�I;�I;�I;H#I;�+I;�4I;c>I;�HI;�SI;�^I;rjI;vI;v�I;p�I;��I;ޟI;��I;�I;��I;9�I;      ��I; �I;��I;Q�I;��I;��I;��I;+�I;.�I;��I;j�I;
�I;�pI;]bI;�TI;�GI;'<I;z1I;�'I;I;^I;gI;w
I;4I;� I;��H;i�H;��H;O�H;K�H;��H;R�H;?�H;�H;��H;��H;~�H;��H;��H;�H;@�H;O�H;��H;M�H;J�H;��H;i�H;��H;� I;.I;~
I;hI;ZI;I;�'I;v1I;'<I;�GI;�TI;\bI;�pI;�I;q�I;��I;*�I;/�I;��I;��I;��I;T�I;��I;��I;      �I;\�I;��I;��I;��I;,�I;��I;G�I; �I;s�I;��I;�I;�I;ڃI;�qI;�`I;QI;�CI;!7I;�+I;'"I;pI;�I;|I;�I;� I;��H;h�H;��H;Q�H;T�H;��H;}�H;��H;��H;��H;o�H;��H;��H;��H;��H;��H;T�H;S�H;��H;f�H;��H;� I;�I;xI;�I;pI;!"I;�+I;%7I;�CI;�QI;�`I;�qI;ڃI;�I;	�I;��I;w�I;�I;A�I;��I;�I;��I;��I;��I;\�I;      a I;N'I;�:I;�XI;�{I;�I;x�I;�I;�I;�I;Q�I;��I;g�I;�I;B�I;�I;�lI;�ZI;_JI;<I;�/I;�$I;I;I;I;I;I;��H;s�H;��H;I�H;U�H;��H;��H;�H;��H;n�H;��H;�H;��H;��H;T�H;L�H;��H;o�H;��H;I;I;I;�I;!I;�$I;�/I;<I;cJI;�ZI;�lI;�I;B�I;�I;i�I;��I;T�I;�I;�I;�I;�I;�I;�{I;�XI;�:I;:'I;      ��F;>�F;��F;Y2G;*�G;&H;T�H;�I;�lI;��I;R�I;q�I;��I;��I;��I;��I;t�I;�wI;�bI; PI;'@I;:2I;U&I;.I;|I;3I;I; I;��H;@�H;w�H;V�H;z�H;&�H;[�H;��H;��H;��H;X�H;&�H;{�H;T�H;z�H;C�H;��H;� I;I;8I;{I;,I;Y&I;<2I;&@I;%PI;�bI;�wI;z�I;��I;��I;��I;��I;l�I;W�I;��I;�lI;�I;Y�H;�%H;4�G;^2G;��F;4�F;      ��?;��?;�@;`tA;��B;J�C;�BE;T�F;j�G;_xH;�I;ˏI;r�I;��I;6�I;��I;�I;.�I;�I;iI;~TI;�BI;�3I;B'I;�I;vI;I;�I;� I;z�H;�H;k�H;]�H;��H;��H;*�H;��H;*�H;��H;��H;`�H;j�H;�H;|�H;� I;�I;I;|I;�I;B'I;�3I;�BI;�TI;iI;�I;+�I;�I;��I;7�I;��I;v�I;ʏI;�I;_xH;f�G;R�F;�BE;<�C; �B;`tA;��@;��?;      ��0;t51;�2;X�4;�07;4#:;�/=;� @;�B;�	E;��F;M%H;	I;N�I;��I;��I;��I;��I;_�I;�I;�mI;BWI;}DI;�4I;>'I;&I;�I;{I;8I;) I;-�H;��H;z�H;��H;c�H;��H;j�H;��H;`�H;��H;~�H;��H;0�H;- I;6I;yI;�I;-I;='I;�4I;�DI;DWI;�mI;��I;e�I;��I;��I;��I;��I;P�I;�	I;M%H;��F;�	E;�B;� @;�/=;)#:;�07;p�4;�2;_51;      D;�; �;��;� ;�&;�\,;ԇ2;98;�/=;�FA;krD;P�F;JH;[9I;-�I;i�I;V�I;��I;~�I;o�I;pI;AXI;�DI;�3I;T&I;I;�I;
I;hI;��H;��H;��H;��H;9�H;H�H;�H;F�H;6�H;��H;��H;��H;��H;oI;|
I;�I;!I;[&I;�3I;�DI;CXI;pI;p�I;��I;��I;R�I;n�I;.�I;[9I;JH;T�F;jrD;�FA;�/=;98;ԇ2;�\,;�&;� ;��;�;�;      <��:��:��:���:���:�P ;�e;�V;H#;e-;��5;�h<;QtA;T	E;�eG;7�H;/�I;�I;��I;�I;�I;�I; pI;GWI;�BI;:2I;�$I;sI;lI;=	I;uI;��H;��H;�H;V�H;/�H;��H;2�H;U�H; �H;��H;��H;yI;C	I;kI;sI;�$I;@2I;�BI;NWI;pI;�I;�I;�I;��I;
�I;/�I;7�H;�eG;T	E;QtA;�h<;��5;e-;M#;�V;�e;�P ;��:��:��:s�:      ��p� �,��!9�ų9��":��u:��:Z��:���:(R;\ ;��,;�6;N)>;�;C;��F;�lH;fkI;o�I;��I;��I;�I;l�I;�mI;yTI;@I;�/I;!"I;VI;�I;�I;�I;r�H;r�H;��H;S�H;��H;T�H;�H;n�H;t�H;�I;�I;�I;UI;""I;�/I;#@I;yTI;�mI;n�I;�I;��I;��I;u�I;fkI;�lH;��F;�;C;P)>;�6;��,;^ ;,R;���:^��:��:��u:��":�ų9`"9 �,�      
p&��!��4���氺�O� =T��t�9��u:�#�:�G�:D;&#;d71;:;;��A;��E;�$H;HVI;�I;��I;�I;~�I;��I;iI;"PI;<I;�+I;I;�I;�I;�I;�I;5�H;��H;��H;�H;��H;��H;.�H;�I;�I;�I;�I;I;�+I;<I;&PI;iI; �I;��I;�I;��I;�I;MVI;�$H;��E;��A;:;;e71;'#;D;�G�:�#�:��u:�t�9�<T�,�O��氺���4��!�      �kٻn�Ի�ǻ����V���n���+�8�Ժ��1���39Dm:��:h�;�;{\,;��8;��@;:]E;�
H;IVI;q�I;��I;��I;`�I;��I;�bI;[JI;"7I;�'I;�I;,I;�
I;6I;9I;i�H;��H;y�H;��H;d�H;6I;6I;�
I;/I;�I;�'I;"7I;bJI;�bI;��I;g�I;��I;��I;r�I;MVI;�
H;8]E;��@;ݍ8;z\,;	�;j�;��:Pm:��39 �1�6�Ժ��+��n��V������ǻj�Ի      7yY��|U�L�I�A�7��� ��!���Ի�᝻��T���#�xu�9���:Kl�:�;�);17;+ @;7]E;�$H;bkI;�I;R�I;��I;+�I;�wI;�ZI;�CI;x1I;I#I;%I;�I;+	I;rI;6I;j�H;��H;k�H;2I;rI;+	I;�I;'I;O#I;w1I;�CI;�ZI;�wI;'�I;��I;S�I;
�I;dkI;�$H;:]E;+ @;17;�);�;Ol�:���:�u�9�#����T��᝻��Ի"��� �B�7�O�I��|U�      ��ü^l��w����R��@ߓ�b�{��M��� �"��̼����B�갺�Io���u:���:�R;/�';17;��@;��E;�lH;.�I;e�I;��I;	�I;s�I;�lI;}QI;'<I;�+I;�I;�I;cI;�I;BI;.I;�I;.I;?I;�I;bI;�I;�I;�+I;&<I;~QI;�lI;t�I;�I;��I;i�I;1�I;�lH;��E;��@;17;/�';�R;���:��u: Io�갺��B�̼�� �컋� ��M�a�{�@ߓ��R��x���]l��      �'��-$�_��Y����
?ټ	w��<���pyY��k� �Ի:��
Y�������#R:���:�R;�);ٍ8;��A;��F;4�H;)�I;��I;��I;��I;�I;�`I;�GI;�4I;�%I;HI;�I;�I;rI;I;EI;I;mI;�I;�I;FI;�%I;�4I;�GI;�`I;�I;��I;��I;��I;*�I;6�H;��F;��A;ڍ8;�);�R;���:�#R:����Y��:�� �Ի�k�qyY�<���	w��
?ټ���Y�`���-$�      Y+����c̀�,l��Q�%�2�B��������@����>�]2��"V���1�����#R:���:�;t\,;4;;�;C;�eG;X9I;��I;0�I;��I;=�I;�qI;�TI;_>I;8-I;0 I;zI;uI;�
I;I;I;I;�
I;qI;zI;- I;6-I;_>I;�TI;�qI;@�I;��I;-�I;��I;X9I;�eG;�;C;8;;t\,;�;���:�#R:ȑ�1�"V��]2����>��@��������B�$�2��Q�-l�c̀���      l�ྲྀhܽo�н^y��`什P ��l��n<�M���>ټ��W|U���������1�������u:Kl�:�;b71;U)>;S	E;JH;T�I;��I;��I;�I;փI;[bI;�HI;'5I;b&I;dI;qI;:I;"I;
I;%I;9I;qI;gI;]&I;$5I;�HI;\bI;׃I;�I;��I;��I;U�I;JH;T	E;L)>;g71;�;Ol�:��u:�����1��������X|U����>ټM���n<�l�P ��`什^y��n�н�hܽ      ��4�g1��&������j�ཅ�������`��'���UR��F�]�~��V���X�� Io����:h�;'#;�6;RtA;R�F;�	I;x�I;��I;i�I;�I;�pI;�SI;�=I;�,I;v I;�I;�I;GI;;I;GI;�I;�I;w I;�,I;�=I;�SI;�pI;�I;k�I;��I;t�I;�	I;T�F;RtA;�6;,#;f�;���:@Ho��X�� V��~��F�]�UR����'��`��������j��������&�g1�      �x���o��ń�HUo���O�*�-�{��hܽ\什Լx���2�tb��VR��X|U�\2��:��&갺`u�9��:D;��,;�h<;drD;N%H;ǏI;e�I;��I;�I;�I;�^I;	FI;S3I;�%I;�I;\I;fI;5I;hI;\I;�I;�%I;R3I;FI;�^I;�I;�I;��I;e�I;��I;N%H;jrD;�h<;��,;D;��:pu�9"갺<��^2��X|U�VR��tb����2�Լx�]什�hܽ{�*�-���O�HUo�ń��o��      w���ྃ�Ѿ(����נ�ń�9�S��#�`O��|n��J̀���2���𛼃�>��Ի��B��#�,m:�G�:_ ;��5;�FA;��F;�I;M�I;M�I;��I;k�I;kjI;�NI;:I;�*I;�I;�I;�I;KI;�I;�I;�I;�*I;:I;�NI;mjI;m�I;��I;P�I;M�I;�I;��F;�FA;��5;U ;�G�:(m:�#���B��Ի��>�������2�J̀�|n��_O���#�9�S�ń��נ�(�����Ѿ��      �3���/��X#��	��A��֌Ⱦ�f��GUo�^1�˰��|n��Լx��'��>ټ�@���k�μ��(����39�#�:.R;e-;�/=;�	E;_xH;�I;�I;m�I; �I;vI;cWI;�@I;�/I;%$I;;I;�I;5I;�I;;I;#$I;�/I;�@I;cWI;vI;�I;p�I;	�I;�I;YxH;�	E;�/=;	e-;$R;�#�:��39$��μ���k��@���>ټ�'�Լx�|n��˰��^1�GUo��f��֌Ⱦ�A���	��X#���/�      ���U���U�v��RZ�[58�͂�q��d���foy�^1�_O��]什�`�M�����pyY�%�컝�T��1���u:���:F#;98;�B;j�G;�lI;�I;��I;.�I;t�I;�_I; GI;�4I;&(I;�I;�I;I;�I;�I;#(I;�4I;GI;�_I;s�I;.�I;�I;�I;�lI;h�G;�B;98;C#;���:��u:$�1���T�$��qyY����M���`�]什_O��^1�foy�d���q��͂�[58��RZ�U�v�U���      	Ŀ6g��&ﱿ���T����U��X#�t��d���HUo��#��hܽ����n<����=����� ��᝻J�Ժ�t�9b��:�V;̇2;� @;W�F;�I;��I;>�I;&�I;g�I;�gI;MI;�9I;�+I;�"I;iI;�I;hI;�"I;�+I;�9I;MI;�gI;i�I;(�I;@�I;��I;�I;R�F;� @;χ2;�V;P��:�t�9N�Ժ�᝻�� �=�������n<�����hܽ�#�HUo�d���t���X#��U�T������'ﱿ6g��      ~x�P9�R��uؿnQ��e_��6�_��X#�r���f��9�S�{�����l�B�	w�� �M���Ի��+�=T���:�e;�\,;�/=;�BE;P�H;v�I;��I;��I;��I;�oI;�RI;>I;\/I;{%I;�I;DI;�I;~%I;\/I;>I;�RI;�oI;��I;��I;��I;w�I;W�H;�BE;�/=;�\,;�e;��: =T��+���Ի�M�	w��B�l�����{�9�S��f��r���X#�6�_�e_��nQ��uؿR��P9�      �X1���,�h���<��5g��e_���U�͂�֌Ⱦ	ń�*�-�j��P ��%�2�?ټb�{�"��n� �O���u:�P ;�&;)#:;:�C;�%H;�I; �I;��I;�I;]vI;�WI;�AI;x2I;(I;A"I;^ I;A"I;(I;x2I;�AI;�WI;YvI;�I;��I;$�I;�I;�%H;<�C;+#:;�&;�P ;t�u: �O��n�"�b�{�?ټ&�2�P ��j��*�-�	ń�֌Ⱦ͂��U�e_��5g��<�h����,�      d��]]�5K��X1�Zf��nQ��T���[58��A���נ���O���`什�Q����@ߓ��� ��V���氺��":и�:� ;�07;�B;,�G;�{I;��I;��I;��I;7|I;4\I;IEI;5I;0*I;1$I;)"I;-$I;3*I;5I;JEI;4\I;4|I;��I;��I;��I;�{I;5�G;�B;�07; ;Ҹ�:܌":�氺�V���� �@ߓ�����Q�`什����O��נ��A��[58�T���nQ���Zf��X1�5K��]]�      N������4z���V��X1��<�uؿ����RZ��	�(���HUo����^y��-l�Z��R��D�7�������ų9���:��;W�4;itA;X2G;�XI;��I;J�I;�I;�I;�_I;�GI;!7I;�+I;�%I;�#I;�%I;�+I;7I;�GI;�_I;�I;�I;H�I;��I;�XI;c2G;gtA;X�4;��;���:�ų9�����D�7��R��Y�-l�^y�����HUo�(����	��RZ����uؿ�<��X1���V��4z�����      �o��e^���ē��4z�5K�h��R��'ﱿU�v��X#���Ѿń��&�o�нc̀�_��v���K�I��ǻ�4�P"9��:2�; �2;��@;��F;�:I;��I;��I;��I;v�I;KbI;�II;�8I;W-I;�&I;�$I;�&I;Z-I;�8I;�II;JbI;p�I;��I;��I;��I;�:I;��F;��@;�2;0�;��:�!9�4��ǻL�I�v���_��c̀�o�н�&�ń���Ѿ�X#�U�v�'ﱿR��h��5K��4z��ē�e^��      q'���X��e^�������]]���,�P9�6g��U�����/����o��g1��hܽ���-$�`l���|U�h�Ի�!� �,�u�:�;�51;��?;1�F;?'I;_�I;�I;<�I;��I;�cI;>KI;x9I;.I;y'I;�%I;v'I; .I;x9I;>KI;�cI;��I;?�I;
�I;b�I;?'I;?�F;��?;51;�;m�: �,��!�j�Ի�|U�_l���-$����hܽg1��o���ྙ�/�U���6g��P9���,��]]�����e^���X��      ����,������T���J�Q�Ǚ$�3�����;�}�H(�A�׾�T���L+���սk����!L���iO���ͻ����m8bo�:Z�;R�1;��?;�uF;f I;e�I;��I;��I;VvI;�WI;�AI;�1I;�'I;�!I;�I;�!I;�'I;�1I;�AI;�WI;TvI;��I;��I;f�I;d I;�uF;��?;O�1;S�;Zo�: m8�����ͻ�iO� L����k����ս�L+��T��A�׾H(�;�}���3���Ǚ$�J�Q�T��������,��      �,��a��#P���{���K��x �����q�����w��$���Ҿg���  (���ѽҷ��(�����K�Hɻ.�� ��8p��:x�;��1;�@;i�F;I;ۿI;�I;��I;�uI;#WI;eAI;�1I;�'I;�!I;�I;�!I;�'I;�1I;fAI;%WI;�uI;��I;�I;޿I;I;t�F;�@;��1;p�;h��: ��8-��Hɻ�K����(�ҷ����ѽ  (�g�����Ҿ�$���w�q��������x ���K��{�#P��a��      ����#P�������d���;�#���㿳���#f�d��ž��z���=�ƽ&0v�U5�2����o@������i��`u9;K�:];�73;�@;��F;FI;��I;M�I;R�I;�sI;�UI;A@I;�0I;�&I;!I;0I;!I;�&I;�0I;?@I;�UI;�sI;V�I;M�I;��I;CI;��F;�@;�73;];3K�:0`u9}i������o@�2���U5�&0v�=�ƽ����z�žd��#f�������#����;���d����#P��      T����{���d��F�Ǚ$�:����ɿ.蒿��K�Q���j���Yb�E�1���s�a����?�����.��d��x�غ���9�Y�:,X;�25;�A;X!G;H7I;q�I;@�I;P�I;�pI;�SI;~>I;y/I;�%I;% I;.I; I;�%I;x/I;~>I;�SI;�pI;R�I;B�I;q�I;F7I;_!G;�A;�25;$X;�Y�:x��9x�غ�d����.�?������s�a�1���E��Yb��j��Q����K�.蒿��ɿ:��Ǚ$��F���d��{�      J�Q���K���;�Ǚ$��;
��޿�����w�q,���澝���'�D������I��$�G�����N��������^�����9:R��:�n!;��7;��B;J�G;�YI;(�I;V�I;��I;�lI;sPI;<I;�-I;$I;�I;�I;�I;$I;�-I;<I;rPI;�lI;��I;V�I;+�I;�YI;P�G;��B;��7;�n!;N��:l�9:\����������N�����$�G��I������'�D��������q,���w�����޿�;
�Ǚ$���;���K�      Ǚ$��x �#��:���޿p���ʅ���F�}�
��~����z��$���ս���@2+���ϼPp�����T�]�,�*���:�;�8';��:;��C;�H;�}I;�I;p�I;ԋI;hgI;�LI;9I;7+I;"I;�I;)I;�I; "I;3+I;9I;�LI;egI;ًI;o�I;�I;�}I;H;��C;��:;�8';�;��:(�*�T�]�����Pp���ϼ@2+������ս�$���z��~��}�
��F�ʅ��p����޿:��#���x �      3��������㿊�ɿ���ʅ����P�d��<�׾�`��T�H����@��R�a���Ρ���D��ɻ� ��ح��W�:�;`I-;4|=;CE;��H;�I;��I;r�I;��I;eaI; HI;�5I;o(I;�I;�I;QI;�I;�I;o(I;�5I;HI;caI;��I;s�I;��I;	�I;��H;CE;4|=;\I-;�;�W�:�ح�� ��ɻ�D�Ρ����R�a��@����T�H��`��<�׾d����P�ʅ�������ɿ�㿳���      ��q�������.蒿��w��F�d��ʰ� ����Yb�)����ѽ�%��D4�ٟ� X�����H���潺���9Br�:��;�93;$Q@;zvF;�H;	�I;��I;��I;�zI;�ZI;CI;�1I;a%I;?I;�I;"I;�I;BI;b%I;�1I;CI;�ZI;�zI;��I;��I;�I;�H;|vF; Q@;�93;��;2r�:���9�潺H����� X��ٟ�D4��%����ѽ)���Yb� ���ʰ�d���F���w�.蒿����q���      ;�}���w�#f���K�q,�}�
�<�׾ �����k���'�fz꽝I���;V�=M�
����iO�nG�toE�̱�0��:A� ;��$;��8;Y�B;��G;,KI;�I;�I;>�I;qI;�SI;�=I;�-I;"I;kI;I;�I;I;mI;"I;�-I;�=I;�SI;	qI;@�I;�I;�I;+KI;��G;X�B;��8;��$;;� ;8��:̱�woE�mG໭iO�
���=M��;V��I��fz���'���k� ���<�׾}�
�q,���K�#f���w�      H(��$�d��Q������~���`���Yb���'��U�H$��C�m�&����ϼ�/��?��������غ88�94��:�F;�G.;|=;GE;�\H;�I;u�I;x�I;��I;gI;�KI;�7I;)I;nI;rI;rI;%I;qI;rI;nI;)I;�7I;LI;gI;��I;y�I;r�I;�I;�\H;DE;|=;�G.;�F;<��:88�9��غ����@���/����ϼ&��C�m�H$���U���'��Yb��`���~�����Q��d���$�      A�׾��Ҿž�j��������z�S�H�)��fz�H$���/v�2+�ݐ�����5��ɻ>4�P(��~��:T��:6o!;P6;lA;��F;p�H;��I;��I;ߦI;F}I;�\I;[DI;2I;p$I;�I;HI;�I;�I;�I;II;�I;p$I;2I;[DI;�\I;J}I;�I;��I;��I;s�H;��F;lA;P6;5o!;f��:~��:h(��<4��ɻ��5���ݐ�2+��/v�H$��fz�)��S�H���z������j��ž��Ҿ      �T��f�����z��Yb�'�D��$�����ѽ�I��C�m�2+�������K�K�ﻛ�p�R������9#T�:�/;q�-;d�<;BzD;YH;�mI;��I;}�I;��I;�oI;�RI;�<I;,I;�I;I;1I;�I;�I;�I;/I;I;�I;�+I;�<I;�RI;�oI;��I;z�I;��I;�mI;YH;FzD;i�<;o�-;�/;#T�:���9L�����p��J�K�������2+�C�m��I����ѽ���$�'�D��Yb���z�f���      �L+�  (���E�������ս�@���%���;V�&��ݐ������MS�N��(���D���n8 q�:�;b�$;�^7;(�A;d�F;��H;_�I;b�I;��I;݃I;RbI;�HI;5I;%&I;/I;>I;�I;�
I;
I;�
I;�I;=I;-I;"&I;5I;�HI;VbI;��I;��I;]�I;b�I;��H;e�F;+�A;�^7;k�$;�;�p�:��n8~D�(��M���MS�����ܐ�&���;V��%���@����ս����E���  (�      ��ս��ѽ<�ƽ1����I�����R�a�D4�=M���ϼ��J�K�O��QG��bf���o���:�B�:�Y;��1;Ol>;�E;�/H;qI;��I;��I;٘I;�rI;�UI;�>I;�-I;b I;�I;�I;�
I;I;0I;I;�
I;�I;�I;^ I;�-I;�>I;�UI;sI;٘I;��I;��I;qI;�/H;�E;Nl>;��1;�Y;�B�:��: �o�df�PG��O��J�K�����ϼ<M�D4�R�a�����I��1���<�ƽ��ѽ      j��ҷ��&0v�s�a�#�G�@2+���؟�	����/����5��)��df��ج���g:3�:�;I-;g;;�NC;SG;�I;ȶI;�I;��I;�I;	cI;}II;�5I;n&I;�I;5I;�I;�I;PI;ZI;NI;�I;�I;5I;�I;r&I;�5I;II;cI;�I;��I;�I;ȶI;�I;
SG;�NC;g;;I-;�;7�:Ԙg:�ج�bf�(�����5��/��	���؟���?2+�$�G�s�a�&0v�ҷ��      
��'�T5���������ϼ͡��X���iO�?���ɻ��p��D���o�ؘg:�_�:AG;n*;o9;��A;�uF;�H;��I;��I;��I;F�I;�pI;1TI;M>I;-I;�I;{I;�I;VI;�I;�I;�I;�I;�I;TI;�I;xI;�I;-I;O>I;5TI;�pI;?�I;��I;��I;��I;�H;�uF;��A;p9;f*;AG;�_�:��g: �o��D⺜�p��ɻ?���iO�X��͡����ϼ������T5�&�      L�����3���?����N��Pp��D����jG�����74�L��� �n8��:;�:GG;�(;��7;Y�@;��E;KQH;mI;��I;��I;��I;#}I;�^I;�FI;�3I;�$I;[I;�I;�	I;I;�I;��H;O�H;��H;�I;I;�	I;�I;^I;�$I;�3I;�FI;�^I;}I;��I;��I;�I;mI;MQH;��E;Z�@;��7;�(;DG;9�:��:��n8J���64�����jG່���D�Pp��N��@���4������      �iO���K��o@���.���������ɻH��qoE���غ8(�����9�p�:�B�:�;l*;��7;�P@;�\E;�H;�II;~�I;f�I;�I;V�I;<hI;�NI;`:I;9*I;xI;�I;�I;I;I;2�H;a�H;��H;^�H;-�H;I;I;�I;�I;{I;6*I;b:I;�NI;7hI;\�I;�I;a�I;�I;�II;�H;�\E;�P@;��7;h*;�;�B�:�p�:���9(����غmoE�H���ɻ���������.��o@�ߔK�      ��ͻNɻ�����d�����B�]�� ��潺���X8�9���:#T�:�;�Y;I-;s9;Y�@;�\E;��G;/5I;��I;C�I;ٵI;R�I;apI;�UI;S@I;2/I;{!I;�I;?I;�I;�I;!�H;��H;�H;��H;�H;��H;�H;�I;�I;AI;�I;x!I;4/I;Q@I;�UI;gpI;S�I;ҵI;E�I;��I;25I;��G;�\E;\�@;o9;I-;�Y;�;)T�:���:H8�9����潺� �J�]�����d������Mɻ      ���1��vi�^�غj����*��׭����98��:<��:f��:�/;e�$;��1;g;;��A;��E;�H;05I;6�I;��I;J�I;��I;�vI;L[I;^EI;�3I;2%I;�I;�I;P	I;�I;|�H;`�H;%�H;��H;l�H;��H;"�H;^�H;|�H;�I;Q	I;�I;�I;5%I;�3I;ZEI;R[I;�vI;��I;L�I;��I;6�I;25I;�H;��E;��A;g;;��1;e�$;�/;h��:<��:<��:���9�׭��*�\���x�غ�i�8��       (m8���8 _u9h��9L�9:��:�W�:Br�:=� ;�F;6o!;n�-;�^7;Nl>;�NC;�uF;MQH;�II;��I;��I;��I;��I;{zI;_I;<II;I7I;a(I;^I;�I;I;�I;) I;p�H;��H; �H;��H;r�H;��H;�H;��H;p�H;% I;�I;I;�I;`I;^(I;G7I;@II;{_I;tzI;��I;��I;��I;��I;�II;MQH;�uF;�NC;Kl>;�^7;n�-;;o!;�F;:� ;6r�:�W�:��:x�9:x��9�_u9@��8      Vo�:���:YK�:�Y�:B��:�;�;��;��$;�G.;P6;f�<;(�A;�E;SG;�H;mI;��I;G�I;M�I;��I;�{I;taI;�KI;�9I;�*I;�I;�I;�I;$I;� I;��H;��H;j�H;��H;�H;��H;�H;��H;j�H;��H;��H;� I;$I;�I;�I;�I;�*I;�9I;�KI;laI;�{I;��I;L�I;E�I;~�I;mI;�H;
SG;�E;(�A;i�<;P6;�G.;��$;��;�;�;r��:�Y�:CK�:z��:      l�;x�;];8X;�n!;�8';jI-;�93;��8;|=;lA;LzD;f�F;�/H;�I;ƔI;��I;h�I;صI;��I;zzI;oaI;uLI;;I;^,I;. I;I;�I;:I;�I;t�H;��H;d�H;l�H;�H;S�H;!�H;N�H;�H;m�H;d�H;��H;w�H;�I;4I;�I;I;. I;b,I;;I;nLI;qaI;zzI;��I;ٵI;d�I;��I;ĔI;�I;�/H;e�F;LzD;lA;|=;��8;�93;fI-;�8';�n!;8X;
];^�;      R�1;��1;�73;�25;{�7;��:;-|=;!Q@;T�B;GE;��F;YH;��H;qI;ƶI;��I;��I;�I;O�I;�vI;{_I;�KI;;I;�,I;� I;I;�I;I;qI;��H;p�H;m�H; �H;��H;m�H;��H;��H;��H;k�H;��H; �H;j�H;u�H;��H;mI;I;�I;I;� I;�,I;;I;�KI;y_I;�vI;L�I;�I;��I;��I;ƶI;qI;��H;YH;��F;EE;V�B;'Q@;+|=;��:;��7;�25;�73;��1;      ��?;�@;�@;�A;��B; �C;&CE;|vF;��G;�\H;w�H;�mI;_�I;�I;�I;��I;��I;_�I;lpI;W[I;GII;�9I;d,I;� I;mI;]I;�I;�I;f�H;��H;��H;+�H;S�H;��H;��H;[�H;1�H;V�H;��H;��H;R�H;&�H;��H;��H;b�H;�I;�I;]I;nI;� I;a,I;�9I;DII;R[I;lpI;\�I;��I;��I;�I;�I;a�I;�mI;x�H;�\H;��G;zvF;#CE;��C;��B;�A;�@;�@;      �uF;w�F;��F;V!G;?�G;H;��H;�H;0KI;"�I;��I;��I;`�I;��I;��I;H�I;&}I;;hI;�UI;[EI;L7I;�*I;- I;I;ZI;�I;DI;��H;��H;��H;#�H;=�H;��H;Z�H;��H;�H;��H;�H;��H;[�H;��H;7�H;#�H;��H;��H;��H;@I;�I;\I;I;) I;�*I;K7I;ZEI;�UI;8hI;'}I;I�I;��I;��I;`�I;��I;��I;!�I;/KI;�H;��H;�H;U�G;i!G;��F;x�F;      t I;)I;@I;I7I;�YI;�}I;�I;�I;�I;u�I;��I;|�I;��I;ژI;�I;�pI;�^I;�NI;V@I;�3I;i(I;�I; I;�I;�I;BI;��H;"�H;��H;1�H;!�H;h�H;�H;�H;�H;�H;��H;��H;|�H;�H;�H;b�H;�H;.�H;��H;�H;��H;EI;�I;�I;I;�I;g(I;�3I;S@I;�NI;�^I;�pI;�I;՘I;��I;|�I;��I;r�I;�I;�I;�I;�}I;�YI;B7I;?I;I;      c�I;�I;��I;w�I;�I;�I;��I;��I;�I;}�I;�I;��I;܃I;sI;cI;3TI;�FI;]:I;3/I;2%I;bI;�I;�I;I;�I;��H;�H;��H;B�H;�H;U�H;��H;��H;��H;X�H;��H;��H;��H;W�H;��H;��H;��H;U�H;�H;=�H;��H;�H;��H;�I;I;�I;�I;`I;1%I;2/I;Y:I;�FI;4TI;cI; sI;܃I;��I;�I;}�I;�I;��I;��I;�I;$�I;{�I;��I;ؿI;      ��I;��I;K�I;S�I;L�I;q�I;w�I;��I;:�I;��I;J}I;�oI;RbI;�UI;II;O>I;�3I;:*I;!I;�I;�I;�I;6I;pI;b�H;��H;��H;B�H;0�H;T�H;��H;��H;��H;��H;y�H;3�H;*�H;-�H;w�H;��H;��H;��H;��H;Q�H;*�H;?�H;��H;��H;d�H;jI;6I;�I;�I;�I;~!I;7*I;�3I;Q>I;�II;�UI;QbI;�oI;M}I;��I;=�I;��I;w�I;i�I;V�I;W�I;I�I;��I;      ��I;��I;`�I;L�I;��I;ԋI;��I;�zI;	qI;	gI;�\I;�RI;�HI;�>I;�5I;-I;�$I;tI;�I;�I;"I; I;�I;��H;��H;��H;1�H;"�H;Z�H;��H;��H;��H;��H;�H;��H;y�H;Y�H;v�H;��H;�H;��H;��H;��H;��H;U�H;!�H;+�H;��H;��H;��H;�I;"I;I;�I;�I;qI;�$I;-I;�5I;�>I;�HI;�RI;�\I;gI;qI;�zI;��I;׋I;��I;W�I;]�I;��I;      UvI;�uI;�sI;�pI;�lI;jgI;faI;�ZI;�SI;LI;`DI;�<I;5I;�-I;u&I;�I;cI;�I;CI;W	I;�I;� I;s�H;t�H;��H;#�H;"�H;\�H;��H;��H;��H;��H;��H;Y�H;�H;��H;��H;��H;	�H;\�H;��H;��H;��H;��H;��H;X�H;�H;$�H;��H;p�H;w�H;� I;�I;P	I;CI;�I;cI;�I;t&I;�-I;5I;�<I;aDI;LI;�SI;�ZI;oaI;agI;�lI;�pI;�sI;�uI;      �WI;-WI;�UI;�SI;ePI;�LI;HI;CI;�=I;�7I;2I;,I;'&I;g I;�I;{I;�I;�I;�I;�I;1 I;��H;��H;j�H;+�H;4�H;e�H;��H;��H;��H;��H;��H;A�H;��H;{�H;?�H;H�H;?�H;x�H;��H;E�H;��H;��H;��H;��H;��H;b�H;6�H;-�H;d�H;��H;��H;* I;�I;�I;�I;�I;}I;�I;g I;'&I;,I;2I;�7I;�=I;CI;'HI;�LI;oPI;�SI;�UI;-WI;      �AI;sAI;C@I;�>I;<I;9I;�5I;�1I;�-I;)I;p$I;�I;-I;�I;7I;�I;�	I;I;�I;��H;}�H;��H;c�H;�H;V�H;��H;�H;��H;��H;��H;��H;D�H;��H;[�H;�H;��H;��H;��H;	�H;\�H;��H;E�H;��H;��H;��H;��H;�H;��H;W�H;�H;e�H;��H;u�H;|�H;�I;I;�	I;�I;9I;�I;/I;�I;u$I;)I;�-I;�1I;�5I;9I;<I;>I;M@I;sAI;      �1I;�1I;�0I;o/I;�-I;*+I;o(I;f%I;"I;uI;�I;I;BI;�I;�I;XI;I;I;#�H;e�H;��H;j�H;j�H;��H;��H;V�H;�H;�H; �H;�H;V�H;��H;\�H;��H;��H;��H;~�H;��H;��H;��H;]�H;��H;U�H;�H;��H;��H;�H;V�H;��H;��H;o�H;g�H;��H;]�H;!�H;I;I;XI;�I;�I;BI;I;�I;uI;"I;b%I;w(I;(+I;�-I;u/I;�0I;�1I;      �'I;�'I;�&I;�%I;$I;"I;�I;II;pI;}I;PI;<I;�I;�
I;�I;�I;�I;/�H;��H;(�H;
�H;��H;�H;c�H;��H;��H;{�H;\�H;��H;��H;�H;{�H;�H;��H;~�H;[�H;U�H;[�H;{�H;��H;�H;|�H;�H;��H;y�H;U�H;z�H;��H;��H;b�H;�H;��H;�H;"�H;��H;2�H;�I;�I;�I;�
I;�I;;I;VI;I;pI;GI;�I;"I;$I;�%I;�&I;�'I;      �!I;�!I;!I; I;�I;�I;�I;�I;I;xI;�I;�I;�
I;I;PI;�I;��H;Z�H;�H;��H;��H;�H;K�H;��H;X�H;�H;�H;�H;:�H;}�H;��H;A�H;��H;��H;_�H;(�H;+�H;+�H;[�H;��H;��H;F�H;��H;x�H;4�H;��H;�H;�H;T�H;��H;O�H;�H;��H;��H;�H;^�H;��H;�I;SI;I;�
I;�I;�I;yI;I;�I;�I;�I;�I;" I;!I;�!I;      �I;�I;>I;+I;�I;!I;TI;(I;�I;'I;�I;�I;
I;7I;`I;�I;V�H;��H;��H;s�H;�H;��H;�H;��H;.�H;��H;��H;��H;1�H;^�H;��H;J�H;��H;z�H;W�H;'�H;�H;(�H;S�H;{�H;��H;K�H;��H;Y�H;,�H;��H;��H;��H;,�H;��H;!�H;��H;w�H;n�H;��H;��H;V�H;�I;aI;;I;
I;�I;�I;'I;�I;&I;ZI;!I;�I;0I;=I;�I;      �!I;�!I;!I; I;�I;�I;�I;�I;I;xI;�I;�I;�
I;I;PI;�I;��H;Z�H;�H;��H;��H;�H;K�H;��H;W�H;�H;�H; �H;:�H;|�H;��H;D�H;��H;��H;a�H;(�H;+�H;+�H;[�H;��H;��H;F�H;��H;v�H;4�H;��H;�H;�H;V�H;��H;O�H;�H;��H;��H;�H;^�H;��H;�I;SI;I;�
I;�I;�I;vI;I;�I;�I;�I;�I;& I;	!I;�!I;      �'I;�'I;�&I;�%I;$I;"I;�I;LI;pI;|I;PI;<I;�I;�
I;�I;�I;�I;/�H;��H;'�H;�H;��H;�H;`�H;��H;��H;z�H;Z�H;~�H;��H;�H;{�H;�H;��H;~�H;\�H;U�H;\�H;}�H;��H;�H;|�H;�H;��H;y�H;T�H;z�H;��H;��H;`�H;�H;��H;�H;!�H;��H;2�H;�I;�I;�I;�
I;�I;<I;VI;|I;pI;MI;�I;"I;$I;�%I;�&I;�'I;      �1I;�1I;�0I;t/I;�-I;/+I;o(I;i%I;"I;tI;�I;I;AI;�I;�I;XI;I;I;"�H;a�H;��H;j�H;h�H;��H;��H;T�H;�H;�H; �H;�H;U�H;��H;\�H;��H;��H;��H;~�H;��H;��H;��H;]�H;��H;U�H;�H;��H;��H;�H;X�H;��H;��H;o�H;h�H;��H;^�H;#�H;I;I;ZI;�I;�I;BI;I;�I;tI;"I;f%I;z(I;-+I;�-I;u/I;�0I;�1I;      �AI;zAI;F@I;~>I;<I;9I;�5I;�1I;�-I;)I;o$I;�I;-I;�I;9I;�I;�	I;I;�I;��H;|�H;��H;`�H;�H;W�H;��H;�H;��H;��H;��H;��H;B�H;��H;[�H;�H;��H;��H;��H;�H;[�H;��H;E�H;��H;��H;��H;��H;�H;��H;U�H;�H;g�H;��H;s�H;�H;�I;I;�	I;�I;7I;�I;2I;�I;u$I;)I;�-I;�1I;�5I;9I;<I;�>I;S@I;tAI;      �WI;2WI;�UI;�SI;ePI;�LI;#HI;CI;�=I;�7I;	2I;,I;%&I;d I;�I;}I;�I;�I;�I;�I;1 I;��H;��H;e�H;-�H;3�H;b�H;��H;��H;��H;��H;��H;B�H;��H;|�H;=�H;H�H;A�H;x�H;��H;D�H;��H;��H;��H;��H;��H;a�H;4�H;*�H;`�H;��H;��H;* I;�I;�I;�I;�I;}I;�I;e I;(&I;
,I;2I;�7I;�=I;CI;&HI;�LI;gPI;�SI;�UI;,WI;      MvI;�uI;�sI;�pI;�lI;hgI;faI;�ZI;�SI;LI;^DI;�<I;5I;�-I;t&I;�I;cI;�I;AI;Q	I;�I;� I;q�H;p�H;��H;�H;�H;Z�H;��H;��H;��H;��H;��H;Z�H;�H;��H;��H;��H;�H;\�H;��H;��H;��H;��H;��H;W�H;�H;#�H;��H;n�H;z�H;� I;�I;Q	I;DI;�I;eI;�I;u&I;�-I;5I;�<I;bDI;LI;�SI;�ZI;oaI;egI;�lI;�pI;�sI;�uI;      ��I;��I;X�I;W�I;��I;��I;��I;�zI;qI;
gI;�\I;�RI;�HI;�>I;�5I;-I;�$I;tI;�I;�I;"I;!I;�I;��H;��H;��H;.�H;!�H;Z�H;��H;��H;��H;��H;�H;��H;x�H;Z�H;y�H;��H;�H;��H;��H;��H;��H;T�H;!�H;.�H;��H;��H;��H;�I;!I;I;�I;�I;qI;�$I;-I;�5I;�>I;�HI;�RI;�\I;gI;	qI;�zI;��I;ҋI;��I;^�I;c�I;��I;      ��I;��I;Z�I;J�I;=�I;v�I;s�I;��I;@�I;�I;G}I;�oI;QbI;�UI;�II;Q>I;�3I;<*I;{!I;�I;�I;�I;2I;nI;c�H;��H;��H;?�H;-�H;Q�H;��H;��H;��H;��H;y�H;1�H;,�H;1�H;w�H;��H;��H;��H;��H;S�H;)�H;=�H;��H;��H;b�H;iI;7I;�I;�I;�I;!I;7*I;�3I;T>I;�II;�UI;RbI;�oI;L}I;�I;=�I;��I;|�I;p�I;N�I;K�I;Z�I;��I;      o�I;׿I;��I;y�I;�I;'�I;��I;��I;�I;|�I;�I;��I;܃I;�rI;	cI;4TI;�FI;]:I;0/I;/%I;aI;�I;�I;I;�I;��H;�H;��H;C�H;�H;T�H;��H;��H;��H;[�H;��H;��H;��H;X�H;�H;��H;��H;X�H;�H;?�H;��H;�H;��H;�I;I;�I;�I;^I;1%I;3/I;Y:I;�FI;4TI;
cI;sI;܃I;��I;�I;�I;�I;��I;��I;�I;#�I;{�I;��I;׿I;      a I;,I;>I;S7I;�YI;�}I;�I;�I;�I;s�I;��I;��I;��I;טI;�I;�pI;�^I;�NI;Q@I;�3I;h(I;�I;I;�I;�I;=I;��H;!�H;��H;-�H;�H;h�H;�H;�H;�H;�H;��H;�H;|�H;�H;�H;i�H;"�H;/�H;��H;�H;��H;DI;�I;�I;!I;�I;d(I;�3I;T@I;�NI;�^I;�pI;�I;֘I;��I;y�I;��I;r�I;�I;�I;�I;�}I;�YI;W7I;>I;I;      �uF;r�F;��F;U!G;C�G;H;��H; �H;/KI; �I;��I;��I;`�I;��I;��I;H�I;#}I;<hI;�UI;WEI;L7I;�*I;& I;I;ZI;�I;AI;��H;��H;��H;#�H;=�H;��H;[�H;��H;�H;��H;�H;��H;[�H;��H;>�H;'�H;��H;��H;��H;DI;�I;ZI;I;, I;�*I;K7I;[EI;�UI;8hI;'}I;K�I;��I;��I;_�I;��I;��I;"�I;)KI;�H;��H;�H;N�G;[!G;��F;i�F;      ��?;�@;�@;�A;��B;�C;!CE;yvF;��G;�\H;t�H;�mI;^�I; �I; �I;��I;��I;_�I;kpI;R[I;DII;�9I;`,I;� I;oI;UI;�I;�I;g�H;��H;��H;.�H;R�H;��H;��H;Z�H;1�H;Z�H;��H;��H;U�H;-�H;��H;��H;c�H;�I;�I;ZI;kI;� I;e,I;�9I;FII;V[I;opI;Z�I;��I;��I;�I; �I;_�I;�mI;u�H;�\H;��G;zvF;&CE;��C;��B;�A;�@;�@;      2�1;��1;�73;�25;w�7;��:;+|=;#Q@;X�B;AE;��F;ZH;��H;qI;ƶI;��I;��I;�I;L�I;�vI;|_I;�KI;;I;�,I;� I;I;�I;I;qI;��H;q�H;q�H;!�H;��H;n�H;��H;��H;��H;j�H;��H;$�H;n�H;u�H;��H;pI;I;�I;I;� I;�,I;;I;�KI;|_I;�vI;R�I;	�I;��I;��I;ƶI;qI;��H;WH;��F;EE;T�B; Q@;0|=;��:;��7;�25;�73;��1;      d�;v�;�\;BX;�n!;�8';bI-;�93;��8;|=;lA;LzD;b�F;�/H;�I;ƔI;��I;h�I;ֵI;��I;wzI;oaI;nLI;;I;a,I;& I;I;�I;;I;�I;v�H;��H;d�H;l�H;
�H;S�H;#�H;R�H;�H;j�H;d�H;�H;z�H;�I;7I;�I; I;, I;^,I;;I;rLI;qaI;{zI;��I;ܵI;c�I;��I;ĔI;�I;�/H;f�F;IzD;lA;|=;��8;�93;dI-;�8';�n!;DX;�\;b�;      To�:���:=K�:�Y�:@��:�;�;��;��$;�G.;P6;j�<;'�A;�E;SG;�H;mI;~�I;A�I;J�I;��I;�{I;maI;�KI;�9I;�*I;�I;�I;�I;!I;� I;��H;��H;j�H;��H;�H;��H;�H;��H;j�H;��H;��H;� I;'I;�I;�I;�I;�*I;�9I;�KI;qaI;�{I;��I;O�I;E�I;{�I;mI;�H;SG;�E;(�A;g�<;P6;�G.;��$;��;�;�;n��:�Y�:;K�:p��:       %m8`��8�_u9x��9H�9:��:�W�::r�:@� ;�F;6o!;n�-;�^7;Kl>;�NC;�uF;KQH;�II;��I;��I;��I;��I;tzI;{_I;?II;B7I;Z(I;^I;�I;I;�I;* I;r�H;��H;�H;��H;t�H;��H;��H;��H;r�H;) I;�I;I;�I;`I;b(I;H7I;<II;_I;wzI;��I;��I;��I;��I;�II;NQH;�uF;�NC;Ll>;�^7;n�-;9o!;�F;=� ;Dr�:�W�:��:��9:���9�`u9���8      ��.��i�^�غp����*� ح�В�9D��::��:f��:�/;d�$;��1;g;;��A;��E;�H;,5I;5�I;��I;J�I;��I;�vI;O[I;WEI;�3I;2%I;�I;�I;P	I;�I;|�H;a�H;%�H;��H;o�H;��H;"�H;]�H;|�H;�I;S	I;�I;�I;4%I;�3I;[EI;L[I;�vI;��I;L�I;��I;6�I;05I;�H;��E;��A;g;;��1;e�$;�/;l��:6��:<��:���9�׭�(�*�\���r�غi�4��      ��ͻNɻ�����d�����C�]�� ��潺���H8�9���:'T�:�;�Y;I-;r9;X�@;�\E;��G;.5I;��I;C�I;յI;N�I;epI;�UI;O@I;0/I;{!I;�I;?I;�I;�I;!�H;��H;�H;��H;�H;��H;�H;�I;�I;CI;�I;z!I;2/I;S@I;�UI;apI;U�I;صI;D�I;��I;25I;��G;�\E;Y�@;o9;I-;�Y;�;'T�:���:H8�9����潺� �F�]�����d������Jɻ      �iO�ޔK��o@���.���������ɻ H��ooE���غ8(�����9�p�:�B�:�;l*;��7;�P@;�\E;�H;�II;|�I;d�I;�I;Y�I;7hI;�NI;_:I;7*I;tI;�I;�I;I;I;/�H;^�H;��H;a�H;,�H;I;I;�I;�I;xI;7*I;`:I;�NI;:hI;U�I;�I;f�I;�I;�II;�H;�\E;�P@;��7;j*;�;�B�:�p�:���9((����غooE�H���ɻ���������.��o@�ޔK�      L�����3���?����N��Pp��D����jG�����74�H�����n8��:;�:GG;�(;��7;U�@;��E;KQH;mI;�I;��I;��I;}I;�^I;�FI;�3I;�$I;\I;�I;�	I;I;�I;��H;R�H;��H;�I;I;�	I;�I;^I;�$I;�3I;�FI;�^I; }I;��I;��I;��I;mI;JQH;��E;X�@;��7;�(;EG;;�:��:��n8L���64�����hG່���D�Pp��N��@���4������      
��'�T5���������ϼ͡��X���iO�@���ɻ��p��D� �o��g:�_�:>G;j*;l9;��A;�uF;�H;��I;��I;��I;B�I;�pI;.TI;O>I;-I;�I;{I;�I;ZI;�I;�I;�I;�I;�I;SI;�I;xI;�I;-I;N>I;3TI;�pI;B�I;��I;��I;ÔI;�H;�uF;��A;l9;h*;AG;�_�:��g:��o��D⺝�p��ɻ@���iO�X��Ρ����ϼ������U5�'�      k��ҷ��&0v�s�a�#�G�?2+���؟�	����/����5��(��bf��ج��g:7�:�;I-;g;;�NC;SG;�I;ƶI;�I;��I;�I;cI;II;�5I;p&I;�I;5I;�I;�I;LI;ZI;NI;�I;�I;5I;�I;n&I;�5I;�II;	cI;�I;��I;�I;ɶI;�I;SG;�NC;g;;I-;�;9�:��g:�ج�bf�*�����5��/��	���؟���?2+�$�G�s�a�&0v�ҷ��      ��ս��ѽ=�ƽ1����I�����R�a�D4�<M���ϼ��J�K�O��PG��_f���o���:�B�:�Y;��1;Ol>;�E;�/H;qI;��I;��I;՘I;�rI;�UI;�>I;�-I;a I;�I;�I;�
I;I;0I;I;�
I;�I;�I;^ I;�-I;�>I;�UI;�rI;טI;��I;��I; qI;�/H;�E;Hl>;��1;�Y;�B�:��:��o�df�PG��O��J�K�����ϼ<M�D4�R�a�����I��1���=�ƽ��ѽ      �L+�  (���E�������ս�@���%���;V�&��ܐ�����MS�N��&��~D� �n8�p�:�;e�$;�^7;(�A;f�F;��H;b�I;]�I;��I;܃I;UbI;�HI;5I;%&I;-I;@I;�I;�
I;
I;�
I;�I;=I;-I;"&I;5I;�HI;UbI;݃I;��I;]�I;^�I;��H;h�F;*�A;�^7;i�$;�;�p�:��n8�D�(��N���MS�����ܐ�&���;V��%���@����ս����E���  (�      �T��f�����z��Yb�'�D��$�����ѽ�I��C�m�2+�������J�K�ﻙ�p�R���p��9#T�:�/;r�-;d�<;EzD;\H;�mI;��I;v�I;��I;�oI;�RI;�<I;,I;�I;I;/I;�I;�I;�I;-I;I;�I; ,I;�<I;�RI;�oI;��I;v�I;��I;�mI;ZH;KzD;d�<;j�-;�/;!T�:x��9P�����p��K�K�������2+�C�m��I����ѽ���$�'�D��Yb���z�f���      A�׾��Ҿž�j��������z�S�H�)��fz�H$���/v�2+�ݐ�����5��ɻ>4�h(��~��:^��:9o!;P6;lA;��F;s�H;��I;��I;ݦI;G}I;�\I;]DI;2I;p$I;�I;FI;�I;�I;�I;FI;�I;p$I;2I;[DI;�\I;I}I;ߦI;��I;��I;n�H;��F;lA;P6;/o!;`��:x��:p(��<4��ɻ��5���ݐ�2+��/v�H$��fz�)��T�H���z������j��ž��Ҿ      H(��$�d��Q������~���`���Yb���'��U�H$��C�m�&����ϼ�/��?��������غ88�9:��:�F;�G.;|=;GE;�\H;�I;q�I;u�I;��I;gI;LI;�7I;)I;pI;oI;oI;%I;qI;qI;nI;)I;�7I; LI;gI;��I;x�I;q�I;�I;�\H;HE;|=;�G.;�F;<��: 8�9��غ����?���/����ϼ&��C�m�H$���U���'��Yb��`���~�����Q��d���$�      ;�}���w�#f���K�q,�}�
�<�׾ �����k���'�fz꽝I���;V�=M�
����iO�mG�woE�̱�6��:B� ;��$;��8;Y�B;��G;)KI;�I;�I;@�I;qI;�SI;�=I;�-I;"I;iI;I;�I;I;jI;"I;�-I;�=I;�SI;qI;@�I;�I;�I;.KI;��G;\�B;��8;��$;:� ;<��:Ա�voE�lG໬iO�
���=M��;V��I��fz���'���k� ���<�׾}�
�q,���K�#f���w�      ��q�������.蒿��w��F�d��ʰ� ����Yb�)����ѽ�%��D4�ٟ� X�����
H���潺���9Dr�:��;�93;%Q@;|vF;�H;�I;��I;��I;�zI;�ZI;CI;�1I;b%I;?I;�I;!I;�I;@I;a%I;�1I;CI;�ZI;�zI;��I;��I;�I;�H;yvF;$Q@;�93;��;2r�:���9�潺H����� X��ٟ�D4��%����ѽ)���Yb� ���ʰ�d���F���w�.蒿����q���      3��������㿊�ɿ���ʅ����P�d��<�׾�`��S�H����@��R�a���Ρ���D��ɻ� �`ح��W�:�;^I-;5|=;CE;��H;�I;��I;s�I;��I;haI;HI;�5I;o(I;�I;�I;PI;�I;�I;o(I;�5I; HI;eaI;��I;r�I;��I;�I;��H;CE;7|=;`I-;�;�W�:`ح�� ��ɻ�D�Ρ����R�a��@����S�H��`��<�׾d����P�ʅ�������ɿ�㿳���      Ǚ$��x �#��:���޿p���ʅ���F�}�
��~����z��$���ս���@2+���ϼPp�����R�]� �*���:�;�8';��:;��C;�H;�}I;�I;p�I;׋I;kgI;�LI;9I;6+I;"I;�I;)I;�I;"I;4+I;9I;�LI;ggI;֋I;o�I;�I;�}I;H;��C;��:;�8';�;��: �*�U�]�����Pp���ϼ@2+������ս�$���z��~��}�
��F�ʅ��p����޿:��#���x �      J�Q���K���;�Ǚ$��;
��޿�����w�q,���澝���'�D������I��$�G�����N��������\�����9:T��:�n!;��7;��B;F�G;�YI;'�I;W�I;��I;�lI;rPI;<I;�-I;$I;�I;�I;�I;$I;�-I;<I;pPI;�lI;��I;W�I;*�I;�YI;P�G;��B;��7;�n!;R��:l�9:X����������N�����$�G��I������'�D��������q,���w�����޿�;
�Ǚ$���;���K�      T����{���d��F�Ǚ$�:����ɿ.蒿��K�Q���j���Yb�E�1���s�a����?�����.��d��t�غ���9�Y�:*X;�25;�A;T!G;E7I;p�I;@�I;O�I;�pI;�SI;|>I;y/I;�%I;" I;/I; I;�%I;v/I;>I;�SI;�pI;S�I;B�I;s�I;F7I;_!G;�A;�25;&X;�Y�:x��9r�غ�d����.�?������s�a�1���E��Yb��j��Q����K�.蒿��ɿ:��Ǚ$��F���d��{�      ����#P�������d���;�#���㿳���#f�d��ž��z���=�ƽ&0v�U5�2����o@������i��`u97K�:];�73;�@;��F;EI;��I;M�I;R�I;�sI;�UI;>@I;�0I;�&I;!I;0I;!I;�&I;�0I;?@I;�UI;�sI;V�I;M�I;��I;EI;��F;�@;�73;];3K�:0`u9|i������o@�2���U5�&0v�=�ƽ����z�žd��#f�������#����;���d����#P��      �,��a��#P���{���K��x �����q�����w��$���Ҿg���  (���ѽҷ��(�����K�Hɻ.�� ��8p��:v�;��1;�@;g�F;I;ۿI;�I;��I;�uI;#WI;eAI;�1I;�'I;�!I;�I;�!I;�'I;�1I;fAI;&WI;�uI;��I;�I;޿I;I;u�F;�@;��1;p�;j��: ��8,��Iɻ�K����(�ҷ����ѽ  (�g�����Ҿ�$���w�q��������x ���K��{�#P��a��      ඕ�S���Ѭ��-�_���7�{�}߿����,b��V�.l¾Gx�d.���Ž��t�*��g����?� N��-�� �x9���:L�;��2;/@@;\fF;5�H;}�I;O�I;|I;�[I;�CI;2I;�%I;[I;�I;0I;�I;ZI;�%I;2I;�CI;�[I;"|I;L�I;~�I;6�H;ifF;.@@;��2;B�;���:Ђx9*�� N����?�g��*����t���Žd.�Gx�.l¾�V��,b����}߿{���7�-�_�Ѭ��S���      S���E���$}��+Y��3�����$ڿ&��Ľ\����(���s��3�6����p�d�V���<<�<������@��9A��:˻;N%3;Ap@;�yF;��H;��I;��I;�{I;K[I;NCI;�1I;Q%I;I;WI;I;SI;I;P%I;�1I;OCI;E[I;�{I;ߛI;��I;��H;�yF;Ap@;J%3;Ļ;7��:��9����<���<<�V��d��p�5����3��s�(�����Ľ\�&���$ڿ����3��+Y�$}�E���      Ѭ��$}�>tf��lG�ע%��p�/�ʿZ����>M����V�����d�ɤ�̷�/�d��
��I���1�j���n�຀��9���:;�U4;��@;ϱF;/�H;׎I;��I;�yI;�YI;7BI;�0I;�$I;�I;�I;I;�I;�I;�$I;�0I;7BI;�YI;�yI;��I;ڎI;,�H;ٱF;��@;�U4;;x��:`��9f��k����1��I���
�/�d�̷�ɤ���d�V�������>M�Z���/�ʿ�p�ע%��lG�>tf�$}�      -�_��+Y��lG�f.�{���꿱���M䂿��5���󾌰��O�N�V��S��"�Q����~���i!��g��x�T	:O
�:��;Z16;��A;6G;�I;5�I;t�I;jvI;HWI;i@I;k/I;�#I;�I;
I;�I;I;�I;�#I;j/I;i@I;DWI;lvI;u�I;3�I;�I;?G;��A;V16;��;I
�:<	:r񳺐g��i!�~������"�Q�S��V��O�N���������5�M䂿�������{�f.��lG��+Y�      ��7��3�ע%�{��<����ſ
���½\�<����Ͼ����`�3��轼z��~�9�`�Ἔ���z��7}��dt� �^:U+�:��#;��8;��B;sG;m%I;��I;�I;rI;TI;�=I;p-I;"I;HI;�I;zI;�I;JI;"I;p-I;�=I;
TI;	rI;�I;��I;k%I;sG;��B;��8;��#;Q+�:��^:�dt��7}��z����`��~�9��z����`�3�������Ͼ<��½\�
�����ſ�<��{�ע%��3�      {�����p������ſ%���Ps���1�1r���d���d�}I�ψŽ��}�`*�KC��!�^��B黃�D�@Gไ �:��;j);7;;%D;/�G;SHI;��I;��I;�lI;�OI;�:I;+I; I;�I;yI;*I;uI;�I; I;+I;�:I;�OI;�lI;��I;��I;NHI;7�G;#D;7;;f);��;v �:0Gไ�D��B�!�^�LC��`*���}�ΈŽ}I��d��d��1r����1��Ps�%����ſ��꿃p����      }߿�$ڿ.�ʿ����
����Ps�PX:����&l¾�ǆ���7����85���Q�����t���75�m�������8�ɼ:��;��.;��=;�EE;�YH;�hI; �I;��I;$fI;KI;"7I;C(I;�I;�I;�I;vI;�I;�I;�I;C(I;!7I;KI;(fI;��I; �I;�hI;�YH;�EE;��=;��.;��;�ɼ: �8���o���75��t������Q�85�������7��ǆ�&l¾���PX:��Ps�
�������.�ʿ�$ڿ      ���&��Z���M䂿½\���1�����J˾青�E�N�x��I������V�'�e�Ҽ��|��z��n��Xx����&:�P�:��;�W4;ˠ@;gF;]�H;�I;�I;.�I;_I;�EI;3I; %I;AI;�I;�I;�I;�I;�I;BI;%I; 3I;�EI;_I;.�I;�I;�I;`�H;!gF;Ơ@;�W4;��;�P�:��&:Xx���n���z���|�e�ҼV�'����I���x��E�N�青��J˾�����1�½\�M䂿Z���&��      �,b�Ľ\��>M���5�<��1r��&l¾青�"&W��3�8Sؽ�z��[G����|I����?���̻��-��
����:��;��&;|9;�C;�dG;GI;=�I;M�I;OvI;{WI;'@I;�.I;�!I;�I;VI;�I;�I;�I;VI;�I;�!I;�.I;&@I;|WI;OvI;P�I;:�I;GI;�dG;�C;|9;��&;��;��:�
����-���̻��?�|I�����[G��z��8Sؽ�3�"&W�青�&l¾1r��<����5��>M�Ľ\�      �V������������Ͼ�d���ǆ�E�N��3��c�[����\�4��*C���o���	�숻`�h��9��:�h;K�/;2�=;CE;�2H;�WI;��I;�I;�kI;�OI; :I;�)I;"I;�I;�I;�I;xI;�I;�I;�I;"I;�)I;!:I;�OI;�kI;��I;��I;�WI;�2H;AE;5�=;L�/;zh;��:h��9d�숻��	��o�*C��3����\�[���cཱ3�E�N��ǆ��d����Ͼ���������      .l¾(��V������������d���7�x��8Sؽ[���d�D*�dkּ.\����'�.���R�h~��h�:�Z;̣#;8=7;$�A;�F;Q�H;k�I;�I;��I;�`I;�GI;�3I;&%I;rI;�I;SI;K
I;J	I;M
I;TI;�I;rI;#%I;�3I;�GI;�`I;��I;�I;h�I;T�H;�F;&�A;8=7;ʣ#;�Z;j�:�~���R�.����'�-\��dkּD*��d�[��8Sؽx����7��d���������V���(��      Gx��s���d�O�N�`�3�}I����H����z����\�D*��ݼJ���1<<��ڻ�V�`dt��&:z��:4C;�</;LD=;ψD;��G;�8I;ØI;��I;tI;$VI;Z?I;�-I;b I;�I;YI;�
I;�I;I;�I;�
I;\I;�I;` I;�-I;^?I;+VI;tI;��I;��I;�8I;��G;ӈD;MD=;�</;>C;z��:�&:Xdt��V��ڻ0<<�J����ݼC*���\��z��H������|I�`�3�O�N���d��s�      c.��3�Ȥ�V����ΈŽ85�����ZG�3��dkּJ���yC��>�p6}����p�x9\��:	;(�&;�;8;��A;��F;��H;.yI;��I;�I;.fI;�KI;I7I;{'I;�I;�I;XI;I;�I;�I;�I;I;WI;�I;�I;'I;P7I;�KI;0fI;�I;��I;2yI;��H;��F;��A;�;8;0�&;	;P��:��x9���p6}��>�yC�J���dkּ3��ZG����85��ΈŽ��V��Ȥ��3�      ��Ž5���̷�S���z����}��Q�V�'����)C��-\��1<<��>n��R��@�"��:"��:�;�'3;��>;�E;bH;]<I;ȗI;��I;�vI;�XI;�AI;t/I;�!I;�I;�I;S	I;cI;#I;tI;#I;bI;S	I;�I;�I;�!I;{/I;�AI;�XI;�vI;��I;͗I;Z<I;dH;�E;��>;�'3;�;��:*��:��R�ຈn���>�0<<�-\��*C�����V�'��Q���}��z��S��̷�5���      ��t��p�/�d�!�Q�}�9�_*����c�Ҽ|I���o���'��ڻq6}�T���9���:Jm�:��;��.;<;�oC;:7G;��H;сI;ќI;хI;fI;;LI;�7I;�'I;�I;rI;LI;HI;�I;� I;P I;� I;�I;HI;NI;qI;�I;�'I;�7I;ALI;fI;˅I;ӜI;ρI;��H;<7G;�oC;<;��.;��;Pm�:��:�9�N��p6}��ڻ��'��o�{I��d�Ҽ���_*�~�9�!�Q�/�d��p�      )��c��
����`��KC���t����|���?���	�,���V�*�������:��:�h;�+;��9;��A;ufF;T�H;p_I;��I;��I;sI;�VI;p@I;�.I;� I;TI;I;�I;jI;O I;~�H;�H;|�H;L I;hI;�I;	I;XI;� I;�.I;u@I;�VI;�rI;��I;��I;p_I;V�H;wfF;��A;��9;�+;�h;��:��:��,����V�+����	���?���|��t��JC��a������
�b�      d��T���I��~������ �^��75��z���̻�눻�R�\dt���x9*��:Rm�:�h;W�*;؍8;��@;ڼE;3(H;b8I;��I;�I;E~I;�`I;�HI;�5I;Y&I;rI;2I;�	I;�I;� I;��H;W�H;��H;S�H;��H;� I;�I;�	I;5I;uI;Y&I;�5I;�HI;�`I;K~I;�I;��I;d8I;5(H;߼E;��@;э8;X�*;�h;Tm�:.��:p�x9Pdt��R��눻��̻�z��75� �^����~����I��R��      ��?��<<��1��h!��z��B�h���n����-�V�`~�� �&:J��:��:��;�+;Ѝ8;:�@;�]E;a�G;@I;�I;L�I;3�I;giI;7PI;<I;�+I;�I;nI;MI;(I;qI;��H;��H;Q�H;��H;N�H;��H;��H;oI;'I;SI;rI;�I;�+I;<I;1PI;kiI;1�I;H�I;�I;BI;f�G;�]E;6�@;ҍ8;�+;��;��:N��:�&:H~��V𳺎�-��n��j���B黶z� i!��1��<<�      N��A��i����g���7}�s�D����Dx���
�����9v�:x��:	;�;��.;��9;��@;�]E;e�G;8I;�I;��I;H�I;�pI;~VI;�AI;z0I;�"I;�I;�I;�I;�I;��H;]�H;v�H;^�H;��H;]�H;s�H;\�H;��H;�I;�I;�I;�I;�"I;y0I;�AI;�VI;�pI;C�I;�I;�I;:I;f�G;�]E;��@;��9;��.;�;	;|��:x�:���9�
��Jx�����y�D��7}��g��i���@��      ,������R��Z��dt�G�@�8��&:��:��:�Z;;C;+�&;�'3;<;��A;ܼE;h�G;9I;T|I;��I;��I;zuI;n[I;FI;�4I;(&I;�I;GI;�	I;�I;9�H;��H;5�H;r�H;|�H;�H;w�H;o�H;4�H;��H;4�H;�I;�	I;DI;�I;'&I;~4I;FI;n[I;vuI;��I;��I;U|I;<I;d�G;޼E;��A;<;�'3;+�&;?C;�Z;��:��:��&:��8�F๬dt�r�l��ʎ��      0�x9���9���94	:��^:~ �:�ɼ:�P�:��;h;̣#;�</;�;8;��>;�oC;xfF;3(H;GI;�I;��I;��I;�wI;k^I;6II;�7I;)I;I;�I;�I;FI;J I;H�H;Q�H;9�H;��H;��H;��H;��H;��H;7�H;P�H;B�H;M I;GI;�I;�I;I;)I;�7I;4II;f^I;�wI;��I;��I;�I;CI;5(H;xfF;�oC;��>;�;8;�</;У#;h;��;�P�:�ɼ:v �:��^:<	:��9ؖ�9      ���:_��:���:e
�:G+�:��;��;��;��&;M�/;:=7;JD=;��A;�E;:7G;X�H;e8I;�I;�I;��I;�wI;�_I;�JI;�9I;�*I;�I;2I;9I;~I;8I;��H;��H;�H;;�H;��H;�H;��H;�H;��H;;�H;�H;��H;��H;8I;{I;9I;/I;�I;�*I;�9I;�JI;�_I;�wI;��I;�I;�I;g8I;V�H;<7G;�E;��A;OD=;<=7;K�/;��&;��;��;��;y+�:U
�:���:K��:      `�;˻;;��;��#;t);��.;�W4;!|9;7�=;+�A;ֈD;��F;kH;��H;u_I;��I;O�I;G�I;zuI;j^I;�JI;!:I;,I;4 I;|I;KI;�I; I;��H;��H;3�H;�H;j�H;b�H;��H;S�H;��H;`�H;k�H;�H;0�H;�H;��H;I;�I;JI;|I;5 I;,I;:I;�JI;k^I;yuI;H�I;J�I;��I;t_I;��H;gH;��F;׈D;1�A;3�=;|9;�W4;��.;n);��#;��;;��;      ��2;V%3;�U4;R16;��8;7;;��=;ɠ@;�C;CE;�F;��G;��H;]<I;΁I;��I;�I;3�I;�pI;j[I;4II;�9I;,I;� I;I;I;PI;�I;G�H;c�H;Z�H;(�H;9�H;��H;��H;^�H;��H;X�H;��H;��H;9�H;&�H;]�H;`�H;C�H;�I;LI;I;I;� I;,I;�9I;2II;g[I;�pI;.�I;�I;��I;΁I;X<I;��H;��G;�F;BE;�C;Ϡ@;��=;7;;��8;S16;�U4;O%3;      P@@;Cp@;��@;��A;��B;0D;�EE;"gF;�dG;�2H;X�H;�8I;/yI;җI;؜I;��I;O~I;qiI;�VI;FI;�7I;�*I;8 I;!I;YI;�I;;I;��H;��H;��H;�H;!�H;��H;n�H;��H;"�H;��H;�H;��H;o�H;��H;�H;�H;��H;��H;��H;6I;�I;ZI;I;5 I;�*I;�7I;FI;�VI;niI;R~I;��I;؜I;їI;0yI;�8I;[�H;�2H;�dG;!gF;�EE;&D;��B;��A;��@;Ap@;      [fF;�yF;ұF;4G;�rG;;�G;�YH;j�H;HI;�WI;n�I;˘I;��I;��I;ЅI;sI;�`I;5PI;�AI;~4I;)I;�I;{I;I;�I;OI;��H;��H;��H;S�H;,�H;e�H;�H;*�H;q�H;�H;�H;	�H;n�H;*�H;�H;_�H;,�H;Q�H;��H;��H;��H;RI;�I;I;xI;�I;)I;|4I;�AI;1PI;�`I;sI;ЅI;��I;��I;ʘI;v�I;�WI;KI;h�H;�YH;0�G;sG;FG;ұF;�yF;      F�H;��H;+�H;�I;c%I;SHI;�hI;�I;@�I;��I;�I;��I;�I;�vI;fI;�VI;�HI;<I;}0I;+&I;I;/I;MI;VI;7I;��H; �H;��H;h�H;0�H;j�H;��H;��H;�H;h�H;�H;�H;�H;e�H;�H;��H;��H;j�H;-�H;b�H;��H;��H;��H;:I;OI;KI;1I;I;'&I;|0I;�;I;�HI;�VI;fI;�vI;�I;��I;�I;��I;<�I;�I;�hI;MHI;x%I;�I;*�H;��H;      ��I;��I;ՎI;:�I;��I;��I;*�I;�I;Q�I;��I;��I;tI;+fI;�XI;:LI;s@I;�5I;�+I;�"I;�I;�I;5I;�I;�I;��H;��H;��H;^�H;E�H;[�H;��H;��H;��H;��H;��H;>�H;#�H;:�H;��H;��H;��H;��H;��H;Z�H;A�H;\�H;��H;��H;��H;�I;�I;6I;�I;�I;�"I;�+I;�5I;u@I;;LI;�XI;-fI;tI;��I;��I;Q�I;�I;*�I;��I;��I;?�I;ӎI;�I;      N�I;ۛI;��I;��I;הI;��I;��I;4�I;IvI;�kI;�`I;+VI;�KI;�AI;�7I;�.I;_&I;�I;�I;JI;�I;xI;I;G�H;��H;��H;_�H;E�H;_�H;��H;��H;��H;��H;#�H;��H;�H;N�H;{�H;��H;#�H;��H;��H;��H;��H;[�H;D�H;\�H;��H;��H;A�H;I;xI;�I;FI;�I;�I;_&I;�.I;�7I;�AI;�KI;+VI;�`I;�kI;LvI;4�I;��I;��I;�I;��I;��I;כI;      |I;�{I;�yI;evI;rI;�lI;'fI;!_I;}WI;�OI;�GI;d?I;N7I;|/I;�'I;� I;wI;iI;�I;�	I;MI;4I;��H;b�H;��H;J�H;0�H;^�H;��H;��H;��H;��H;��H;�H;�H;��H;��H;��H;	�H;�H;��H;��H;��H;��H;��H;\�H;*�H;N�H;��H;]�H;��H;6I;GI;�	I;�I;hI;xI;� I;�'I;y/I;O7I;a?I;�GI;�OI;}WI;_I;+fI;�lI;rI;ovI;�yI;�{I;      �[I;`[I;�YI;PWI;
TI;�OI;KI;�EI;-@I;':I;�3I;�-I;�'I;�!I;�I;XI;9I;QI;�I;�I;T I;��H;��H;]�H;�H;*�H;m�H;��H;��H;��H;}�H;��H;U�H;��H;u�H;Y�H;R�H;V�H;r�H;��H;W�H;��H;~�H;��H;��H;��H;j�H;,�H;�H;Z�H;�H;��H;P I;�I;�I;QI;;I;[I;�I;�!I;�'I;�-I;�3I;(:I;.@I;�EI;#KI;�OI;TI;SWI;�YI;`[I;      �CI;UCI;6BI;a@I;�=I;�:I;7I;3I;�.I;�)I;#%I;g I;�I;�I;rI;I;�	I;)I;�I;=�H;P�H;��H;0�H;'�H;!�H;\�H;��H;��H;��H;��H;��H;B�H;��H;M�H;�H;��H;��H;��H;�H;N�H;��H;@�H;��H;��H;��H;��H;��H;_�H;"�H;�H;3�H;��H;I�H;7�H;�I;,I;
I;I;uI;�I;�I;e I;+%I;�)I;�.I;3I;*7I;�:I;�=I;i@I;=BI;UCI;      2I;�1I;�0I;k/I;m-I;
+I;>(I;%I;�!I;I;rI;�I;�I;�I;LI;�I;�I;qI;��H;��H;^�H;�H;�H;7�H;��H;�H;��H;��H;��H; �H;S�H;��H;2�H;��H;��H;}�H;m�H;}�H;��H;��H;2�H;��H;P�H;��H;��H;��H;��H;�H;��H;6�H;�H;�H;U�H;��H;��H;qI;�I;�I;OI;�I;�I;�I;xI; I;�!I;%I;C(I;+I;s-I;j/I;�0I;�1I;      �%I;M%I;�$I;�#I;	"I; I;�I;GI;�I;�I;�I;aI;]I;X	I;KI;kI;� I;��H;a�H;;�H;A�H;<�H;g�H;��H;l�H;%�H;�H;�H;)�H;��H;��H;O�H;��H;��H;\�H;6�H;$�H;6�H;[�H;��H;��H;O�H;��H;}�H;"�H;��H;�H;&�H;l�H;��H;k�H;;�H;;�H;4�H;^�H;��H;� I;nI;NI;X	I;]I;aI;�I;�I;�I;DI;�I; I;"I;�#I;�$I;Z%I;      NI;4I;�I;�I;TI;�I;�I;�I;YI;�I;\I;�
I;I;jI;�I;P I;��H;��H;v�H;v�H;��H;��H;]�H;��H;��H;g�H;c�H;��H;��H;�H;n�H;�H;��H;[�H;�H;�H;�H;�H;�H;\�H;��H;�H;m�H;	�H;��H;��H;c�H;i�H;��H;��H;`�H;��H;��H;o�H;t�H;��H;��H;S I;�I;jI;I;�
I;_I;�I;[I;�I;�I;�I;QI;�I;�I;5I;      �I;ZI;�I;I;�I;pI;�I;�I;�I;�I;O
I;�I;�I;&I;� I;{�H;V�H;K�H;a�H;|�H;��H;�H;��H;P�H;�H;�H;�H;A�H;��H;��H;V�H;��H;��H;8�H;�H;��H;��H;��H;�H;<�H;��H;��H;U�H;��H;��H;<�H;�H;�H;�H;P�H;��H;�H;��H;w�H;`�H;O�H;Z�H;~�H;� I;(I;�I;�I;T
I;�I;�I;�I;�I;rI;�I;I;�I;hI;      6I;�I;�I;�I;rI;"I;xI;�I;�I;vI;S	I;I;�I;{I;V I;�H;��H;��H;��H; �H;��H;��H;P�H;��H;��H;�H;�H;*�H;V�H;��H;M�H;��H;o�H; �H;�H;��H;��H;��H;�H;!�H;q�H;��H;M�H;��H;O�H;&�H;�H;	�H;��H;��H;S�H;��H;��H;�H;��H;��H;��H;�H;W I;|I;�I;I;W	I;xI;�I;�I;~I;"I;pI;�I;�I;	I;      �I;]I;�I;I;�I;sI;�I;�I;�I;�I;N
I;�I;�I;(I;� I;{�H;V�H;K�H;`�H;{�H;��H;�H;��H;O�H;�H;�H;�H;?�H;��H;��H;V�H;��H;��H;8�H;�H;��H;��H;��H;�H;;�H;��H;��H;U�H;��H;��H;;�H;�H;�H;�H;P�H;��H;
�H;��H;w�H;`�H;O�H;W�H;~�H;� I;%I;�I;�I;T
I;�I;�I;�I;�I;rI;�I;	I;�I;dI;      FI;6I;�I;�I;TI;�I;�I;�I;YI;�I;[I;�
I;I;iI;�I;P I;��H;��H;v�H;u�H;��H;��H;\�H;��H;��H;d�H;c�H;��H;��H;�H;m�H;�H;��H;[�H;�H;�H;�H;�H;�H;\�H;��H;�H;m�H;�H;��H;��H;e�H;j�H;��H;��H;`�H;��H;��H;o�H;t�H;��H;��H;S I;�I;jI;I;�
I;_I;�I;YI;�I;�I;�I;TI;�I;�I;8I;      �%I;N%I;�$I;�#I;	"I; I;�I;II;�I;�I;�I;`I;[I;W	I;MI;kI;� I;��H;`�H;8�H;@�H;;�H;e�H;��H;n�H;#�H;�H; �H;)�H;��H;��H;O�H;��H;��H;^�H;5�H;$�H;8�H;[�H;��H;��H;O�H;��H;}�H;"�H;��H;�H;(�H;n�H;��H;k�H;;�H;9�H;5�H;`�H;��H;� I;nI;NI;X	I;[I;`I;�I;�I;�I;HI;�I; I;"I;�#I;�$I;P%I;      2I;�1I;�0I;h/I;l-I;+I;<(I;!%I;�!I;I;qI;�I;�I;�I;OI;�I;�I;qI;��H;��H;\�H;�H;�H;4�H;��H;�H;��H;��H;��H;��H;P�H;��H;0�H;��H;��H;~�H;m�H;~�H;��H;��H;0�H;��H;P�H;��H;��H;��H;��H;�H;��H;3�H;	�H;�H;T�H;��H;��H;pI;�I;�I;OI;�I;�I;�I;uI;I;�!I;%I;E(I;	+I;p-I;o/I;�0I;�1I;      �CI;YCI;'BI;a@I;�=I;�:I;&7I;3I;�.I;�)I;'%I;g I;�I;�I;tI;I;�	I;,I;�I;:�H;P�H;��H;/�H;!�H;!�H;\�H;��H;��H;��H;��H;��H;A�H;��H;K�H;�H;��H;��H;��H;�H;M�H;��H;A�H;��H;��H;��H;��H;��H;^�H;�H;�H;6�H;��H;I�H;9�H;�I;)I;�	I;I;uI;�I;�I;g I;*%I;�)I;�.I;3I;(7I;�:I;�=I;l@I;.BI;SCI;      �[I;`[I;�YI;KWI;TI;�OI;KI;�EI;*@I;$:I;�3I;�-I;�'I;�!I;�I;YI;;I;SI;�I;�I;T I;��H;��H;Z�H;�H;&�H;h�H;��H;��H;��H;}�H;��H;V�H;��H;x�H;X�H;R�H;[�H;r�H;��H;W�H;��H;}�H;��H;��H;��H;j�H;,�H;�H;Y�H;�H; �H;O I;�I;�I;PI;<I;YI;�I;�!I;�'I;�-I;�3I;':I;.@I;�EI;"KI;�OI;TI;VWI;�YI;a[I;      (|I;�{I;�yI;qvI;�qI;�lI;%fI;#_I;}WI;�OI;�GI;a?I;L7I;y/I;�'I;� I;wI;kI;�I;�	I;MI;5I;��H;]�H;��H;G�H;,�H;\�H;��H;��H;��H;��H;��H;�H;�H;��H;��H;��H;
�H;�H;��H;��H;��H;��H;��H;\�H;-�H;M�H;��H;\�H;��H;6I;GI;�	I;�I;gI;wI;� I;�'I;{/I;N7I;^?I;�GI;�OI;{WI;"_I;+fI;�lI;rI;xvI;�yI;�{I;      Y�I;ۛI;��I;~�I;ɔI;��I;��I;2�I;OvI;�kI;�`I;+VI;�KI;�AI;�7I;�.I;]&I;�I;�I;FI;�I;wI;I;D�H;��H;��H;\�H;D�H;_�H;��H;��H;��H;��H;%�H;��H;�H;O�H;��H;��H;#�H;��H;��H;��H;��H;[�H;B�H;_�H;��H;��H;@�H;I;zI;�I;FI;�I;�I;]&I;�.I;�7I;�AI;�KI;(VI;�`I;�kI;MvI;5�I;��I;��I;ڔI;��I;��I;қI;      ��I;�I;ŎI;:�I;��I;��I;*�I;#�I;N�I;��I;��I;tI;-fI;�XI;<LI;u@I;�5I;�+I;�"I;�I;�I;5I;�I;�I;��H;��H;��H;[�H;G�H;X�H;��H;��H;��H;��H;��H;<�H;'�H;>�H;��H;��H;��H;��H;��H;[�H;B�H;[�H;��H;��H;��H;�I;�I;5I;�I;�I;�"I;�+I;�5I;u@I;<LI;�XI;-fI;tI;��I;��I;M�I;�I;*�I;��I;��I;?�I;ҎI;�I;      6�H;��H;'�H;
I;n%I;THI;�hI;�I;?�I;��I;�I;��I;�I;�vI;fI;�VI;�HI;<I;y0I;$&I;I;/I;GI;TI;7I;��H;��H;��H;f�H;-�H;i�H;��H;��H;�H;i�H;�H;�H;�H;e�H;�H;��H;��H;m�H;0�H;c�H;��H;��H;��H;9I;PI;OI;1I;	I;(&I;}0I; <I;�HI;�VI;fI;�vI;�I;��I;�I;��I;<�I;�I;�hI;NHI;u%I;I;(�H;��H;      QfF;�yF;رF;4G;sG;D�G;�YH;l�H;KI;�WI;q�I;˘I;��I;��I;ЅI;sI;�`I;5PI;�AI;|4I;)I;�I;wI;I;�I;KI;��H;��H;��H;P�H;,�H;e�H;�H;*�H;r�H;�H;�H;�H;n�H;*�H;�H;f�H;0�H;S�H;��H;��H;��H;OI;�I;I;|I;�I;)I;~4I;�AI;3PI;�`I;sI;҅I;��I;��I;ȘI;t�I;�WI;DI;d�H;�YH;0�G;sG;6G;��F;�yF;      M@@;>p@;~�@;��A;��B;4D;�EE;!gF;�dG;�2H;W�H;�8I;.yI;ΗI;ٜI;��I;O~I;qiI;�VI;FI;�7I;�*I;3 I;I;ZI;�I;4I;��H;��H;��H;�H;"�H;��H;n�H;��H;!�H;��H;!�H;��H;o�H;��H;"�H; �H;��H;��H;��H;:I;�I;YI;I;: I;�*I;�7I;FI;�VI;liI;R~I;��I;ٜI;ΗI;/yI;�8I;W�H;�2H;�dG;"gF;�EE;&D;��B;��A;}�@;@p@;      �2;=%3;�U4;_16;��8;$7;;��=;ˠ@;�C;?E;�F;��G;��H;W<I;ρI;��I;�I;2�I;�pI;e[I;2II;�9I;,I;� I;I;I;JI;�I;G�H;_�H;\�H;+�H;9�H;��H;��H;[�H; �H;^�H;��H;��H;;�H;+�H;a�H;c�H;F�H;�I;PI;I;I;� I;,I;�9I;4II;j[I;�pI;.�I;�I;��I;΁I;X<I;��H;��G;�F;AE;�C;Ơ@;��=;7;;��8;t16;�U4;(%3;      P�;ƻ;;�;��#;l);��.;�W4;$|9;6�=;'�A;׈D;��F;iH;��H;u_I;��I;L�I;D�I;wuI;i^I;�JI;:I;,I;5 I;uI;GI;�I;!I;��H;��H;6�H;�H;j�H;c�H;��H;U�H;��H;`�H;h�H;�H;6�H;�H;��H;I;�I;OI;zI;4 I;,I; :I;�JI;k^I;zuI;J�I;H�I;��I;u_I;��H;fH;��F;ԈD;*�A;6�=;!|9;�W4;��.;n);��#; �;;��;      v��:Y��:���:U
�:G+�:��;��;��;��&;I�/;9=7;PD=;��A;�E;<7G;W�H;b8I;�I;��I;��I;�wI;�_I;�JI;�9I;�*I;�I;.I;9I;|I;5I;��H;��H;�H;;�H;��H;�H;��H;�H;��H;9�H;�H;��H;�H;;I;|I;9I;5I;�I;�*I;�9I;�JI;�_I;�wI;��I;�I;�I;e8I;W�H;<7G;�E;��A;MD=;<=7;I�/;��&;��;��;w�;s+�:?
�:���:C��:      p�x9X��9��9<	:��^:� �:�ɼ:�P�:��;zh;ͣ#;�</;�;8;��>;�oC;xfF;3(H;CI;�I;��I;��I;�wI;d^I;2II;�7I;�(I; I;�I;�I;CI;J I;I�H;Q�H;;�H;��H;��H;��H;��H;��H;9�H;S�H;H�H;O I;II;�I;�I;I; )I;�7I;5II;i^I;�wI;��I;��I;�I;BI;6(H;zfF;�oC;��>;�;8;�</;У#;~h;��;�P�:�ɼ:~ �:�^:H	:���9薒9      ������d��T��dt��F���8��&:��:��:�Z;>C;+�&;�'3;<;��A;ܼE;d�G;6I;R|I;��I;��I;tuI;j[I;FI;z4I;!&I;�I;GI;�	I;�I;9�H;��H;6�H;r�H;x�H;�H;{�H;o�H;2�H;��H;:�H;�I;�	I;GI;�I;)&I;~4I;FI;o[I;zuI;��I;��I;U|I;:I;d�G;޼E;��A;<;�'3;)�&;;C;�Z;��:��:��&:��80G๬dt�j�f����      N��B��j����g���7}�r�D����Fx���
�����9r�:|��:	;
�;��.;��9;��@;�]E;b�G;8I;�I;��I;C�I;�pI;�VI;�AI;u0I;�"I;�I;�I;�I;�I;��H;]�H;v�H;^�H;��H;^�H;s�H;\�H;��H;�I;�I;�I;�I;�"I;z0I;�AI;~VI;�pI;F�I; �I;�I;:I;e�G;�]E;��@;��9;��.;
�;	;z��:r�:x��9�
��Bx�����v�D��7}��g��l���>��      ��?��<<�	�1� i!��z��B�h���n����-�V�P~���&:J��:��:��;�+;Ѝ8;6�@;�]E;c�G;?I;�I;J�I;/�I;jiI;0PI;�;I;�+I;�I;iI;PI;)I;pI;��H;��H;N�H;��H;R�H;��H;��H;qI;)I;SI;nI;�I;�+I;<I;1PI;giI;2�I;K�I;�I;@I;f�G;�]E;6�@;Ѝ8;�+;��;��:J��: �&:H~��Z𳺏�-��n��h���B黸z� i!��1��<<�      d��T���I��}������ �^��75��z���̻�눻�R�Ldt���x9(��:Xm�:�h;X�*;ҍ8;��@;ۼE;3(H;a8I;��I;�I;J~I;�`I;�HI;�5I;[&I;pI;2I;�	I;�I;� I;��H;V�H;��H;V�H;��H;� I;�I;�	I;5I;rI;[&I;�5I;�HI;�`I;E~I;�I;��I;d8I;2(H;߼E;��@;ҍ8;X�*;�h;Tm�:*��:��x9Xdt��R��눻��̻�z��75��^����~����I��S��      )��c��
����`��JC���t����|���?���	�,���V�*�������:��:�h;�+;��9;��A;wfF;T�H;p_I;��I;��I;�rI;�VI;o@I;�.I;� I;UI;I;�I;kI;O I;{�H;�H;~�H;J I;gI;�I;	I;UI;� I;�.I;r@I;�VI;�rI;��I;��I;r_I;V�H;sfF;��A;��9;�+;�h;��:��:��,����V�,����	���?���|��t��JC��a�����	�
�c�      ��t��p�/�d�!�Q�}�9�_*����c�Ҽ|I���o���'��ڻq6}�N�ະ9���:Lm�:��;��.;<;�oC;97G;��H;΁I;ҜI;ͅI;fI;:LI;�7I;�'I;�I;rI;LI;JI;�I;� I;P I;� I;�I;HI;LI;qI;�I;�'I;�7I;<LI;fI;ͅI;ϜI;сI;��H;<7G;�oC;<;��.;��;Rm�:��:�9�R��s6}��ڻ��'��o�|I��d�Ҽ���_*�~�9�!�Q�/�d��p�      ��Ž5���̷�S���z����}��Q�U�'����*C��-\��0<<��>n��F�຀�&��:��:	�;�'3;��>;�E;cH;]<I;͗I;��I;�vI;�XI;�AI;t/I;�!I;�I;�I;Q	I;aI;!I;tI;#I;^I;S	I;�I;�I;�!I;x/I;�AI;�XI;�vI;��I;ǗI;^<I;iH;�E;��>;�'3;	�; ��:*��:��R�ຈn���>�0<<�-\��*C�����V�'��Q���}��z��S��̷�5���      c.��3�ɤ�V����ΈŽ85�����ZG�3��dkּJ���yC��>�l6}������x9R��:	;+�&;�;8;��A;��F;��H;0yI;��I;�I;+fI;�KI;K7I;|'I;�I;�I;ZI;I;�I;�I;�I;I;WI;�I;�I;|'I;L7I;�KI;-fI;��I;��I;,yI;��H;��F;��A;�;8;/�&;	;P��:��x9"���o6}��>�yC�J���dkּ3��ZG����85��ΈŽ��V��ɤ��3�      Gx��s���d�O�N�`�3�}I����H����z����\�C*��ݼJ���0<<��ڻ�V�hdt���&:z��::C;�</;JD=;҈D;��G;�8I;ØI;��I;tI;%VI;W?I;�-I;a I;�I;\I;�
I;�I;I;�I;�
I;ZI;�I;` I;�-I;Z?I;(VI;tI;��I;ØI;�8I;��G;ԈD;JD=;�</;=C;x��: �&:`dt��V��ڻ1<<�J����ݼD*���\��z��H������}I�`�3�O�N���d��s�      .l¾(��V������������d���7�x��8Sؽ[���d�D*�dkּ.\����'�.���R��~��h�:�Z;Σ#;6=7;&�A;�F;T�H;k�I;�I;��I;�`I;�GI;�3I;&%I;rI;�I;SI;K
I;J	I;K
I;SI;�I;rI;#%I;�3I;�GI;�`I;��I;�I;k�I;Q�H;�F;'�A;5=7;ţ#;�Z;b�:�~���R�.����'�.\��dkּD*��d�[��8Sؽx����7��d���������V���(��      �V������������Ͼ�d���ǆ�E�N��3��c�[����\�3��*C���o���	�숻h�x��9	��:�h;K�/;3�=;BE;�2H;�WI;��I;�I;�kI;�OI;!:I;�)I;"I;�I;�I;�I;xI;�I;�I;�I;"I;�)I;!:I;�OI;�kI;�I;��I;�WI;�2H;BE;6�=;I�/;wh;��:P��9d�숻��	��o�*C��4����\�[���cཱ3�E�N��ǆ��d����Ͼ���������      �,b�Ľ\��>M���5�<��1r��&l¾青�"&W��3�8Sؽ�z��ZG����|I����?���̻��-��
��
��:��;��&;|9;�C;�dG;FI;:�I;L�I;OvI;yWI;)@I;�.I;�!I;�I;TI;�I;�I;�I;UI;�I;�!I;�.I;'@I;yWI;MvI;M�I;:�I;HI;�dG;�C;|9;��&;�;��:�
����-���̻��?�|I�����[G��z��8Sؽ�3�"&W�青�&l¾1r��<����5��>M�Ľ\�      ���&��Z���M䂿½\���1�����J˾青�E�N�x��I������V�'�e�Ҽ��|��z��n��Tx����&:�P�:��;�W4;̠@;!gF;Z�H;�I;�I;-�I;_I;�EI;3I;%I;AI;�I;�I;�I;�I;�I;AI; %I;3I;�EI;_I;-�I;�I;�I;^�H;gF;ˠ@;�W4;��;�P�:��&:Zx���n���z���|�e�ҼV�'����I���x��E�N�青��J˾�����1�½\�M䂿Z���&��      }߿�$ڿ.�ʿ����
����Ps�PX:����&l¾�ǆ���7����85���Q�����t���75�o����� �8�ɼ:��;��.;��=;�EE;�YH;�hI;�I;��I;%fI;KI;"7I;C(I;�I;�I;�I;tI;�I;�I;�I;C(I;"7I;KI;'fI;��I;!�I;�hI;�YH;�EE;��=;��.;��;�ɼ:`�8���n���75��t������Q�85�������7��ǆ�&l¾���PX:��Ps�
�������.�ʿ�$ڿ      {�����p������ſ%���Ps���1�1r���d���d�}I�ψŽ��}�`*�KC��!�^��B黃�D�(Gไ �:��;j);7;;#D;,�G;QHI;��I;��I;�lI;�OI;�:I;+I; I;�I;vI;*I;vI;�I; I;+I;�:I;�OI;�lI;��I;��I;PHI;6�G;#D;7;;h);��;z �:(Gไ�D��B� �^�KC��`*���}�ΈŽ}I��d��d��1r����1��Ps�%����ſ��꿃p����      ��7��3�ע%�{��<����ſ
���½\�<����Ͼ����`�3��轼z��~�9�`�Ἔ���z��7}��dt���^:U+�:��#;��8;��B;sG;k%I;��I;�I;rI;TI;�=I;o-I;"I;DI;�I;yI;�I;GI;"I;o-I;�=I;TI;	rI;�I;��I;n%I;sG;��B;��8;��#;U+�:��^:�dt��7}��z����`��~�9��z����`�3�������Ͼ<��½\�
�����ſ�<��{�ע%��3�      -�_��+Y��lG�f.�{���꿱���M䂿��5���󾌰��O�N�V��S��"�Q����~���i!��g��r�T	:M
�:��;X16;��A;4G;�I;3�I;t�I;hvI;IWI;h@I;h/I;�#I;�I;	I;�I;I;�I;�#I;k/I;k@I;GWI;nvI;t�I;5�I;�I;?G;��A;X16;��;I
�:8	:r񳺐g��i!�~������"�Q�S��V��O�N���������5�M䂿�������{�f.��lG��+Y�      Ѭ��$}�>tf��lG�ע%��p�/�ʿZ����>M����V�����d�ɤ�̷�/�d��
��I���1�j���h�຀��9~��:;�U4;��@;αF;.�H;َI;��I;�yI;�YI;7BI;�0I;�$I;�I;�I;I;�I;�I;�$I;�0I;7BI;�YI;�yI;��I;܎I;.�H;رF;��@;�U4;;x��:`��9d��k����1��I���
�/�d�̷�ɤ���d�V�������>M�Z���/�ʿ�p�ע%��lG�>tf�$}�      S���E���$}��+Y��3�����$ڿ&��Ľ\����(���s��3�6����p�d�V���<<�<������H��9A��:˻;N%3;Ap@;�yF;��H;��I;��I;�{I;K[I;NCI;�1I;Q%I;I;VI;I;SI;I;Q%I;�1I;OCI;E[I;�{I;ߛI;��I;��H;�yF;@p@;K%3;Ļ;7��:��9����=���<<�V��d��p�6����3��s�(�����Ľ\�&���$ڿ����3��+Y�$}�E���      �Aq���i���U�G:�@�����;���v���{A�d5�� ��^Z�����A���]�����d��M",��5����Ѻ���9���:�;XY4;B�@;HVF;~�H;�GI;�bI;OI;:I;�)I;I;{I;�I;�I;�I;~I;�I;{I;I;�)I;:I;OI;�bI;�GI;~�H;TVF;C�@;VY4;�;���:���9��Ѻ�5��L",��d������]��A�����^Z�� ��d5�{A�v���;�������@�G:���U���i�      ��i���b�Z�O�.5�2i�������������q<�����e��`
V�GE	�!���IY�j9�F�����(��R���ȺH�:G��:ޔ;<�4;8�@;hF;��H;
II;vbI;�NI;�9I;�)I;�I;ZI;�I;`I;ZI;[I;�I;ZI;�I;�)I;�9I;�NI;vbI;II;��H;#hF;:�@;9�4;֔;A��:0�:�Ⱥ�R����(�F���j9��IY�!��GE	�`
V��e������q<������������2i�.5�Z�O���b�      ��U�Z�O�H-?�.�'���M�ῴ欿`�{�fa/���뾝���I����d���ZN�]5������>H�h ��x���h�":��:x�;��5;�`A;��F;H�H;MI;�aI;�MI;�8I;�(I;@I;�I;7I;I;I;I;9I;�I;@I;�(I;�8I;�MI;�aI;MI;H�H;��F;�`A;��5;p�;}�:X�":n���j ��>H�����]5���ZN�d������I�������fa/�`�{��欿M����.�'�H-?�Z�O�      G:�.5�.�'��������jȿ���k$_���W�Ҿܕ���6�����*���`=�>�漯)��KG�*6������Q:��:�/";�7;X&B;��F;��H;�RI;�`I;vKI;7I;�'I;;I;I;�I;oI;n
I;jI;�I;I;;I;�'I;7I;yKI;�`I;�RI;��H;��F;X&B;�7;�/";��:��Q:���,6��KG��)��?���`=��*������6�ܕ��W�Ҿ��k$_����jȿ�������.�'�.5�      @�2i�������I�ѿk��� ���q<��:��a����q����Wн罅���'�Vb̼�zl��.��T�X������:��;ˎ&;ë9;C;8MG;��H;5YI;�^I;�HI;�4I;�%I;�I;I;�I;�
I;�	I;�
I;�I;I;�I;�%I;�4I;�HI;�^I;6YI;��H;?MG;C;��9;ǎ&;��;��:p��W�X��.���zl�Vb̼��'�罅��Wн����q��a���:��q<� ��k���I�ѿ������2i�      �������M��jȿk���������O���{]׾{����I�����A��?�d�n�֮�RH��jλW�$�@)�i��:BN;��+;�<;�3D;��G;�I;|^I;h[I;�DI;2I;�#I;CI;�I;]I;�	I;�I;�	I;]I;�I;BI;�#I;2I;�DI;h[I;�^I;�I;��G;�3D;�<;��+;@N;W��:)�X�$��jλRH��֮�n�>�d��A������I�{���z]׾����O�����k���jȿM�Ῡ��      ;��������欿��� ����O��x����� ���l���"��ܽ���`=����x���k"�0R��Nۺ���9�?�:ZL;{�0;��>;�ME;G#H;�%I;�aI;�VI;�@I;�.I;<!I;>I; I;
I;MI;�I;JI;
I;I;=I;;!I;�.I;�@I;�VI;�aI;�%I;K#H;�ME;��>;x�0;WL;r?�:���9Rۺ0R���k"�x������`=����ܽ��"��l�� ����뾁x���O� ������欿����      v�������`�{�k$_��q<�������}��w��	�6�����!���h����㷾�� d��.���^e�I[���Z:X��:�, ;��5;�A;�VF;��H;�@I;kbI;�QI;�;I;:+I;kI;I;5I;}	I;�I;,I;�I;	I;7I;I;iI;9+I;�;I;�QI;pbI;�@I;��H;�VF;�A;��5;�, ;J��:��Z: I[��^e��.��� d�ⷾ�����h�!������	�6�w���}��������q<�k$_�`�{�����      {A��q<�fa/����:�z]׾� ��w��>�DE	�����ڽ����3�_�꼚���",��W��d��@Q�o��:�M
;�f);��:;#@C;�?G;M�H;GTI;�_I;$KI;�6I;K'I;eI;�I;<I;�I;oI;�I;lI;�I;;I;�I;eI;L'I;�6I;'KI;�_I;BTI;M�H;�?G; @C;��:;�f);�M
;w��:@Q�j���W��",�����_�꼙�3�ڽ������DE	�>�w��� ��z]׾�:���fa/��q<�      d5�������W�Ҿ�a��{����l�	�6�DE	���Ƚk���aG����f֮��W����t�k�6���c,:��:��;��1;:�>;<E;�G;I;$_I;>ZI;3DI;�1I;-#I;CI;�I;
I;	I;�I;!I;�I;	I;
I;�I;?I;/#I;�1I;6DI;AZI;"_I;I;"�G;7E;<�>;��1;�;���:�c,:@��q�k�����W�f֮�����aG�k����ȽDE	�	�6��l�{����a��W�Ҿ������      � ���e�����ܕ����q��I���"���������k���ZN�\�"¼R�y��$��Q���� � tX���:0;!�&;�w8;j B;��F;ΐH;R@I;�aI;hRI;=I;,I;�I;�I;[I;�I;5I;I;cI;I;5I;�I;ZI;�I;�I;,I;=I;jRI;�aI;P@I;ԐH;��F;k B;�w8;�&;0;��: �X��� ��Q���$�P�y�"¼[��ZN�k������������"��I���q�ܕ������e��      ~^Z�`
V��I��6�������ܽ!��ڽ���aG�[��ȼ�)��~�(�k��QG5������Z:�:S;'1;��=;��D;+�G;��H;�XI;^I;|II;�5I;�&I;�I;�I;�
I;�I;KI;` I;��H;` I;KI;�I;�
I;~I;�I;�&I;�5I;|II;^I;�XI;��H;+�G;��D;��=;'1;S;�:��Z:���OG5�l��}�(��)��
�ȼ[��aG�ڽ��!���ܽ������6��I�`
V�      ���GE	��������Wн�A�����h���3����!¼�)��3x/��һy�X�x#����9F��:�>;)f);e`9;[&B;��F;c}H;�6I;NaI;�UI;^@I;�.I;� I;DI;'I;�I;LI;P I;��H;��H;��H;O I;LI;�I;$I;HI;!I;�.I;a@I;�UI;IaI;�6I;d}H;��F;]&B;``9;3f);�>;<��:��9x#��w�X��һ3x/��)��"¼�����3��h��󑽢A���Wн��콺��GE	�      �A��!��d���*��潅�?�d��`=����_��e֮�P�y�~�(��һ�]e�􄮺0�f9���:6�;C1";�4;�m?;�E;��G;d�H;�WI;}^I;
KI;o7I;�'I;�I;"I;�
I;#I;I;k�H;��H;:�H;��H;j�H;I; I;�
I;%I;�I;�'I;r7I;KI;w^I;�WI;c�H;��G;�E;�m?;�4;C1";0�;���:�f9򄮺�]e��һ~�(�P�y�f֮�^�꼗���`=�>�d�罅��*��d��!��      �]��IY��ZN��`=���'�n����᷾������W��$�l��|�X������9p��:Q��:m�;��0;��<;P�C;G;��H;�?I;#aI;�TI;<@I;/I;T!I;�I;I;xI;�I;��H;|�H;�H;��H;�H;z�H;��H;�I;uI;I;�I;W!I;/I;<@I;�TI;'aI;�?I;��H; G;N�C;��<;��0;e�;W��:n��:�9򄮺y�X�j���$��W�����᷾����n���'��`=��ZN��IY�      ���j9�\5��=��Ub̼֮�v��� d�",�����Q��SG5��#��0�f9n��:��:�;��-;��:;�KB;8VF;KH;�I;�\I;\I;�HI;6I;'I;I;�I;
I;BI;��H;��H;��H;X�H;��H;W�H;��H;��H;��H;?I;
I;�I;I;'I;6I;�HI;\I;�\I;�I;KH;8VF;�KB;��:;��-;
�;��:p��:�f9�#��OG5��Q�����",�� d�w��~֮�Vb̼=��\5��i9�      �d��D��������)���zl�RH��k"�z.���W��j�k��� ������9���:]��:�;�-;ɫ9;?aA;��E;#�G;r�H;�RI;`I;�OI;�<I;�,I;�I;-I;I;zI;TI;��H;��H;��H;��H;`�H;��H;��H;��H;��H;QI;{I;I;-I;�I;�,I;~<I;�OI;`I;�RI;u�H;#�G;��E;BaA;«9;�-;�;_��:���:��9����� �l�k��W��|.���k"�RH��zl��)������C���      E",���(�>H�HG��.���jλ*R���^e�d��2�� tX�l�Z:8��:.�;i�;��-;��9;tA;�cE;�G;��H;LGI;�`I;�UI;7BI;�1I;�#I;�I;�I;�I;�I;��H;H�H;��H;
�H;�H;��H;�H;�H;��H;D�H;|�H;�I;�I;�I;�I;�#I;�1I;;BI;�UI;�`I;OGI;��H;�G;�cE;pA;ë9;��-;i�;.�;:��:��Z: \X�.��]���^e�+R���jλ�.��HG�<H���(�      �5���R��h ��(6��W�X�F�$�8ۺ�H[��Q��c,:��:�:�>;@1";��0;��:;?aA;�cE;�G;p�H;�=I;(`I;kYI;�FI;�5I;�'I;�I;�I;�
I;�I;��H;�H;�H;��H;�H;��H;<�H;��H;}�H;��H;�H; �H;��H;�I;�
I;�I;�I;�'I;�5I;�FI;iYI;*`I;�=I;s�H;��G;�cE;BaA;��:;��0;A1";�>;�:��:�c,:�Q��H[�>ۺL�$�T�X�,6��g ���R��      ��Ѻ�Ⱥ^����������(��9��Z:y��:���:!0;S;,f);�4;��<;�KB;��E; �G;p�H;Y:I;L_I;|[I;JI; 9I;�*I;�I;�I;�I;[I;I;��H;��H;�H;/�H;��H;7�H;��H;0�H;��H;-�H;�H;��H;��H;I;XI;�I;�I;�I;�*I; 9I;JI;|[I;O_I;[:I;u�H;�G;��E;�KB;��<;�4;.f);S;!0;���:y��:��Z:ؓ�9p(�d�����t���(�Ⱥ      ���9 �:�":��Q:��:_��:n?�:R��:�M
;��; �&;'1;]`9;�m?;M�C;:VF;!�G;��H;�=I;J_I;\I;�KI;;I;�,I;� I;�I;�I;�I;GI;��H;3�H;x�H;5�H;��H;��H;��H;��H;��H;��H;��H;1�H;q�H;6�H;��H;CI;�I;�I;�I;� I;�,I;;I;�KI;\I;K_I;�=I;��H;#�G;<VF;P�C;�m?;_`9;'1;!�&;��;�M
;L��:z?�:U��:��:��Q:8�":�:      ���:k��:��:��:��;BN;WL;�, ;�f);��1;�w8;��=;Z&B;�E; G;KH;u�H;QGI;+`I;[I;�KI;�;I;�-I;."I;*I;I;	I;aI;��H;��H;��H;i�H;y�H;�H;D�H;��H;d�H;��H;B�H;�H;v�H;e�H;��H;��H;��H;aI;	I;I;-I;+"I;�-I;�;I;�KI;~[I;,`I;NGI;v�H;KH; G;�E;[&B;��=;�w8;��1;�f);�, ;^L;>N;��;��:��:W��:      .�;ݔ;p�;�/";��&;��+;��0;��5;��:;A�>;s B;��D;��F;��G;��H;�I;�RI;�`I;kYI;JI;;I;�-I;�"I;�I;�I;�	I;'I;G�H;o�H;W�H;��H;��H;��H;��H;��H;��H;`�H;��H;��H;��H;��H;��H;��H;T�H;h�H;I�H;&I;�	I;�I;�I;"I;�-I;;I;JI;mYI;�`I;�RI;�I;��H;��G;��F;��D;y B;<�>;��:;��5;��0;��+;Ύ&;�/";o�;ɔ;      XY4;F�4;��5; �7;��9;�<;��>;�A;@C;<E;��F;(�G;_}H;c�H;�?I;�\I;`I;�UI;�FI;�8I;�,I;%"I;�I; I;U
I;�I;��H;��H;��H;��H;��H;��H;��H;��H;��H;��H;f�H;��H;��H;��H;��H;��H;��H;��H;��H;��H;��H;�I;Y
I;I;�I;("I;�,I;�8I;�FI;�UI;`I;�\I;�?I;a�H;_}H;,�G;��F;:E;!@C;�A;��>;�<;��9; �7;��5;<�4;      d�@;<�@;�`A;S&B;C;4D;�ME;�VF;�?G;#�G;ؐH;��H;�6I;�WI;)aI;&\I;�OI;BBI;�5I;�*I;� I;.I;�I;`
I;�I; I;-�H;��H;!�H;��H;��H;��H;K�H;z�H;��H;��H;e�H;��H;��H;z�H;G�H;��H;��H;��H;�H;��H;)�H; I;�I;]
I;�I;1I;� I;�*I;�5I;<BI;�OI;'\I;)aI;�WI;�6I;��H;ڐH;#�G;�?G;�VF;�ME;�3D;$C;X&B;�`A;;�@;      FVF;*hF;��F;��F;-MG;��G;K#H;��H;L�H;I;V@I;�XI;OaI;�^I;�TI;�HI;�<I;�1I;�'I;�I;�I;
I;�	I;�I; I;;�H;�H;X�H;��H;��H;w�H;H�H;=�H;x�H;�H;��H;|�H;��H;�H;x�H;<�H;D�H;w�H;��H;��H;U�H;�H;?�H; I;�I;�	I;I;�I;�I;�'I;�1I;�<I;�HI;�TI;~^I;OaI;�XI;^@I;I;O�H;��H;M#H;��G;EMG;��F;��F;'hF;      ��H;��H;E�H;��H;��H;�I;�%I;�@I;GTI;&_I;�aI;^I;�UI;	KI;;@I;6I;�,I;�#I;�I;�I;�I;	I;'I;��H;)�H;�H;F�H;�H;+�H;n�H;&�H;�H;5�H;��H;7�H;��H;��H;��H;4�H;��H;6�H;�H;%�H;k�H;%�H;�H;A�H;�H;,�H;��H;'I;	I;�I;�I;�I;�#I;�,I;6I;;@I;KI;�UI;^I;�aI;"_I;DTI;�@I;�%I;�I;��H;��H;E�H;��H;      �GI;II;MI;�RI;(YI;�^I;�aI;obI;�_I;DZI;oRI;�II;]@I;t7I;/I;'I;�I;�I;�I;�I;�I;\I;B�H;��H;��H;O�H;�H;�H;y�H;&�H;��H;�H;b�H;��H;t�H;=�H;2�H;9�H;r�H;��H;d�H;�H;��H;"�H;v�H;�H;�H;U�H;��H;��H;B�H;^I;�I;�I;�I;�I;�I;'I;/I;t7I;[@I;�II;qRI;HZI;�_I;obI;�aI;u^I;3YI;�RI;MI;II;      �bI;rbI;�aI;�`I;�^I;k[I;WI;�QI; KI;6DI;=I;�5I;�.I;�'I;U!I;I;2I;�I;�
I;]I;KI;��H;j�H;��H;�H;��H;$�H;z�H;�H;��H;��H;8�H;��H;)�H;��H;��H;��H;��H;��H;*�H;��H;5�H;��H;��H;�H;w�H;!�H;��H;�H;��H;k�H;��H;JI;YI;�
I;�I;4I;I;X!I;�'I;�.I;�5I;=I;7DI;$KI;�QI;WI;c[I;�^I;�`I;�aI;nbI;      OI;�NI;�MI;qKI;�HI;�DI;�@I;�;I;�6I;�1I;,I;�&I; !I;�I;�I;�I;I;�I;�I;I;��H;��H;S�H;��H;��H;��H;k�H;(�H;��H;��H;#�H;|�H;��H;��H;A�H;�H;�H;�H;@�H;��H;��H;{�H;#�H;��H;��H;#�H;g�H;��H;��H;��H;V�H;��H;��H;	I;�I;�I;I;�I;�I;�I; !I;�&I;,I;�1I;�6I;�;I;�@I;�DI;�HI;yKI;�MI;�NI;      :I;�9I;�8I;!7I;�4I;2I;�.I;E+I;P'I;6#I;�I;�I;MI;,I;I;
I;�I;�I;��H;��H;<�H;��H;��H;��H;��H;u�H;&�H;�H;��H;)�H;��H;��H;Y�H;	�H;��H;��H;��H;��H;��H;�H;\�H;��H;��H;&�H;��H;�H;%�H;w�H;��H;��H;��H;��H;9�H;��H;��H;�I;�I; 
I;I;+I;OI;�I;�I;9#I;U'I;B+I;�.I;2I;�4I;#7I;�8I;�9I;      �)I;�)I;�(I;�'I;�%I;�#I;9!I;nI;hI;EI;�I;�I;'I;�
I;vI;CI;XI;��H;
�H;��H;}�H;i�H;��H;��H;��H;@�H;	�H;�H;:�H;}�H;��H;t�H;��H;��H;t�H;L�H;6�H;L�H;p�H;��H;��H;t�H;��H;|�H;5�H;	�H;�H;B�H;��H;��H;��H;i�H;x�H;��H;�H;��H;ZI;FI;{I;�
I;(I;�I;�I;HI;jI;mI;C!I;�#I;�%I;�'I;�(I;�)I;      "I;�I;JI;>I;�I;8I;:I;	I;�I;�I;[I;�
I;�I;&I;�I;��H;��H;H�H; �H;�H;?�H;{�H;��H;��H;I�H;9�H;6�H;i�H;��H;��H;V�H;��H;��H;S�H;�H; �H;�H;��H;	�H;U�H;��H;��H;V�H;��H;��H;g�H;6�H;:�H;L�H;��H;��H;x�H;9�H;�H; �H;I�H;��H; I;�I;&I;�I;�
I;_I;�I;�I;	I;>I;2I;�I;;I;QI;�I;      sI;WI;�I;I; I;�I;I;9I;:I;
I;�I;�I;RI; I;��H;��H;��H;��H;��H;4�H;��H;�H;��H;��H;u�H;q�H;��H;��H;,�H;��H;�H;��H;U�H;�H;��H;��H;��H;��H;��H;�H;W�H;��H;�H;��H;&�H;��H;��H;v�H;w�H;��H;��H;�H;��H;+�H;��H;��H;��H;��H;��H;!I;RI;�I;�I;
I;<I;6I;I;�I;I;I;�I;bI;      �I;�I;;I;�I;�I;TI;I;�	I;�I;I;<I;VI;X I;t�H;��H;��H;��H;	�H;~�H;��H;��H;B�H;��H;��H;��H;��H;1�H;r�H;��H;D�H;��H;v�H;�H;��H;��H;��H;��H;��H;��H;��H;�H;w�H;��H;?�H;��H;o�H;3�H; �H;��H;��H;��H;@�H;��H;��H;~�H;
�H;��H;��H;��H;u�H;[ I;VI;BI;I;�I;�	I;I;VI;�I;�I;=I;�I;      zI;`I;I;mI;�
I;}	I;QI;�I;jI;�I;!I;d I;��H;��H;�H;U�H;��H;�H;��H;7�H;��H;��H;��H;x�H;��H;��H;��H;>�H;��H;"�H;��H;P�H;�H;��H;��H;z�H;y�H;}�H;��H;��H;�H;P�H;��H;�H;��H;;�H;��H;��H;��H;x�H;��H;��H;��H;2�H;��H;�H;��H;Z�H;�H;��H;��H;b I;$I;�I;mI;�I;[I;	I;�
I;mI;�I;nI;      �I;SI;I;n
I;�	I;�I;�I;0I;�I;I;lI;��H;��H;A�H;��H;��H;h�H;��H;>�H;��H;��H;g�H;]�H;]�H;c�H;r�H;��H;7�H;��H;"�H;��H;8�H;�H;��H;��H;u�H;~�H;u�H;��H;��H;�H;;�H;��H;�H;��H;3�H;��H;v�H;b�H;\�H;`�H;d�H;��H;��H;>�H;��H;h�H;��H;��H;A�H;��H;��H;pI;I;�I;0I;�I;�I;�	I;t
I;I;`I;      zI;aI;�I;jI;�
I;	I;PI;�I;jI;�I; I;e I;��H;��H;�H;U�H;��H;�H;��H;6�H;��H;��H;��H;x�H;��H;��H;��H;>�H;��H;!�H;��H;P�H;�H;��H;��H;z�H;y�H;}�H;��H;��H;�H;P�H;��H;�H;��H;:�H;��H;��H;��H;w�H;��H;��H;��H;2�H;��H;�H;��H;X�H;�H;��H;��H;b I;%I;�I;mI;�I;WI;	I;�
I;nI;I;hI;      �I;�I;9I;�I;�I;QI;I;�	I;�I;I;;I;VI;X I;t�H;��H;��H;��H;
�H;~�H;��H;��H;C�H;��H;��H;��H;��H;1�H;r�H;��H;C�H;��H;v�H;�H;��H;��H;��H;��H;��H;��H;��H;�H;v�H;��H;=�H;��H;n�H;3�H;�H;��H;��H;��H;B�H;��H;��H;~�H;
�H;��H;��H;��H;t�H;Z I;VI;AI;I;�I;�	I;I;QI;�I;�I;>I;�I;      sI;XI;�I;I; I;�I; I;<I;<I;
I;�I;�I;PI; I;��H;��H;��H;��H;��H;1�H;��H;�H;��H;��H;x�H;s�H;��H;��H;-�H;��H;�H;��H;U�H;�H;��H;��H;��H;��H;��H;�H;W�H;��H;�H;��H;&�H;��H;��H;v�H;u�H;��H;��H;�H;��H;-�H;��H;��H;��H;��H;��H; I;PI;�I;�I;
I;<I;:I;
I;�I;I;I;�I;ZI;       I;�I;MI;<I;�I;;I;9I;I;�I;�I;ZI;�
I;�I;&I;�I;��H;��H;H�H;�H;�H;?�H;y�H;��H;��H;K�H;3�H;6�H;i�H;��H;��H;U�H;��H;��H;S�H;�H;�H;�H; �H;�H;T�H;��H;��H;V�H;��H;��H;e�H;6�H;9�H;I�H;��H;��H;x�H;5�H;�H;�H;G�H;��H;  I;�I;$I;�I;�
I;^I;�I;�I;I;@I;6I;�I;BI;UI;�I;      �)I;�)I;�(I;�'I;�%I;�#I;@!I;jI;eI;EI;�I;�I;(I;�
I;yI;CI;XI;��H;�H;��H;�H;i�H;��H;��H;��H;>�H;	�H;�H;<�H;|�H;��H;t�H;��H;��H;w�H;G�H;6�H;L�H;p�H;��H;��H;t�H;��H;{�H;5�H;�H;	�H;B�H;��H;��H;��H;i�H;v�H;��H;�H;��H;ZI;FI;yI;�
I;(I;�I;�I;EI;gI;jI;B!I;�#I;�%I;�'I;�(I;�)I;      :I;�9I;�8I;7I;�4I;2I;�.I;E+I;N'I;3#I;�I;�I;MI;)I;I;
I;�I;�I;��H;��H;=�H;��H;��H;��H;��H;p�H;"�H;�H;��H;'�H;��H;��H;[�H;�H;��H;��H;��H;��H;��H;�H;\�H;��H;��H;%�H;��H;��H;&�H;w�H;��H;��H;��H;��H;6�H;��H;��H;�I;�I;
I;I;+I;MI;�I;�I;4#I;R'I;G+I;�.I;2I;�4I;(7I;�8I;�9I;      #OI;�NI;�MI;|KI;yHI;�DI;�@I;�;I;�6I;�1I;,I;�&I;� I;�I;�I;�I;I;�I;�I;I;��H;��H;O�H;��H;��H;��H;h�H;%�H;��H;��H;#�H;}�H;��H;��H;C�H;�H;�H;�H;@�H;��H;��H;�H;#�H;��H;��H;%�H;k�H;��H;��H;��H;W�H;��H;��H;	I;�I;�I;I;�I;�I;�I;� I;�&I;,I;�1I;�6I;�;I;�@I;�DI;�HI;�KI;�MI;�NI;      �bI;qbI;�aI;�`I;{^I;n[I;�VI;�QI;'KI;2DI;=I;�5I;�.I;�'I;X!I;I;1I;�I;�
I;YI;KI;��H;e�H;��H;�H;��H;!�H;y�H;�H;��H;��H;:�H;��H;)�H;��H;��H;��H;��H;��H;)�H;��H;:�H;��H;��H;�H;w�H;$�H;��H;�H;��H;m�H;��H;HI;YI;�
I;�I;1I;I;X!I;�'I;�.I;�5I;=I;2DI;"KI;�QI;WI;h[I;�^I;�`I;�aI;jbI;      �GI;II;�LI;�RI;$YI;�^I;�aI;ubI;�_I;CZI;lRI;�II;[@I;r7I;/I;'I;�I;�I;�I;�I;�I;]I;>�H;��H;��H;K�H;
�H;�H;z�H;"�H;��H;�H;b�H;��H;u�H;;�H;4�H;>�H;q�H;��H;e�H;�H;�H;%�H;w�H;�H;�H;Q�H;��H;��H;E�H;]I;�I;�I;�I;�I;�I;'I;/I;q7I;[@I;II;oRI;EZI;�_I;nbI;�aI;z^I;2YI;�RI;	MI;II;      ��H;��H;A�H;��H;��H;�I;�%I;�@I;GTI;#_I;�aI;^I;�UI;KI;:@I;6I;�,I;�#I;�I;�I;�I;	I;"I;��H;*�H;	�H;C�H;�H;+�H;k�H;%�H;�H;5�H;��H;8�H;��H;��H;��H;4�H;��H;6�H;�H;(�H;n�H;(�H;�H;G�H;�H;*�H;��H;,I;	I;�I;�I;�I;�#I;�,I;6I;<@I;KI;�UI;^I;�aI;"_I;DTI;�@I;�%I;�I;��H;��H;C�H;��H;      <VF;&hF;��F;��F;4MG;��G;J#H;��H;O�H;I;V@I;�XI;OaI;~^I;�TI;�HI;�<I;�1I;�'I;�I;�I;I;�	I;�I; I;7�H;�H;Y�H;��H;��H;v�H;H�H;:�H;x�H;�H;��H;}�H;��H;�H;x�H;=�H;I�H;z�H;��H;��H;X�H;�H;;�H; I;�I;�	I;I;�I;�I;�'I;�1I;�<I;�HI;�TI;}^I;NaI;�XI;[@I;I;H�H;��H;J#H;��G;>MG;��F;�F;hF;      a�@;7�@;�`A;X&B;C;4D;�ME;�VF;�?G;"�G;ԐH;��H;�6I;�WI;,aI;'\I;�OI;ABI;�5I;�*I;� I;0I;�I;_
I;�I; I;)�H;��H; �H;��H;��H;��H;G�H;x�H;��H;��H;f�H;��H;��H;{�H;I�H;��H;�H;��H;�H;��H;-�H; I;�I;\
I;�I;0I;� I;�*I;�5I;;BI;�OI;'\I;*aI;�WI;�6I;��H;֐H;"�G;�?G;�VF;�ME;�3D; C;X&B;�`A;8�@;      2Y4;+�4;��5;�7;��9;�<;��>;�A;#@C;7E;��F;+�G;_}H;`�H;�?I;�\I;`I;�UI;�FI;�8I;�,I;$"I;�I;I;Y
I;�I;��H;��H;��H;��H;��H;��H;��H;��H;��H;��H;i�H;��H;��H;��H;��H;��H;��H;��H;��H;��H;��H;�I;V
I;I;�I;%"I;�,I;�8I;�FI;�UI;`I;�\I;�?I;`�H;_}H;*�G;��F;9E;@C;�A;��>;�<;ū9;!�7;��5;�4;      �;֔;b�;�/";��&;��+;�0;��5;��:;?�>;n B;��D;��F;��G;��H;�I;�RI;�`I;iYI;JI;;I;�-I;|"I;�I;�I;�	I;%I;H�H;m�H;S�H;��H;��H;��H;��H;��H;��H;c�H;��H;��H;��H;��H;��H;��H;X�H;k�H;H�H;,I;�	I;�I;�I;�"I;�-I;;I;JI;nYI;�`I;�RI;�I;��H;��G;��F;��D;r B;?�>;��:;��5;�0;��+;��&;�/";c�;;      ���:c��:��:��:��;HN;[L;�, ;�f);��1;�w8;��=;Z&B;�E;"G;KH;t�H;OGI;(`I;|[I;�KI;�;I;�-I;+"I;.I;I;	I;aI;��H;��H;��H;j�H;v�H;�H;C�H;��H;e�H;��H;B�H;�H;y�H;l�H;��H;��H;��H;aI;	I;I;,I;."I;�-I;�;I;�KI;[I;,`I;LGI;u�H;KH; G;�E;Z&B;��=;�w8;��1;�f);�, ;WL;2N;��;��:��:O��:      ���9T�:<�":�Q:��:i��:t?�:T��:�M
;�; �&;'1;]`9;�m?;P�C;:VF;"�G;��H;�=I;J_I;\I;�KI;
;I;�,I;� I;�I;�I;�I;DI;��H;3�H;x�H;2�H;��H;��H;��H;��H;��H;��H;��H;5�H;x�H;7�H;��H;DI;�I;�I;�I;� I;�,I;;I;�KI;\I;L_I;�=I;��H;#�G;<VF;P�C;�m?;_`9;'1;#�&;��;�M
;X��:|?�:_��:��: �Q:p�":�:      ��Ѻ�Ⱥl���������p(����9��Z:��:���:0;S;.f);�4;��<;�KB;��E;�G;o�H;Y:I;L_I;|[I;JI;�8I;�*I;�I;�I;�I;YI;I;��H;��H;�H;/�H;��H;3�H;��H;6�H;��H;-�H;�H;��H;��H;I;[I;�I;�I;�I;�*I;9I;JI;|[I;N_I;[:I;s�H;�G;��E;�KB;��<;�4;,f);S;!0;���:y��:��Z:���9)�h�����n����Ⱥ      �5���R��h ��'6��[�X�H�$�>ۺ�H[�@Q��c,:��:�:�>;>1";��0;��:;?aA;�cE;�G;p�H;�=I;(`I;jYI;�FI;�5I;�'I;�I;�I;�
I;�I;��H;�H;�H;��H;}�H;��H;;�H;��H;z�H;��H;�H;�H;��H;�I;�
I;�I;�I;�'I;�5I;�FI;mYI;*`I;�=I;s�H;��G;�cE;AaA;��:;��0;@1";�>;�:��:�c,: Q��H[�@ۺJ�$�Z�X�'6��j ���R��      I",���(�?H�HG��.���jλ(R���^e�`��4�� pX�t�Z:4��:,�;l�;��-;«9;pA;�cE;�G;��H;NGI;�`I;�UI;8BI;�1I;�#I;�I;�I;�I;�I;~�H;D�H;��H;	�H;�H;��H;�H;�H;��H;G�H;��H;�I;�I;�I;�I;�#I;�1I;5BI;�UI;�`I;OGI;��H;�G;�cE;qA;«9;��-;k�;,�;4��:l�Z: pX�6��c���^e�*R���jλ�.��HG�BH���(�      �d��D��������)���zl�RH��k"�|.���W��l�k��� ������9���:_��:�;�-;ū9;>aA;��E;%�G;t�H;�RI;`I;�OI;}<I;�,I;�I;+I;I;zI;QI;��H;��H;��H;��H;a�H;��H;��H;��H;��H;SI;|I;I;.I;�I;�,I;~<I;�OI;`I;�RI;t�H;�G;��E;?aA;ë9;�-;�;_��:���:��9����� �n�k��W��|.���k"�RH��zl��)������D���      ���j9�\5��<��Vb̼~֮�w��� d�",�����Q��OG5��#�� �f9t��:��:	�;��-;��:;�KB;<VF;KH;�I;�\I;\I;�HI;�5I;'I;I;�I;
I;?I;��H;��H;��H;W�H;��H;W�H;��H;��H;��H;AI;
I;�I;I;'I;6I;�HI;\I;�\I;�I;KH;4VF;�KB;��:;��-;
�;��:p��:�f9�#��UG5��Q�����",�� d�w��~֮�Wb̼=��^5��j9�      �]��IY��ZN��`=���'�n����᷾������W��$�k��y�X������9n��:W��:h�;��0;��<;R�C;G;��H;�?I;#aI;�TI;7@I;/I;U!I;�I;I;vI;�I;��H;|�H;�H;��H;�H;y�H;��H;�I;vI;I;I;X!I;/I;:@I;�TI;"aI;�?I;��H; G;J�C;��<;��0;e�;Y��:j��:�9􄮺}�X�k���$��W�����᷾����n���'��`=��ZN��IY�      �A��!��d���*��潅�>�d��`=����^��f֮�P�y�}�(��һ�]e�섮�@�f9���:.�;@1";�4;�m?;�E;��G;c�H;�WI;|^I;KI;k7I;�'I;�I;%I;�
I; I;I;k�H;��H;:�H;��H;i�H;I; I;�
I;"I;�I;�'I;o7I;KI;y^I;�WI;e�H;��G;�E;�m?;�4;=1";.�;���:�f9�����]e��һ}�(�P�y�f֮�^�꼗���`=�>�d�罅��*��d��!��      ���GE	��������Wн�A�����h���3����!¼�)��3x/��һs�X�x#��x�9@��:�>;.f);f`9;[&B;��F;c}H;�6I;KaI;�UI;[@I;�.I;� I;GI;%I;�I;OI;P I;��H;��H;��H;O I;LI;�I;"I;FI;� I;�.I;]@I;�UI;IaI;�6I;c}H;��F;Z&B;]`9;2f);�>;:��:��9|#��w�X��һ3x/��)��"¼�����3��h��󑽢A���Wн��콺��GE	�      ~^Z�`
V��I��6�������ܽ!��ڽ���aG�[�
�ȼ�)��~�(�j��OG5����d�Z:�:
S;'1;��=;��D;+�G;��H;�XI;^I;xII;�5I;�&I;�I;I;�
I;�I;KI;^ I;��H;` I;JI;�I;�
I;I;�I;�&I;�5I;{II;^I;�XI;��H;,�G;��D;��=;'1;S;�:x�Z:���RG5�j��~�(��)���ȼ[��aG�ڽ��!���ܽ������6��I�`
V�      � ���e�����ܕ����q��I���"���������k���ZN�[�"¼Q�y��$��Q���� � �X���:0;$�&;�w8;l B;��F;АH;S@I;�aI;iRI;=I;,I;�I;�I;[I;�I;3I;I;cI;I;3I;�I;[I;�I;�I;,I;=I;lRI;�aI;P@I;ΐH;��F;n B;�w8;�&;0;��: xX��� ��Q���$�Q�y�"¼\��ZN�k������������"��I���q�ܕ������e��      d5�������W�Ҿ�a��{����l�	�6�DE	���Ƚk���aG����f֮��W����s�k�B���c,:���:��;��1;;�>;:E;�G;I; _I;=ZI;5DI;�1I;0#I;AI;�I;
I;I;�I;I;�I;I;
I;�I;?I;/#I;�1I;5DI;@ZI;_I;I;�G;:E;?�>;��1;�;���:�c,:@��q�k�����W�f֮�����aG�k����ȽDE	�	�6��l�{����a��W�Ҿ������      {A��q<�fa/����:�z]׾� ��w��>�DE	�����ڽ����3�_�꼚���",��W��j���Q�s��:�M
;�f);��:; @C;�?G;K�H;BTI;�_I;&KI;�6I;N'I;dI;�I;;I;�I;lI;�I;jI;�I;;I;�I;dI;L'I;�6I;'KI;�_I;BTI;M�H;�?G;$@C;��:;�f);�M
;y��: Q�g���W��",�����_�꼙�3�ڽ������DE	�>�w��� ��z]׾�:���fa/��q<�      v�������`�{�k$_��q<�������}��w��	�6�����!���h����ⷾ�� d��.���^e�I[���Z:Z��:�, ;��5;�A;�VF;��H;�@I;kbI;�QI;�;I;;+I;kI;I;6I;{	I;�I;+I;�I;}	I;5I;I;iI;;+I;�;I;�QI;nbI;�@I;��H;�VF;�A;��5;�, ;F��:��Z:(I[��^e��.��� d�㷾�����h�!������	�6�w���}��������q<�k$_�`�{�����      ;��������欿��� ����O��x����� ���l���"��ܽ���`=����x���k"�0R��Nۺ���9|?�:XL;z�0;��>;�ME;C#H;�%I;�aI;�VI;�@I;�.I;<!I;=I;I;I;JI;�I;II;	I; I;=I;;!I;�.I;�@I;�VI;�aI;�%I;M#H;�ME;��>;}�0;UL;n?�:���9Tۺ0R���k"�x������`=����ܽ��"��l�� ����뾁x���O� ������欿����      �������M��jȿk���������O���z]׾{����I�����A��?�d�n�֮�RH��jλV�$� )�c��:@N;��+;�<;�3D;��G;�I;|^I;g[I;�DI;"2I;�#I;BI;�I;[I;�	I;�I;�	I;[I;�I;CI;�#I;2I;�DI;h[I;�^I;�I;��G;�3D;�<;��+;<N;[��:)�Z�$��jλRH�֮�n�>�d��A������I�{���z]׾����O�����k���jȿM�Ῡ��      @�2i�������I�ѿk��� ���q<��:��a����q����Wн罅���'�Vb̼�zl��.��T�X�t����:��;Ȏ&;��9; C;2MG;��H;2YI;�^I;�HI;�4I;�%I;�I;I;�I;�
I;�	I;�
I;�I;I;�I;�%I;�4I;�HI;�^I;6YI;��H;>MG; C;��9;ǎ&;��;��:t��W�X��.���zl�Vb̼��'�罅��Wн����q��a���:��q<� ��k���I�ѿ������2i�      G:�.5�.�'��������jȿ���k$_���W�Ҿܕ���6�����*���`=�>�漯)��KG�*6������Q:��:�/";�7;X&B;��F;��H;�RI;�`I;uKI;7I;�'I;:I;I;�I;nI;p
I;kI;I;I;<I;�'I;7I;zKI;�`I;�RI;��H;��F;Z&B;�7;�/";��:��Q:���,6��JG��)��>���`=��*������6�ܕ��W�Ҿ��k$_����jȿ�������.�'�.5�      ��U�Z�O�H-?�.�'���M�ῴ欿`�{�fa/���뾝���I����d���ZN�]5������?H�h ��t���p�":��:w�;��5;�`A;��F;G�H;MI;�aI;�MI;�8I;�(I;?I;�I;6I;I;I;I;9I;�I;BI;�(I;�8I;�MI;�aI;MI;H�H;��F;�`A;��5;o�;{�:X�":l���j ��>H�����]5���ZN�d������I�������fa/�`�{��欿M����.�'�H-?�Z�O�      ��i���b�Z�O�.5�2i�������������q<�����e��`
V�GE	�!���IY�j9�F�����(��R���ȺH�:G��:ޔ;<�4;:�@;hF;��H;
II;vbI;�NI;�9I;�)I;�I;ZI;�I;^I;\I;ZI;�I;ZI;�I;�)I;�9I;�NI;vbI;II;��H;$hF;:�@;:�4;֔;A��:0�:�Ⱥ�R����(�F���j9��IY�!��GE	�`
V��e������q<������������2i�.5�Z�O���b�      �>���8���*�O������˿p��E�b�C\�4m־^��R�:��J�)��F�B�>��������4/��`���̑>:]t�:
p ;�J6;�DA;WIF;�NH;��H;�!I;�I;�I;|I;NI;�I;J I;��H;�H;��H;H I;�I;NI;|I;�I;�I;�!I;��H;�NH;aIF;�DA;�J6;p ;Yt�:��>:Z���6/���������>��F�B�)���J�R�:�^��4m־C\�E�b�p���˿����O���*���8�      ��8��4��g&�6��<����<ƿ񲗿�>]�®�P�Ѿ�p���*7����%W��MR?�}�s8����"���䅍�p�G:g �:�!;�6;�kA;bYF;�TH;B�H;�!I;�I;�I;gI;(I;�I;; I;��H;��H;��H;; I;�I;(I;gI;�I;�I;�!I;C�H;�TH;lYF;�kA;�6;�!;c �:l�G:ޅ��"�����r8��}�MR?�%W�����*7��p��P�Ѿ®��>]�񲗿�<ƿ<���6���g&��4�      ��*��g&��#�t�U[�pL�������M�r5��>ľ����,��D�钐��5�3�ݼ���q
� �x�<uk���b:l�:�#;��7;P�A;��F;�dH;�I;!"I;�I;DI;I;�I;�I;��H;[�H;��H;T�H;��H;�I;�I;I;>I;�I;!"I;�I;�dH;��F;O�A;��7;�#;l�:��b:,uk�$�x��q
���3�ݼ�5�蒐��DὪ�,����>ľr5���M����pL��U[�t��#��g&�      O�6��t����˿@1��6�y�Î6��z �����1�l�+��ͽ$�����&���˼B�k�(�����X�� �h��:3�;�&;z9;f�B;��F;�}H;�	I;/"I;I;�I;yI;TI;"I;��H;�H;a�H;��H;��H;"I;QI;xI;I;I;/"I;�	I;�}H;��F;f�B;v9;�&;0�;`��:� ���X�(���B�k���˼��&�$����ͽ+�1�l������z �Î6�6�y�@1���˿���t�6��      ����<���U[忶˿�T���{�R�����E۾ӗ����M���	������j��3�d����O�?�׻��/����1��:� 
;�*;K;;�jC;z'G;ӛH;�I;�!I;�I;vI;�
I;�I;�I;"�H;��H;��H;��H;!�H;�I;�I;�
I;pI;�I;�!I;�I;ԛH;�'G;�jC;G;;�*;� 
;%��:p����/�?�׻��O�d���3���j������	���M�ӗ���E۾���{�R���T���˿U[�<���      �˿�<ƿpL��@1����>]���)��$��ֳ���{���,�r��(��R`I��J���,���3/�,�� � ��,69�4�:΄;�o.;.=;9aD;��G;P�H;�I;!I;<I;'I;�	I;�I;� I;��H;��H;B�H;��H;~�H;� I;�I;�	I;%I;AI;!I;�I;M�H;��G;8aD;
.=;�o.;ʄ;�4�:�,69 � �,���3/��,���J��R`I�'��r�齤�,���{�ֳ��$����)��>]��@1��pL���<ƿ      p��񲗿���6�y�{�R���)�nv��>ľ^���I�Xl����������&�ծҼ�}�3B�Ю��,���`�!:�*�:z;T3;Dj?;l\E;��G;��H;GI;|I;iI;�I;VI;�I;��H;��H;C�H;��H;A�H;��H;��H;�I;SI;�I;nI;{I;EI;��H;��G;m\E;Dj?;T3;z;�*�:l�!:*���Ү��3B��}�ծҼ��&��������Xl��I�^���>ľnv���)�{�R�6�y����񲗿      E�b��>]���M�Î6�����$���>ľ"q��y�Z�+�R9ݽ!W����L����#F���G��׻;�ho�rȊ:zi;�O$;��7;P�A;�IF;�BH;��H;� I;AI;TI;�I;I;I;��H;��H;t�H;��H;r�H;��H;��H;|I;I;�I;ZI;@I;� I;��H;CH;�IF;L�A;��7; P$;ti;zȊ:xo�;��׻�G�"F�������L�!W��R9ݽ+�y�Z�"q���>ľ�$�����Î6���M��>]�      C\����r5��z ��E۾ֳ�^��y�Z�L?#����A����j�&��Eϼ�����ε���lۺ89�9X4�:=�;A�,;P�;;�C;zG;�H;I;�!I;�I;"I;I;qI;$I;��H;��H;��H;�H;��H;��H;��H; I;pI;I;'I;�I;�!I;|I;�H;}G;�C;R�;;C�,;4�;`4�:(9�9�lۺε�������Eϼ&����j��A�����L?#�y�Z�^��ֳ��E۾�z �r5����      4m־P�Ѿ�>ľ����ӗ����{��I�+�����V���{�?�/�&���,��B=�F�һu�@�T� ���k:��:�a;��3;j?;M2E;��G;<�H;I;K I;�I;�I;�I;�I;��H;��H;��H;��H;8�H;��H;��H;��H;��H;�I;�I;�I;�I;K I;I;;�H;��G;J2E;j?;��3;�a;��:��k:d� �r�@�F�һB=��,��&��?�/��{��V�����+��I���{�ӗ�������>ľP�Ѿ      ^���p����1�l���M���,�Xl�Q9ݽ�A���{���5��J��
;���T[�#?�����jP���O�9��:��;*;�9;0kB;��F;RNH;Q�H;�I;eI;�I;�I;�I; I;C�H;��H;��H;��H;I�H;��H;��H;��H;A�H;I;�I;I;�I;fI;�I;P�H;VNH;��F;1kB; �9;*;��;��:�O�9dP������$?��T[�
;���J����5��{��A��Q9ݽXl���,���M�1�l����p��      Q�:��*7���,�+���	�r�齂���!W����j�?�/��J���I���k�n�.��l��x���Ȋ:!o�:�;@r3;��>;��D;J�G;!�H;�I;!I;�I;cI;_
I;�I;> I;��H;x�H;��H;��H;@�H;��H;��H;{�H;��H;< I;�I;d
I;jI;�I;!I;�I;$�H;J�G;�D;��>;?r3;�;#o�:�Ȋ:P��l��.��n��k��I���J��?�/���j�!W������q�齃�	�+���,��*7�      �J�����D��ͽ���'�������L�&��%��
;���k����pI����/��/��>:��:�B;9�,;��:;
�B;fxF;r<H;��H;�I;pI;�I;I;�I;�I;k�H;W�H;�H;N�H;~�H;M�H;~�H;N�H;�H;U�H;j�H;�I;�I;I;�I;oI;�I;��H;r<H;ixF;�B;��:;D�,;�B;��:�>:�/���/�nI������k�
;��&��%����L����'������ͽ�D����      (��%W��蒐�$�����j�R`I���&����Dϼ�,���T[�n�rI��k;��nk�\:�4�:�;�&;��6;�!@;2E;��G;~�H;�I;� I;0I;�I;�
I;I;O I;��H;��H;��H;@�H;t�H;'�H;t�H;?�H;��H;��H;��H;S I;I;�
I;�I;.I;� I;�I;|�H;��G;2E;�!@;��6;�&;|;�4�:X:�nk�h;�oI��n��T[��,��Dϼ�����&�R`I���j�$���蒐�%W��      E�B�MR?��5���&��3��J��ԮҼ!F����@=�"?�.����/��nk����9׳:��;!;63;��=;��C;��F;�cH;��H;kI;�I;�I;�I;�I;�I;�H;��H;r�H;_�H; �H;d�H;�H;b�H;�H;`�H;r�H;��H;!�H;�I;�I;I;�I;�I;nI;��H;�cH;��F;��C;��=;:3;!;��;׳:���9�nk���/�.��"?�A=���!F��ԮҼ�J���3���&��5�MR?�      ;�� }�2�ݼ��˼d���,���}��G����F�һ����m���/�X:׳:�;Kb;��0;j<;~�B;�IF;HH;��H;�I;J I;�I;I;6
I;�I;  I;�H;5�H;��H;�H;�H;\�H;�H;Z�H;��H;�H;��H;2�H;�H; I;�I;9
I;I;�I;O I;�I;�H;KH;�IF;��B;m<;��0;Lb;�;׳:X:�/�k������E�һ����G��}��,��d����˼2�ݼ�|�      ����q8����B�k���O��3/�0B��׻ʵ��k�@�ZP��`���>:�4�:��;Pb;|�/;;;�A;a�E;��G;έH;�
I;C I;�I;�I;�I;�I;�I;e�H;�H;��H;x�H;��H;��H;O�H;�H;K�H;��H;��H;w�H;��H;�H;h�H;�I;�I;�I;�I;�I;D I;�
I;ѭH;��G;k�E;�A;
;;}�/;Ob;��;�4�:�>:P��ZP��m�@�ʵ���׻1B��3/���O�D�k���p8��      ������q
� ���8�׻ ,��ʮ��;��lۺL� ��O�9�Ȋ:��:z;!;��0;;;��A;�pE;J�G;��H;��H;�I;I;,I;�I;�I;RI;��H;"�H;W�H;��H;��H;��H;��H;F�H;�H;C�H;��H;��H;��H;��H;Z�H;(�H;��H;RI;�I;�I;2I;I;�I;��H;��H;P�G;�pE;��A;
;;��0;!;|;	��:�Ȋ:P�9@� ��lۺ;�ͮ���+��4�׻"����q
���      (/��(��� �x���X���/�� ����0o�p9�9��k:��:o�:�B;�&;:3;k<;�A;�pE;<tG;�|H;�H;I;LI; I;�I;J
I;�I;0 I;*�H;�H;��H;^�H;��H;��H;��H;X�H;C�H;V�H;��H;��H;��H;Z�H;��H;�H;)�H;1 I;�I;F
I;�I;"I;JI;I;�H;�|H;?tG;�pE;�A;i<;<3;�&;�B;!o�:��:��k:p9�9@o����� ���/���X��x�(���      X���셍�uk�ș �����,69��!:rȊ:b4�:��:��;�;?�,;��6;��=;��B;h�E;S�G;�|H;p�H;SI;�I;\I;6I;�I;I;fI;&�H;��H;�H;��H;��H;��H;��H;��H;o�H;S�H;h�H;��H;��H;��H;��H;��H;�H;��H;(�H;cI;�I;�I;6I;[I;�I;WI;q�H;�|H;O�G;k�E;��B;��=;��6;A�,;�;��;��:f4�:|Ȋ:��!:0-69h��� �,uk�����      D�>:,�G:X�b:X��:��:�4�:�*�:xi;7�;�a;*;9r3;��:;�!@;��C;�IF;��G;��H;�H;OI;�I;I;I;�I;�I;7I;��H;k�H;��H;X�H;*�H;��H;z�H;��H;��H;��H;c�H;��H;��H;��H;y�H;��H;-�H;Z�H;��H;j�H;��H;6I;�I;�I;I;I;�I;QI;�H;��H;��G;�IF;��C;�!@;��:;<r3;
*;�a;4�;ti;�*�:�4�:+��:^��:��b:8�G:      Yt�:� �:9l�:A�;� 
;Є;z;�O$;H�,;��3;�9;��>;
�B;2E;��F;KH;ѭH;��H;I;�I;I;YI;I;�I;�I;��H;�H;.�H;��H;x�H;��H;��H;o�H;��H;�H;��H;��H;��H;�H;��H;o�H;��H;��H;y�H;��H;.�H;��H;��H;�I;�I;I;ZI;!I;�I;I;��H;խH;LH;��F;2E;�B; �>;�9;��3;G�,;P$;"z;ʄ;� 
;8�;%l�:s �:       p ;�!;�#;�&;�*;�o.;_3;��7;Y�;;
j?;8kB;�D;ixF;��G;�cH;�H;�
I;�I;LI;^I;I;I;�I;7I;�H;n�H;n�H;	�H;��H;��H;��H;c�H;r�H;��H;6�H;�H;��H;��H;5�H;��H;r�H;`�H;��H;��H;��H;�H;k�H;o�H;�H;3I;�I;I;I;^I;NI;�I;�
I;�H;�cH;��G;jxF;�D;>kB;j?;[�;;��7;^3;�o.;�*;�&;�#;�!;      �J6;�6;��7;v9;=;;.=;Aj?;P�A;�C;N2E;��F;H�G;n<H;{�H;��H;�I;A I;I;"I;3I;�I;�I;2I;,�H;��H;��H;@�H;�H;�H;��H;g�H;T�H;t�H;	�H;��H;S�H;*�H;M�H;��H;	�H;t�H;Q�H;j�H;��H;�H;�H;<�H;��H;��H;)�H;/I;�I;�I;0I; I;I;D I;�I;��H;{�H;n<H;J�G;��F;P2E;�C;X�A;Bj?;�-=;L;;v9;��7;�6;      �DA;�kA;J�A;a�B;�jC;JaD;y\E;�IF;�G;��G;]NH;(�H;��H;�I;qI;V I;�I;6I;�I;�I;�I;�I;�H;��H;��H;\�H;�H;/�H;��H;x�H;M�H;e�H;��H;A�H;��H;��H;��H;��H;��H;A�H;��H;_�H;O�H;x�H;��H;.�H;�H;]�H;��H;��H;�H;�I;�I;�I;�I;2I;�I;V I;qI;�I;��H;.�H;^NH;��G;�G;�IF;y\E;@aD;�jC;g�B;L�A;�kA;      WIF;pYF;��F;��F;r'G;��G;��G;CH;�H;B�H;T�H;�I;�I;� I;�I;�I;�I;�I;G
I;I;:I;��H;k�H;��H;[�H;7�H;A�H;��H;y�H;\�H;F�H;��H;�H;|�H;6�H;�H;�H;�H;3�H;|�H;�H;��H;F�H;Y�H;v�H;��H;?�H;;�H;]�H;��H;k�H;��H;:I;�I;G
I;�I;�I;�I;�I;� I;�I;�I;]�H;C�H;�H;CH;��G;��G;�'G;��F;��F;oYF;      �NH;�TH;�dH;�}H;ɛH;P�H;��H;��H;�I;I;�I;!I;lI;.I;�I;I;�I;�I;�I;hI;�H;��H;l�H;D�H;�H;?�H;��H;}�H;K�H;L�H;��H;��H;U�H;��H;��H;��H;w�H;��H;��H;��H;U�H;��H;��H;J�H;G�H;|�H;��H;D�H;�H;@�H;l�H;��H;�H;cI;�I;�I;�I;I;�I;+I;mI;!I;  I;I;�I;��H;��H;L�H;�H;�}H;�dH;uTH;      ��H;F�H;�I;�	I;�I;�I;RI;� I;�!I;T I;kI;�I;�I;�I;�I;9
I;�I;OI;0 I;&�H;k�H;)�H;�H;�H;(�H;��H;{�H;\�H;B�H;s�H;��H;2�H;��H;q�H;0�H;�H;��H;��H;0�H;r�H;��H;/�H;��H;r�H;?�H;[�H;x�H;��H;,�H;�H;�H;,�H;k�H;&�H;. I;NI;�I;<
I;�I;�I;�I;�I;mI;U I;�!I;� I;RI;�I;�I;�	I;�I;;�H;      �!I;�!I;!"I;B"I;�!I;!I;�I;EI;�I;�I;�I;lI;I;�
I;�I;�I;�I;��H;.�H;��H;��H;��H;��H;�H;��H;r�H;D�H;D�H;��H;��H;�H;��H;=�H;��H;��H;��H;��H;��H;��H;��H;A�H;��H;"�H;��H;��H;B�H;@�H;t�H;��H;�H;��H;��H;��H;��H;.�H;��H;�I;�I;�I;�
I;I;lI;�I;�I;�I;EI;�I;!I;�!I;D"I;"I;�!I;      �I;�I;�I;I;�I;:I;kI;ZI;%I;�I;I;i
I;�I;I;�I;  I;j�H;�H;��H;�H;^�H;t�H;��H;��H;t�H;Q�H;G�H;u�H;��H;�H;��H;<�H;��H;��H;_�H;@�H;/�H;?�H;\�H;��H;��H;9�H;��H;�H;��H;s�H;C�H;V�H;x�H;��H;��H;u�H;[�H;�H;�H;�H;l�H; I;�I;I;�I;f
I;I;�I;(I;XI;pI;:I;�I;I;�I;�I;      �I;�I;KI;�I;qI;'I;�I;�I;	I;	I;�I;�I;�I;X I;%�H;�H;"�H;[�H;��H;��H;3�H;��H;��H;j�H;M�H;C�H;��H;��H;&�H;��H;�H;��H;l�H;1�H;�H;��H;��H;��H; �H;4�H;m�H;��H;�H;��H;"�H;��H;��H;G�H;O�H;g�H;��H;��H;0�H;��H;��H;[�H;$�H;�H;'�H;Z I;�I;�I;�I;	I;
I;�I;�I; I;~I;�I;II;�I;      }I;nI;I;nI;�
I;�	I;VI;	I;wI;�I; I;C I;n�H;��H;��H;8�H;��H;��H;b�H;��H;��H;��H;a�H;R�H;c�H;��H;��H;3�H;��H;=�H;��H;M�H;�H;��H;��H;��H;��H;��H;��H;��H;�H;J�H;��H;:�H;��H;0�H;��H;��H;e�H;K�H;e�H;��H;��H;��H;a�H;��H;��H;;�H;��H;��H;p�H;B I;'I;�I;vI;I;^I;�	I;�
I;vI;I;lI;      UI;3I;�I;UI;�I;�I;�I;{I;I;��H;D�H;��H;V�H;��H;s�H;��H;~�H;�H;��H;��H;��H;t�H;r�H;t�H;��H;�H;U�H;��H;F�H;��H;i�H;�H;��H;��H;��H;d�H;^�H;d�H;~�H;��H;��H;�H;h�H;��H;A�H;��H;V�H;�H;��H;s�H;w�H;r�H;��H;��H;��H;�H;�H;��H;v�H;��H;Z�H;��H;J�H;��H; I;{I;�I;�I;�I;RI;�I;0I;      �I;�I;�I;I;~I;� I;��H;��H;��H;��H;��H;�H;�H;��H;d�H;�H;��H;��H;��H;��H;��H;��H;��H;�H;<�H;x�H;��H;u�H;��H;��H;-�H;��H;��H;e�H;P�H;A�H;4�H;A�H;O�H;g�H;��H;��H;.�H;�H;��H;q�H;��H;y�H;>�H;�H;��H;��H;��H;��H;��H;��H;��H;�H;d�H;��H;�H;�H;��H;��H;��H;��H;  I;� I;�I;I;�I;�I;      B I;M I;��H;��H;,�H;u�H;��H;��H;��H;��H;��H;��H;V�H;G�H;'�H;�H;��H;��H;��H;��H;��H;�H;4�H;��H;��H;,�H;��H;2�H;��H;c�H;��H;��H;��H;O�H;-�H;�H;"�H;�H;)�H;P�H;��H;��H;��H;\�H;��H;.�H;��H;/�H;��H;��H;8�H;�H;��H;��H;��H;��H;��H;�H;'�H;H�H;Y�H;��H;��H;��H;��H;��H;��H;x�H;-�H;��H;��H;P I;      ��H;��H;T�H;��H;�H;��H;H�H;u�H;��H;��H;��H;��H;�H;w�H;d�H;Y�H;Q�H;@�H;X�H;m�H;��H;��H;��H;E�H;��H;�H;��H;�H;��H;F�H;��H;��H;i�H;B�H;#�H;�H;�H;�H;�H;F�H;l�H;��H;��H;@�H;��H;��H;��H;�H;��H;E�H;��H;��H;��H;h�H;W�H;F�H;R�H;\�H;d�H;x�H;�H;��H;��H;��H;��H;u�H;S�H;��H;��H;��H;O�H;��H;      �H;��H;��H;c�H;��H;:�H;��H;��H;�H;5�H;Q�H;H�H;T�H;.�H;�H;�H;�H;�H;F�H;Y�H;m�H;��H;��H;#�H;��H;��H;t�H;��H;��H;5�H;��H;��H;a�H;1�H;#�H;�H;�H;�H; �H;3�H;e�H;��H;��H;/�H;��H;��H;w�H; �H;��H;"�H;��H;��H;g�H;U�H;F�H;�H;�H;�H;�H;.�H;T�H;G�H;V�H;6�H;�H;��H;��H;;�H;��H;h�H;��H;��H;      ��H;��H;N�H;��H;��H;��H;H�H;u�H;��H;��H;��H;��H;��H;x�H;d�H;Y�H;Q�H;@�H;X�H;m�H;��H;��H;��H;E�H;��H;�H;��H;�H;��H;D�H;��H;��H;k�H;C�H;#�H;�H;�H;�H;�H;E�H;l�H;��H;��H;?�H;��H;��H;��H;�H;��H;C�H;��H;��H;��H;g�H;W�H;D�H;Q�H;\�H;d�H;v�H;�H;��H;��H;��H;��H;x�H;P�H;��H;��H;�H;T�H;��H;      7 I;P I;��H;��H;-�H;t�H;��H;��H;��H;��H;��H;��H;Y�H;G�H;'�H;�H;��H;��H;��H;��H;��H;�H;2�H;��H;��H;*�H;��H;0�H;��H;b�H;��H;��H;��H;O�H;,�H;�H;"�H; �H;*�H;P�H;��H;��H;��H;\�H;��H;,�H;��H;0�H;��H;��H;8�H;�H;��H;��H;��H;��H;��H;�H;$�H;G�H;V�H;��H;��H;��H;��H;��H;��H;u�H;3�H;��H;  I;Q I;      �I;�I;�I;I;I;� I;��H;��H;��H;��H;��H;�H;�H;��H;d�H;�H;��H;��H;��H;��H;��H;��H;��H;�H;>�H;x�H;��H;t�H;��H;��H;-�H;��H;��H;e�H;S�H;?�H;4�H;A�H;O�H;g�H;��H;��H;-�H;��H;��H;q�H;��H;{�H;>�H;��H;��H;��H;��H;��H;��H;��H;��H;�H;d�H;��H;�H;~�H;��H;��H;��H;��H;  I;� I;�I;I;�I;�I;      SI;7I;�I;RI;�I;�I;�I;�I;I;��H;C�H;��H;Y�H;��H;v�H;��H;~�H;�H;��H;��H;��H;t�H;n�H;s�H;��H;�H;S�H;��H;G�H;��H;f�H;�H;��H;��H;��H;e�H;^�H;e�H;��H;��H;��H;�H;h�H;��H;?�H;��H;V�H;�H;��H;q�H;x�H;q�H;}�H;��H;��H;��H;~�H;��H;s�H;��H;Z�H;��H;G�H;��H;I;~I;�I;�I;�I;XI;�I;3I;      oI;nI;I;oI;�
I;�	I;[I;I;qI;�I;$I;E I;p�H;��H;��H;9�H;��H;��H;a�H;��H;��H;��H;a�H;O�H;e�H;��H;��H;2�H;��H;<�H;��H;J�H;�H;��H;��H;��H;��H;��H;��H;��H;�H;L�H;��H;:�H;��H;/�H;��H;��H;c�H;J�H;e�H;��H;��H;��H;`�H;��H;��H;9�H;��H;��H;p�H;B I;"I;�I;tI;I;[I;�	I;�
I;vI;I;hI;      �I;�I;GI;�I;wI;&I;�I;�I;	I;	I;�I;�I;�I;X I;'�H;�H;$�H;[�H;��H;��H;3�H;��H;��H;h�H;N�H;@�H;��H;��H;&�H;��H;�H;��H;l�H;2�H;�H;��H;��H;��H;�H;5�H;m�H;��H;�H;��H;!�H;��H;��H;G�H;M�H;d�H;��H;��H;/�H;��H;��H;[�H;%�H;�H;(�H;X I;�I;�I;�I;	I;
I;�I;�I;"I;�I;�I;NI;�I;      �I;�I;�I;I;�I;EI;kI;^I;(I;�I;I;g
I;�I;I;�I; I;j�H;�H;��H;�H;^�H;u�H;��H;��H;v�H;O�H;F�H;s�H;��H;�H;��H;<�H;��H;��H;b�H;?�H;/�H;B�H;^�H;��H;��H;=�H;��H;�H;��H;s�H;G�H;V�H;u�H;��H;��H;u�H;Z�H;�H;�H;�H;j�H; I;�I;I;�I;f
I;I;�I;'I;[I;pI;7I;�I;!I;�I;I;      �!I;�!I;-"I;<"I;�!I;!I;I;DI;�I;�I;�I;jI;I;�
I;�I;�I;�I;��H;*�H;��H;��H;��H;��H;�H;��H;n�H;A�H;C�H;��H;��H;!�H;��H;?�H;��H;��H;��H;��H;��H;��H;��H;@�H;��H;"�H;��H;��H;@�H;D�H;r�H;��H;�H;��H;��H;��H;��H;0�H;��H;�I;�I;�I;�
I;I;hI;�I;�I;�I;EI;�I;!I;�!I;<"I;-"I;�!I;      ��H;<�H;uI;�	I;�I;�I;SI;� I;�!I;R I;hI;�I;�I;�I;�I;7
I;�I;OI;, I;#�H;k�H;*�H;�H;�H;+�H;��H;x�H;[�H;C�H;r�H;��H;2�H;��H;q�H;3�H;��H;��H;�H;0�H;r�H;��H;2�H;��H;s�H;@�H;Y�H;{�H;��H;'�H;�H;	�H;*�H;j�H;&�H;0 I;KI;�I;9
I;I;�I;�I;�I;lI;T I;�!I;� I;SI;�I;�I;�	I;�I;<�H;      �NH;�TH;�dH;�}H;؛H;S�H;��H;��H;�I;I;�I;!I;jI;+I;�I;I;�I;�I;�I;cI;�H;��H;g�H;D�H;�H;<�H;��H;}�H;K�H;I�H;��H;��H;S�H;��H;��H;��H;w�H;��H;��H;��H;U�H;��H;��H;L�H;H�H;|�H;��H;C�H;�H;@�H;p�H; �H;��H;fI;�I;�I;�I;I;�I;+I;jI;!I;�I;I;I;��H;��H;O�H;ߛH;�}H;�dH;TH;      MIF;lYF;��F;��F;y'G;ÈG;��G;CH;�H;A�H;X�H;�I;�I;� I;�I;�I;�I;�I;G
I;�I;:I;��H;g�H;��H;[�H;3�H;?�H;��H;{�H;Y�H;F�H;��H;�H;}�H;6�H;�H;	�H;�H;3�H;|�H;�H;��H;I�H;[�H;v�H;��H;D�H;8�H;[�H;��H;n�H;��H;9I;�I;H
I;�I;�I;�I;�I;� I;�I;�I;[�H;C�H;�H;CH;��G;��G;�'G;��F;��F;_YF;      �DA;�kA;F�A;d�B;�jC;MaD;w\E;�IF;�G;��G;[NH;+�H;��H;�I;rI;V I;�I;5I;�I;�I;�I;�I;�H;��H;��H;U�H;�H;.�H;��H;v�H;M�H;e�H;��H;A�H;��H;��H;��H;��H;��H;C�H;��H;f�H;T�H;y�H;��H;.�H;�H;\�H;��H;��H;�H;�I;�I;�I;�I;2I;�I;W I;tI;�I;��H;(�H;ZNH;��G;~G;�IF;y\E;?aD;�jC;f�B;E�A;�kA;      �J6;��6;��7;�9;7;;.=;Ej?;Q�A;�C;J2E;��F;I�G;m<H;w�H;��H;�I;A I;I;I;/I;�I;�I;,I;*�H;��H;��H;<�H;�H;�H;��H;h�H;U�H;v�H;	�H;��H;Q�H;,�H;S�H;��H;�H;z�H;X�H;n�H;��H;�H;�H;A�H;��H;��H;*�H;0I;�I;�I;2I;"I;I;D I;�I;��H;y�H;m<H;I�G;��F;M2E;�C;L�A;Dj?;.=;O;;�9;��7;�6;      p ;�!;�#;�&;�*;�o.;[3;��7;_�;;	j?;2kB;�D;fxF;��G;�cH;�H;�
I;�I;KI;[I;I;I;�I;3I;�H;e�H;i�H;�H;��H;��H;��H;e�H;q�H;��H;9�H;�H;��H;�H;4�H;��H;u�H;h�H;��H;��H;��H;�H;r�H;n�H;�H;4I;�I;I;I;^I;OI;�I;�
I;�H;�cH;��G;jxF;�D;5kB;	j?;\�;;��7;[3;�o.;�*;�&;�#;�!;      Ot�:� �:l�::�;� 
;ք; z;P$;G�,;��3;�9;�>;	�B;2E;��F;KH;ЭH;��H;I;�I;I;WI;I;�I;�I;��H;��H;.�H;��H;t�H;��H;��H;o�H;��H;�H;��H;��H;��H;�H;��H;u�H;��H;��H;{�H;��H;.�H;�H;��H;�I;�I;I;YI;!I;�I;I;��H;ҭH;LH;��F;2E;	�B;��>;�9;��3;G�,; P$;z;��;� 
;,�;l�:s �:      �>:��G:��b:f��:��:�4�:�*�:zi;:�;�a;	*;=r3;��:;�!@;��C;�IF;��G;��H;�H;PI;�I;I;I;�I;�I;0I;��H;i�H;��H;T�H;)�H;��H;z�H;��H;��H;��H;f�H;��H;��H;��H;}�H;��H;0�H;[�H;��H;k�H;��H;6I;�I;�I;I;I;�I;SI;�H;��H;��G;�IF;��C;�!@;��:;9r3;*;�a;6�;zi;�*�:�4�:=��:b��:��b:D�G:      2���慍�,uk��� ����0-69��!:�Ȋ:l4�:��:��;�;@�,;��6;��=;��B;h�E;P�G;�|H;p�H;TI;�I;ZI;2I;�I;�I;_I;$�H;��H;�H;��H;��H;��H;��H;��H;k�H;V�H;m�H;��H;��H;��H;��H;��H;�H;��H;'�H;hI;I;�I;7I;aI;�I;TI;q�H;�|H;O�G;k�E;��B;��=;��6;?�,;�;��;��:b4�:|Ȋ:��!:�,69h���� �,uk��      '/��(���!�x���X���/�� ����0o�p9�9��k:��:o�:�B;�&;=3;m<;�A;�pE;;tG;�|H;�H;I;KI;I;�I;C
I;�I;- I;)�H;��H;��H;]�H;��H;��H;��H;V�H;C�H;W�H;��H;��H;��H;^�H;��H;�H;*�H;0 I;�I;F
I;�I;#I;NI;I;�H;�|H;<tG;�pE;�A;j<;<3;�&;�B;o�:��:��k:p9�9(o����� ���/���X�'�x�&���      ������q
� ���8�׻�+��ʮ�� ;��lۺL� ��O�9�Ȋ:��:z;!;��0;;;��A;�pE;M�G;��H;��H;�I;I;,I;�I;�I;OI;��H;�H;X�H;��H;��H;��H;��H;D�H;�H;F�H;��H;��H;��H;��H;Z�H;"�H;��H;SI;�I;�I;+I;I;�I;��H;��H;P�G;�pE;��A;	;;��0;!;z;��:�Ȋ: P�9T� ��lۺ;�̮�� ,��7�׻"����q
���      ����q8����A�k���O��3/�1B��׻ʵ��m�@�\P��H���>:�4�:��;Rb;}�/;;;�A;f�E;��G;έH;�
I;A I;�I;�I;�I;�I;�I;b�H;�H;��H;x�H;��H;��H;N�H;�H;N�H;��H;��H;w�H;��H;�H;e�H;�I;�I;�I;�I;�I;C I;�
I;έH;��G;j�E;�A;
;;|�/;Ob;��;�4�:�>:`��ZP��n�@�ɵ���׻1B��3/���O�C�k���p8��      ;���|�2�ݼ��˼d���,���}��G����H�һ����k���/�L:׳:�;Ib;��0;i<;�B;�IF;IH;�H;�I;L I;�I;I;2
I;�I;��H;�H;5�H;��H;�H;�H;Y�H;�H;Y�H;��H;�H;��H;4�H;�H;  I;�I;6
I;I;�I;I I;�I;�H;KH;�IF;��B;i<;��0;Lb;�;׳:X:�/�o������F�һ����G��}��,��d����˼4�ݼ }�      E�B�MR?��5���&��3��J��ծҼ!F����A=�#?�.����/��nk����9׳:��;!;83;��=;��C;��F;�cH;��H;kI;�I;�I;�I;�I;�I;!�H;��H;r�H;b�H; �H;b�H;�H;d�H;�H;`�H;r�H;��H;!�H;�I;�I;�I;�I;�I;jI;��H;�cH;��F;��C;��=;63;!;��;׳:���9�nk���/�.��"?�B=���!F��ծҼ�J���3���&��5�MR?�      (��%W��蒐�$�����j�R`I���&����Dϼ�,���T[�m�pI��j;��nk�d:�4�:z;�&;��6;�!@;2E;��G;{�H;�I;� I;+I;�I;�
I;I;S I;��H;��H;��H;?�H;s�H;&�H;v�H;:�H;��H;��H;��H;P I;I;�
I;�I;)I;� I;�I;~�H;��G;2E;�!@;��6;�&;|;�4�:X:�nk�k;�rI��n��T[��,��Dϼ�����&�R`I���j�$���蒐�%W��      �J�����D��ͽ���'�������L�&��&��
;���k����pI����/��/��>:��:�B;?�,;��:;	�B;ixF;r<H;��H;�I;jI;�I;I;�I;�I;m�H;W�H;�H;N�H;~�H;M�H;~�H;L�H;�H;U�H;j�H;�I;�I;I;�I;lI;�I;��H;q<H;mxF;	�B;��:;C�,;�B;	��:�>:�/���/�pI������k�
;��&��%����L����'������ͽ�D����      Q�:��*7���,�+���	�r�齂���!W����j�?�/��J���I���k�n�.��k��x���Ȋ:!o�:�;Cr3;��>;�D;J�G;"�H;�I;
!I;�I;eI;]
I;�I;< I;��H;{�H;��H;��H;A�H;��H;��H;z�H;��H;< I;�I;b
I;hI;�I;!I;�I;�H;J�G;�D;��>;9r3;�;o�:�Ȋ:h��m��.��n��k��I���J��?�/���j�!W������q�齂�	�+���,��*7�      ^���p����1�l���M���,�Xl�Q9ݽ�A���{���5��J��
;���T[�#?�����nP���O�9��:��;*; �9;2kB;��F;SNH;S�H;�I;cI;�I;�I;�I; I;C�H;��H;��H;��H;J�H;��H;��H;��H;C�H;I;�I; I;�I;eI;�I;Q�H;PNH;��F;2kB;��9; *;��;��:�O�9dP������$?��T[�
;���J����5��{��A��R9ݽXl���,���M�1�l����p��      4m־P�Ѿ�>ľ����ӗ����{��I�+�����V���{�?�/�&���,��A=�F�һr�@�p� ���k:��:�a;��3;j?;M2E;��G;<�H;I;J I;�I;�I;�I;�I;��H;��H;��H;��H;8�H;��H;��H;��H;��H;�I;�I;�I;�I;K I;I;<�H;��G;J2E;j?;��3;�a;��:|�k:d� �r�@�F�һB=��,��&��?�/��{��V�����+��I���{�ӗ�������>ľP�Ѿ      C\����r5��z ��E۾ֳ�^��y�Z�L?#����A����j�&��Eϼ�����е���lۺ89�9^4�:;�;@�,;Q�;;�C;}G;�H;|I;�!I;�I;"I;I;qI;#I;��H;��H;��H;�H;��H;��H;��H; I;sI;I;$I;�I;�!I;|I;�H;zG;�C;R�;;@�,;4�;`4�:(9�9�lۺε�������Eϼ&����j��A�����L?#�y�Z�^��ֳ��E۾�z �r5����      E�b��>]���M�Î6�����$���>ľ"q��y�Z�+�R9ݽ!W����L����"F���G��׻;�ho�vȊ:zi;�O$;��7;Q�A;�IF;�BH;��H;� I;@I;TI;�I;I;I;��H;��H;q�H;��H;q�H;��H;��H;~I;I;�I;ZI;@I;� I;��H;CH;�IF;M�A;��7;�O$;ri;zȊ:�o�;��׻�G�#F�������L�!W��R9ݽ+�y�Z�"q���>ľ�$�����Î6���M��>]�      p��񲗿���6�y�{�R���)�nv��>ľ^���I�Xl����������&�ծҼ�}�3B�Ү��*���l�!:�*�:z;R3;Dj?;l\E;��G;��H;EI;|I;jI;�I;VI;�I;��H;��H;A�H;��H;A�H;��H;��H;�I;WI;�I;nI;~I;GI;��H;��G;k\E;Dj?;W3;z;�*�:t�!:,���Ю��2B��}�ծҼ��&��������Xl��I�^���>ľnv���)�{�R�6�y����񲗿      �˿�<ƿpL��@1����>]���)��$��ֳ���{���,�r��'��R`I��J���,���3/�,��� ��,69�4�:ʄ;�o.;
.=;9aD;��G;L�H;�I;!I;?I;,I;�	I;�I;� I;�H;��H;B�H;��H;~�H;� I;�I;�	I;'I;BI;!I;�I;O�H;��G;8aD;
.=;�o.;Ȅ;�4�:�,69#� �,���3/��,���J��R`I�'��r�齤�,���{�ֳ��$����)��>]��@1��pL���<ƿ      ����<���U[忶˿�T���{�R�����E۾ӗ����M���	������j��3�d����O�@�׻��/����1��:� 
;�*;I;;�jC;w'G;ћH;�I;�!I;�I;vI;�
I;�I;�I;�H;��H;��H;��H;�H;I;�I;�
I;sI;�I;�!I;�I;֛H;�'G;�jC;I;;�*;� 
;%��:p����/�?�׻��O�d���3���j������	���M�ӗ���E۾���{�R���T���˿U[�<���      O�6��t����˿@1��6�y�Î6��z �����1�l�+��ͽ$�����&���˼B�k�(�����X�� �l��:1�;�&;w9;f�B;��F;�}H;�	I;/"I;I;�I;xI;QI;"I;��H;�H;a�H;��H;��H; I;RI;yI;�I;I;/"I;�	I;�}H;��F;d�B;y9;�&;0�;b��:� ���X�&���B�k���˼��&�$����ͽ+�1�l������z �Î6�6�y�@1���˿���t�6��      ��*��g&��#�t�U[�pL�������M�r5��>ľ����,��D�钐��5�3�ݼ���q
� �x�8uk���b:l�:�#;7;P�A;��F;�dH;�I;!"I;�I;DI;I;�I;�I;��H;X�H;��H;T�H;��H;�I;�I;I;@I;�I;!"I;�I;�dH;��F;O�A;��7;�#;l�:��b:(uk�"�x��q
���3�ݼ�5�钐��DὪ�,����>ľr5���M����pL��U[�t��#��g&�      ��8��4��g&�6��<����<ƿ񲗿�>]�®�P�Ѿ�p���*7����%W��MR?�}�s8����"�������x�G:g �:�!;�6;�kA;aYF;�TH;B�H;�!I;�I;�I;gI;(I;�I;; I;��H;��H;��H;; I;�I;(I;hI;�I;�I;�!I;C�H;�TH;lYF;�kA;�6;�!;c �:l�G:څ��#�����s8��}�MR?�%W�����*7��p��P�Ѿ®��>]�񲗿�<ƿ<���6���g&��4�      ��$������꿯�ſ�ޞ�%3s��2�=����� j���yHͽŸ����'�C<ͼt�n�j���IQ^�..�b��:fW;ZS%;ao8;��A;DF;�H;y�H;��H;��H;�H;�H;!�H;��H;��H;��H;
�H;��H;��H;��H;!�H;�H;�H;��H;��H;y�H;�H;DF;��A;^o8;QS%;cW;^��:..�KQ^�h���t�n�C<ͼ��'�Ÿ��zHͽ�� j���=����2�%3s��ޞ���ſ������$�      $�������忇�����cm�V�-�����Qh��Vde�"-�תɽ�v��)�$���ɼ}mj�<���X�@���ņ:`x;�%;,�8;?B;RF;�H;�H;�H;��H;C�H;�H;�H;u�H;��H;��H;�H;��H;��H;u�H;�H;�H;>�H;��H;�H;�H;�H;%RF;?B;*�8;��%;]x;�ņ:4��X�<���}mj���ɼ(�$��v��תɽ"-�Vde�Qh������V�-�cm��������忝����      ����������ԿLw�����:�\�"����k��Z0X�����;����w����������]�$���F�(���ɒ:��;��';��9;�oB;|zF;�!H;p�H;��H; �H;n�H;�H;�H;}�H;��H;��H;��H;��H;��H;}�H;�H;�H;h�H;�H;��H;n�H;�!H;�zF;�oB;��9;��';��;�ɒ:����F�$�黮�]����������w��;�����Z0X�k�����"�:�\����Lw���Կ��𿝏�      ������Կp���ޞ�`F�h�C�-E�"�;�I��D���"��g�c�}��֯���J��ѻآ)�P�K���:�
;�M*;i�:;�C;øF;�8H;*�H;G�H;W�H;��H;�H;�H;�H;��H;��H;��H;��H;��H;}�H;�H;�H;��H;[�H;F�H;&�H;�8H;ʸF;�C;e�:;�M*;�
;��:�K�ڢ)��ѻ��J��֯�}�g�c�"����D��I��"�;-E�h�C�`F��ޞ�p���Կ��      ��ſ���Lw���ޞ�����>�W�5�%�����hɰ��|x�g{+�ұ����J��  �ж��\�1�,���&+��
9��:��;ڷ-;��<;W�C;�G;�TH;!�H;��H;��H;��H;+�H;�H;d�H;��H;t�H;��H;o�H;��H;a�H;�H;'�H;��H;��H;��H; �H;�TH;�G;V�C;~�<;շ-;��;��:�
9)+�,���]�1�ж���  ��J���ұ�g{+��|x�hɰ�����5�%�>�W������ޞ�Lw�����      �ޞ�������_F�>�W�W�-���?Kɾ�G����O����ƽǸ��΄-���ۼㄼ84� ǐ�϶��\:��:x;v�1;�c>;>�D;r\G;)sH;s�H;3�H;A�H;��H;H�H;
�H;G�H;j�H;]�H;��H;Y�H;h�H;D�H;	�H;G�H;��H;F�H;0�H;s�H;'sH;y\G;=�D;�c>;r�1;v;ؤ�:]:϶� ǐ�84�ㄼ��ۼ΄-�Ǹ��ƽ�����O��G��?Kɾ��W�-�>�W�_F�������      %3s�cm�:�\�h�C�5�%����TҾj��
 j��C(����_P����[�}������Y�?��lX���<���k:(��:�� ;Ο5;+R@;1uE;ʲG;�H;�H;��H;��H;�H;D�H;�H;@�H;L�H;7�H;k�H;4�H;K�H;@�H;�H;A�H;�H;��H;��H;�H;�H;ѲG;1uE;*R@;̟5;�� ;��:��k:��<�mX�>����Y����}���[�_P����콪C(�
 j�j���TҾ��5�%�h�C�:�\�cm�      �2�V�-�"�-E�����?Kɾj����s�8�5���v㻽�v��
z0��;��+���*����96��CS�9M�:I�	;j�(;�9;�/B;CDF;H;��H;X�H;��H;��H;I�H;b�H;��H;�H;�H;�H;9�H;�H;�H;�H;��H;_�H;G�H;��H;��H;X�H;��H;H;DDF;�/B;�9;j�(;A�	;AM�: DS�96�����*��+���;�
z0��v��v㻽��8�5���s�j��?Kɾ����-E�"�V�-�      =����������"�;hɰ��G��
 j�8�5��	�ϪɽY����J�t���沼��]�����	x�b	�� n:z��:�v;��/;]-=;��C;�F;�HH;z�H;��H;��H;��H;x�H;d�H;��H;��H;��H;��H;�H;��H;��H;��H;��H;d�H;x�H;�H;��H;��H;w�H;�HH;�F;��C;a-=;��/;�v;���: n:j	���	x������]��沼t���J�Y���Ϫɽ�	�8�5�
 j��G��hɰ�"�;��徶���      ��Qh��k���I���|x���O��C(���Ϫɽ����RDX�I��(<ͼ
ㄼ�X!��s���W�0vK���:�y;��#;�H6;R@;�PE;b�G;V�H;��H;�H;��H;z�H;��H;R�H;��H;��H;��H;��H;��H;��H;��H;��H;��H;N�H;��H;��H;��H;�H;��H;V�H;g�G;�PE;R@;�H6;�#;�y;��:`vK��W��s���X!�
ㄼ(<ͼI��RDX�����Ϫɽ���C(���O��|x��I��k��Qh��       j�Vde�Z0X�D�g{+�������v㻽Z���RDX������ۼ̾����;�J>ۻ)X���y��>":���:��;��-;~�;;��B;izF;�H;Z�H;T�H;��H;��H;��H;��H;K�H;��H;z�H;q�H;��H;[�H;��H;r�H;|�H;��H;G�H;��H;��H;��H;��H;T�H;Y�H;�H;ezF;��B;~�;;��-;��;���:�>":|�y�)X�K>ۻ��;�̾����ۼ���RDX�Y���v㻽��콂��g{+�D�Z0X�Vde�      ��"-������ұ�ƽ^P���v���J�I����ۼ��f�J������+���rѺ�'
9�M�:��;l $;��5;��?;X�D;<\G;�eH;��H;��H;��H;��H;��H;��H;0�H;R�H;9�H;2�H;D�H;�H;D�H;2�H;<�H;O�H;.�H;��H;�H;��H;��H;��H;��H;�eH;<\G;\�D;��?;��5;v $;��;�M�:�'
9�rѺ�+������f�J�����ۼI���J��v��^P��ƽұ轄����"-�      yHͽתɽ�;��"����Ǹ����[�	z0�s��'<ͼ̾��f�J�����j���*��ب�:0b�:2�;��/;zL<;�C;�lF;k�G;סH;��H;��H;��H;�H;.�H;��H;�H;�H;��H;��H;��H;��H;��H;��H;��H;�H;�H;��H;5�H;�H;��H;��H;��H;ݡH;k�G;mF;�C;zL<;��/;5�;$b�:ਂ: ��*��j�����e�J�̾��'<ͼs��	z0���[�Ǹ����"���;��תɽ      Ÿ���v����w�g�c��J�τ-�|��;缆沼	ㄼ��;������j���5�����>Q:$��:Ii;�M*;`�8;a�@;�PE;�uG;iH;��H;��H;��H;��H;��H;S�H;��H;��H;��H;��H;��H;��H;��H;��H;��H;��H;��H;��H;��H;[�H;��H;��H;��H;��H;��H;iH;�uG;�PE;`�@;h�8;�M*;Gi;0��:�>Q:��깬5��j��������;�	ㄼ�沼�;�|�΄-��J�g�c���w��v��      ��'�)�$����}��  ���ۼ����+����]��X!�H>ۻ�+���*���깬�>:���:��;�%;ʟ5;s�>;(D;��F;P!H;�H;'�H;��H;��H;��H;��H;I�H;��H;��H;i�H;m�H;I�H;4�H;N�H;2�H;G�H;p�H;i�H;��H;��H;P�H;��H;��H;��H;��H;*�H;�H;R!H;��F;(D;z�>;Ο5;�%;��;���:��>:��깅*��+��G>ۻ�X!���]��+�������ۼ�  �}����)�$�      @<ͼ��ɼ�����֯�϶��ㄼ��Y��*�����s��$X��rѺ0��>Q:���:��
;.�#;K�3;nc=;�#C;DF;��G;�H;��H;��H;�H;��H;3�H;��H;C�H;l�H;C�H;�H;1�H;��H;��H;��H;��H;��H;1�H;�H;@�H;p�H;G�H;��H;5�H;��H;�H;��H;��H;�H;��G;DF;�#C;qc=;F�3;/�#;��
;���:�>Q:@��rѺ X��s������*���Y�ㄼж���֯�����~�ɼ      o�n�zmj���]���J�[�1�64�9������	x��W�`�y��'
9⨂:0��:��;2�#;5�2;�<;GpB;��E;��G;�eH;��H;�H;��H;��H;��H;��H;�H;'�H;�H;��H;��H;��H;��H;��H;��H;��H;��H;��H;��H;��H;�H;*�H;�H;��H;��H;��H;��H;�H;��H;�eH;��G;�E;JpB;߆<;7�2;2�#;��;2��:ܨ�:�'
9\�y��W��	x����<��64�\�1���J���]�xmj�      \���7���#���ѻ&���ǐ�dX�26�d	���uK��>":�M�:b�:Di;�%;D�3;ۆ<;&0B;��E;O\G;�HH;�H;s�H;;�H;��H;�H;�H;��H;��H;��H;��H;��H;��H;B�H;5�H;5�H;�H;4�H;4�H;C�H;��H;��H;��H; �H;��H;��H;�H;�H;��H;9�H;s�H; �H;�HH;U\G;��E;#0B;݆<;D�3;�%;Ei;"b�:�M�:�>":�uK�V	��26�hX�ǐ�"����ѻ ��8���      4Q^�!X��F�Ԣ)�++��ζ�`�<�@BS�n:��:���:��;2�;�M*;Ο5;pc=;GpB;��E;�JG;)8H;F�H;a�H;��H;�H;`�H;��H;p�H;��H;��H;��H;s�H;Z�H;5�H;��H;��H;��H;��H;��H;��H;��H;4�H;W�H;v�H;��H;��H;��H;n�H;��H;d�H;�H;��H;d�H;J�H;-8H;�JG;��E;KpB;mc=;Ο5;�M*;5�;��;���:��:n:@BS�l�<�϶�(+�ޢ)��F�!X�      ..�\�����K��
9]:�k:9M�:���:�y;��;t $;��/;d�8;|�>;�#C;�E;Y\G;,8H;��H;��H;��H;i�H;�H;c�H;0�H;��H;��H;��H;b�H;�H;��H;��H;��H;|�H;u�H;\�H;o�H;y�H;��H;��H;��H;�H;`�H;��H;��H;��H;,�H;h�H;�H;f�H;��H;��H;��H;/8H;U\G;�E;�#C;}�>;d�8;��/;x $;��;�y;���:GM�:�k:,]:�
9�K��김��      ���:�ņ:�ɒ:���:��:��:��:F�	;�v;��#;��-;��5;vL<;^�@;~(D;DF;��G;�HH;G�H;��H;��H;$�H;��H;:�H;��H;k�H;��H;��H;?�H;�H;��H;��H;S�H;G�H;�H;�H;�H;�H;�H;G�H;P�H;��H;��H;�H;<�H;��H;��H;i�H;��H;9�H;��H;'�H;��H;��H;J�H;�HH;��G;DF;�(D;]�@;wL<;��5;��-;��#;�v;D�	;$��:ؤ�:��:���:�ɒ:�ņ:      eW;ox;��;�
;��;};�� ;j�(;��/;�H6;��;;��?;�C;�PE;��F;��G;�eH;#�H;d�H;��H;*�H;��H;�H;��H;>�H;a�H;i�H;I�H;��H;��H;��H;-�H;��H;��H;��H;��H;��H;��H;��H;��H;��H;(�H;��H;��H;��H;I�H;d�H;b�H;A�H;��H;�H;��H;+�H;��H;e�H;!�H;�eH;��G;��F;�PE;�C;��?;��;;�H6;��/;p�(;�� ;v;��;
�
;��;dx;      rS%;�%;��';�M*;ӷ-;��1;ڟ5;��9;h-=;R@;��B;^�D;mF;�uG;T!H;�H;��H;w�H;��H;g�H;��H;�H;��H;E�H;^�H;V�H;�H;��H;��H;y�H;�H;��H;��H;�H;m�H;X�H;9�H;R�H;k�H;��H;��H;��H;
�H;x�H;��H;��H;�H;W�H;a�H;C�H;��H;�H;��H;g�H;��H;s�H;��H;�H;U!H;�uG;mF;b�D;��B;R@;j-=;��9;؟5;z�1;�-;�M*;��';��%;      ^o8;4�8;��9;f�:;u�<;�c>;+R@;�/B;��C;�PE;fzF;:\G;i�G;iH;�H;��H;�H;?�H;�H;�H;9�H;��H;A�H;P�H;H�H;'�H;��H;��H;R�H;��H;��H;��H;D�H;�H;�H;�H;��H;�H;�H;�H;C�H;��H;��H;��H;N�H;��H;��H;*�H;J�H;M�H;>�H;��H;:�H;�H;�H;9�H;�H;��H;�H;iH;i�G;=\G;mzF;�PE;��C;�/B;+R@;�c>;��<;e�:;��9;*�8;      ��A;?B;�oB;�C;P�C;P�D;=uE;GDF;�F;i�G;�H;�eH;ݡH;��H;-�H;��H;��H;��H;k�H;n�H;�H;B�H;a�H;P�H;�H;��H;��H;W�H;��H;��H;_�H;0�H;��H;��H;��H;��H;��H;��H;��H;��H;��H;+�H;b�H;��H;��H;V�H;��H;��H;�H;M�H;a�H;C�H;�H;j�H;k�H;��H;��H;��H;.�H;��H;ߡH;�eH;�H;k�G;�F;HDF;=uE;F�D;a�C;�C;�oB;?B;      DF;)RF;�zF;¸F;�G;\G;ѲG;)H;�HH;]�H;]�H;��H;��H;��H;��H;�H;��H;�H;��H;,�H;l�H;^�H;S�H;-�H;��H;r�H;G�H;��H;��H;R�H;�H;��H;��H;��H;e�H;T�H;a�H;N�H;b�H;��H;��H;��H;�H;Q�H;��H;��H;B�H;v�H;��H;,�H;S�H;`�H;l�H;*�H;��H;�H;��H;�H;��H;��H;��H;��H;e�H;_�H;�HH;)H;ҲG;u\G;�G;͸F;�zF;'RF;      �H;�H;�!H;�8H;�TH;*sH;�H;��H;{�H;��H;W�H;��H;��H;��H;��H;��H;��H;�H;r�H;��H;��H;e�H;�H;��H;��H;D�H;��H;w�H;:�H;�H;��H;��H;T�H;6�H; �H;��H;�H;��H;�H;8�H;T�H;��H;��H;�H;6�H;t�H;��H;I�H;��H;��H;�H;g�H;��H;��H;p�H;�H;��H;��H;��H;��H;��H;��H;X�H;��H;x�H;��H;�H;%sH;�TH;�8H;�!H;�H;      ~�H;�H;m�H;1�H;�H;x�H;)�H;\�H;�H;�H;��H;��H;��H;��H;��H;4�H;��H;��H;��H;��H;��H;C�H;��H;��H;P�H;��H;t�H;H�H;��H;��H;f�H;<�H;�H;��H;��H;��H;��H;��H;��H;��H;�H;8�H;f�H;��H;��H;F�H;p�H;��H;S�H;��H;��H;E�H;��H;��H;��H;��H;��H;7�H;��H;��H;��H;��H;�H;�H;�H;]�H;*�H;l�H;$�H;2�H;m�H;��H;      ��H;�H;��H;X�H;��H;3�H;��H;��H;��H;��H;��H;��H;�H;��H;��H;�H;�H;��H;��H;��H;E�H;��H;��H;O�H;��H;��H;3�H;��H;��H;_�H;(�H;��H;��H;��H;��H;��H;u�H;��H;��H;��H;��H;��H;*�H;^�H;��H;��H;/�H;��H;��H;L�H;��H;��H;C�H;��H;��H;��H;�H;�H;��H;��H;�H;��H;��H;��H;��H;��H;��H;,�H;��H;[�H;��H;�H;      ��H;��H;�H;N�H;��H;?�H;��H;��H;�H;��H;��H;�H;4�H;[�H;J�H;D�H;+�H;��H;��H;b�H;�H;��H;r�H;��H;��H;G�H;�H;��H;_�H;!�H;��H;��H;��H;~�H;^�H;C�H;5�H;A�H;Z�H;~�H;��H;��H;��H;�H;^�H;��H;��H;M�H;��H;��H;v�H;��H;�H;`�H;��H;��H;.�H;I�H;J�H;X�H;5�H;�H;��H;��H;�H;��H;��H;?�H;��H;T�H;�H;��H;      #�H;Z�H;v�H;��H;��H;��H;!�H;P�H;~�H;��H;��H;��H;��H;��H;��H;s�H;�H;��H;w�H;"�H;��H;��H;�H;��H;]�H;�H;��H;j�H;.�H;��H;��H;|�H;n�H;7�H;�H;�H;�H;�H;�H;8�H;p�H;z�H;��H;��H;*�H;h�H;��H;�H;`�H;��H;�H;��H;��H;�H;w�H;��H; �H;v�H;��H;��H;��H;��H;��H;��H;��H;P�H;+�H;��H;��H;��H;v�H;X�H;      �H;�H;�H;�H;!�H;A�H;D�H;c�H;i�H;Q�H;J�H;5�H;�H;��H;��H;F�H;��H;��H;]�H;��H;��H;,�H;��H;��H;.�H;��H;�H;=�H;��H;��H;u�H;Z�H;8�H;�H;��H;��H;��H;��H;��H;�H;<�H;X�H;s�H;��H;��H;<�H;�H;��H;/�H;��H;��H;/�H;��H;��H;]�H;��H;��H;I�H;��H;��H;�H;5�H;Q�H;U�H;j�H;f�H;M�H;C�H;/�H;�H;�H;�H;      ,�H;!�H;%�H;�H;�H; �H;�H;��H;��H;��H;��H;U�H;�H;��H;j�H;�H;��H;��H;:�H;��H;]�H; �H;��H;D�H;��H;��H;T�H;�H;��H;��H;k�H;;�H;��H;��H;��H;��H;��H;��H;��H;��H;��H;<�H;i�H;��H;��H;�H;T�H;��H;��H;C�H;��H;��H;Y�H;��H;:�H;��H;��H;�H;l�H;��H;�H;V�H;��H;��H;��H;��H;�H;��H;�H;�H;-�H;�H;      v�H;r�H;}�H;t�H;`�H;:�H;A�H;�H;��H;��H;��H;@�H;�H;��H;s�H;6�H;��H;E�H;��H;��H;N�H;��H;|�H;�H;��H;�H;2�H;��H;��H;��H;1�H;�H;��H;��H;��H;��H;��H;��H;��H;��H;��H;�H;1�H;|�H;��H;��H;4�H;��H;��H;�H;��H;��H;I�H;��H;��H;H�H;��H;6�H;t�H;��H;�H;@�H;��H;��H;��H;�H;G�H;9�H;h�H;v�H;��H;|�H;      ��H;��H;��H;��H;��H;]�H;R�H;�H;��H;��H;z�H;=�H;��H;��H;P�H;��H;��H;5�H;��H;��H;�H;��H;i�H;�H;��H;[�H;�H;��H;��H;a�H;�H;��H;��H;��H;��H;��H;��H;��H;��H;��H;��H;��H;�H;Z�H;��H;��H;�H;^�H;��H;�H;n�H;��H;�H;y�H;��H;8�H;��H;��H;P�H;��H;�H;=�H;|�H;��H;��H;!�H;W�H;`�H;��H;��H;��H;��H;      ��H;��H;��H;��H;d�H;R�H;=�H;�H;��H;��H;��H;H�H;��H;��H;4�H;��H;��H;3�H;��H;t�H;�H;��H;O�H;��H;��H;G�H;��H;��H;��H;H�H;�H;��H;��H;��H;��H;��H;��H;��H;��H;��H;��H;��H;�H;B�H;��H;��H;��H;J�H;��H;�H;V�H;��H;�H;o�H;��H;7�H;��H;��H;4�H;��H;��H;G�H;��H;��H;��H;�H;G�H;U�H;h�H;��H;��H;��H;      �H;��H;�H;��H;��H;��H;o�H;:�H;�H;��H;c�H;!�H;��H;��H;W�H;��H;��H;�H;��H;c�H;�H;��H;9�H;��H;��H;Z�H;	�H;��H;z�H;>�H;�H;��H;��H;��H;��H;��H;x�H;��H;��H;��H;��H;��H;�H;8�H;u�H;��H;�H;\�H;��H;��H;=�H;��H;�H;^�H;��H;�H;��H;��H;U�H;��H;��H; �H;f�H;��H;�H;;�H;x�H;��H;��H;��H;�H;�H;      ��H;��H;��H;��H;e�H;U�H;;�H;�H;��H;��H;��H;H�H;��H;��H;4�H;��H;��H;3�H;��H;t�H;�H;��H;N�H;��H;��H;G�H;��H;��H;��H;F�H;�H;��H;��H;��H;��H;��H;��H;��H;��H;��H;��H;��H;�H;A�H;��H;��H;��H;L�H;��H;��H;U�H;��H;�H;o�H;��H;7�H;��H;��H;4�H;��H;��H;G�H;��H;��H;��H;�H;A�H;R�H;h�H;��H;��H;��H;      ��H;��H;��H;��H;��H;\�H;R�H;"�H;��H;��H;x�H;=�H;��H;��H;Q�H;��H;��H;7�H;��H;��H;�H;��H;g�H;�H;��H;[�H;�H;��H;��H;`�H;�H;��H;��H;��H;��H;��H;��H;��H;��H;��H;��H;��H;�H;Z�H;��H;��H;�H;_�H;��H;	�H;n�H;��H;�H;y�H;��H;8�H;��H;��H;M�H;��H;��H;?�H;z�H;��H;��H;&�H;Y�H;\�H;��H;��H;��H;��H;      y�H;r�H;|�H;y�H;c�H;>�H;@�H;�H;��H;��H;��H;?�H;�H;��H;t�H;6�H;��H;H�H;��H;��H;N�H;��H;{�H;�H;��H;�H;4�H;��H;��H;��H;1�H;�H;��H;��H;��H;��H;��H;��H;��H;��H;��H;�H;0�H;}�H;��H;��H;4�H;��H;��H;�H;��H;��H;G�H;��H;��H;F�H;��H;8�H;t�H;��H;��H;?�H;��H;��H;��H;�H;H�H;;�H;j�H;y�H;��H;t�H;      *�H;&�H;(�H;�H;�H;�H;�H;��H;��H;��H;��H;X�H;�H;��H;l�H;�H;��H;��H;;�H;��H;]�H; �H;��H;C�H;��H;��H;S�H;�H;��H;��H;i�H;:�H;��H;��H;��H;��H;��H;��H;��H;��H;��H;<�H;i�H;��H;��H;�H;T�H;��H;��H;A�H;��H;��H;V�H;��H;;�H;��H;��H;�H;j�H;��H;�H;T�H;��H;��H;��H;��H;
�H;��H;�H;�H;0�H;!�H;      �H;�H;	�H;�H; �H;K�H;J�H;b�H;g�H;R�H;N�H;6�H;�H;��H;��H;I�H;��H;��H;]�H;��H;��H;/�H;��H;��H;/�H;��H;}�H;=�H;��H;��H;s�H;W�H;8�H;�H;��H;��H;��H;��H;��H;�H;;�H;X�H;r�H;��H;��H;;�H;~�H;��H;.�H;��H;��H;/�H;��H;��H;]�H;��H;��H;G�H;��H;��H;�H;6�H;O�H;R�H;g�H;b�H;M�H;@�H;"�H;�H;�H;�H;      �H;X�H;s�H;��H;��H;��H;#�H;Q�H;~�H;��H;��H;��H;��H;��H;��H;v�H; �H;��H;v�H;�H;��H;��H;�H;��H;`�H;�H;��H;h�H;/�H;��H;��H;|�H;n�H;8�H;�H;�H;�H;�H;�H;:�H;p�H;}�H;��H;��H;(�H;h�H;��H;�H;\�H;��H;�H;��H;��H;�H;y�H;��H;!�H;t�H;��H;��H;��H;��H;��H;��H;~�H;S�H;'�H;��H;��H;��H;y�H;W�H;      ��H;��H;�H;[�H;��H;J�H;��H;��H;�H;��H;��H;�H;4�H;Z�H;M�H;F�H;-�H;��H;��H;a�H;�H;��H;o�H;��H;��H;F�H;��H;��H;_�H;#�H;��H;��H;��H;~�H;^�H;B�H;5�H;C�H;[�H;~�H;��H;��H;��H; �H;\�H;��H;�H;K�H;��H;��H;y�H;��H;�H;`�H;��H;��H;-�H;G�H;L�H;Z�H;2�H; �H;��H;��H;�H;��H;��H;<�H;��H;a�H;�H;��H;      ��H;�H;�H;U�H;��H;7�H;��H;��H;��H;��H;��H;��H;�H;��H;��H;�H;�H;��H;��H;��H;E�H;��H;��H;O�H;��H;~�H;/�H;��H;��H;^�H;(�H;��H;��H;��H;��H;��H;u�H;��H;��H;��H;��H;��H;*�H;_�H;��H;��H;3�H;��H;��H;H�H;��H;��H;B�H;��H;��H;��H;�H;�H;��H;��H;�H;��H;��H;��H;��H;��H;��H;0�H;��H;T�H;�H;�H;      ��H;��H;`�H;2�H;�H;��H;*�H;c�H;��H;�H;��H;��H;��H;��H;��H;5�H;��H;��H;��H;��H;��H;E�H;��H;��H;S�H;��H;p�H;F�H;��H;��H;f�H;<�H;�H;��H;��H;��H;��H;��H;��H;��H;�H;<�H;h�H;��H;��H;F�H;t�H;��H;O�H;��H;��H;F�H;~�H;��H;��H;��H;��H;7�H;��H;��H;��H;��H;�H;�H;��H;]�H;)�H;q�H;!�H;2�H;j�H;��H;      �H;H;�!H;�8H;�TH;.sH;�H;��H;{�H;��H;W�H;��H;��H;��H;��H;��H;��H;�H;o�H;��H;��H;g�H;�H;��H;��H;A�H;��H;u�H;9�H;�H;��H;��H;S�H;6�H;!�H;��H;�H;��H;�H;8�H;T�H;��H;��H;�H;6�H;u�H;��H;H�H;��H;��H;�H;h�H;��H;��H;p�H;�H;��H;��H;��H;��H;��H;��H;U�H;��H;x�H;��H;!�H;)sH;�TH;�8H;�!H;�H;      �CF;%RF;�zF;��F;�G;�\G;ͲG;,H;�HH;\�H;c�H;��H;��H;��H;��H;�H;��H;�H;��H;'�H;l�H;]�H;O�H;,�H;��H;n�H;B�H;��H;��H;Q�H;�H;��H;��H;��H;f�H;P�H;c�H;S�H;b�H;��H;��H;��H;	�H;R�H;��H;��H;H�H;t�H;��H;*�H;V�H;^�H;k�H;*�H;��H;�H;��H;�H;��H;��H;��H;��H;a�H;]�H;�HH;#H;ͲG;u\G;�G;��F;rzF;RF;      ��A;;B;�oB;�C;R�C;R�D;<uE;GDF;�F;i�G;�H;�eH;ۡH;��H;0�H;��H;��H;��H;i�H;h�H; �H;B�H;]�H;O�H;�H;��H;��H;V�H;��H;��H;_�H;0�H;��H;��H;��H;��H;��H;��H;��H;��H;��H;2�H;d�H;��H;��H;U�H;��H;��H;�H;M�H;d�H;C�H;�H;k�H;m�H;��H;��H;��H;0�H;��H;ޡH;�eH;�H;k�G;�F;HDF;;uE;E�D;Z�C;�C;�oB;;B;      9o8;�8;��9;q�:;p�<;�c>;.R@;�/B;��C;�PE;izF;=\G;h�G;iH;�H;��H;�H;>�H;�H;	�H;9�H;��H;;�H;O�H;I�H;"�H;��H;��H;P�H;��H;��H;��H;D�H;�H;�H;�H;��H;�H;�H;�H;H�H;��H;��H;��H;P�H;��H;��H;)�H;H�H;O�H;A�H;��H;:�H;�H;�H;9�H;�H;��H;�H;iH;f�G;:\G;hzF;�PE;��C;�/B;-R@;�c>;��<;��:;��9;�8;      ZS%;��%;�';�M*;ͷ-;v�1;ԟ5;��9;o-=;R@;��B;b�D; mF;�uG;U!H;�H;��H;w�H;��H;e�H;��H;
�H;��H;C�H;`�H;O�H;�H;��H;��H;t�H;	�H;��H;��H;�H;n�H;X�H;<�H;X�H;m�H;�H;��H;��H;�H;{�H;��H;��H;�H;V�H;^�H;B�H;��H;�H;��H;g�H;��H;s�H;��H;�H;W!H;�uG;mF;\�D;��B;R@;k-=;��9;ԟ5;x�1;з-;�M*;�';��%;      `W;ox;��;�
;��;�;�� ;p�(;��/;�H6;��;;��?;�C;�PE;��F;��G;�eH;!�H;a�H;��H;(�H;��H;�H;��H;A�H;Z�H;g�H;I�H;��H;��H;��H;-�H;��H;��H;��H;��H;��H;��H;��H;��H;��H;/�H;��H;��H;��H;I�H;k�H;b�H;>�H;��H;�H;��H;*�H;��H;d�H; �H;�eH;��G;��F;�PE;�C;��?;��;;�H6;��/;p�(;�� ;h;��;��
;��;ex;      ���:�ņ:�ɒ:��:��:��:$��:F�	;�v;�#;��-;��5;vL<;\�@;�(D;DF;��G;�HH;F�H;��H;��H;%�H;��H;9�H;��H;d�H;��H;~�H;>�H;��H;��H;��H;R�H;H�H;�H;�H;�H;�H;�H;G�H;U�H;��H;��H;�H;>�H;��H;��H;i�H;��H;:�H;��H;$�H;��H;��H;I�H;�HH;��G;DF;�(D;]�@;wL<;��5;��-;��#;�v;H�	;(��:��:��:��:�ɒ:�ņ:      �-.�L�� ���~K�p
9,]:�k:QM�:���:�y;��;x $;��/;b�8;}�>;�#C;�E;V\G;*8H;��H;��H;��H;f�H;�H;g�H;)�H;��H;��H;��H;[�H;�H;��H;��H;��H;}�H;r�H;^�H;t�H;{�H;��H;��H;��H;�H;a�H;��H;��H;��H;,�H;d�H;�H;j�H;��H;��H;��H;-8H;U\G;�E;�#C;|�>;b�8;��/;v $;��;�y;���:CM�:�k:]:�
9�K����X��      3Q^� X��F�Ѣ)�/+��ζ�p�<�@BS�n:��:���:��;2�;�M*;П5;pc=;GpB;��E;�JG;*8H;J�H;c�H;��H;�H;c�H;��H;l�H;��H;��H;��H;s�H;X�H;4�H;��H;��H;��H;��H;��H;��H;��H;5�H;Z�H;v�H;��H;��H;��H;p�H;��H;`�H;�H;��H;a�H;I�H;-8H;�JG;��E;HpB;nc=;Ο5;�M*;2�;��;���:��:n:�AS�t�<�϶�-+�Ӣ)��F�X�      c���2���&���ѻ$���ǐ�bX�+6�Z	���uK��>":�M�:b�:Bi;�%;E�3;܆<;#0B;��E;R\G;�HH; �H;t�H;9�H;��H;�H;�H;��H;��H;��H;��H;��H;��H;C�H;5�H;4�H;�H;7�H;3�H;C�H;��H;��H;��H;��H;��H;��H;�H;�H;��H;9�H;v�H;�H;�HH;U\G;��E;#0B;܆<;D�3;�%;Di;b�:�M�:�>": vK�Z	��06�eX�ǐ�$����ѻ*��4���      o�n�zmj���]���J�Z�1�64�:������	x��W�h�y��'
9ܨ�:.��:��;3�#;7�2;߆<;FpB; �E;��G;�eH;��H;�H;��H;��H;��H;��H;�H;$�H;�H;��H;��H;��H;��H;��H;��H;��H;��H;��H;��H;��H;�H;(�H;�H;��H;��H;��H;��H;�H;��H;�eH;��G;�E;GpB;݆<;7�2;2�#;��;0��:ਂ:�'
9`�y��W��	x����<��64�]�1���J���]�ymj�      @<ͼ��ɼ�����֯�϶��ㄼ��Y��*�����s��#X��rѺ0��>Q:���:��
;,�#;E�3;mc=;�#C;DF;��G;�H;��H;��H;�H;��H;0�H;��H;B�H;o�H;C�H;�H;5�H;��H;��H;��H;��H;��H;1�H;�H;C�H;o�H;D�H;��H;4�H;��H;�H;��H;��H;�H;��G;�CF;�#C;mc=;D�3;.�#;��
;���:�>Q:0��rѺ#X��s������*���Y�ㄼж���֯�������ɼ      ��'�(�$����|��  ���ۼ����+����]��X!�H>ۻ�+���*������>:���:��;�%;ʟ5;w�>;�(D;��F;W!H;
�H;&�H;��H;��H;��H;��H;I�H;��H;��H;i�H;p�H;I�H;1�H;N�H;2�H;G�H;p�H;h�H;��H;��H;J�H;��H;��H;��H;��H;&�H;�H;U!H;��F;{(D;z�>;ʟ5;�%;��;���:��>:��깈*��+��H>ۻ�X!���]��+�������ۼ�  �}����)�$�      Ÿ���v����w�g�c��J�΄-�|��;缆沼	ㄼ��;������j���5�����>Q:.��:Ei;�M*;b�8;e�@;�PE;�uG;iH;��H;��H;��H;��H;��H;T�H;��H;��H;��H;��H;��H;��H;�H;��H;��H;��H;��H;��H;��H;X�H;��H;��H;��H;��H;��H;iH;�uG;�PE;\�@;f�8;�M*;Ei;.��:�>Q:��깮5��j��������;�	ㄼ�沼�;�}�΄-��J�g�c���w��v��      yHͽתɽ�;��"����Ǹ����[�	z0�s��'<ͼ˾��e�J�����j���*� �ڨ�:$b�:2�;��/;}L<;�C;mF;l�G;ڡH;��H;��H;��H;�H;/�H;��H;�H;�H;��H;��H;��H;��H;��H;��H;��H;�H;�H;��H;4�H;�H;��H;��H;��H;סH;i�G;mF;�C;sL<;��/;/�;"b�:ܨ�: ��*��j�����f�J�̾��(<ͼs��	z0���[�Ǹ����"���;��תɽ      ��"-������ұ�ƽ^P���v���J�I����ۼ��f�J������+���rѺ�'
9�M�:��;r $;��5;��?;\�D;<\G;�eH;��H;��H;��H;��H;��H;��H;/�H;U�H;<�H;2�H;A�H;�H;D�H;0�H;:�H;Q�H;/�H;��H;��H;��H;��H;��H;��H;�eH;<\G;^�D;��?;��5;v $;��;�M�:�'
9�rѺ�+������f�J�����ۼI���J��v��^P��ƽұ轄����"-�       j�Vde�Z0X�D�g{+�������v㻽Z���RDX������ۼ̾����;�J>ۻ)X���y��>":���:��;��-;�;;��B;fzF;�H;[�H;S�H;��H;��H;��H;��H;K�H;��H;|�H;p�H;��H;[�H;��H;p�H;{�H;��H;H�H;��H;��H;��H;��H;Q�H;Y�H;�H;hzF;��B;{�;;��-;��;���:�>":��y�)X�K>ۻ��;�̾����ۼ���RDX�Y���v㻽��콂��g{+�D�Z0X�Vde�      ��Qh��k���I���|x���O��C(���Ϫɽ����RDX�I��(<ͼ
ㄼ�X!��s���W�`vK���:�y;��#;�H6;R@;�PE;e�G;X�H;��H;�H;��H;|�H;��H;Q�H;��H;��H;��H;��H;��H;��H;��H;��H;��H;O�H;��H;~�H;��H;�H;��H;V�H;a�G;�PE;R@;�H6;��#;�y;��:`vK��W��s���X!�
ㄼ(<ͼI��RDX�����Ϫɽ���C(���O��|x��I��k��Qh��      =����������"�;hɰ��G��
 j�8�5��	�ϪɽY����J�s���沼��]�����	x�j	��n:~��:�v;��/;`-=;��C;�F;�HH;w�H;��H;��H;��H;{�H;d�H;��H;��H;��H;��H;�H;��H;��H;��H;��H;f�H;x�H; �H;��H;��H;x�H;�HH;�F;��C;c-=;��/;�v;���:�m:h	���	x������]��沼t���J�Y���Ϫɽ�	�8�5�
 j��G��hɰ�"�;��徶���      �2�V�-�"�-E�����?Kɾj����s�8�5���v㻽�v��
z0��;��+���*����=6��CS�;M�:H�	;h�(;�9;�/B;DDF;H;��H;V�H;��H;�H;J�H;b�H;��H;�H;�H;�H;9�H;�H;�H;�H;��H;`�H;I�H;��H;��H;X�H;��H;H;ADF;�/B;�9;h�(;A�	;AM�:�DS�96�����*��+���;�
z0��v��v㻽��8�5���s�j��?Kɾ����-E�"�V�-�      %3s�cm�:�\�h�C�5�%����TҾj��
 j��C(����_P����[�}������Y�>��oX���<���k:$��:�� ;̟5;*R@;/uE;ʲG;�H;�H;��H;��H; �H;D�H;�H;@�H;I�H;4�H;k�H;3�H;K�H;>�H;�H;D�H;�H;��H;��H;�H;�H;ϲG;.uE;+R@;Ο5;�� ;��:��k:��<�mX�>����Y����}���[�_P����콪C(�
 j�j���TҾ��5�%�h�C�:�\�cm�      �ޞ�������_F�>�W�W�-���?Kɾ�G����O����ƽǸ��΄-���ۼㄼ74� ǐ�϶�]:��:u;t�1;�c>;>�D;q\G;'sH;s�H;1�H;D�H;��H;K�H;	�H;G�H;h�H;Z�H;��H;Z�H;g�H;E�H;	�H;K�H;��H;F�H;3�H;v�H;*sH;{\G;=�D;�c>;t�1;s;ޤ�:]:϶� ǐ�84�ㄼ��ۼ΄-�Ǹ��ƽ�����O��G��?Kɾ��W�-�>�W�_F�������      ��ſ���Lw���ޞ�����>�W�5�%�����hɰ��|x�g{+�ұ����J��  �϶��\�1�.���(+��
9��:��;׷-;�<;W�C;�G;�TH;�H;��H;��H;��H;)�H;�H;e�H;��H;r�H;��H;n�H;��H;a�H;�H;(�H;��H;��H;��H;#�H;�TH;�G;T�C;��<;շ-;��;��:�
9)+�,���]�1�϶���  ��J���ұ�g{+��|x�hɰ�����5�%�>�W������ޞ�Lw�����      ������Կp���ޞ�`F�h�C�-E�"�;�I��D���"��g�c�}��֯���J��ѻע)� �K���:�
;�M*;f�:;�C;��F;�8H;'�H;F�H;U�H;��H;�H;�H;}�H;��H;��H;��H;��H;��H;{�H;�H;�H;��H;\�H;G�H;(�H;�8H;̸F;�C;f�:;�M*;��
;��:�K�ڢ)��ѻ��J��֯�}�g�c�"����D��I��"�;-E�h�C�`F��ޞ�p���Կ��      ����������ԿLw�����:�\�"����k��Z0X�����;����w����������]�&���F����ɒ:��;��';��9;�oB;zzF;�!H;p�H;��H; �H;o�H;�H;�H;|�H;��H;��H;��H;��H;��H;|�H;�H;�H;i�H;�H;��H;q�H;�!H;�zF;�oB;��9;��';��;�ɒ:����F�$�黮�]����������w��;�����Z0X�k�����"�:�\����Lw���Կ��𿝏�      $�������忇�����cm�V�-�����Qh��Vde�"-�תɽ�v��(�$���ɼ}mj�>���X�<���ņ:`x;�%;,�8;AB;RF;�H;�H;�H;��H;B�H;�H;�H;u�H;��H;��H;�H;��H;��H;u�H;�H;�H;>�H;��H;�H;�H;�H;'RF;>B;*�8;��%;]x;�ņ:0��X�<���~mj���ɼ(�$��v��תɽ"-�Vde�Qh������V�-�cm��������忝����      dܿ3�ֿ�aǿ=^��/���Yo���7����iþ�(���-=��` �A���_�0]�0p����I�V�ѻ��)��R���:*�
;�*;�:;��B;�HF;#�G;�lH;�H;q�H;7�H;��H;|�H;I�H;y�H;�H;��H;�H;x�H;I�H;{�H;��H;6�H;{�H;�H;�lH;&�G;�HF;��B;�:;�*;&�
;��:��R���)�V�ѻ��I�0p��0]��_�A���` ��-=��(���iþ����7�Yo�/���=^���aǿ3�ֿ      2�ֿCpѿ�¿������_Xi�Е3��
�VD��Fl��@�9��.���R��!\� �fx��2�E��ͻ%�$�� �ˍ�:8�;E�*;1�:;�B;�TF;��G;#nH;��H;��H;g�H;��H;��H;X�H;|�H;�H;��H;�H;}�H;V�H;��H;��H;b�H;ķH;��H;#nH;��G;�TF;�B;+�:;>�*;5�;Ǎ�:� �%�$��ͻ2�E�fx�� �!\��R���.��@�9�Fl��VD���
�Е3�_Xi��������¿Cpѿ      �aǿ�¿����������"Y��f'�����7o���.}��k/����%ڟ�"<Q�.#�ע��(;�4���@�� q7���:�;l,;��;;�C;�vF;�G;�rH;�H;��H;�H;��H;��H;��H;��H;J�H;��H;B�H;��H;��H;��H;��H;�H;��H;�H;�rH;�G;�vF;�C;|�;;e,;�;��: j7�B��4����(;�ע�.#�"<Q�%ڟ�����k/��.}�7o�������f'��"Y�����������¿      =^������k���Yo���@�)�$�޾����9ce�0����ڽ󻒽g@������R���O*�NG��"����B^9��:�;Vd.;��<;��C;�F;��G;�yH;��H;�H;�H;��H;h�H;��H;��H;�H;�H;z�H;��H;��H;e�H;��H;�H;�H;��H;�yH;��G;��F;��C;��<;Md.;�;��:`C^9(���MG���O*��R������g@�󻒽��ڽ0��9ce�����$�޾)���@�Yo�k�������      /����������Yo��!J�K�#��\��VD������zPH�����b�� C��� +���ټ*����񿐻"���8�:��:=�;�Y1;>;�0D;x�F;]H;A�H;��H;�H;W�H;��H;	�H;_�H;H�H;��H;\�H;��H;F�H;_�H;�H;��H;Q�H;�H;��H;?�H;^H;|�F;�0D;�>;�Y1;=�;��:T�:&���񿐻��*����ټ� +� C���b�����zPH�����VD���\��K�#��!J�Yo��������      Yo�_Xi��"Y���@�K�#��
��о�A���i���(�~��wr���_��5��ɺ�r�`��<��n�d���\�,�X:�P�:�`;±4;��?;��D;q8G;i0H;��H;i�H;p�H;��H;��H;��H;��H;��H;�H;��H;�H;��H;��H;��H;��H;��H;u�H;g�H;��H;g0H;w8G;��D;��?;��4;�`;�P�:<�X:��\�m�d��<��s�`��ɺ��5��_�vr��~����(��i��A���о�
�K�#���@��"Y�_Xi�      ��7�Е3��f'�)��\���о�����.}��-=�{
���Ľ\��,:����������7�&GĻʃ$�@O�����:�{;D&;�+8;JA;�E;��G;yLH;�H;t�H;/�H;��H;��H;��H;��H;�H;��H;�H;|�H;�H;��H;��H;��H;��H;5�H;r�H;��H;tLH;��G;�E;JA;�+8;~D&;�{;���:HO��˃$�%GĻ�7���������,:�\����Ľ{
��-=��.}������о�\��)��f'�Е3�      ���
�����$�޾VD���A���.}�(�D�ht���ڽ�!��\����\�ļ�
v�>��ο���Iɺ�R�9���:(;�-;}�;;��B;bIF;��G;fH;��H;�H;)�H;��H;c�H;��H;Y�H;��H;��H;d�H;��H;��H;Z�H;��H;_�H;��H;0�H;�H;��H;fH;��G;cIF;��B;}�;;�-;(;���:�R�9�Iɺο��>���
v�\�ļ���\��!����ڽht�(�D��.}��A��VD��$�޾�����
�      �iþVD��7o�����������i��-=�ht� ���R��iys�z +����z񗼖(;�.�ѻ�s@��!��3j:�P�:��;�D3;,�>;FD;��F;�	H;5|H;��H;o�H;0�H;��H;��H;��H;�H;+�H;m�H;��H;j�H;,�H;�H;��H;��H;��H;6�H;o�H;��H;5|H;�	H;��F;FD;-�>;�D3;��;�P�:�3j:�!��s@�.�ѻ�(;�z����z +�iys��R�� ��ht��-=��i���������7o��VD��      �(��Fl���.}�9ce�zPH���(�|
���ڽ�R�� �{�C�6�� �.p��`�`�Ϩ��,��VIҺ�K^9���:ԣ;�~(;(�8;�IA;�{E;jG;�=H;>�H;ѬH;�H;Y�H;"�H;h�H;��H;��H;��H;��H;H�H;��H;��H;��H;��H;e�H;"�H;`�H;�H;ѬH;<�H;�=H;jG;�{E;�IA;)�8;�~(;٣;���:�K^9TIҺ�,��Ψ�`�`�.p��� �C�6� �{��R����ڽ{
���(�zPH�9ce��.}�Fl��      �-=�@�9��k/�0�����~��Ľ�!��iys�C�6�%#��ɺ��vz����D^��o�$��$�r:���:��;�Y1;�H=; xC;!wF;�G;�eH;E�H;~�H;��H;��H;L�H;��H;��H;��H;c�H;w�H;��H;y�H;d�H;��H;��H;��H;M�H;��H;��H;�H;F�H;�eH;�G;!wF;#xC;�H=;�Y1;��;���:$�r:�~�o�$�D^������vz��ɺ�%#�C�6�iys��!����Ľ~���0���k/�@�9�      �` ��.�����ڽ�b��wr��[��\�z +�� ��ɺ�A��O*�Jͻ�5R� ǅ���:��:~�;�);�t8;_�@;S*E;g8G;8$H;9�H;@�H;�H;�H;��H;h�H;`�H; �H;M�H;��H;��H;�H;��H;��H;O�H;��H;]�H;k�H;��H;&�H;�H;;�H;9�H;=$H;g8G;W*E;b�@;�t8;�);�;��:��: ǅ��5R�Iͻ�O*�@��ɺ�� �z +�\�[��vr���b����ڽ��.��      A���R��%ڟ�����C���_�+:�������-p���vz��O*��4ֻk�<�����09 �:1;J� ;�D3;B�=;��C;�kF;��G;�\H;��H;I�H;��H;6�H;��H;t�H;��H;��H;�H;��H;T�H;��H;S�H;��H;�H;��H;��H;w�H;��H;;�H;��H;H�H;��H;�\H;��G;�kF;��C;A�=;�D3;O� ;1;(�:��096���k��4ֻ�O*��vz�-p����輤��,:��_� C������%ڟ��R��      �_� \�!<Q�g@�� +��5�����[�ļz�_�`����Lͻk�Iɺ �6�0�:�P�:%�;�d.;@�:;�A;$|E;sNG;@'H;��H;åH;Z�H;��H;!�H;G�H;W�H;2�H;��H;��H;�H;��H;��H;��H;	�H;��H;��H;/�H;Z�H;Q�H;(�H;��H;X�H;��H;��H;@'H;xNG;'|E;�A;I�:;�d.;"�;�P�:0�: �6�
Iɺk�Jͻ���_�`�y�[�ļ�����5�� +�g@�!<Q� \�      /]� �.#�������ټ�ɺ������
v��(;�Ψ�B^���5R�>��� �6����:���:�;#�*;�+8;|!@;T�D;]�F;��G;�eH;{�H;��H;��H;��H;��H;��H;�H;r�H;��H;a�H;x�H;)�H;V�H;(�H;w�H;b�H;��H;n�H; �H;��H;��H;��H;��H;��H;~�H;�eH;��G;`�F;U�D;�!@;�+8;�*;��;���:���: �6�:����5R�@^��Ψ��(;��
v������ɺ���ټ����.#� �      -p��ex��ע��R��)��r�`� �7�<��.�ѻ�,��k�$� ǅ���090�:���:z;�~(;�Z6;~�>;ŨC;�HF;נG;�DH;D�H;��H;��H;�H;&�H;�H;��H;��H;��H;��H;�H;��H;��H;��H;�H;��H;�H;��H;��H;��H;��H;�H;)�H;�H;��H;��H;D�H;�DH;٠G;�HF;̨C;�>;�Z6;�~(;|;���:0�:��09ǅ�h�$��,��+�ѻ<���7�p�`�*���R��ע�dx��      ��I�0�E��(;��O*����<��!GĻʿ���s@�DIҺ�~�:*�:�P�:�;�~(;�5;�>;3C;*�E;tcG;6$H;�{H;4�H;�H;��H;��H;9�H;��H;�H;T�H;��H;M�H;��H;?�H;��H;��H;��H;<�H;��H;J�H;��H;W�H;�H;��H;9�H;��H;��H;�H;5�H;�{H;8$H;wcG;2�E;3C;�>;�5;�~(;��;�P�:*�:��:�~�BIҺ�s@�ȿ��#GĻ�<�����O*��(;�.�E�      I�ѻ�ͻ2���HG��쿐�k�d���$��Iɺ�!� L^90�r:��:�0;!�;�*;�Z6;�>;8�B;��E;�8G;�	H;�mH;�H;C�H;��H;`�H;��H;��H;E�H;��H;�H;u�H;��H;��H;��H;�H;!�H;�H;��H;��H;��H;q�H;��H;�H;E�H;��H;��H;]�H;��H;E�H;�H;�mH;�	H;�8G;��E;2�B;�>;�Z6;�*;!�; 1;��:H�r:@L^9؅!��IɺŃ$�f�d�运�JG��.����ͻ      t�)�2�$�A�����*���H�\��N���R�9 4j:���:��:x�;M� ;�d.;�+8;|�>;3C;��E;�)G;��G;dH;{�H;��H;Y�H;��H;0�H;��H;��H;��H;��H;��H;H�H;z�H;_�H;��H;6�H;I�H;3�H;��H;]�H;w�H;C�H;��H;��H;��H;��H;��H;0�H;��H;\�H;��H;~�H;dH;��G;�)G;��E;4C;{�>;�+8;�d.;O� ;~�;��:���:4j:�R�9O��\�\�&���0���@��2�$�      ��R� � c7�PD^9@�:D�X:Ϳ�:���:�P�:ۣ;��;�);�D3;E�:;�!@;ɨC;1�E;�8G;��G;�`H;j�H;�H;�H;u�H;5�H;-�H;I�H;[�H;��H;��H;��H;�H;��H;��H;,�H;m�H;c�H;g�H;*�H;��H;��H;�H;��H;��H;��H;]�H;H�H;-�H;;�H;v�H;�H;�H;o�H;�`H;��G;�8G;.�E;˨C;�!@;C�:;�D3;�);��;ܣ;�P�:���:ÿ�:`�X:T�:PC^9 k7�� �      ��:���:��:��:���:�P�:�{;(;��;�~(;�Y1;�t8;=�=;�A;T�D;�HF;tcG;�	H;dH;h�H;B�H;ѶH;.�H;��H;��H;7�H;E�H;��H; �H;��H;|�H;��H;R�H;��H;E�H;��H;��H;��H;G�H;��H;Q�H;��H;}�H;��H;�H;��H;A�H;6�H;��H;��H;+�H;ӶH;G�H;j�H;dH;�	H;tcG;�HF;T�D;�A;?�=;�t8;�Y1;�~(;��;(;�{;�P�:��:
��:��:���:      &�
;C�;��;;<�;�`;|D&;�-;�D3;/�8;I=;_�@;��C;)|E;`�F;٠G;8$H; nH;�H;�H;ӶH;��H;3�H;�H;d�H;��H;��H;r�H;f�H;�H;�H;��H;��H;�H;d�H;��H;��H;��H;`�H;�H;��H;��H;�H;�H;d�H;p�H;��H;��H;g�H;�H;0�H;��H;ֶH;�H;�H;�mH;;$H;٠G;c�F;$|E;��C;c�@;I=;+�8;�D3;�-;�D&;�`;R�;;�;6�;      �*;D�*;e,;dd.;�Y1;α4;�+8;��;;7�>;�IA;-xC;Z*E;�kF;�NG;��G;�DH;�{H;�H;��H;�H;,�H;2�H;��H;��H;��H;[�H;�H;��H;��H;��H;��H;m�H;��H;9�H;��H;��H;��H;��H;��H;:�H;��H;g�H;��H;��H;��H;��H;�H;\�H;��H;��H;��H;5�H;/�H;�H;��H;�H;�{H;�DH;��G;}NG;�kF;^*E;1xC;�IA;7�>;��;;�+8;ȱ4;�Y1;bd.;e,;-�*;      �:;5�:;y�;;��<;�>;��?;JA;��B;FD;|E;!wF;g8G;��G;B'H;�eH;H�H;7�H;I�H;\�H;r�H;��H;�H;��H;��H;�H;��H;��H;2�H;u�H;m�H;�H;��H;�H;\�H;}�H;��H;��H;��H;y�H;\�H;�H;��H;�H;l�H;o�H;2�H;��H;��H;�H;��H;��H;�H;��H;q�H;Y�H;C�H;7�H;H�H;�eH;?'H;��G;j8G;(wF;|E;FD;��B;JA;��?;>;��<;|�;;*�:;      ̣B;�B;�C;��C;�0D;��D;��E;fIF;��F;jG; �G;A$H;�\H;�H;��H;��H;!�H;��H;��H;A�H;��H;g�H;��H;�H;��H;o�H;��H;B�H;(�H;��H;��H;��H;*�H;q�H;��H;��H;��H;��H;��H;q�H;)�H;��H;��H;��H;$�H;A�H;��H;p�H;��H;�H;��H;j�H;��H;<�H;��H;��H;$�H;��H;��H;�H;�\H;F$H;!�G;jG;��F;fIF;��E;��D;�0D;��C;�C;�B;      �HF;�TF;�vF;�F;q�F;|8G;��G;��G;�	H;�=H;�eH;?�H;��H;ʥH;��H;��H;��H;`�H;0�H;,�H;:�H;��H;X�H;��H;j�H;��H; �H;�H;��H;C�H;��H;�H;3�H;n�H;��H;��H;��H;��H;��H;n�H;2�H;�H;��H;@�H;��H;�H;�H;��H;o�H;��H;W�H;��H;:�H;*�H;0�H;^�H;��H;��H;��H;ĥH;��H;@�H;fH;�=H;�	H;��G;��G;q8G;��F;�F;�vF;�TF;      5�G;��G;�G;��G;VH;j0H;�LH;fH;4|H;?�H;F�H;;�H;G�H;Z�H;��H;�H;��H;��H;��H;I�H;I�H;��H;�H;��H;��H;�H;��H;��H;N�H;��H;��H;/�H;L�H;q�H;��H;��H;��H;�H;��H;t�H;O�H;,�H;��H;��H;J�H;��H;��H;#�H;��H;��H;�H;��H;K�H;F�H;��H;��H;��H;�H;��H;W�H;H�H;@�H;I�H;>�H;4|H;fH;}LH;c0H;kH;��G;�G;��G;      �lH;&nH;�rH;�yH;7�H;��H;�H;��H;��H;جH;��H;��H;��H;��H;��H;(�H;7�H;��H;��H;X�H;��H;l�H;��H;2�H;;�H;�H;��H;3�H;��H;��H;�H;;�H;^�H;d�H;|�H;��H;�H;��H;{�H;d�H;]�H;4�H;�H;��H;��H;/�H;��H;�H;?�H;/�H;��H;n�H;��H;W�H;��H;��H;9�H;)�H;��H;��H;��H;��H;��H;٬H;��H;��H;�H;��H;B�H;�yH;�rH;nH;      �H;��H;�H;��H;��H;i�H;{�H;�H;h�H;�H;��H;#�H;:�H;%�H;��H;�H;��H;I�H;��H;��H;&�H;c�H;��H;r�H;#�H;��H;F�H;��H;��H;�H;)�H;K�H;]�H;c�H;a�H;m�H;j�H;g�H;`�H;d�H;^�H;E�H;)�H;	�H;��H;��H;C�H;��H;$�H;n�H;��H;b�H;#�H;��H;��H;G�H;��H;�H;��H;%�H;9�H;"�H;��H;�H;l�H;�H;y�H;b�H;��H;��H;�H;��H;      u�H;��H;��H;�H;
�H;m�H;1�H;*�H;3�H;]�H;��H;��H;��H;O�H;��H;��H;�H;��H;��H;��H;��H; �H;��H;j�H;��H;9�H;��H;��H;�H;!�H;>�H;B�H;L�H;a�H;K�H;Y�H;n�H;V�H;G�H;a�H;N�H;=�H;=�H;�H;	�H;��H;��H;?�H;��H;h�H;��H; �H;��H;��H;��H;��H; �H;��H;��H;M�H;��H;��H;��H;c�H;6�H;,�H;4�H;m�H;�H;�H;��H;��H;      =�H;|�H;�H;�H;S�H;��H;��H;��H;��H;(�H;Q�H;t�H;{�H;^�H;#�H;��H;]�H;��H;��H;��H;��H;�H;��H;�H;��H;��H;��H;
�H;-�H;D�H;U�H;N�H;=�H;=�H;^�H;L�H;,�H;H�H;Z�H;>�H;>�H;K�H;S�H;@�H;)�H;�H;��H;��H;��H;�H;��H;�H;~�H;��H;��H;��H;^�H;��H;#�H;]�H;~�H;u�H;T�H;*�H;��H;��H;��H;��H;a�H; �H;�H;|�H;      ��H;��H;��H;��H;��H;��H;��H;d�H;��H;f�H;��H;b�H;��H;9�H;r�H;��H;��H;v�H;L�H;�H;��H;��H;i�H;��H;��H;�H;*�H;;�H;I�H;D�H;H�H;U�H;:�H;6�H;H�H;)�H;"�H;)�H;E�H;7�H;>�H;S�H;E�H;B�H;E�H;6�H;)�H;�H;��H;��H;p�H;��H;��H;�H;I�H;x�H;��H;��H;r�H;6�H;��H;d�H;��H;j�H;��H;f�H;�H;��H;��H;��H;��H;��H;      ��H;��H;��H;g�H;�H;��H;��H;��H;��H;��H;��H;�H;��H;��H;��H;��H;S�H; �H;~�H;��H;\�H;��H;��H;�H;*�H;/�H;N�H;e�H;d�H;S�H;:�H;>�H;A�H;;�H;�H;�H;I�H;�H;�H;=�H;B�H;>�H;9�H;N�H;^�H;`�H;L�H;0�H;-�H;�H;��H;��H;Y�H;��H;}�H; �H;T�H;��H;��H;��H; �H;�H;��H;��H;��H;��H;��H;��H;�H;d�H;
�H;��H;      B�H;T�H;��H;��H;a�H;��H;��H;Y�H;�H;��H;��H;T�H;�H;��H;h�H;�H;��H;��H;b�H;��H;��H;�H;4�H;U�H;n�H;k�H;o�H;e�H;d�H;e�H;9�H;:�H;;�H;&�H;�H;�H;#�H;�H;�H;&�H;>�H;9�H;9�H;a�H;a�H;a�H;o�H;k�H;q�H;S�H;=�H;�H;��H;��H;`�H;�H;��H;�H;h�H;��H;�H;T�H;��H;��H;�H;Z�H;��H;��H;i�H;��H;��H;`�H;      u�H;��H;��H;��H;T�H;��H;�H;��H;.�H;��H;j�H;��H;��H;�H;��H;��H;D�H;��H;��H;0�H;K�H;`�H;��H;o�H;��H;��H;��H;}�H;d�H;O�H;W�H;L�H;�H;�H;!�H;�H;��H;�H;�H;�H;�H;N�H;V�H;H�H;`�H;y�H;��H;��H;��H;q�H;��H;`�H;G�H;*�H;��H;��H;H�H;��H;��H;�H;��H;��H;o�H;��H;3�H;��H;&�H;��H;T�H;��H;��H;��H;      �H;�H;G�H;{�H;��H;�H;��H;��H;g�H;��H;z�H;��H;W�H;��H;+�H;��H;��H;�H;6�H;j�H;��H;��H;��H;��H;��H;��H;�H;��H;o�H;^�H;I�H;0�H;�H;�H;�H;�H;�H;�H;�H;�H;"�H;0�H;H�H;Y�H;k�H;��H;��H;��H;��H;��H;��H;��H;��H;e�H;4�H;�H;��H;��H;+�H;��H;U�H;��H;��H;��H;m�H;��H;��H;�H;��H;x�H;D�H;(�H;      ��H;��H;��H;�H;X�H;��H;�H;g�H;��H;H�H;��H;&�H;��H;�H;_�H;��H;��H;&�H;L�H;j�H;��H;��H;��H;��H;��H;��H;��H;��H;o�H;x�H;*�H;)�H;N�H;"�H;��H;�H;��H;�H;��H;#�H;S�H;*�H;*�H;r�H;k�H;��H;��H;��H;��H;��H;��H;��H;��H;d�H;L�H;(�H;��H;��H;]�H;�H;��H;'�H;��H;J�H;��H;h�H;�H;��H;[�H;�H;��H;��H;      �H;�H;C�H;z�H;��H;�H;��H;��H;h�H;��H;z�H;��H;W�H;��H;+�H;��H;��H;�H;6�H;j�H;��H;��H;��H;��H;��H;��H;�H;��H;q�H;]�H;I�H;2�H;�H;�H;�H;�H;�H;�H;�H;�H;"�H;0�H;H�H;Y�H;k�H;��H;��H;��H;��H;��H;��H;��H;��H;e�H;4�H;�H;��H;��H;+�H;��H;U�H;��H;~�H;��H;k�H;��H;��H;�H;��H;~�H;I�H;&�H;      h�H;��H;��H;��H;V�H;��H; �H;��H;/�H;��H;h�H;��H;��H;�H;��H;��H;D�H;��H;��H;0�H;L�H;c�H;��H;q�H;��H;��H;��H;|�H;d�H;N�H;V�H;K�H;�H;�H;"�H;�H;��H;�H;�H;�H;"�H;L�H;V�H;H�H;`�H;y�H;��H;��H;��H;o�H;��H;a�H;E�H;*�H;��H;��H;G�H;��H;~�H;�H;��H;��H;k�H;��H;0�H;��H;&�H;��H;Z�H;��H;��H;��H;      C�H;T�H;��H;��H;b�H;��H;��H;\�H;�H;��H;��H;R�H;�H;��H;i�H;�H;��H;��H;b�H;��H;��H;�H;7�H;W�H;r�H;h�H;n�H;d�H;e�H;e�H;9�H;9�H;;�H;&�H;�H;�H;#�H;�H;�H;&�H;@�H;:�H;7�H;a�H;`�H;c�H;q�H;m�H;o�H;P�H;=�H;�H;��H;��H;b�H;��H;��H;�H;h�H;��H;�H;R�H;��H;��H;�H;]�H;��H;��H;i�H;��H;��H;V�H;      ��H;��H;�H;e�H;�H;��H;��H;��H;��H;��H;��H;�H;��H;��H;��H;��H;S�H;��H;}�H;��H;[�H;��H;��H;�H;-�H;*�H;K�H;a�H;d�H;R�H;9�H;:�H;@�H;;�H;�H;�H;I�H;�H;�H;=�H;B�H;@�H;9�H;O�H;^�H;`�H;N�H;2�H;*�H;�H;��H;��H;U�H;��H;~�H;��H;S�H;��H;��H;��H; �H;�H;��H;��H;��H;��H;��H;��H;�H;l�H;�H;��H;      v�H;��H;��H;��H;�H;��H;�H;c�H;��H;f�H;��H;b�H;��H;6�H;u�H;��H;��H;x�H;I�H;�H;��H;��H;i�H;��H;��H;�H;(�H;9�H;I�H;A�H;D�H;S�H;9�H;6�H;I�H;)�H;"�H;,�H;E�H;6�H;>�H;U�H;E�H;A�H;G�H;7�H;)�H;�H;��H;��H;q�H;��H;��H;�H;J�H;x�H;��H;��H;r�H;6�H;��H;b�H;��H;h�H;��H;c�H;�H;��H;��H;��H;��H;��H;      5�H;~�H;�H;�H;Z�H;��H;��H;��H;��H;(�H;S�H;t�H;}�H;`�H;$�H;��H;]�H;��H;��H;��H;��H;�H;��H;�H;��H;��H;��H;�H;,�H;B�H;R�H;L�H;;�H;>�H;`�H;K�H;,�H;L�H;\�H;A�H;@�H;N�H;S�H;A�H;(�H;�H;��H;��H;��H;�H;��H; �H;~�H;��H;��H;��H;a�H;��H;#�H;]�H;{�H;t�H;Q�H;(�H;��H;��H;��H;��H;f�H;&�H;�H;{�H;      ��H;��H;��H;�H;�H;x�H;2�H;1�H;7�H;`�H;��H;��H;��H;N�H;��H;��H;�H;��H;��H;��H;��H;�H;��H;h�H;��H;7�H;��H;��H;�H;!�H;=�H;@�H;I�H;a�H;K�H;W�H;n�H;Y�H;I�H;c�H;P�H;B�H;>�H;�H;	�H;��H;��H;?�H;��H;e�H;��H;�H;��H;��H;��H;��H;�H;��H;��H;N�H;��H;��H;��H;`�H;3�H;0�H;5�H;i�H;�H;�H;��H;��H;      ��H;��H;&�H;��H;��H;n�H;x�H;�H;p�H;�H;��H;#�H;:�H;&�H;��H;�H;��H;K�H;��H;��H;&�H;c�H;��H;p�H;$�H;��H;C�H;��H;��H;	�H;&�H;I�H;]�H;c�H;a�H;k�H;k�H;m�H;a�H;d�H;`�H;I�H;)�H;�H;��H;��H;F�H;��H;!�H;k�H;��H;c�H;#�H;��H;��H;G�H;��H;�H;��H;#�H;:�H;!�H;��H;�H;m�H;�H;|�H;g�H;��H;��H;'�H;|�H;      �lH;nH;�rH;�yH;3�H;��H;�H;��H;��H;٬H;��H;��H;��H;��H;��H;(�H;7�H;��H;��H;W�H;��H;l�H;��H;2�H;>�H;��H;��H;/�H;��H;��H;�H;7�H;Z�H;c�H;|�H;��H;��H;��H;|�H;e�H;a�H;:�H;�H;��H;��H;/�H;��H;�H;;�H;-�H;��H;l�H;��H;W�H;��H;��H;9�H;(�H;��H;��H;��H;��H;��H;جH;��H;��H;�H;��H;A�H;�yH;�rH;nH;      (�G;��G;�G;��G;dH;n0H;�LH;fH;7|H;?�H;H�H;@�H;E�H;X�H;��H;�H;��H;��H;��H;E�H;H�H;��H;��H;��H;��H;�H;��H;��H;M�H;��H;��H;/�H;K�H;r�H;��H;��H;��H;��H;��H;u�H;O�H;2�H;��H;��H;J�H;��H;��H;#�H;��H;��H;�H;��H;G�H;I�H;��H;��H;��H;�H;��H;W�H;G�H;>�H;F�H;>�H;4|H;fH;�LH;g0H;lH;��G;�G;��G;      �HF;�TF;�vF;�F;v�F;�8G;��G;��G;�	H;�=H;fH;C�H;��H;ƥH;��H;��H;��H;b�H;.�H;(�H;:�H;��H;S�H;��H;m�H;��H;�H;�H;��H;@�H;��H;!�H;2�H;o�H;��H;��H;��H;��H;��H;q�H;4�H;"�H;��H;D�H;��H;�H;�H;��H;l�H;��H;Z�H;��H;9�H;*�H;0�H;[�H;��H;��H;��H;ĥH;��H;?�H; fH;�=H;�	H;��G;��G;q8G;��F;�F;�vF;�TF;      ǣB;�B;�C;��C;�0D;��D;��E;hIF;��F;jG; �G;F$H;�\H;��H;��H;��H;�H;��H;��H;;�H;��H;g�H;��H;�H;��H;h�H;��H;A�H;'�H;��H;��H;��H;)�H;r�H;��H;��H;��H;��H;��H;u�H;-�H;��H;��H;��H;&�H;?�H;��H;p�H;��H;�H;��H;i�H;��H;<�H;��H;��H;"�H;��H;��H;��H;�\H;B$H;�G;jG;��F;eIF;��E;��D;�0D;��C;�C;�B;      �:;�:;r�;;��<;�>;��?;JA;��B;FD; |E;$wF;k8G;��G;<'H;�eH;H�H;4�H;G�H;X�H;o�H;��H;�H;��H;��H;�H;��H;��H;2�H;r�H;j�H;�H;��H;�H;\�H;}�H;��H;��H;��H;{�H;]�H;�H;��H;�H;p�H;u�H;2�H;��H;��H;�H;��H;��H;�H;��H;t�H;[�H;E�H;7�H;H�H;�eH;@'H;��G;i8G;$wF; |E;FD;��B;JA;��?;	>;�<;q�;;�:;      �*;9�*;Y,;kd.;|Y1;ı4;�+8;��;;:�>;�IA;'xC;[*E;�kF;{NG;��G;�DH;�{H;�H;��H;�H;+�H;0�H;��H;��H;��H;T�H;�H;��H;��H;��H;��H;m�H;��H;9�H;��H;��H;��H;��H;��H;:�H;��H;p�H;��H;��H;��H;��H;�H;[�H;��H;��H;��H;2�H;.�H;�H;��H;�H;�{H;�DH;��G;zNG;�kF;Z*E;*xC;�IA;:�>;��;;�+8;±4;}Y1;ld.;Z,;"�*;      "�
;C�;�;;>�;�`;�D&;�-;�D3;(�8;�H=;c�@;��C;#|E;`�F;۠G;8$H;�mH;|�H;�H;նH;��H;.�H;�H;g�H;��H;��H;r�H;f�H;�H;�H;��H;��H;�H;a�H;��H;��H;��H;a�H;�H;��H;��H;!�H;�H;g�H;r�H;��H;��H;d�H;�H;3�H;��H;նH;�H;~�H;�mH;:$H;۠G;a�F;$|E;��C;_�@;�H=;&�8;�D3;�-;{D&;�`;R�;�;�;;�;      ��:ݍ�:��:��:���:�P�:�{;(;��;�~(;�Y1;�t8;?�=;�A;U�D;�HF;scG;�	H;dH;g�H;B�H;ѶH;(�H;��H;��H;2�H;@�H;��H;�H;��H;|�H;��H;Q�H;��H;G�H;��H;��H;��H;E�H;��H;R�H;��H;��H;��H;�H;��H;G�H;6�H;��H;��H;,�H;϶H;E�H;j�H;dH;�	H;tcG;�HF;T�D;�A;?�=;�t8;�Y1;�~(;��;(;�{;�P�: ��:��:��:���:      ��R�� � l7��D^9D�:d�X:Ͽ�:���:�P�:ܣ;��;�);�D3;C�:;�!@;̨C;.�E;�8G;��G;�`H;l�H;�H;�H;t�H;:�H;)�H;C�H;X�H;��H;��H;��H;�H;��H;��H;-�H;h�H;c�H;j�H;*�H;��H;��H;�H;��H;��H;��H;[�H;I�H;,�H;7�H;y�H;�H;�H;k�H;�`H;��G;�8G;1�E;̨C;�!@;B�:;�D3;�);��;٣;�P�:���:ÿ�:<�X:\�:�C^9 j7�  �      s�)�1�$�C�����2���D�\�O���R�94j:���:���:~�;N� ;�d.;�+8;~�>;1C;��E;�)G;��G;dH;{�H;��H;X�H;��H;,�H;��H;��H;��H;��H;��H;F�H;z�H;_�H;��H;4�H;I�H;4�H;��H;_�H;z�H;H�H;��H;��H;��H;��H;��H;/�H;��H;\�H;��H;|�H;dH;��G;�)G;��E;1C;{�>;�+8;�d.;M� ;|�;��:���:4j:S�9 O��`�\�.������I��-�$�      P�ѻ�ͻ6���FG��꿐�a�d���$��Iɺ�!� L^98�r:��: 1;�; �*;�Z6;�>;4�B;��E;�8G;�	H;�mH;�H;B�H;��H;]�H;��H;��H;D�H;��H;��H;t�H;��H;��H;��H;�H;!�H;�H;��H;��H;��H;t�H;��H; �H;E�H;��H;��H;[�H;��H;C�H;�H;�mH;�	H;�8G;��E;2�B;�>;�Z6; �*;�;�0;��:D�r: L^9�!��IɺÃ$�i�d�꿐�HG��:����ͻ      ��I�0�E��(;��O*����<��#GĻȿ���s@�DIҺ�~�:*�:�P�:��;�~(;�5;�>;0C;+�E;vcG;4$H;�{H;3�H;�H;��H;��H;3�H;��H;�H;V�H;��H;M�H;��H;@�H;��H;��H;��H;<�H;��H;J�H;��H;W�H;�H;��H;6�H;��H;��H;�H;4�H;�{H;6$H;scG;/�E;0C;�>;�5;�~(;��;�P�:*�:��:�~�HIҺ�s@�ʿ��$GĻ�<�����O*��(;�.�E�      -p��ex��ע��R��)��p�`� �7�<��.�ѻ�,��k�$�ǅ���09,�:���:~;�~(;�Z6;{�>;ȨC;�HF;ؠG;�DH;D�H;��H;��H;�H;#�H;�H;��H;��H;��H;��H;�H;��H;�H;��H;�H;��H;�H;��H;��H;��H;��H;�H;&�H;�H;��H;��H;D�H;�DH;ؠG;�HF;̨C;x�>;�Z6;�~(;z;���:0�:��09ǅ�j�$��,��.�ѻ<���7�p�`�*���R��ע�ex��      0]� �.#�������ټ�ɺ������
v��(;�Ψ�B^���5R�:��� �6����:���:�;�*;�+8;!@;V�D;^�F;��G;�eH;}�H;��H;��H;��H;��H;��H;�H;o�H;��H;d�H;z�H;'�H;V�H;(�H;w�H;b�H;��H;n�H;�H;��H;��H;��H;��H;��H;z�H;�eH;��G;^�F;N�D;�!@;�+8;�*;�;���:���: �6�>����5R�B^��Ψ��(;��
v������ɺ���ټ����.#� �      �_� \�"<Q�g@�� +��5�����[�ļz�`�`����Iͻk�Iɺ �6�:�:�P�:!�;�d.;B�:;!�A;$|E;xNG;@'H;��H;åH;W�H;��H;%�H;H�H;Y�H;0�H;��H;��H;�H;��H;��H;��H;�H;��H;��H;/�H;V�H;K�H;#�H;��H;V�H;��H;��H;@'H;{NG;#|E;�A;F�:;�d.;�;�P�:0�: �6�
Iɺk�Iͻ���`�`�y�Z�ļ�����5�� +�g@�!<Q� \�      A���R��%ڟ�����C���_�,:�������-p���vz��O*��4ֻk�2�����09&�:1;K� ;�D3;E�=;��C;�kF;��G;�\H;��H;G�H;��H;:�H;��H;v�H;��H;��H;�H;��H;S�H;��H;Q�H;��H;�H;��H;��H;t�H;��H;:�H;��H;E�H;��H;�\H;��G;�kF;��C;=�=;�D3;H� ; 1;"�:��098���k��4ֻ�O*��vz�.p����輤��,:��_� C������&ڟ��R��      �` ��.�����ڽ�b��vr��[��\�z +�� ��ɺ�@��O*�Jͻ�5R�ǅ���:��:~�;�);�t8;`�@;X*E;i8G;=$H;;�H;;�H;�H;�H;��H;m�H;]�H;�H;M�H;��H;��H;�H;��H;��H;M�H;��H;]�H;j�H;��H;"�H;�H;:�H;8�H;8$H;g8G;Z*E;]�@;�t8;�);{�;��:��:"ǅ��5R�Jͻ�O*�@��ɺ�� �z +�\�\��vr���b����ڽ��.��      �-=�@�9��k/�0�����~��Ľ�!��iys�C�6�%#��ɺ��vz����C^��n�$� ��r:���:��;�Y1;�H=;'xC;"wF;�G;�eH;B�H;�H;��H;��H;N�H;��H;��H;��H;`�H;v�H;��H;v�H;`�H;��H;��H;��H;L�H;��H;��H;~�H;B�H;�eH;�G;!wF;&xC;�H=;�Y1;��;���: �r:�~�p�$�D^������vz��ɺ�%#�C�6�iys��!����Ľ~���0���k/�@�9�      �(��Fl���.}�9ce�zPH���(�{
���ڽ�R�� �{�C�6�� �.p��`�`�Ψ��,��TIҺ�K^9���:գ;�~(;(�8;�IA;�{E;	jG;�=H;<�H;ѬH;�H;\�H;#�H;f�H;��H;��H;��H;��H;I�H;��H;��H;��H;��H;e�H;#�H;_�H;�H;ѬH;<�H;�=H;jG;�{E;�IA;&�8;�~(;أ;|��:�K^9TIҺ�,��Ψ�`�`�.p��� �C�6� �{��R����ڽ|
���(�zPH�9ce��.}�Fl��      �iþVD��7o�����������i��-=�ht� ���R��iys�z +����z񗼖(;�.�ѻ�s@��!��3j:�P�:��;�D3;-�>;FD;��F;�	H;5|H;��H;p�H;2�H;��H;��H;��H;�H;)�H;h�H;��H;h�H;+�H;�H;��H;��H;��H;3�H;p�H;��H;7|H;�	H;��F;FD;0�>;�D3;��;�P�:�3j: �!��s@�.�ѻ�(;�z����z +�iys��R�� ��ht��-=��i���������7o��VD��      ���
�����$�޾VD���A���.}�(�D�ht���ڽ�!��\����\�ļ�
v�>��ο���Iɺ�R�9���:(;�-;�;;��B;cIF;��G;fH;��H;�H;)�H;��H;c�H;��H;Y�H;��H;��H;d�H;��H;��H;V�H;��H;`�H;��H;0�H;�H;��H;fH;��G;`IF;��B;�;;�-;(;���:�R�9�IɺͿ��?���
v�\�ļ���\��!����ڽht�(�D��.}��A��VD��$�޾�����
�      ��7�Е3��f'�)��\���о�����.}��-=�{
���Ľ\��,:����������7�&GĻ΃$�XO�����:�{;~D&;�+8;JA;�E;��G;tLH;�H;t�H;/�H;��H;��H;��H;��H;�H;|�H;�H;{�H;�H;��H;��H;��H;��H;5�H;t�H;�H;wLH;��G;�E;JA;�+8;zD&;�{;���:`O��̓$�%GĻ�7���������,:�\����Ľ{
��-=��.}������о�\��)��f'�Е3�      Yo�_Xi��"Y���@�K�#��
��о�A���i���(�~��wr���_��5��ɺ�r�`��<��p�d���\�8�X:�P�:�`;��4;��?;��D;n8G;f0H;��H;i�H;r�H;�H;��H;��H;��H;��H;�H;��H;�H;��H;��H;��H;��H;��H;u�H;j�H;��H;j0H;w8G;��D;��?;��4;�`;�P�:<�X:��\�p�d��<��r�`��ɺ��5��_�wr��~����(��i��A���о�
�K�#���@��"Y�_Xi�      /����������Yo��!J�K�#��\��VD������zPH�����b�� C��� +���ټ*����򿐻"���H�:��:=�;�Y1;>;�0D;r�F;[H;?�H;��H;�H;W�H;��H;�H;a�H;B�H;��H;[�H;��H;C�H;\�H;�H;��H;T�H;�H;��H;A�H;bH;}�F;�0D;>;�Y1;<�;��:P�:&���𿐻��)����ټ� +� C���b�����zPH�����VD���\��K�#��!J�Yo��������      =^������k���Yo���@�)�$�޾����9ce�0����ڽ󻒽g@������R���O*�NG�� ��� C^9��:�;Rd.;��<;��C;�F;��G;�yH;��H;�H;�H;��H;g�H;��H;��H;~�H;�H;{�H;��H;��H;h�H;��H;�H;�H;��H;�yH;��G;��F;��C;��<;Pd.;�;��:pC^9(���LG���O*��R������g@�󻒽��ڽ0��9ce�����$�޾)���@�Yo�k�������      �aǿ�¿����������"Y��f'�����7o���.}��k/����%ڟ�"<Q�.#�ע��(;�4���@�� o7���:�;h,;��;;�C;�vF;�G;�rH;�H;��H;�H;��H;��H;��H;��H;G�H;��H;C�H;��H;��H;��H;��H;
�H;��H;�H;�rH;�G;�vF;�C;�;;e,;�;��: j7�A��4����(;�ע�.#�"<Q�%ڟ�����k/��.}�7o�������f'��"Y�����������¿      3�ֿCpѿ�¿������_Xi�Е3��
�VD��Fl��A�9��.���R��!\� �fx��2�E��ͻ#�$�� �ύ�:6�;E�*;1�:;�B;�TF;��G;#nH;��H;��H;g�H;��H;��H;W�H;}�H;�H;��H;�H;}�H;W�H;��H;��H;b�H;ķH;��H;#nH;��G;�TF;�B;-�:;>�*;4�;Ǎ�:p �&�$��ͻ3�E�fx�� �!\��R���.��@�9�Fl��VD���
�Е3�_Xi��������¿Cpѿ      �?��|h��=v��� ��7�X��O/�/y�A�;ఖ��+X����ѽ����_n;�]�������B(�ߚ��f��Оe9�:�;�Y.;P�<;aWC;�ZF;��G;�/H;/jH;4�H;B�H;~�H;%�H;��H;V�H;��H;��H;��H;P�H;��H;"�H;z�H;>�H;<�H;/jH;�/H;��G;�ZF;\WC;L�<;�Y.;�;
�:�e9h��ޚ���B(�����]��_n;������ѽ���+X�ఖ�A�;/y��O/�7�X�� ��=v��|h��      |h��/���a�����y�VvS�pM+��v�9ɾ�����T� ]�\ν����y\8�����x��%�R�������9a-�:a�;��.;�<;�nC;�dF;�G;�1H;�jH;��H;��H;ǵH;f�H;��H;a�H;��H;��H;��H;a�H;��H;c�H;ƵH;��H;��H;�jH;�1H;�G;�dF;�nC;�<;��.;_�;[-�:0�9���R���%��x�����y\8�����\ν ]��T�����9ɾ�v�pM+�VvS���y�a���/���      =v��b���W ��`�h�6E�W��i���|㼾}���nH�ӈ�y�ý�Ȅ��s/��o��#�����)J��:к	�9Hg�:�l;0;]=;ӲC;ҀF;j�G;6H;mH;"�H;��H;{�H;��H;;�H;��H;�H;��H;��H;��H;:�H;��H;z�H;��H;)�H;mH;6H;m�G;݀F;ҲC;]=;0;�l;Dg�:0	�9>к(J������#���o��s/��Ȅ�y�ýӈ��nH�}��|㼾i���W��6E�`�h�W ��a���      � ����y�`�h���N��O/����B�߾B���*|��6�p}�䳽jSt�=�!�prμDF{��_��X��ޓ��:��:�Z;�2;�O>;iD;#�F;v�G;=H;�pH;��H;D�H;ȷH;��H;��H;Z�H;y�H;[�H;r�H;Z�H;��H;��H;ƷH;>�H;��H;�pH;=H;v�G;,�F;eD;�O>;�2;�Z;��:<:�����X���_�DF{�prμ=�!�jSt�䳽p}��6��*|�B��B�߾����O/���N�`�h���y�      7�X�VvS�6E��O/��S�GW����������LS\��� ���:����Y�{��҃����]�����,�b���Y��Y:��:\`;1�4;�?;4�D;��F;�G; FH;AuH;��H;��H;�H;�H;��H;�H;�H;��H;�H;�H;��H;�H;}�H;��H;��H;@uH; FH;	�G;��F;2�D;�?;+�4;\`;��:,�Y:ȇY�,�b�������]�҃��{���Y�:����彑� �LS\���������GW���S��O/�6E�VvS�      �O/�pM+�W�����GW��9ɾA���Mw�� :�j��x�ý�L��\n;�_���tv���E<��˻��-�p��Ty�:�^;�%;v�7;q�@;5E;�"G;�G;3PH;�zH;��H;T�H;v�H;��H;��H;�H;��H;��H;��H;�H;��H;��H;v�H;O�H;��H;�zH;3PH;�G;�"G;5E;m�@;v�7;�%;�^;\y�:x����-��˻�E<�tv��^���\n;��L��w�ýi��� :��Mw�A��9ɾGW�����X��pM+�      /y��v�i���B�߾����A��?����nH���CὝu����d�0O�jrμJ"�����
	������q89F;�:Y�;�+;K|:;t7B;��E;�aG;mH;�ZH;_�H;&�H;��H;�H;E�H;A�H;�H;��H;o�H;��H; �H;A�H;A�H;�H;��H;*�H;^�H;�ZH;kH;�aG;��E;q7B;J|:;�+;T�;R;�:�q89���		�����J"��jrμ0O���d��u��C����nH�?���A������B�߾i����v�      @�;9ɾ|㼾B�������Mw��nH�����Z�䳽˕��r\8�o#������^N�Q���b�$Ix�5:ˮ�:)�;��0;]=;:�C;�[F;ΞG;�)H;�eH;n�H; �H;7�H;��H;�H;��H;&�H;��H;h�H;��H;'�H;��H;�H;|�H;6�H;&�H;n�H;�eH;�)H;ҞG;�[F;5�C;]=;��0;#�;ٮ�: 5:$Ix��b�Q��^N�����o#��r\8�˕��䳽�Z񽰯��nH��Mw�����B��|㼾9ɾ      ఖ�����}���*|�LS\�� :����Z�l$�������K�v���Oļ����������I&�`��5/�:�^;��#;�G6;0�?;�D;@�F;��G;�?H;�pH;ڏH;p�H;�H;H�H;-�H;i�H;m�H;��H;t�H;��H;m�H;g�H;'�H;G�H;�H;t�H;ُH;�pH;�?H;��G;B�F;�D;2�?;�G6;��#;�^;9/�:���J&������������Oļv���K�����l$���Z���� :�LS\��*|�}������      �+X��T��nH��6��� �j��C�䳽�����mR����ټ�����E<��?ݻ?d\������ :�d�:��;"�,;s�:;O7B;��E;gLG;'H;USH;�{H;x�H;�H;�H;:�H;Q�H;�H;��H;��H;��H;��H;��H;�H;N�H;7�H;�H;�H;|�H;�{H;VSH;(H;mLG;��E;P7B;s�:;�,;��;�d�:� :����>d\��?ݻ�E<�����ټ����mR�����䳽C�i���� ��6��nH��T�      �� ]�ӈ�p}���x�ý�u��˕���K�����o�kv���&R�!��Z^����� �>����:UB;2";`�4;��>;6D;��F;�G;�)H;`dH;m�H;�H;[�H;"�H;*�H;~�H;��H;�H;	�H;��H;
�H;�H;��H;|�H;'�H;%�H;c�H;	�H;n�H;adH;�)H;�G;��F;:D;��>;_�4;9";WB;���: �>����Z^�� ���&R�jv���o�����K�˕���u��w�ý��p}�ӈ� ]�       �ѽ\νy�ý䳽9����L����d�r\8�v��ټjv����Y��_����F���[�x�Y:I��:Cm;�r-;�:;f�A;%oE;�"G;D�G;TGH;�sH;ސH;�H;�H;�H;�H;��H;t�H;{�H;%�H;��H;%�H;{�H;x�H;��H;�H;#�H;�H;��H;ߐH;�sH;TGH;I�G;�"G;)oE;i�A;�:;�r-;Cm;I��:��Y:�[�D������_���Y�iv��ټv��q\8���d��L��:���䳽y�ý\ν      ���������Ȅ�kSt��Y�\n;�0O�n#���Oļ�����&R��_������N3��Y��3:��:ί;�?&;�G6;zX?;�D;xF;��G;'!H;�^H;�H;�H;��H;8�H;��H;��H;��H;�H;��H;M�H;�H;M�H;��H;�H;��H;��H;��H;B�H;ƭH;�H;��H;~^H;-!H;��G;"xF;�D;zX?;�G6;�?&;ʯ;��:�3:��Y��N3������_��&R������Oļn#��0O�\n;��Y�kSt��Ȅ�����      ^n;�y\8��s/�=�!�z��`���jrμ��������E<�������N3�tHx�x�9��:�^;K ;#2;Z�<;�B;��E;5G;��G;$FH;sqH;��H;;�H;��H;C�H;��H;��H;��H;��H;�H;k�H; �H;k�H;�H;��H;��H;��H;��H;M�H;��H;>�H;��H;rqH;)FH;��G;$5G;��E;�B;b�<;'2;I ;�^;��:��9dHx��N3�������E<��������jrμ_���{��=�!��s/�x\8�      [������o�prμу��tv��J"��^N�����?ݻX^��K���Y�p�9��:Ŧ�:��;H�.;w|:;�>A;��D;�F;��G;�)H;aH;�H;q�H;׬H;(�H;�H;,�H;T�H;��H;�H;M�H;��H;��H;��H;K�H;�H;��H;P�H;/�H;�H;/�H;ެH;q�H;�H;aH;�)H;��G; �F;��D;�>A;z|:;D�.;��;Ŧ�:��:��9 �Y�F��V^���?ݻ���^N�J"��sv��Ӄ��prμ�o����      �����x���#��BF{���]��E<����N�뻬���=d\�����[��3:��:ɦ�:p[;Z�,;��8;!@;�0D;l[F;{G;�
H;8PH;vH;אH;4�H;�H;�H;[�H;o�H;��H;��H;q�H;m�H;��H;��H;��H;j�H;q�H;��H;��H;q�H;`�H; �H;�H;4�H;ӐH;vH;8PH;�
H;{G;n[F;�0D;!@;��8;^�,;p[;Ϧ�:��:�3:�[����:d\�����L�뻤���E<���]�BF{��#���x��      �B(�%�����_������˻	���b�B&����� �>�|�Y:��:�^;��;_�,;`8;[�?;��C;fF;�FG;<�G;�?H;kH;�H;��H;�H;I�H;��H;_�H;h�H;�H;r�H;��H;��H;{�H;��H;w�H;}�H;��H;o�H;�H;l�H;c�H;��H;J�H;�H;��H;�H;kH;�?H;?�G;�FG;nF;��C;U�?;`8;_�,;��;�^;��:��Y: �>�����A&�
�b�	���˻�����_����%�      њ��M���(J���X��"�b���-����Ix�`��� :���:;��:ǯ;I ;D�.;��8;P�?;�C;��E;$#G;��G;�1H;�aH;=�H;g�H;j�H;��H;��H;P�H;�H;%�H;-�H;��H;�H;�H;2�H;��H;/�H;}�H;�H;��H;)�H;)�H;�H;R�H;��H;��H;h�H;m�H;<�H;�aH;�1H;��G;+#G;��E;��C;S�?;��8;F�.;I ;ȯ;G��:���:� :��Ix������-��b��X��$J��M���      :�����>кؓ��ЇY����r8985:?/�:�d�:^B;?m;�?&;&2;x|:;!@;��C;��E;lG;��G;H(H;�ZH;]zH;,�H;ŤH;��H;W�H;��H;��H;S�H;��H;��H;A�H;#�H;A�H;��H;t�H;��H;?�H;#�H;>�H;��H;��H;W�H;��H;��H;V�H;��H;ʤH;.�H;ZzH;�ZH;L(H;��G;lG;��E;��C;!@;z|:;&2;�?&;Cm;aB;�d�:C/�:85:`r898��ȇY��>к���      ��e9��9X	�9d:�Y:`y�:h;�:Ѯ�:�^;��;9";�r-;�G6;_�<;�>A;�0D;mF;0#G;��G;�$H;OWH;�vH;f�H;1�H;3�H;k�H;�H;�H;n�H;-�H;��H;u�H;��H; �H;�H;��H;��H;��H;�H;�H;��H;q�H;��H;,�H;k�H;�H;��H;i�H;8�H;2�H;c�H;�vH;RWH;�$H;��G;+#G;mF;�0D;�>A;]�<;�G6;�r-;>";��;�^;߮�:`;�:jy�: �Y::	�9��9      H�:C-�:g�: ��:��:�^;T�;#�;��#; �,;`�4;��:;xX?;�B;��D;n[F;�FG;��G;J(H;KWH;YuH;|�H;	�H;�H;�H;��H;��H;��H;��H;��H;��H;��H;��H;��H;��H;P�H;J�H;I�H;��H;��H;��H;��H;��H;��H;��H;��H;��H;��H;�H;�H;�H;}�H;\uH;MWH;K(H;��G;�FG;n[F;��D;�B;zX?;�:;c�4; �,;��#;"�;Z�;�^;��:��:&g�:;-�:      �;k�;�l;�Z;Z`;�%;�+;��0;�G6;x�:;��>;f�A;�D;��E;"�F;{G;@�G;�1H;�ZH;�vH;~�H;<�H;��H;��H;z�H;F�H;��H;��H;��H;��H;0�H;1�H;��H;��H;b�H;��H;��H;��H;`�H;��H;��H;+�H;2�H;��H;��H;��H;��H;G�H;|�H;��H;��H;<�H;��H;�vH;�ZH;�1H;B�G;{G;%�F;��E;�D;l�A;��>;u�:;�G6;��0;�+;�%;p`;�Z;�l;_�;      �Y.;��.;0;�2;'�4;��7;[|:;!]=;<�?;Z7B;BD;,oE;$xF;/5G;��G;�
H;�?H;�aH;^zH;b�H;�H;��H;<�H;��H;X�H;��H;��H;��H;�H;��H;��H;U�H;O�H;>�H;��H;�H;=�H;�H;��H;?�H;K�H;O�H;��H;��H;�H;��H;��H;��H;\�H;��H;8�H;��H;�H;c�H;^zH;�aH;�?H;�
H;��G;+5G;&xF;/oE;ED;V7B;<�?;!]=;Y|:;��7;6�4;�2;0;��.;      J�<;�<;]=;�O>;ہ?;u�@;t7B;:�C;�D;��E;��F;�"G;��G; �G;�)H;;PH;kH;C�H;.�H;.�H;�H;��H;��H;+�H;&�H;)�H;;�H;��H;�H;3�H;��H;�H;�H;��H;<�H;x�H;��H;q�H;;�H;��H; �H;�H;��H;0�H;�H;��H;7�H;,�H;)�H;(�H;��H;��H;�H;-�H;+�H;<�H;kH;=PH;�)H;��G;��G;�"G;��F;��E;�D;A�C;u7B;d�@;�?;�O>;]=;�<;      �WC;�nC;βC;cD;.�D;#5E;��E;�[F;H�F;oLG;��G;M�G;-!H;0FH;aH;vH;��H;t�H;ѤH;<�H;�H;|�H;\�H;/�H;��H;��H;7�H;��H;��H;��H;��H;��H;��H;.�H;��H;��H;��H;��H;��H;1�H;��H;��H;��H;��H;��H;��H;3�H;��H;��H;,�H;[�H;~�H;�H;8�H;ѤH;o�H;��H;vH;aH;-FH;.!H;Q�G;��G;qLG;K�F;�[F;��E;5E;;�D;bD;ϲC;�nC;      �ZF;�dF;׀F;"�F;��F;�"G;�aG;ݞG;��G;/H;�)H;[GH;�^H;|qH;�H;ڐH;��H;j�H;��H;e�H;��H;C�H;��H;,�H;��H;�H;��H;��H;e�H;��H;��H;��H;�H;q�H;��H;�H;�H;�H;��H;q�H;�H;��H;��H;��H;b�H;��H;�H;�H;��H;)�H;��H;D�H;��H;g�H;��H;f�H;��H;ؐH;�H;vqH;�^H;[GH;�)H;0H;��G;ݞG; bG;�"G;��F;'�F;݀F;�dF;      	�G;�G;j�G;w�G;��G;�G;xH;�)H;�?H;YSH;cdH;�sH;�H;��H;p�H;5�H;�H;��H;W�H;��H;��H;��H;��H;>�H;4�H;��H;�H;8�H;{�H;��H;]�H;��H;o�H;��H;�H;5�H;O�H;,�H;��H;��H;o�H;��H;Z�H;��H;w�H;5�H;|�H;��H;6�H;:�H;��H;��H;��H;��H;W�H;��H;�H;6�H;p�H;��H;��H;�sH;fdH;VSH;�?H;�)H;uH;��G;�G;i�G;i�G;֪G;      �/H;�1H;6H;=H;�EH;7PH;�ZH;�eH;�pH;�{H;n�H;�H;�H;A�H;جH;�H;H�H;��H;��H;}�H;��H;��H;��H;��H;��H;��H;5�H;r�H;Z�H;F�H;��H;a�H;��H;�H;@�H;T�H;?�H;O�H;=�H;�H;��H;[�H;��H;C�H;V�H;p�H;2�H;��H;��H;��H;��H;��H;��H;{�H;��H;��H;I�H;�H;׬H;A�H;�H;�H;r�H;�{H;�pH;�eH;�ZH;*PH;FH;=H;6H;�1H;      )jH;�jH;mH;�pH;2uH;�zH;f�H;n�H;ԏH;y�H;	�H;��H;ĭH;��H;*�H; �H;��H;U�H;��H;n�H;��H;��H;�H;�H;��H;^�H;r�H;\�H;O�H;��H;L�H;��H;��H;.�H;]�H;d�H;U�H;`�H;[�H;/�H;��H;��H;L�H;��H;L�H;W�H;n�H;^�H;��H;�H;�H;��H;��H;j�H;��H;R�H;��H; �H;*�H;��H;ĭH;��H;�H;|�H;ԏH;n�H;f�H;�zH;>uH;�pH;mH;�jH;      5�H;��H;,�H;��H;��H;��H;)�H;!�H;t�H;�H;a�H;�H;>�H;L�H;�H;[�H;c�H;	�H;N�H;*�H;��H;��H;��H;-�H;��H;��H;}�H;F�H;��H;B�H;��H;��H;,�H;V�H;b�H;w�H;��H;u�H;_�H;U�H;,�H;��H;��H;=�H;��H;F�H;{�H;��H;��H;,�H;��H;��H;��H;'�H;N�H;�H;c�H;]�H;�H;I�H;>�H;�H;b�H;�H;t�H;!�H;,�H;��H;H;��H;/�H;��H;      I�H;��H;��H;E�H;��H;S�H;��H;:�H;�H;�H;*�H;)�H;�H;��H;3�H;s�H;p�H;,�H;��H;��H;��H;3�H;��H;��H;��H;��H;X�H;��H;N�H;��H;��H;"�H;V�H;f�H;�H;~�H;x�H;{�H;|�H;g�H;Y�H; �H;��H;��H;J�H;��H;V�H;��H;��H;��H;��H;2�H;��H;��H;��H;*�H;s�H;t�H;2�H;��H;�H;,�H;,�H;�H;�H;;�H;��H;I�H;��H;E�H;��H;��H;      {�H;εH;x�H;��H;x�H;k�H;�H;��H;L�H;:�H;*�H;�H;��H;��H;W�H;��H;�H;0�H;��H;x�H;��H;1�H;Q�H;�H;��H;��H;��H;b�H;��H;��H;�H;:�H;`�H;~�H;��H;��H;��H;��H;��H;�H;d�H;7�H;�H;��H;��H;^�H;��H;��H;��H;��H;V�H;1�H;��H;u�H;��H;2�H;�H;��H;W�H;��H;��H;�H;/�H;=�H;L�H;��H;��H;o�H;��H;��H;��H;еH;      (�H;p�H;�H;��H;�H;�H;C�H;�H;%�H;O�H;��H;��H;��H;��H;��H;��H;u�H;��H;E�H;��H;��H;��H;K�H;��H;��H;�H;l�H;��H;��H;2�H;U�H;d�H;t�H;��H;��H;��H;��H;��H;��H;��H;w�H;d�H;T�H;+�H;��H;��H;m�H;�H;��H;��H;P�H;��H;��H;��H;E�H;��H;z�H;��H;��H;��H;��H;��H;��H;R�H;)�H;�H;F�H;w�H;�H;��H;�H;n�H;      ��H;��H;>�H;��H;��H;��H;E�H;��H;j�H;�H;��H;}�H;�H;��H;�H;v�H;��H;�H;$�H;$�H;��H;��H;8�H;��H;(�H;j�H;��H;�H;,�H;Y�H;b�H;��H;��H;�H;��H;��H;��H;��H;��H;�H;��H;��H;b�H;V�H;+�H;�H;��H;l�H;+�H;��H;A�H;��H;��H;�H;$�H;�H;��H;x�H;�H;��H;�H;|�H;��H;�H;n�H;��H;I�H;��H;��H;��H;D�H;��H;      P�H;r�H;��H;\�H;(�H;��H;
�H;(�H;q�H;��H;�H;��H;��H;�H;T�H;o�H;��H;}�H;A�H;�H;��H;`�H;��H;1�H;��H;��H;��H;?�H;`�H;f�H;z�H;��H;��H;��H;��H;��H;��H;��H;��H;��H;��H;��H;x�H;`�H;Y�H;:�H;��H;��H;��H;1�H;��H;^�H;��H; �H;@�H;��H;��H;r�H;T�H;�H;��H;��H;$�H;��H;w�H;+�H;�H;��H;(�H;^�H;��H;s�H;      ��H;��H;��H;u�H;�H;��H;��H;��H;��H;��H;�H;)�H;N�H;q�H;��H;��H;{�H;/�H;��H;��H;Q�H;��H;�H;i�H;��H;�H;+�H;T�H;g�H;~�H;|�H;��H;��H;��H;��H;��H;��H;��H;��H;��H;��H;��H;{�H;x�H;d�H;R�H;/�H;�H;��H;j�H;�H;��H;O�H;��H;��H;3�H;��H;��H;��H;p�H;S�H;)�H;�H;��H;��H;��H;��H;��H;�H;p�H;��H;��H;      ��H;��H;��H;[�H;��H;��H;v�H;i�H;x�H;��H;��H;��H;�H;
�H;��H;��H;��H;��H;u�H;��H;S�H;��H;<�H;��H;��H;�H;H�H;G�H;[�H;��H;u�H;��H;��H;��H;��H;��H;��H;��H;��H;��H;��H;��H;u�H;��H;V�H;D�H;M�H;�H;��H;��H;C�H;��H;O�H;��H;v�H;��H;��H;��H;��H;	�H;�H;��H;��H;��H;{�H;n�H;|�H;��H;��H;\�H;��H;��H;      ��H;��H;��H;s�H;�H;��H;��H;��H;��H;��H;�H;)�H;N�H;q�H;��H;��H;z�H;.�H;��H;��H;Q�H;��H;�H;i�H;��H;�H;+�H;R�H;i�H;|�H;|�H;��H;��H;��H;��H;��H;��H;��H;��H;��H;��H;��H;{�H;w�H;d�H;Q�H;/�H;	�H;��H;i�H;�H;��H;O�H;��H;��H;3�H;�H;��H;��H;n�H;P�H;)�H;�H;��H;��H;��H;��H;��H;�H;u�H;�H;��H;      C�H;u�H;��H;U�H;)�H;��H;�H;+�H;q�H;��H; �H;��H;��H;�H;U�H;r�H;��H;~�H;A�H;�H;��H;a�H;��H;1�H;��H;��H;��H;=�H;_�H;d�H;x�H;��H;��H;��H;��H;��H;��H;��H;��H;��H;��H;��H;x�H;_�H;\�H;:�H;��H;��H;��H;/�H;��H;`�H;��H; �H;@�H;��H;��H;r�H;R�H;�H;��H;��H;!�H;��H;r�H;2�H;�H;��H;/�H;Z�H;��H;v�H;      ��H;��H;;�H;��H;��H;��H;B�H;��H;k�H;�H;��H;{�H;�H;��H;�H;x�H;��H;�H;$�H;"�H;��H;��H;;�H;��H;+�H;l�H;��H;�H;.�H;Y�H;`�H;��H;��H;�H;��H;��H;��H;��H;��H;��H;��H;��H;`�H;V�H;(�H;�H;��H;o�H;*�H;��H;A�H;��H;��H; �H;&�H;�H;��H;x�H;�H;��H;�H;{�H;��H;�H;k�H;��H;K�H;��H;��H;��H;D�H;��H;      )�H;r�H;�H;��H;�H;��H;A�H;�H;&�H;R�H;��H;��H;��H;��H;��H;��H;w�H;��H;D�H;��H;��H;��H;I�H; �H;��H;�H;j�H;��H;��H;2�H;T�H;b�H;r�H;��H;��H;��H;��H;��H;��H;��H;u�H;d�H;T�H;,�H;��H;��H;m�H;�H;��H;��H;R�H;��H;��H;��H;D�H;��H;w�H;��H;��H;��H;��H;��H;��H;Q�H;'�H;�H;I�H;~�H;�H;��H;�H;m�H;      o�H;͵H;p�H;��H;w�H;{�H;��H;��H;K�H;:�H;+�H;�H;��H;��H;Z�H;��H;�H;2�H;��H;x�H;��H;2�H;Q�H;�H;��H;��H;��H;_�H;��H;��H;�H;7�H;`�H;|�H;��H;��H;��H;��H;��H;�H;c�H;9�H;�H;��H;��H;^�H;��H;��H;��H;��H;X�H;2�H;��H;u�H;��H;/�H;�H;��H;V�H;��H;��H;�H;+�H;:�H;N�H;��H;��H;n�H;x�H;��H;u�H;ǵH;      >�H;��H;��H;B�H;��H;S�H;��H;;�H;�H;�H;)�H;,�H;�H;��H;5�H;t�H;r�H;*�H;��H;��H;��H;3�H;��H;��H;��H;��H;V�H;��H;P�H;��H;��H;"�H;U�H;f�H;��H;|�H;x�H;�H;~�H;i�H;[�H;"�H;��H;��H;J�H;��H;W�H;��H;��H;��H;��H;4�H;��H;��H;��H;*�H;u�H;t�H;3�H;��H;�H;*�H;)�H;�H;�H;@�H;��H;P�H;��H;L�H;��H;��H;      A�H;��H;(�H;��H;��H;��H;*�H;'�H;w�H;�H;a�H;�H;?�H;J�H;�H;\�H;b�H;�H;N�H;*�H;��H;��H;�H;,�H;��H;��H;}�H;F�H;��H;@�H;��H;��H;)�H;X�H;c�H;w�H;��H;x�H;`�H;X�H;.�H;��H;��H;?�H;��H;C�H;}�H;��H;��H;'�H;��H;��H;��H;'�H;P�H;�H;c�H;]�H;�H;J�H;>�H;�H;b�H;�H;t�H;&�H;,�H;��H;H;��H;0�H;��H;      6jH;�jH;&mH;�pH;,uH;�zH;e�H;n�H;ڏH;x�H;
�H;��H;ƭH;��H;,�H; �H;��H;V�H;��H;k�H;��H;��H;�H;�H;��H;[�H;p�H;W�H;P�H;��H;J�H;��H;��H;/�H;]�H;d�H;V�H;d�H;\�H;/�H;��H;��H;M�H;��H;L�H;V�H;p�H;a�H;��H;�H;�H;��H;��H;k�H;��H;R�H;��H;!�H;,�H;��H;ĭH;��H;
�H;x�H;ُH;s�H;i�H;�zH;:uH;�pH;'mH;�jH;      	0H;�1H;	6H;=H;�EH;APH;�ZH;�eH;�pH;�{H;q�H;�H;�H;A�H;۬H;�H;H�H;��H;��H;{�H;��H;��H;��H;��H;��H;��H;2�H;p�H;Z�H;C�H;��H;_�H;��H;�H;?�H;R�H;A�H;T�H;=�H;	�H;��H;_�H;��H;F�H;W�H;p�H;4�H;��H;��H;��H;��H;��H;��H;{�H;��H;��H;I�H;�H;۬H;>�H;�H;�H;r�H;�{H;�pH;�eH;�ZH;0PH;FH;=H;6H;�1H;      ��G;��G;d�G;~�G;�G;	�G;xH;�)H; @H;WSH;ddH;�sH;�H;��H;q�H;5�H;�H;��H;V�H;��H;��H;��H;��H;?�H;4�H;��H;|�H;6�H;z�H;��H;X�H;��H;m�H;��H;�H;0�H;O�H;0�H;��H;��H;p�H;��H;]�H;��H;w�H;5�H;}�H;��H;3�H;:�H;��H;��H;��H;��H;Y�H;��H;�H;6�H;r�H;��H;~�H;�sH;cdH;VSH;�?H;�)H;zH;�G;�G;}�G;i�G;ߪG;      �ZF;�dF;ހF;�F;��F;�"G;�aG;��G;��G;.H;�)H;\GH;�^H;xqH;�H;ڐH;��H;l�H;��H;d�H;��H;C�H;��H;,�H;��H;�H;��H;��H;e�H;��H;��H;��H;�H;s�H;��H;�H;�H;�H;��H;s�H;�H;��H;��H;��H;a�H;��H;��H;�H;��H;)�H;��H;C�H;��H;g�H;��H;f�H;��H;ڐH;�H;xqH;�^H;YGH;�)H;/H;��G;ٞG;�aG;�"G;��F;�F;ȀF;}dF;      }WC;�nC;ȲC;aD;1�D;#5E;��E;�[F;K�F;oLG;��G;P�G;-!H;+FH;aH;vH;��H;r�H;ФH;8�H;�H;|�H;Z�H;/�H;��H;��H;3�H;��H;��H;��H;��H;��H;��H;/�H;��H;��H;��H;��H;��H;1�H;��H;��H;��H;��H;��H;��H;7�H;��H;��H;,�H;^�H;~�H;�H;;�H;ӤH;o�H;��H;vH;aH;-FH;.!H;P�G;��G;qLG;G�F;�[F;��E;5E;7�D;bD;ʲC;�nC;      '�<;�<;	]=;�O>;Ӂ?;y�@;v7B;<�C;��D;��E;��F;�"G;��G;��G;�)H;;PH;kH;A�H;)�H;+�H;�H;��H;��H;+�H;(�H;#�H;8�H;��H;�H;.�H;��H;�H;�H;��H;=�H;x�H;��H;z�H;<�H;��H;�H;	�H;��H;3�H;�H;��H;<�H;*�H;(�H;+�H;��H;��H;�H;/�H;.�H;=�H;kH;;PH;�)H;��G;��G;�"G;��F;��E;�D;8�C;t7B;n�@;�?;�O>;	]=;��<;      �Y.;��.;0;�2;$�4;z�7;R|:;!]=;>�?;V7B;=D;,oE;"xF;)5G;��G;�
H;�?H;�aH;\zH;`�H;�H;��H;8�H;��H;[�H;��H;��H;��H;�H;��H;��H;U�H;L�H;>�H;��H;�H;@�H;�H;��H;<�H;O�H;V�H;��H;��H;�H;��H;��H;��H;Z�H;��H;;�H;��H;�H;d�H;^zH;�aH;�?H;�
H;��G;(5G;#xF;,oE;>D;V7B;>�?;$]=;T|:;z�7;$�4;�2;	0;~�.;      �;k�;�l;�Z;\`;�%;�+;��0;�G6;s�:;��>;l�A;�D;��E;#�F;{G;?�G;�1H;�ZH;�vH;~�H;:�H;��H;��H;|�H;A�H;��H;��H;��H;��H;0�H;/�H;��H;��H;`�H;��H;��H;��H;`�H;��H;��H;1�H;6�H;��H;��H;��H;��H;G�H;{�H;¸H;��H;<�H;~�H;�vH;�ZH;�1H;@�G;{G;#�F;��E;�D;j�A;��>;u�:;�G6;��0;�+;�%;r`;�Z;�l;a�;      2�:s-�:2g�:��:��:�^;Y�;&�;��#;�,;b�4;�:;xX?;�B;��D;o[F;�FG;��G;H(H;KWH;XuH;}�H;�H;�H;�H;��H;��H;��H;��H;��H;��H;��H;��H;��H;��H;L�H;L�H;M�H;��H;��H;��H;��H;��H;��H;��H;��H;��H;��H;�H;�H;�H;z�H;[uH;OWH;K(H;��G;�FG;n[F;��D;�B;xX?; �:;e�4;�,;��#;)�;Z�;�^;��:��:Jg�:K-�:      ��e9�9	�9p:�Y:jy�:j;�:��:�^;��;=";�r-;�G6;]�<;�>A;�0D;lF;-#G;��G;�$H;PWH;�vH;c�H;/�H;7�H;g�H;��H;}�H;m�H;'�H;��H;u�H;��H;!�H;�H;��H;��H;��H;�H;�H;��H;u�H;��H;-�H;n�H;��H;�H;k�H;4�H;5�H;c�H;�vH;PWH;�$H;��G;+#G;nF;�0D;�>A;^�<;�G6;�r-;>";��;�^;ٮ�:`;�:Zy�:$�Y:<:(	�9��9      :�����Bкғ����Y���@r8985:?/�:�d�:[B;Cm;�?&;#2;||:;!@;��C;��E;iG;��G;K(H;�ZH;]zH;+�H;ɤH;��H;U�H;��H;��H;Q�H;��H;��H;@�H;#�H;C�H;��H;t�H;��H;A�H;!�H;@�H;��H;��H;U�H;��H;��H;Y�H;��H;ƤH;.�H;]zH;�ZH;J(H;��G;kG;��E;��C;!@;{|:;#2;�?&;Bm;^B;�d�:C/�:D5:0r890��܇Y�ؓ��Jк���      ؚ��H���+J���X���b���-�����Hx�0��� :���:C��:ȯ;D ;H�.;��8;Q�?;�C;��E;'#G;��G;�1H;�aH;<�H;k�H;f�H;��H;��H;P�H;�H;(�H;,�H;��H;�H;~�H;0�H;��H;2�H;{�H;�H;��H;*�H;(�H;�H;P�H;��H;��H;h�H;e�H;<�H;�aH;�1H;��G;*#G;��E;��C;Q�?;��8;H�.;F ;ů;C��:���:� :0��Ix������-� �b��X��0J��I���      �B(�%�����_������˻	���b�D&����� �>���Y:��:�^;��;b�,;`8;W�?;��C;jF;�FG;=�G;�?H;kH;�H;��H;�H;E�H;��H;[�H;k�H;�H;r�H;��H;��H;z�H;��H;z�H;}�H;��H;n�H;�H;k�H;_�H;��H;F�H;�H;�H;�H;kH;�?H;9�G;�FG;lF;��C;U�?;`8;_�,;��;�^;��:��Y: �>�����A&�
�b�		���˻�����_����%�      �����x���#��@F{���]��E<����L�뻬���>d\�����[��3:��:Ѧ�:t[;[�,;��8;!@;�0D;p[F;{G;�
H;7PH;vH;֐H;/�H;�H;�H;Y�H;o�H;��H;��H;s�H;n�H;��H;��H;��H;j�H;p�H;��H;��H;o�H;\�H;�H;�H;.�H;АH;vH;4PH;�
H;{G;g[F;�0D;!@;��8;]�,;p[;˦�:��:�3:�[����>d\�����M�뻥���E<���]�BF{��#���x��      \������o�prμу��sv��J"��^N�����?ݻX^��G���Y���9��:˦�:��;F�.;w|:;�>A;��D; �F;��G;�)H;aH;�H;n�H;׬H;,�H;�H;.�H;T�H;��H;�H;M�H;��H;��H;��H;M�H;�H;��H;P�H;,�H;�H;-�H;׬H;k�H;��H;
aH;�)H;��G;�F;��D;�>A;u|:;A�.;��;æ�:��:��9�Y�H��X^���?ݻ���^N�J"��sv��Ӄ��qrμ�o����      ^n;�x\8��s/�=�!�z��_���jrμ��������E<�������N3�hHx���9��:�^;G ;#2;]�<;�B;��E;$5G;��G;)FH;vqH;��H;:�H;��H;D�H;��H;��H;��H;��H;�H;j�H; �H;m�H;�H;��H;��H;��H;��H;I�H;��H;;�H;��H;oqH;#FH;��G;(5G;��E;�B;_�<; 2;G ;�^;��:��9dHx��N3�������E<��������jrμ_���{��=�!��s/�x\8�      ���������Ȅ�jSt��Y�\n;�0O�n#���Oļ�����&R��_������N3���Y��3:��:˯;�?&;�G6;~X?;�D;$xF;��G;,!H;^H;}�H;�H;ƭH;;�H;��H;��H;��H;	�H;��H;L�H;�H;L�H;��H;�H;��H;��H;��H;>�H;ĭH;�H;~�H;{^H;&!H;��G;$xF;�D;sX?;�G6;�?&;ǯ;��:�3:��Y��N3������_��&R������Oļn#��0O�\n;��Y�kSt��Ȅ�����      �ѽ\νy�ý䳽:����L����d�q\8�v��ټiv����Y��_����D���[�|�Y:A��:Cm;�r-;�:;i�A;,oE;�"G;I�G;TGH;�sH;ݐH;��H;�H;#�H;�H;��H;u�H;z�H;"�H;��H;#�H;x�H;t�H;��H;�H;!�H;�H;��H;ݐH;sH;PGH;C�G;�"G;,oE;f�A;��:;�r-;Am;A��:��Y:�[�D������_���Y�jv��ټv��q\8���d��L��:���䳽y�ý\ν      �� ]�ӈ�p}���x�ý�u��˕���K�����o�jv���&R�!��Y^����� �>����:UB;5";e�4;��>;>D;��F;�G;�)H;`dH;k�H;�H;\�H;%�H;(�H;~�H;��H;�H;	�H;��H;	�H;�H;��H;z�H;&�H;"�H;a�H;	�H;k�H;^dH;�)H;�G;��F;=D;��>;Y�4;5";TB;���: �>����Z^��!���&R�jv���o�����K�˕���u��w�ý��p}�ӈ� ]�      �+X��T��nH��6��� �j��C�䳽�����mR����ټ�����E<��?ݻ>d\������ :�d�:��;$�,;s�:;V7B;��E;kLG;)H;USH;�{H;{�H;�H;�H;9�H;Q�H;�H;��H;��H;��H;��H;��H;�H;M�H;6�H;�H;�H;{�H;�{H;SSH;'H;gLG;��E;U7B;q�:;�,;��;�d�:� :����@d\��?ݻ�E<�����ټ����mR�����䳽C�j���� ��6��nH��T�      ఖ�����}���*|�LS\�� :����Z�l$�������K�v���Oļ����������J&����3/�:�^;��#;�G6;4�?;�D;E�F;��G;�?H;�pH;ڏH;q�H;�H;H�H;,�H;i�H;k�H;��H;v�H;��H;k�H;g�H;'�H;H�H;�H;t�H;ڏH;�pH;�?H;��G;B�F;��D;5�?;�G6;��#;�^;-/�:���I&������������Oļv���K�����l$���Z���� :�LS\��*|�}������      @�;9ɾ|㼾B�������Mw��nH�����Z�䳽˕��r\8�o#������^N�Q���b�8Ix� 5:ͮ�:)�;��0;]=;9�C;�[F;ϞG;�)H;�eH;n�H;�H;9�H;��H;�H;��H;$�H;��H;h�H;��H;&�H;��H;�H;~�H;7�H;&�H;p�H;�eH;�)H;ўG;�[F;8�C;]=;��0; �;ծ�:5:(Ix��b�Q��^N�����p#��r\8�˕��䳽�Z񽰯��nH��Mw�����B��|㼾9ɾ      /y��v�i���B�߾����A��?����nH���CὝu����d�0O�jrμJ"�����
	������q89L;�:Y�;�+;H|:;r7B;��E;�aG;jH;�ZH;a�H;'�H;��H;�H;C�H;A�H;�H;��H;o�H;��H; �H;@�H;A�H;�H;��H;-�H;b�H;�ZH;nH;�aG;��E;t7B;N|:;�+;R�;R;�:�q89���	�����J"��jrμ0O���d��u��C����nH�?���A������B�߾j����v�      �O/�pM+�X�����GW��9ɾA���Mw�� :�j��x�ý�L��\n;�_���tv���E<��˻��-�h��Vy�:�^;�%;v�7;n�@;5E;�"G;�G;1PH;�zH;��H;V�H;x�H;��H;��H;�H;��H;��H;��H;�H;��H;��H;x�H;Q�H;��H;�zH;4PH;�G;�"G;5E;o�@;w�7;�%;�^;\y�:�����-��˻�E<�tv��^���\n;��L��w�ýj��� :��Mw�A��9ɾGW�����X��pM+�      7�X�VvS�6E��O/��S�GW����������LS\��� ���:����Y�{��҃����]�����0�b�ȇY� �Y:��:\`;.�4;�?;4�D;��F;�G; FH;AuH;��H;��H;~�H;�H;��H;�H;�H;��H;�H;�H;��H;�H;~�H;��H;œH;CuH;FH;�G;��F;4�D;�?;.�4;Z`;��:$�Y:ȇY�+�b�������]�҃��{���Y�:����彑� �LS\���������GW���S��O/�6E�VvS�      � ����y�`�h���N��O/����B�߾B���*|��6�p}�䳽jSt�=�!�prμDF{��_��X��ܓ��$:��:�Z;�2;�O>;fD; �F;s�G;=H;�pH;��H;E�H;ȷH;��H;��H;Z�H;v�H;\�H;s�H;W�H;��H;��H;ɷH;B�H;��H;�pH;=H;w�G;,�F;eD;�O>;�2;�Z;��:<:�����X���_�CF{�prμ=�!�jSt�䳽p}��6��*|�B��B�߾����O/���N�`�h���y�      =v��b���W ��`�h�6E�W��j���|㼾}���nH�ӈ�y�ý�Ȅ��s/��o��#�����)J��:к	�9Jg�:�l;0;]=;ղC;ЀF;i�G;6H;mH;"�H;��H;|�H;��H;:�H;��H;�H;��H;��H;��H;9�H;��H;z�H;��H;)�H;mH;6H;n�G;݀F;ҲC;]=;0;�l;Dg�:8	�9>к(J������#���o��s/��Ȅ�y�ýӈ��nH�}��|㼾j���W��6E�`�h�W ��b���      |h��/���b�����y�VvS�pM+��v�9ɾ�����T� ]�\ν����y\8�����x��%�R�������9g-�:a�;��.;�<;�nC;�dF;�G;�1H;�jH;��H;��H;ɵH;f�H;��H;b�H;��H;��H;��H;`�H;��H;c�H;ǵH;��H;��H;�jH;�1H;�G;�dF;�nC;�<;��.;_�;[-�:8�9���R���%��x�����y\8�����\ν ]��T�����9ɾ�v�pM+�VvS���y�b���/���      EEb�`]��N��7����s� ���˾��)�j��!,�p���L��Cm�,��9,˼��x�^���1�� ���4�:b�:�;
�1;0,>;_�C;NwF;�G;i H;�>H;�hH;'�H;>�H;�H;�H;��H;�H;i�H;�H;��H;�H;�H;;�H;#�H;�hH;�>H;i H;�G;\wF;^�C;/,>;�1;�;`�:@�: ����1��^����x�9,˼,��Dm�L��p����!,�)�j�����˾s� �����7��N�`]�      `]�d�W��TI�v3��D�������Ǿv����f�8)�%��s;���Fi��k���Ǽ�[t�P�	�0Ȅ�.X����:���:��;$J2;LZ>;!	D;6F;4�G;�H;�?H;siH;��H;��H;O�H;�H;��H;3�H;��H;,�H;��H;�H;L�H;��H;��H;xiH;�?H;�H;7�G;BF; 	D;LZ>; J2;��;���:��:.X��/Ȅ�P�	��[t���Ǽ�k��Fi�s;��%��8)��f�v�����Ǿ�����D�v3��TI�d�W�      �N��TI���;�/�'�l��쾀���x󐾳Z��K ��s�A����&^���"����g����ڨu�!���2<:��:�
;1g3;��>;PBD;p�F;ڔG;gH;BH;YkH;)�H;��H;�H;��H;?�H;��H; �H;��H;>�H;��H;�H;��H;"�H;`kH;BH;eH;ޔG;}�F;PBD;��>;-g3;�
;��:�2<:!��ڨu������g��"����&^�A����s潥K ��Z�x󐾀�����l�/�'���;��TI�      �7�v3�/�'����s� ��{Ծ ���H���y�F�����ӽ���_�L�Jv��뮼TT����PV���=�4)i:f��:�z ;w$5;��?;�D;��F;�G;oH;aFH;pnH;^�H;H�H;H�H;��H;�H;.�H;��H;(�H;�H;��H;F�H;F�H;W�H;tnH;_FH;kH;�G;��F;�D;��?;r$5;�z ;`��:D)i:��=��PV���TT��뮼Jv�_�L�����ӽ���y�F�H��� ����{Ծs� ����/�'�v3�      ����D�l�s� �V�ݾj���V͓��f��>/�����'���섽P�6��t�w��a�:�,Tʻ�.�x۷�,t�:�;��$;|Y7;K�@;�	E;��F;&�G;�H;LH;�rH;��H;��H;��H;�H;�H;!�H;��H;�H;�H;�H;��H;��H;�H;�rH;LH;�H;'�G;��F;�	E;I�@;yY7;��$;�;6t�:�۷��.�,Tʻa�:�w���t�P�6��섽�'������>/��f�V͓�j���V�ݾs� �l��D�      s� ��������{Ծj���v���Z�x��SC��^��޽@���y�e�(��D�Ѽ&G������R������ܤ8���:�Y;>�);��9;��A;��E;yG;	�G;<!H;SH;�wH;G�H;V�H;�H;��H;H�H;S�H;��H;N�H;G�H;��H;�H;V�H;A�H;�wH;SH;:!H;�G;�G;��E;��A;��9;=�);�Y;���:�ܤ8����R�����%G��D�Ѽ(��x�e�@����޽�^��SC�Z�x�v���j����{Ծ�쾠���      ��˾��Ǿ���� ���V͓�Z�x���J��K �m���������?����뮼-�[�#���!3|��W��h�:)�:�';Y/;5g<;C;?F;�NG;��G;-H;7[H;�}H;��H;��H;��H;|�H;��H;��H;��H;��H;��H;|�H;��H;��H;��H;�}H;7[H;-H;��G;�NG;@F;}C;5g<;Y/;�';3�:`�:�W�� 3|�$���-�[��뮼���?������m����K ���J�Z�x�V͓� ���������Ǿ      ��v���x�H����f��SC��K �nn����Ž����Z��k�}ռ.X��cy-�1���|.����P�:x+�:u�;4;
�>;�D;�wF;��G;��G;�9H;#dH;P�H;|�H;/�H;E�H;��H;{�H;(�H;B�H;%�H;|�H;��H;A�H;+�H;w�H;V�H;#dH;�9H;��G;��G;�wF;�D;�>;4;q�;�+�:�P�:���|.�0���cy-�.X��}ռ�k��Z������Žnn���K ��SC��f�H���x�v���      (�j��f��Z�y�F��>/��^�m�����ŽF ���Fi��Q+�}t�oT��p�W�����1��<Ⱥ�W�9cP�:xY;{�(;��8;�A;�E;��F;2�G;mH;�FH;�mH;g�H;��H;�H;F�H;��H;]�H;��H;��H;��H;]�H;��H;A�H;�H;��H;k�H;�mH;�FH;lH;4�G;��F;�E;�A;��8;w�(;�Y;gP�:�W�9:Ⱥ�1�����o�W�oT��|t�Q+��Fi�F ����Žm����^��>/�y�F��Z��f�      �!,�8)��K ��������޽������Fi��0����鷼��x�����.��[�(� ���*i:j��:�;��0;0�<;hC;�E;�<G;��G;�$H;5TH;�wH;ĒH;�H;�H;U�H;�H;b�H;q�H;K�H;o�H;c�H;�H;S�H;�H;�H;ʒH;�wH;8TH;�$H;��G;�<G;~�E;mC;4�<;��0;$�;j��:�*i:��[�(��.�������x�鷼����0��Fi�������޽�������K �8)�      p���%��s��ӽ�'��@�������Z��Q+�����"��G��»0���׻ӕb�NW���X�9���:`;w*';�Y7;�#@;��D;ۖF;�G;��G;8H;�aH;ɁH;0�H;v�H;F�H;h�H;t�H;V�H;"�H;
�H;#�H;W�H;v�H;g�H;C�H;w�H;9�H;΁H;�aH;8H;��G;�G;ۖF; �D;�#@;�Y7;*';`;���:�X�9LW��ҕb���׻»0�G���"������Q+��Z����@����'���ӽ�s�%��      K��s;��A�������섽y�e��?��k�}t�鷼G���e7����Ȅ��0㺀�t�u�:�+�:f;e1;;�<;B�B;��E;�G;��G;+H;MJH;/oH;͋H;��H;�H;k�H;��H;��H;g�H;��H;��H;��H;g�H;��H;��H;g�H;�H;��H;֋H;2oH;MJH;,H;��G;�G; �E;H�B;>�<;p1;f;�+�:u�: �t��0�Ȅ���껆e7�G��鷼|t��k��?�x�e��섽���A���s;��      Dm��Fi��&^�`�L�O�6�(����}ռoT����x���0����������ط��n`:p�:�;�*;�8;�@;�D;>�F;�}G;u�G;g1H;�[H;?|H;��H;��H;V�H;��H;��H;[�H;e�H;��H;B�H;��H;d�H;[�H;��H;��H;Z�H;��H;��H;B|H;�[H;e1H;z�G;�}G;A�F;�D;��@; �8;�*;�;z�:�n`:�ط���
��������0���x�nT��}ռ��(��Q�6�`�L��&^��Fi�      +���k��Kv�}t�F�Ѽ�뮼-X��p�W������׻Ȅ�"��h���4<:E��:�Y;�t%;�$5;�Z>;�`C;��E;*G;=�G;�H;�GH;AlH;ňH;ўH;��H;��H;m�H;��H;��H;G�H;C�H;��H;B�H;F�H;��H;��H;i�H;��H;��H;ٞH;ǈH;BlH;�GH;�H;=�G;*G;��E;�`C;�Z>;�$5;~t%;�Y;C��:�4<:X����Ȅ���׻���n�W�-X���뮼D�Ѽ�t�Kv���k�      7,˼��Ǽ�"���뮼w��%G��-�[�ay-�����.��Еb��0� ٷ��4<:�L�:�\;h�!;�J2;{g<;&0B;	CE;�F; �G;��G;[4H;r\H;�{H;|�H;t�H;,�H;��H;�H;g�H;!�H;"�H;��H;~�H;��H;"�H;#�H;e�H;�H;��H;3�H;y�H;��H;�{H;o\H;_4H;��G;!�G;
�F;CE;10B;g<;�J2;n�!;�\;�L�:�4<:�ط��0�͕b��.�����ay-�-�[�$G��w���뮼�"����Ǽ      ��x��[t���g�RT�a�:�������.����1��Z�(�HW��@�t��n`:C��:�\;�z ;}�0;J;;�<A;�D;�wF;�cG;'�G;�!H;}MH;SoH;G�H;W�H;��H;b�H;6�H;��H;,�H;A�H;��H;j�H;��H;h�H;��H;A�H;)�H;��H;9�H;h�H;��H;Z�H;F�H;OoH;�MH;�!H;)�G;�cG;�wF;��D;�<A;F;;�0;�z ;�\;C��:�n`:@�t�DW��Y�(��1��-��� ������d�:�RT���g��[t�      [��N�	������*Tʻ�R��3|�w.�2Ⱥ ���X�9u�:z�:�Y;l�!;��0;Ε:;��@;�BD;^2F;S8G;��G;�H;<@H;�cH;��H;H�H;�H;�H;�H;b�H;��H;��H;?�H;��H;��H;W�H;��H;}�H;@�H;��H;��H;f�H;"�H;�H;�H;E�H;��H;�cH;>@H;�H;��G;V8G;f2F;�BD;��@;ѕ:;��0;p�!;�Y;v�:u�:�X�9��.Ⱥu.�3|��R��,Tʻ�����M�	�      �1��,Ȅ�ۨu��PV�{.�����W������W�9�*i:ġ�:�+�:
�;~t%;�J2;C;;��@;VD;�F;�G;Q�G;aH;S5H;RZH; xH;�H;��H;�H;�H;*�H;<�H;��H;��H;��H;�H;0�H;��H;.�H;�H;��H;��H;��H;@�H;2�H;�H;�H;��H;�H;xH;QZH;P5H;dH;T�G;G;�F;SD;��@;@;;�J2;|t%;�;�+�:Ρ�:�*i:X�9���W�����w.��PV�Ԩu�+Ȅ�      ����LX��!����=��۷� ޤ8��:�P�:iP�:j��:`;b;�*;�$5;g<;�<A;�BD;�F;�G;Q�G;:�G;s-H;�RH;(qH;��H;��H;P�H;�H;�H;��H;��H;��H;$�H;��H;q�H;h�H;��H;e�H;n�H;��H;!�H;��H;��H;��H;�H;�H;L�H;��H;��H;+qH;�RH;v-H;>�G;U�G;�G;�F;�BD;�<A;�g<;�$5;�*;f; `;j��:oP�:�P�:|�:`ݤ8�۷���=�!��LX��      �:��:�2<:t)i:"t�:���:E�:x+�:|Y;$�;�*';m1;�8;�Z>;10B;��D;c2F;G;S�G;��G;R)H;WNH;FlH;�H;4�H;S�H;m�H; �H;W�H;��H;	�H;��H; �H;.�H;��H;��H;��H;��H;��H;.�H; �H;��H;	�H;��H;U�H; �H;k�H;Q�H;8�H;�H;ClH;YNH;U)H;��G;V�G;G;c2F;��D;30B;�Z>;�8;o1;�*';%�;|Y;�+�:A�:Ň�:.t�:$)i:�2<:\�:      ��:���:���:J��:�;�Y;�';q�;z�(;��0;�Y7;7�<;�@;�`C;CE;�wF;S8G;[�G;<�G;P)H;�LH;�iH;�H;+�H;t�H;��H;��H;4�H;��H;��H;��H;,�H;��H;o�H;��H;{�H;��H;t�H;��H;n�H;��H;%�H;��H;��H;��H;4�H;��H;��H;x�H;(�H;�H;�iH;�LH;P)H;=�G;U�G;T8G;�wF;CE;�`C;��@;;�<;�Y7;��0;v�(;m�;�';�Y;�;J��:���:���:      �;��;�
;�z ;��$;>�);Y/;4;��8;6�<;�#@;B�B;�D;��E;	�F;�cG;��G;gH;v-H;YNH;�iH;�H;��H;��H;��H;��H;v�H;u�H;�H;��H;G�H;�H;�H;��H;��H;D�H;��H;?�H;��H;��H;�H; �H;H�H;��H;�H;s�H;q�H;��H;��H;~�H;~�H;�H;�iH;YNH;v-H;dH;��G;�cG;�F;��E;�D;H�B;�#@;4�<;��8;4;[/;6�);��$;�z ;�
;��;      !�1;"J2;*g3;�$5;uY7;��9;Gg<;�>;�A;qC;	�D;�E;B�F;*G;#�G;+�G;�H;X5H;�RH;BlH;�H;��H;��H;��H;Y�H;:�H;/�H;�H;��H;~�H;^�H;��H;[�H;��H;��H;�H;I�H;��H;�H;��H;Z�H;��H;a�H;}�H;��H;�H;,�H;;�H;\�H;��H;��H;��H;�H;BlH;�RH;S5H;�H;+�G;$�G;*G;D�F;�E;
�D;nC;�A;�>;Fg<;��9;�Y7;�$5;)g3;J2;      *,>;TZ>;��>;��?;B�@;��A;�C;�D;�E;��E;ݖF;�G;�}G;A�G;��G;�!H;?@H;YZH;*qH;�H;(�H;|�H;��H;�H;��H;��H;�H;��H;��H;��H;9�H;�H;~�H;x�H;=�H;��H;��H;��H;:�H;x�H;}�H;
�H;<�H;��H;��H;��H;�H;��H;��H;�H;��H;}�H;(�H;�H;'qH;RZH;>@H;�!H;��G;=�G;�}G;�G;��F;��E;�E;�D;�C;��A;M�@;��?;��>;JZ>;      ��C;	D;LBD;ߚD;�	E;��E;KF;�wF;��F;�<G;�G;��G;z�G;�H;a4H;�MH;�cH;xH;��H;=�H;|�H;��H;]�H;��H;�H;��H;��H;L�H;S�H;��H;��H;W�H;u�H;0�H;��H;;�H;>�H;5�H;��H;2�H;t�H;Q�H;��H;��H;P�H;J�H;��H;��H; �H;��H;\�H;��H;|�H;8�H;��H;xH;�cH;�MH;a4H;�H;|�G;��G;�G;�<G;��F;�wF;MF;��E;�	E;ښD;MBD;	D;      JwF;?F;u�F;��F;��F;�G;�NG;	�G;5�G;��G;��G;3H;i1H;�GH;s\H;VoH;��H;�H;��H;P�H;��H;��H;5�H;��H;��H;<�H;�H;�H;��H;v�H;�H;F�H;%�H;��H;g�H;��H;��H;��H;b�H;��H;&�H;@�H;�H;v�H;��H;
�H;�H;A�H;��H;��H;5�H;��H;��H;M�H;��H;�H;��H;UoH;p\H;�GH;h1H;3H;��G;��G;4�G;�G;�NG;yG;��F;��F;z�F;>F;      ��G;:�G;ڔG;�G;�G;�G;��G;��G;kH;�$H;8H;KJH;�[H;ClH;�{H;G�H;I�H;��H;P�H;m�H;��H;s�H;/�H;�H;��H;
�H;��H;U�H;>�H;��H;'�H;�H;��H;}�H;��H;��H;	�H;��H;��H;~�H;��H;��H;%�H;��H;:�H;T�H;��H;�H;��H;�H;/�H;t�H;��H;j�H;M�H;��H;I�H;H�H;�{H;?lH;�[H;PJH;8H;�$H;hH;��G;��G;��G;4�G;أG;ڔG;&�G;      g H;�H;aH;sH;�H;<!H;-H;�9H;�FH;>TH;�aH;6oH;A|H;ɈH;|�H;W�H;�H;�H;�H;��H;4�H;p�H;�H;��H;F�H;�H;T�H;L�H;��H;��H;��H;��H;n�H;��H;�H;W�H;Z�H;Q�H;�H;��H;l�H;��H;��H;��H;��H;K�H;P�H;
�H;J�H;��H;�H;o�H;3�H;��H;�H;�H;�H;Y�H;y�H;ɈH;A|H;7oH;�aH;>TH;�FH;�9H;-H;2!H;�H;pH;bH;�H;      �>H;u?H;BH;mFH;�KH;SH;>[H;"dH;�mH;�wH;ЁH;֋H;��H;՞H;v�H;��H;�H;�H;�H;W�H;��H;�H;��H;��H;N�H;{�H;6�H;��H;�H;��H;��H;b�H;��H;-�H;f�H;��H;��H;��H;e�H;.�H;��H;]�H;��H;��H;�H;��H;3�H;}�H;O�H;��H;��H;�H;��H;S�H;
�H;�H;�H;��H;u�H;ӞH;��H;ԋH;сH;�wH;�mH;"dH;;[H; SH;LH;mFH;BH;y?H;      �hH;jiH;ckH;gnH;�rH;�wH;�}H;P�H;k�H;ʒH;7�H;��H;��H;��H;/�H;b�H;!�H;*�H;��H;��H;��H;��H;w�H;��H;��H;m�H;��H;��H;��H;��H;h�H;��H;�H;t�H;��H;��H;��H;��H;��H;s�H;�H;��H;g�H;��H;��H;��H;��H;q�H;��H;��H;z�H;��H;��H;��H;��H;(�H;!�H;d�H;.�H;��H;��H;��H;9�H;̒H;k�H;T�H;�}H;�wH;�rH;jnH;dkH;iiH;      0�H;ԈH;0�H;a�H;��H;E�H;��H;}�H;��H;�H;}�H;�H;^�H;��H;��H;<�H;i�H;A�H;��H;�H;��H;G�H;[�H;7�H;��H;�H;$�H;��H;��H;n�H;��H;'�H;~�H;��H;��H;��H;��H;��H;��H;��H;��H;$�H;��H;i�H;��H;��H;"�H;�H;��H;7�H;a�H;F�H;��H;�H;��H;?�H;k�H;=�H;��H;��H;`�H;�H;~�H;�H;��H;��H;��H;=�H;��H;^�H;2�H;ԈH;      >�H;��H;��H;=�H;��H;L�H;��H;/�H;�H;�H;H�H;p�H;��H;t�H;�H;��H;��H;��H;��H; �H;/�H;�H;��H;�H;T�H;=�H;��H;��H;a�H;��H;!�H;t�H;��H;��H;��H;��H;�H;��H;��H;��H;��H;q�H;�H;��H;]�H;��H;��H;@�H;W�H;�H;��H;�H;*�H;��H;��H;��H;��H;��H;�H;q�H;��H;p�H;N�H;!�H;�H;3�H;��H;O�H;��H;@�H;��H;��H;      �H;Z�H;�H;G�H; �H;�H;��H;@�H;=�H;U�H;l�H;��H;��H;��H;i�H;0�H;��H;�H;(�H;�H;��H;�H;X�H;z�H;u�H;!�H;��H;r�H;��H;�H;}�H;��H;��H;��H;�H;�H;��H;�H;�H;��H;��H;��H;z�H;�H;��H;n�H;��H;#�H;x�H;z�H;^�H;�H;��H;�H;(�H;�H;��H;3�H;i�H;��H;��H;��H;o�H;X�H;A�H;A�H;��H;�H;�H;A�H;�H;Z�H;      �H;�H;��H;��H;��H;��H;��H;��H;��H;�H;��H;��H;b�H;��H;(�H;E�H;C�H;��H;��H;0�H;t�H;��H;��H;m�H;,�H;��H;v�H;��H;-�H;w�H;��H;��H;��H;��H;%�H;/�H;�H;.�H;$�H;��H;��H;��H;��H;s�H;(�H;��H;w�H;��H;0�H;m�H;��H;��H;o�H;,�H;��H;�H;I�H;G�H;(�H;��H;d�H;��H;��H;�H;��H;��H;��H;~�H;��H;��H;��H;�H;      ��H;��H;I�H;	�H;�H;=�H;��H;|�H;a�H;k�H;`�H;r�H;r�H;O�H;)�H;��H;��H;�H;p�H;��H;��H;��H;z�H;-�H;��H;Z�H;��H;�H;h�H;��H;��H;��H;�H;'�H;�H;$�H;C�H;%�H;�H;)�H;�H;��H;��H;��H;e�H;	�H;��H;]�H;��H;/�H;��H;��H;��H;��H;n�H;�H;��H;��H;*�H;Q�H;s�H;u�H;d�H;n�H;g�H;��H;��H;@�H;�H;�H;J�H;��H;       �H;0�H;��H;*�H;�H;G�H;��H;)�H;��H;w�H;*�H;��H;��H;I�H;��H;h�H;��H;,�H;g�H;��H;{�H;?�H;��H;��H;3�H;��H;��H;U�H;��H;��H;��H;��H;�H;2�H;'�H;�H;/�H;�H;'�H;6�H;�H;��H;��H;��H;��H;T�H;��H;��H;5�H;��H; �H;?�H;x�H;~�H;g�H;0�H;��H;m�H;��H;J�H;��H;��H;/�H;z�H;��H;.�H;��H;I�H;�H;$�H;��H;>�H;      o�H;��H;7�H;��H;��H;��H;��H;B�H;��H;O�H;�H;��H;N�H;�H;��H;��H;^�H;��H;��H;��H;��H;��H;E�H;��H;;�H;��H;�H;a�H;��H;��H;��H;�H;��H;�H;F�H;.�H;�H;/�H;C�H;�H;�H;�H;��H;��H;��H;\�H;�H;��H;>�H;��H;L�H;��H;��H;��H;��H;��H;a�H;��H;��H;�H;O�H;��H;�H;R�H;��H;G�H;��H;��H;��H;��H;7�H;��H;      �H;3�H;��H;(�H;�H;L�H;��H;)�H;��H;w�H;)�H;��H;��H;J�H;��H;h�H;��H;,�H;g�H;��H;}�H;@�H;��H;��H;3�H;��H;��H;U�H;��H;��H;��H;��H;�H;5�H;)�H;�H;/�H;�H;'�H;5�H;�H;��H;��H;��H;��H;T�H;��H;��H;4�H;��H; �H;=�H;x�H;~�H;g�H;0�H;��H;m�H;��H;H�H;��H;��H;/�H;w�H;��H;.�H;��H;I�H; �H;+�H;��H;:�H;      ��H;��H;C�H;�H;�H;;�H;��H;��H;a�H;k�H;`�H;r�H;p�H;Q�H;,�H;��H;��H;�H;p�H;��H;��H;��H;z�H;/�H;��H;X�H;��H;�H;f�H;��H;��H;��H;�H;(�H;	�H;%�H;C�H;%�H;	�H;)�H;�H;��H;��H;��H;e�H;	�H;��H;]�H;��H;-�H;�H;��H;��H;��H;n�H;�H;��H;��H;)�H;O�H;s�H;u�H;a�H;k�H;b�H;��H;��H;;�H;�H;�H;I�H;��H;      �H;�H;��H;��H;��H;��H;��H;��H;��H;�H;��H;��H;b�H;��H;*�H;G�H;F�H; �H;��H;/�H;r�H;��H;��H;p�H;/�H;��H;v�H;��H;-�H;w�H;��H;��H;��H;��H;'�H;.�H;�H;.�H;%�H;��H;��H;��H;��H;s�H;(�H;��H;w�H;��H;-�H;i�H;��H;��H;k�H;,�H;��H; �H;G�H;H�H;(�H;��H;b�H;��H;��H;�H;��H;��H;��H;��H;��H;��H;��H;
�H;      �H;^�H;�H;D�H;��H;�H;��H;D�H;?�H;W�H;l�H;��H;��H;��H;l�H;0�H;��H;�H;'�H;�H;��H;�H;W�H;{�H;x�H;�H;��H;p�H;��H;�H;z�H;��H;��H;��H;�H;�H;��H;�H;�H;��H;��H;��H;{�H;�H;��H;n�H;��H;"�H;u�H;w�H;`�H;�H;��H;�H;(�H; �H;��H;2�H;i�H;��H;��H;��H;l�H;U�H;A�H;D�H;��H;�H;�H;J�H;�H;X�H;      2�H;��H;��H;?�H;��H;\�H;��H;0�H;�H;�H;J�H;p�H;��H;r�H;�H;��H;��H;��H;��H;��H;0�H;�H;��H;�H;W�H;?�H;��H;��H;b�H;��H;�H;s�H;��H;��H;��H;��H;�H;��H;��H;��H;��H;s�H;�H;��H;^�H;��H;��H;A�H;T�H; �H;��H;�H;(�H;��H;��H;��H;��H;��H;�H;q�H;��H;p�H;H�H; �H;�H;2�H;��H;P�H;��H;@�H;��H;��H;      #�H;ӈH;0�H;]�H;��H;G�H;��H;~�H;��H;�H;~�H;�H;^�H;��H;��H;=�H;j�H;A�H;��H;	�H;��H;H�H;[�H;9�H;��H;�H;!�H;��H;��H;l�H;��H;&�H;�H;��H;��H;��H;��H;��H;��H;��H;��H;'�H;��H;k�H;��H;��H;!�H;�H;��H;3�H;b�H;H�H;��H;	�H;��H;?�H;m�H;=�H;��H;��H;^�H;�H;}�H;�H;��H;��H;��H;D�H;��H;g�H;6�H;шH;      �hH;miH;^kH;tnH;�rH;�wH;�}H;W�H;n�H;̒H;7�H;��H;��H;��H;0�H;d�H;!�H;*�H;��H;��H;��H;��H;v�H;��H;��H;m�H;��H;��H;��H;��H;g�H;��H;�H;t�H;��H;��H;��H;��H;��H;t�H;�H;��H;h�H;��H;��H;��H;��H;t�H;��H;��H;~�H;��H;��H;��H;��H;(�H;!�H;e�H;/�H;��H;��H;��H;9�H;̒H;k�H;W�H;�}H;�wH;�rH;xnH;hkH;iiH;      �>H;u?H;BH;kFH;�KH;SH;;[H;"dH;�mH;�wH;΁H;֋H;��H;֞H;y�H;��H;�H;�H;�H;T�H;��H;�H;��H;��H;O�H;x�H;2�H;��H;�H;��H;��H;a�H;��H;.�H;h�H;��H;��H;��H;f�H;.�H;��H;a�H;��H;��H;�H;��H;4�H;~�H;L�H;��H;��H;�H;��H;T�H;�H;�H;�H;��H;x�H;ӞH;��H;ӋH;ЁH;�wH;�mH;'dH;@[H;SH;�KH;kFH;BH;s?H;      t H;�H;WH;rH;~H;G!H;-H;�9H;�FH;>TH;�aH;6oH;B|H;ɈH;}�H;Y�H;�H;�H;�H;��H;4�H;r�H; �H;��H;I�H;�H;P�H;K�H;��H;��H;��H;��H;i�H;��H;�H;T�H;\�H;U�H;�H;��H;o�H;��H;��H;��H;��H;H�H;S�H;
�H;F�H;��H;�H;r�H;2�H;��H;�H;�H;�H;W�H;}�H;ǈH;A|H;6oH;�aH;>TH;�FH;�9H;-H;9!H;�H;pH;aH;�H;      �G;D�G;ՔG;�G;+�G;�G;��G;��G;lH;�$H;8H;PJH;�[H;AlH;�{H;G�H;I�H;��H;N�H;i�H;��H;t�H;*�H;�H;��H;�H;��H;T�H;=�H;��H;$�H;�H;��H;~�H;��H;��H;�H;��H;��H;~�H;��H;�H;(�H;��H;:�H;T�H;��H;�H;��H;�H;2�H;v�H;��H;m�H;N�H;��H;I�H;H�H;�{H;?lH;�[H;NJH;8H;�$H;iH;��G;��G;�G;2�G;�G;ؔG;/�G;      =wF;>F;}�F;��F;��F;�G;�NG;
�G;8�G;��G;��G;6H;k1H;�GH;r\H;VoH;��H;�H;��H;M�H;��H;��H;3�H;��H;��H;8�H;�H;�H;��H;u�H;�H;D�H;#�H;��H;e�H;��H;��H;��H;b�H;��H;&�H;D�H;�H;v�H;�H;
�H;�H;A�H;��H;��H;8�H;��H;��H;N�H;��H;�H;��H;VoH;u\H;�GH;i1H;3H;��G;��G;/�G;�G;�NG;{G;��F;��F;g�F;0F;      ~�C;	D;GBD;ܚD;�	E;��E;MF;�wF;��F;�<G;�G;��G;y�G;�H;b4H;�MH;�cH;xH;��H;9�H;{�H;��H;Z�H;��H; �H;��H;��H;J�H;S�H;��H;��H;W�H;r�H;0�H;��H;:�H;?�H;:�H;��H;3�H;u�H;W�H;��H;��H;P�H;I�H;��H;��H;�H;��H;`�H;��H;|�H;9�H;��H;xH;�cH;�MH;c4H;�H;|�G;��G;�G;�<G;��F;�wF;JF;��E;�	E;ښD;GBD;	D;      ,>;<Z>;��>;��?;;�@;��A;�C;�D;�E;�E;ߖF;�G;�}G;=�G;��G;�!H;>@H;XZH;(qH;�H;)�H;|�H;��H;�H;��H;��H;�H;��H;��H;��H;:�H;�H;~�H;w�H;:�H;��H;��H;��H;9�H;u�H;��H;�H;?�H;��H;��H;��H;�H;��H;��H;�H;��H;}�H;)�H;�H;*qH;TZH;?@H;�!H;��G;>�G;�}G;�G;ߖF;�E;�E;�D;�C;��A;R�@;��?;��>;$Z>;      �1;J2;g3;�$5;qY7;��9;Bg<;�>;�A;oC;�D;�E;A�F;*G;%�G;-�G;�H;X5H;�RH;AlH;�H;��H;��H;��H;\�H;3�H;,�H;�H;��H;x�H;`�H;��H;Z�H;��H;��H;�H;K�H;�H;�H;��H;[�H;��H;d�H;��H;��H;�H;2�H;;�H;Z�H;��H;��H;��H;�H;BlH;�RH;S5H;�H;+�G;'�G;*G;B�F;�E;�D;oC;�A;�>;@g<;��9;rY7;�$5;g3;J2;      �;��;�
;�z ;��$;C�);]/;	4;��8;2�<;�#@;I�B;�D;��E;�F;�cG;��G;gH;t-H;YNH;�iH;�H;��H;~�H;��H;��H;s�H;r�H;�H;��H;G�H;�H;�H;��H;��H;@�H;��H;C�H;��H;��H;�H;�H;K�H;��H;�H;u�H;w�H;��H;��H;��H;��H;�H;�iH;ZNH;v-H;dH;��G;�cG;�F;��E;�D;G�B;�#@;2�<;��8;4;V/;-�);��$;�z ;�
;��;      ��:��:���:^��:�;�Y;�';r�;z�(;��0;�Y7;:�<;�@;�`C;CE;�wF;S8G;X�G;=�G;P)H;�LH;�iH;�H;)�H;w�H;��H;��H;2�H;��H;��H;��H;*�H;��H;n�H;��H;w�H;��H;x�H;��H;k�H;��H;)�H;��H;��H;��H;4�H;��H;��H;u�H;+�H;�H;�iH;�LH;Q)H;=�G;U�G;T8G;�wF;CE;�`C;��@;:�<;�Y7;��0;z�(;u�;�';�Y;�;V��:��:���:      p�:��:�2<:x)i:&t�:Ç�:I�:�+�:�Y;%�;�*';m1;�8;�Z>;10B;��D;b2F;G;S�G;��G;U)H;YNH;ClH;�H;6�H;N�H;i�H;��H;X�H;��H;	�H;��H;�H;/�H;��H;��H;��H;��H;��H;+�H; �H;��H;�H;��H;X�H; �H;n�H;T�H;5�H;�H;ClH;WNH;T)H;��G;U�G;G;e2F;��D;30B;�Z>;�8;m1;�*';"�;~Y;�+�:A�:���:2t�:H)i:�2<:��:      ����HX��!����=��۷� ޤ8|�:�P�:kP�:j��:`;f;�*;�$5;�g<;�<A;�BD;�F;�G;R�G;>�G;t-H;�RH;'qH;��H;��H;L�H;�H;�H;��H;��H;��H;$�H;��H;q�H;g�H;��H;g�H;n�H;��H;"�H;��H;��H;��H;�H;�H;P�H;��H;��H;*qH;�RH;s-H;<�G;S�G;�G;�F;�BD;�<A;�g<;�$5;�*;f;`;d��:kP�:�P�:x�:�ݤ8�۷���=�!��@X��      �1��'Ȅ��u��PV�x.�����W��h�� X�9�*i:ơ�:�+�:
�;|t%;�J2;D;;��@;RD;�F; G;T�G;cH;U5H;QZH;xH;�H;��H;�H;�H;)�H;?�H;��H;��H;��H;�H;/�H;��H;/�H;�H;��H;��H;��H;?�H;0�H;�H;�H;��H;�H;�wH;QZH;T5H;aH;P�G;G;�F;RD;��@;C;;�J2;|t%;�;�+�:̡�:�*i:�W�9���W�����{.��PV��u�'Ȅ�      \��N�	������(Tʻ�R��3|�t.�6Ⱥ���X�9u�:v�:�Y;p�!;��0;Е:;��@;�BD;b2F;W8G;��G;�H;>@H;�cH;��H;E�H;�H;�H;�H;d�H;��H;��H;@�H;��H;��H;X�H;��H;}�H;?�H;��H;��H;d�H; �H;�H;�H;E�H;��H;�cH;<@H;�H;��G;P8G;c2F;�BD;��@;Е:;��0;p�!;�Y;v�:u�:�X�9��.Ⱥw.�!3|��R��.Tʻ�����L�	�      ��x��[t���g�QT�a�:�������,����1��Z�(�DW�� �t��n`:C��:�\;�z ;|�0;F;;�<A;��D;�wF;�cG;+�G;�!H;�MH;SoH;D�H;V�H;��H;b�H;9�H;��H;,�H;D�H;��H;h�H;��H;h�H;��H;>�H;(�H;��H;7�H;d�H;��H;W�H;D�H;OoH;zMH;�!H;+�G;�cG;�wF;��D;�<A;C;;�0;�z ;�\;C��:�n`:��t�HW��Z�(��1��.���"������d�:�RT���g��[t�      8,˼��Ǽ�"���뮼w��$G��-�[�ay-�����.��ϕb��0��ط��4<:�L�:�\;l�!;�J2;}g<;*0B;CE;	�F;'�G;��G;_4H;s\H;�{H;|�H;x�H;,�H;��H;�H;g�H;$�H;#�H;��H;|�H;��H; �H;!�H;d�H;�H;��H;.�H;x�H;z�H;�{H;l\H;X4H;��G;$�G;	�F;CE;-0B;{g<;�J2;l�!;�\;�L�:�4<: ٷ��0�Еb��.�����ay-�-�[�%G��w���뮼�"����Ǽ      +���k��Kv�~t�D�Ѽ�뮼-X��o�W������׻Ȅ� ��X���4<:G��:�Y;|t%;�$5;�Z>;�`C;��E;*G;@�G;�H;�GH;AlH;ňH;՞H;��H;��H;m�H;��H;��H;G�H;A�H;��H;C�H;C�H;��H;��H;i�H;��H;��H;ӞH;ÈH;>lH;�GH;�H;>�G;*G;��E;�`C;�Z>;�$5;|t%;�Y;?��:�4<:`��!��Ȅ���׻���o�W�-X���뮼E�Ѽ�t�Kv���k�      Dm��Fi��&^�`�L�O�6�(����}ռoT����x���0����
������ط��n`:t�:�;�*;�8;��@;�D;D�F;�}G;y�G;h1H;�[H;?|H;��H;��H;Y�H;��H;��H;]�H;e�H;��H;A�H;��H;b�H;Z�H;��H;��H;V�H;��H;��H;?|H;�[H;a1H;s�G;�}G;D�F;�D;�@;�8;�*;
�;t�:�n`:�ط�����������0���x�oT��}ռ��(��Q�6�`�L��&^��Fi�      L��s;��A�������섽x�e��?��k�}t�鷼G���e7����Ȅ��0���t�u�:�+�:f;l1;A�<;E�B;�E;�G;��G;-H;KJH;-oH;ҋH;��H;�H;i�H;��H;��H;g�H;��H;��H;��H;d�H;��H;��H;g�H;�H;��H;ӋH;-oH;JJH;)H;��G;�G;�E;D�B;7�<;m1;d;�+�:u�:��t��0�Ȅ���껆e7�G��鷼|t��k��?�x�e��섽���A���r;��      o���%��s��ӽ�'��@�������Z��Q+�����"��G��»0���׻ҕb�LW���X�9���:`;{*';�Y7;�#@;�D;ۖF;�G;��G;8H;�aH;ˁH;2�H;y�H;F�H;h�H;v�H;T�H;"�H;
�H;"�H;T�H;u�H;e�H;C�H;v�H;6�H;́H;�aH;8H;��G;�G;ܖF;�D;�#@;�Y7;|*';`;���:�X�9PW��ԕb���׻û0�G���"������Q+��Z����@����'���ӽ�s�%��      �!,�8)��K ��������޽������Fi��0����鷼��x�����.��[�(����*i:f��:!�;��0;2�<;mC;�E;�<G;��G;�$H;4TH;�wH;ŒH;�H;�H;U�H;�H;b�H;m�H;K�H;m�H;`�H;�H;S�H;�H;�H;ȒH;�wH;5TH;�$H;��G;�<G;~�E;nC;.�<;�0;$�;b��:�*i:��\�(��.�������x�鷼����0��Fi�������޽�������K �8)�      (�j��f��Z�y�F��>/��^�m�����ŽF ���Fi��Q+�|t�oT��p�W�����1��<Ⱥ�W�9cP�:zY;{�(;��8;�A;�E;��F;2�G;lH;�FH;�mH;h�H;��H;�H;F�H;��H;[�H;��H;��H;��H;[�H;��H;A�H;�H;��H;j�H;�mH;�FH;mH;2�G;��F;�E;�A;��8;t�(;�Y;]P�:�W�9<Ⱥ�1�����p�W�oT��|t�Q+��Fi�F ����Žm����^��>/�y�F��Z��f�      ��v���x�H����f��SC��K �nn����Ž����Z��k�}ռ.X��cy-�0���|.����P�:z+�:x�;4;�>;�D;�wF;��G;��G;�9H;"dH;P�H;}�H;/�H;E�H;��H;{�H;%�H;A�H;%�H;{�H;��H;B�H;,�H;|�H;W�H;%dH;�9H;��G;��G;�wF;�D;�>;4;p�;�+�:�P�:���z.�2���cy-�.X�� }ռ�k��Z������Žnn���K ��SC��f�H���x�v���      ��˾��Ǿ���� ���V͓�Z�x���J��K �m���������?����뮼.�[�#��� 3|��W��\�:-�:�';Z/;5g<;C;@F;�NG;��G;-H;7[H;�}H;��H;��H;��H;|�H;��H;��H;��H;��H;��H;|�H;��H;��H;��H;�}H;:[H;-H;��G;�NG;?F;�C;9g<;W/;�';3�:X�:�W�� 3|�$���-�[��뮼���?������m����K ���J�Z�x�V͓� ���������Ǿ      s� ��������{Ծj���v���Z�x��SC��^��޽@���y�e�(��D�Ѽ&G������R������ܤ8���:�Y;;�);��9;��A;��E;yG;�G;<!H;SH;�wH;H�H;W�H;�H;��H;G�H;P�H;��H;P�H;G�H;��H;�H;W�H;D�H;�wH;SH;=!H;	�G;�G;��E;��A;��9;:�);�Y;���:`ܤ8����R�����%G��D�Ѽ(��y�e�@����޽�^��SC�Z�x�v���j����{Ծ�쾠���      ����D�l�s� �V�ݾj���V͓��f��>/�����'���섽P�6��t�w��a�:�,Tʻ�.��۷�.t�:�;��$;{Y7;I�@;�	E;��F;#�G;�H;LH;�rH;��H;��H;��H;�H;��H;!�H;��H;�H;�H;�H;��H;��H;��H;�rH;LH;�H;*�G;��F;�	E;K�@;yY7;��$;�;4t�:�۷��.�-Tʻa�:�w���t�P�6��섽�'������>/��f�V͓�j���V�ݾs� �l��D�      �7�v3�/�'����s� ��{Ծ ���H���y�F�����ӽ���^�L�Kv��뮼TT����PV���=�<)i:l��:�z ;t$5;��?;�D;��F;�G;lH;aFH;nnH;`�H;H�H;G�H;��H;�H;-�H;��H;(�H;�H;��H;G�H;H�H;]�H;xnH;aFH;nH;�G;��F;�D;��?;s$5;�z ;`��:L)i:��=��PV���ST��뮼Kv�_�L�����ӽ���z�F�H��� ����{Ծs� ����/�'�v3�      �N��TI���;�/�'�l��쾀���x󐾳Z��K ��s�A����&^���"����g����ۨu�!���2<:��:�
;0g3;��>;PBD;n�F;ڔG;eH;BH;ZkH;+�H;��H;�H;��H;>�H;��H;�H;��H;>�H;��H;�H;��H;'�H;`kH;BH;gH;ߔG;}�F;PBD;��>;+g3;�
;��:�2<:
!��ڨu������g��"����&^�A����s潥K ��Z�x󐾀�����l�/�'���;��TI�      `]�d�W��TI�v3��D�������Ǿv����f�8)�%��s;���Fi��k���Ǽ�[t�P�	�0Ȅ�.X����:���:��;$J2;LZ>;!	D;4F;4�G;�H;�?H;siH;��H;��H;O�H;�H;��H;1�H;��H;,�H;��H;�H;L�H;��H;��H;ziH;�?H;�H;8�G;DF;	D;LZ>; J2;��;���:��:0X��/Ȅ�P�	��[t���Ǽ�k��Fi�s;��%��8)��f�v�����Ǿ�����D�v3��TI�d�W�      1�$��� ����#��?��'�þ�*��1Dx���=�����Pν���$'K��c� ��s�V����E^���S�Xw[:���:
e;!�4;=`?;�mD;M�F;HvG;�G;9H;^OH;�sH;��H;x�H;|�H;�H;P�H;!�H;K�H;�H;|�H;w�H;��H;�sH;hOH;7H;�G;LvG;Y�F;�mD;:`?;�4;e;���:hw[:��S�E^����r�V� ���c�$'K�����Pν�����=�1Dx��*��(�þ?��#������� �      �� ����R��O��/������0��4�s�׀:�g9��ʽ1Z����G��8�.���5S����	0X���D�FBd:�B�:� ;��4;È?;�~D;�F;	yG;��G;J H;'PH;tH;�H;ʢH;ðH;(�H;n�H;1�H;j�H;(�H;°H;ȢH; �H;tH;.PH;I H;��G;yG;�F;�~D;��?;��4;� ;�B�:ZBd:��D�0X���껰5S�.���8���G�1Z���ʽg9�׀:�4�s��0�����/��O��R�����      ���R��8�
������Yؾ���ޥ����f���0�Z[�N8��ϐ���>�����LȤ��6H�f�ܻrF�����}:���:\";&�5;��?;O�D;��F;�G;��G;,#H;]RH;�uH;C�H;��H;s�H;��H;�H;��H;�H;��H;q�H;��H;B�H;�uH;dRH;*#H;��G;�G;��F;M�D;��?;�5;X";���:��}:���rF�g�ܻ�6H�KȤ������>�ϐ��N8��Z[���0���f�ޥ������Yؾ����8�
�Q��      #��O������>I�(�þ�R��;���tS��Q"��s������}��0��켊�����6�K�ƻB}*�X�����:tx;R%;�l7;ҳ@;��D;��F;��G;�G;�'H;�UH;ZxH;K�H;C�H;��H;��H;��H;u�H;��H;��H;��H;@�H;H�H;TxH;�UH;�'H;|�G;��G;��F;��D;ҳ@;�l7;N%;sx;��:`���B}*�L�ƻ��6��������0���}�����s��Q"�tS�;����R��(�þ>Iᾣ���O��      ?��/�待Yؾ(�þĪ�|쏾�k�׀:�~�{�ؽ�����c�^y���Ҽ����F� �o�4�� (71�:��
;��(;y_9;��A;a\E;g�F;��G;��G;.H;�ZH;�{H;�H;G�H;M�H;�H;��H;t�H;��H;�H;M�H;D�H;�H;�{H;�ZH;.H;��G;��G;o�F;a\E;��A;s_9;��(;��
;;�: (74��o�F� �������Ҽ^y��c�����|�ؽ~�׀:��k�|쏾Ī�(�þ�Yؾ/��      '�þ��� ����R��|쏾5�s��H�����������ΐ����D��c�����?�f�V,�����P�� �9���:�;j-;E�;;n�B;��E;TG;��G;��G;|6H;�`H;T�H;I�H;ҩH;K�H;��H;O�H;��H;K�H;��H;H�H;ΩH;H�H;Q�H;�`H;{6H;��G;��G;\G;��E;k�B;B�;;j-;�;���: �9�P�����V,�>�f������c���D�ΐ�������������H�5�s�|쏾�R�� ������      �*���0��ޥ��;����k��H��#%�Z[��Pνt��a�f�3/%���伇���w�=��?ػ�FL���D�D�R:��:,�;,2;��=;��C;_0F;@GG;��G;H;�?H;�gH;��H;)�H;��H;��H;}�H;��H;p�H;��H;}�H;��H;��H;&�H;~�H;�gH;�?H;H;��G;FGG;a0F;��C;��=;,2;(�;��:@�R:��D��FL��?ػw�=��������3/%�a�f�t���PνZ[��#%��H��k�;���ޥ���0��      0Dx�4�s���f�tS�׀:����Z[��7ս�榽��}���;��8�V�����r����@G����@ά���:�;�}$;��6;��?;�D;��F;�pG;��G;�H;JH;;oH;9�H;s�H;��H;3�H;��H;��H;#�H;��H;��H;4�H;��H;o�H;4�H;BoH; JH;�H;��G;�pG;ÔF;�D;��?;��6;�}$;�;��:@ά���@G�������r�V����8���;���}��榽�7սZ[����׀:�tS���f�4�s�      ��=�ր:���0��Q"�~������Pν�榽@����G�2����Ҽ ��KE:�B�ܻ�D^�ʸ��<i:-��:�;2|,;��:;D�A;;iE;��F;�G;z�G;�(H;-UH;xwH;l�H;�H;��H;�H;��H;��H;�H;��H;��H;�H;��H;�H;j�H;}wH;1UH;�(H;{�G;�G;��F;8iE;G�A;��:;0|,;�;3��:8i:ʸ���D^�@�ܻKE:� ����Ҽ2����G�@���榽�Pν����~��Q"���0�ր:�      ���g9�Z[��s�{�ؽ���t����}���G������2c��Y�V�H,��*���������:��:I ;\�3;�0>;��C;�F;�8G;$�G;eH;�7H;�`H;�H;�H;��H;H�H;��H;E�H;��H;�H;��H;E�H;��H;B�H;�H;�H;�H;�`H;�7H;fH;$�G;�8G;�F;��C;�0>;Y�3;P ;��:�:p������*��H,�Y�V�1c���������G���}�t�����|�ؽ�s�Z[�g9�      �Pν�ʽO8���������ϐ��b�f���;�2�����DȤ�6�f�,��Rߵ�_o5� �D��-:4��:�>;�+;�_9;�A;^�D;�F;�vG;��G;H;qGH;VlH;��H;��H;��H;)�H;��H;��H;�H;!�H;�H;��H;��H;(�H;�H;��H;ÈH;[lH;tGH;H;��G;�vG;�F;b�D;�A;�_9;�+;�>;2��:�-:��D�^o5�Pߵ�+��5�f�CȤ����2����;�b�f�ΐ���������O8���ʽ      ���1Z��ϐ����}��c���D�2/%��8���Ҽ2c��5�f�����ƻ�/X�n���H��9��:3�;�";��3;6>;:YC;m�E;�G;�G;_�G;�,H;�VH;xH;��H;+�H;�H;�H;��H;.�H;B�H;,�H;A�H;.�H;��H;�H;�H;.�H;��H;xH; WH;�,H;^�G;�G;�G;t�E;AYC;8>;��3;�";3�;��:H��9j����/X��ƻ���4�f�2c����Ҽ�8�3/%���D��c���}�ϐ��1Z��      $'K���G��>��0�]y��c����U��� ��Y�V�+���ƻ�od���º r(7y4�:���:��;�P.;ʡ:;zA;%�D;¨F;HnG;4�G;�H;�@H; fH;Y�H;)�H;��H;ѸH;��H;��H;��H;z�H;5�H;x�H;��H;��H;��H;͸H;��H;0�H;^�H;!fH;�@H;�H;9�G;HnG;ŨF;*�D;zA;֡:;�P.;��;���:}4�: u(7��º�od��ƻ+��Y�V� ��U�����伖c�^y��0��>���G�      �c��8���������Ҽ����������r�KE:�G,�Oߵ��/X���º Ȭ�D�}:� �:�;A�);m7;�?;��C;F;Q)G;�G;A�G;�)H;�SH;�tH;X�H;x�H;�H;��H;��H;��H;�H;��H;I�H;��H;�H;��H;��H;��H;�H;��H;b�H;�tH;�SH;�)H;F�G;
�G;V)G;F;��C;�?;!m7;?�);�;� �:L�}:�Ǭ���º�/X�Nߵ�G,�IE:���r�����������Ҽ�켸����8�      ��.��LȤ���������>�f�w�=����B�ܻ�*��[o5�z��� r(7H�}:�n�:#�;�>&;��4;��=;��B;�E;�F;��G;��G;'H;}AH;�eH;7�H;͘H;U�H;ַH;d�H;�H;��H;h�H;��H;M�H;��H;g�H;��H;�H;`�H;ڷH;[�H;ԘH;=�H;�eH;xAH;+H;��G;��G;�F;�E;��B;��=;��4;�>&;"�;�n�:P�}: t(7p���Xo5��*��>�ܻ���w�=�<�f� �������LȤ�.��      m�V��5S��6H���6�F� �W,��?ػ=G���D^������D�8��9u4�:� �:"�;�%;��3;�<;OB;�E;��F;�XG;��G;A H;d0H;HWH;UvH;�H;w�H;��H;��H;��H;l�H;K�H;��H;��H;5�H;��H;��H;K�H;i�H;��H;��H;��H;{�H;�H;VvH;BWH;h0H;A H;��G;�XG;��F;�E;RB;�<;��3;�%;%�;� �:s4�:H��9��D�����D^�;G���?ػT,�I� ���6��6H��5S�      ��ﻲ��l�ܻN�ƻl󩻾���FL���ĸ����(�-:��:���:�;�>&;��3;K9<;�A;԰D;:ZF;5G;��G;��G;e!H;(JH;*kH;��H;��H;^�H;��H;��H;��H;��H;��H;��H;b�H;��H;^�H;��H;��H;��H;��H;��H;��H;c�H;��H;��H;&kH;,JH;f!H;��G;��G;5G;BZF;װD;
�A;N9<;��3;�>&;�;���:��:4�-:���������FL����o�Q�ƻq�ܻ���      E^�0X�rF�9}*�)���P����D��ͬ�@i:��::��:,�;��;>�);��4;�<;�A;�D;o9F;�G;h�G;?�G;8H;?H;UaH;}H;x�H;q�H;��H;ݾH;��H;_�H;|�H;�H;��H;%�H;��H;"�H;��H;�H;x�H;[�H;��H;�H;��H;q�H;v�H;}H;ZaH;?H;4H;@�G;k�G;�G;p9F;�D;	�A;�<;��4;>�);��;/�;D��:��:Pi:`ͬ���D��P��&��B}*�rF�0X�      h�S���D����@��� (7P�9h�R:��:3��:��:�>;�";�P.; m7;��=;QB;԰D;w9F;G;�G;N�G;�H;�6H;eYH;�uH;�H;�H;��H;��H;��H;�H;��H;�H;5�H;^�H;��H;��H;��H;\�H;4�H;�H;��H;�H;��H;��H;��H;�H;�H;�uH;fYH;�6H;�H;Q�G;�G;G;p9F;ذD;LB;��=; m7;�P.;�";�>;��:7��:��:d�R:(�9 (7���������D�      Lw[:6Bd:�}:��:%�:���:��:�;�;P ;�+;��3;ҡ:;�?;��B;�E;AZF;�G;�G;i�G;:H;N1H;�SH;[pH;ӇH;D�H;�H;v�H;��H;��H;��H;��H;o�H;�H;��H;�H;Y�H;�H;��H;�H;n�H;��H;��H;��H;��H;x�H;ߪH;A�H;ׇH;]pH;�SH;P1H;=H;k�G;�G;�G;?ZF;�E;��B;
�?;ҡ:;��3;�+;P ;�;�;��:˳�:1�:��:��}:�Ad:      ��:�B�:���:dx;z�
;�;)�;�}$;.|,;[�3;�_9;1>;zA;��C;�E;��F;5G;q�G;P�G;8H;�/H;�PH;�lH;C�H;��H;��H;i�H;��H;��H;�H;Y�H;��H;��H;��H;i�H;I�H;��H;A�H;g�H;��H;��H;��H;\�H;�H;��H;��H;e�H;��H;��H;B�H;�lH;�PH;�/H;8H;Q�G;k�G;5G;��F;�E;��C;zA;6>;�_9;[�3;,|,;�}$;-�;�;��
;dx;���:zB�:      �d; ;f";\%;��(;j-;*2;��6;��:;�0>;�A;:YC;)�D;F;�F;�XG;��G;E�G;�H;P1H;�PH;�kH;p�H;w�H;-�H;(�H;ӼH;��H;��H;	�H;j�H;��H;s�H;m�H;��H;^�H;��H;X�H;��H;m�H;r�H;��H;j�H;	�H;��H;�H;μH;)�H;1�H;v�H;i�H;�kH;�PH;N1H;�H;@�G;��G;�XG;�F;F;)�D;?YC;�A;�0>;��:;��6;.2;j-;��(;P%;[";� ;      7�4;��4;�5;�l7;r_9;M�;;��=;�?;O�A;ƚC;j�D;t�E;ƨF;[)G;��G;��G;��G;?H;�6H;�SH;�lH;n�H;��H;�H;��H;K�H; �H;/�H;��H;~�H;�H;��H;/�H;��H;��H;_�H;��H;Z�H;��H;��H;/�H;��H;�H;{�H;��H;/�H;�H;L�H;��H;�H;��H;n�H;�lH;�SH;�6H;8H;��G;��G;��G;V)G;ƨF;x�E;l�D;C;N�A;�?;��=;I�;;�_9;�l7;�5;��4;      ;`?;ʈ?;��?;̳@;��A;o�B;��C;�D;3iE;�F;�F;�G;HnG;�G;��G;D H;f!H;?H;fYH;WpH;A�H;q�H;�H;?�H;��H;"�H;@�H;�H;��H;p�H;P�H;��H;��H;��H;��H;:�H;K�H;3�H;��H;��H;��H;��H;S�H;n�H;��H;�H;:�H;#�H;��H;;�H;��H;s�H;?�H;VpH;cYH;?H;e!H;D H;��G;
�G;EnG;�G; �F;�F;8iE;�D;��C;^�B;��A;ɳ@;��?;��?;      �mD;�~D;I�D;��D;Z\E;��E;l0F;��F;��F;�8G;�vG;�G;;�G;L�G;-H;l0H;2JH;baH;�uH;ۇH;��H;1�H;��H;��H;��H;��H;g�H;�H;��H;��H;[�H;>�H;��H;��H;��H;��H;(�H;��H;��H;��H;��H;9�H;\�H;��H;��H;�H;`�H;��H;��H;��H;��H;1�H;��H;ׇH;�uH;^aH;2JH;n0H;-H;H�G;;�G;�G;�vG;�8G;��F;ÔF;m0F;��E;f\E;��D;L�D;�~D;      D�F;�F;��F;��F;e�F;_G;JGG;�pG;�G;0�G;��G;e�G;�H;*H;}AH;KWH;,kH;}H;�H;>�H;��H;$�H;G�H;!�H;��H;,�H;��H;|�H;��H;�H;�H;��H;��H;��H;9�H;��H;��H;��H;6�H;��H;��H;��H;
�H;�H;��H;{�H;��H;/�H;��H;�H;G�H;$�H;��H;=�H;�H;}H;,kH;HWH;{AH;�)H;�H;e�G;��G;-�G;�G;�pG;JGG;TG;y�F;��F;��F;�F;      ]vG;yG;�G;��G;��G;��G;��G;��G;z�G;hH;H;�,H;�@H;�SH;�eH;XvH;��H;|�H;�H;ߪH;l�H;мH;�H;@�H;d�H;��H;a�H;[�H;��H;��H;]�H;��H;��H;>�H;��H;%�H;"�H;�H;��H;A�H;��H;��H;]�H;��H;��H;X�H;Z�H;��H;g�H;<�H;�H;мH;l�H;ܪH;�H;u�H;��H;YvH;�eH;�SH;�@H;�,H;H;fH;x�G;��G;��G;��G;ĝG;y�G;�G;�xG;      �G;��G;��G;��G;��G;��G;-H;�H;�(H;�7H;uGH;WH; fH;�tH;7�H;�H;��H;q�H;��H;t�H;��H;}�H;)�H;�H;�H;{�H;[�H;��H;��H;b�H;��H;��H;S�H;��H;M�H;��H;��H;��H;L�H;��H;V�H;��H;��H;b�H;��H;��H;T�H;{�H;�H;��H;,�H;{�H;��H;r�H;��H;m�H;��H;�H;7�H;�tH; fH;WH;xGH;�7H;�(H;�H;-H;|�G;��G;�G;��G;��G;      4H;? H;&#H;�'H;q.H;�6H;�?H;JH;*UH;�`H;]lH;xH;]�H;]�H;јH;{�H;e�H;��H;��H;��H;��H;��H;��H;��H;��H;��H;��H;��H;0�H;��H;��H;N�H;��H;r�H;��H;��H;��H;��H;��H;s�H;��H;H�H;��H;��H;0�H;��H;��H;��H;��H;��H;��H;~�H;��H;��H;��H;��H;e�H;|�H;јH;\�H;\�H;xH;^lH;�`H;*UH;JH;�?H;{6H;{.H;�'H;(#H;C H;      ^OH; PH;gRH;�UH;�ZH;�`H;�gH;;oH;|wH;
�H;ÈH;��H;/�H;��H;V�H;��H;��H;ݾH;��H;��H;�H;�H;v�H;i�H;��H;�H;��H;b�H;��H;�H;I�H;��H;d�H;��H;��H;�H;2�H;�H;��H;��H;e�H;��H;G�H;~�H;��H;a�H;��H;�H;��H;g�H;z�H;�H;�H;��H;��H;ܾH;��H;��H;U�H;�H;/�H;��H;ÈH;�H;{wH;AoH;�gH;�`H;�ZH;�UH;jRH;PH;      �sH;)tH;�uH;[xH;�{H;T�H;��H;7�H;o�H;�H;��H;5�H;��H;��H;޷H;��H;��H;��H; �H;��H;^�H;j�H;�H;O�H;X�H;
�H;]�H;��H;��H;N�H;��H;k�H;��H;�H;W�H;b�H;Z�H;^�H;T�H;�H;��H;g�H;��H;K�H;��H;��H;X�H;�H;\�H;N�H;�H;i�H;\�H;��H;�H;��H;��H;��H;޷H;��H;��H;6�H;��H;�H;p�H;;�H;��H;L�H;�{H;ZxH;�uH;*tH;      ��H;�H;B�H;@�H;�H;>�H;0�H;s�H;$�H;��H;��H;�H;׸H;��H;d�H;��H;��H;b�H;��H;��H;��H;��H;��H;��H;;�H;��H;��H;��H;K�H;��H;d�H;��H;�H;X�H;��H;~�H;��H;~�H;�H;Z�H;�H;��H;b�H;��H;I�H;��H;��H;��H;>�H;��H;��H;��H;��H;��H;��H;c�H;��H;��H;d�H;��H;ָH;�H;��H;��H;$�H;w�H;5�H;A�H;�H;C�H;J�H;�H;      |�H;֢H;ȣH;B�H;L�H;ͩH;��H;��H;��H;I�H;0�H;�H;��H;��H; �H;q�H;��H;�H;�H;u�H;��H;u�H;+�H;��H;��H;��H;��H;Y�H;��H;k�H;��H;�H;P�H;��H;��H;��H;��H;��H;��H;��H;Q�H;�H;��H;e�H;��H;W�H;��H;��H;��H;��H;2�H;s�H;��H;p�H;�H;�H;��H;s�H;!�H;��H;��H;�H;0�H;K�H;��H;��H;��H;ƩH;P�H;=�H;ԣH;֢H;      w�H;��H;t�H;��H;O�H;@�H;��H;7�H;�H;��H;��H;��H;��H;��H;��H;R�H;��H;�H;8�H;#�H;��H;k�H;��H;��H;��H;��H;:�H;��H;o�H;��H;�H;X�H;��H;��H;��H;��H;��H;��H;��H;��H;��H;X�H;�H;��H;l�H;��H;;�H;��H;��H;��H;��H;k�H;��H;�H;6�H;�H;��H;R�H;��H;��H;��H;��H;��H;��H;��H;;�H;��H;?�H;W�H;��H;}�H;ɰH;      �H;9�H;κH;��H;�H;��H;��H;��H;��H;N�H;��H;8�H;��H;�H;o�H;��H;��H;��H;]�H;��H;k�H;��H;��H;��H;��H;/�H;��H;M�H;��H;�H;S�H;��H;��H;��H;��H;��H;��H;��H;��H;��H;��H;��H;P�H;��H;��H;J�H;��H;0�H;��H;��H;��H;��H;g�H;��H;\�H;��H;��H;��H;o�H;�H;��H;:�H;��H;O�H;��H;��H;��H;��H;�H;��H;ϺH;?�H;      K�H;m�H;�H;��H;��H;B�H;��H;��H;��H;��H;�H;H�H;~�H;��H;��H;��H;b�H;"�H;��H;�H;K�H;Z�H;U�H;(�H;��H;��H;�H;��H;��H;#�H;_�H;��H;��H;��H;��H;��H;��H;��H;��H;��H;��H;��H;^�H;�H;��H;��H; �H;��H;��H;)�H;\�H;X�H;G�H;�H;��H;%�H;e�H;��H;��H;��H;�H;H�H;�H;��H;��H;��H;�H;G�H;��H;��H;�H;{�H;      (�H;/�H;��H;r�H;o�H;��H;w�H;%�H;�H;�H;0�H;;�H;@�H;W�H;V�H;;�H;��H;��H;��H;_�H;��H;��H;��H;@�H;&�H;��H;�H;��H;��H;<�H;W�H;��H;��H;��H;��H;��H;��H;��H;��H;��H;��H;��H;X�H;6�H;��H;��H; �H;��H;&�H;A�H;��H;��H;��H;Y�H;��H;��H;��H;>�H;V�H;W�H;A�H;:�H;2�H;�H;�H;)�H;|�H;��H;r�H;t�H;��H;9�H;      L�H;o�H;�H;��H;��H;H�H;��H;��H;��H;��H;�H;H�H;�H;��H;��H;��H;a�H;"�H;��H;�H;L�H;[�H;U�H;(�H;��H;��H;�H;��H;��H;!�H;_�H;��H;��H;��H;��H;��H;��H;��H;��H;��H;��H;��H;_�H;�H;��H;��H;�H;��H;��H;(�H;\�H;W�H;G�H;�H;��H;%�H;c�H;��H;��H;��H;~�H;H�H;�H;��H;��H;��H;��H;G�H;��H;��H;�H;x�H;      ۹H;=�H;ȺH;��H;�H;��H;��H;��H;��H;O�H;��H;8�H;��H;�H;q�H;��H;��H;��H;]�H;��H;m�H;��H;��H;��H;��H;/�H;��H;O�H;��H; �H;Q�H;��H;��H;��H;��H;��H;��H;��H;��H;��H;��H;��H;Q�H;��H;��H;I�H;��H;2�H;��H;��H;��H;��H;f�H;��H;\�H;��H;��H;��H;n�H;�H;��H;;�H;��H;O�H;��H;��H;��H;��H;�H;��H;̺H;?�H;      z�H;��H;s�H;��H;P�H;D�H;��H;:�H;��H;��H;��H;��H;��H;��H;��H;R�H;��H;�H;8�H;!�H;��H;n�H;��H;��H;��H;��H;:�H;��H;p�H;��H;�H;X�H;��H;��H;��H;��H;��H;��H;��H;��H;��H;Z�H;�H;��H;k�H;��H;:�H;��H;��H;��H;��H;m�H;��H;�H;8�H;�H;��H;T�H;��H;��H;��H;��H;��H;��H;��H;=�H;��H;A�H;W�H;��H;~�H;��H;      ~�H;ڢH;ˣH;?�H;H�H;ЩH;��H;��H;��H;K�H;/�H;�H;��H;��H;"�H;q�H;��H;}�H;�H;s�H;��H;u�H;)�H;��H;��H;��H;��H;\�H;��H;k�H;��H;�H;N�H;��H;��H;��H;��H;��H;��H;��H;P�H;�H;��H;e�H;��H;V�H;��H;��H;��H;��H;3�H;s�H;��H;r�H;�H;}�H;��H;s�H;!�H;��H;��H;�H;/�H;I�H;��H;��H;��H;˩H;N�H;F�H;ԣH;բH;      ��H;	�H;4�H;A�H;�H;M�H;3�H;w�H;!�H;��H;��H;�H;ָH;��H;f�H;��H;��H;b�H;��H;��H;��H;��H;��H;��H;>�H;��H;��H;��H;O�H;��H;b�H;��H;�H;W�H;��H;�H;��H;��H;�H;Z�H;�H;��H;b�H;��H;I�H;��H;��H;��H;;�H;��H;��H;��H;��H;��H;��H;b�H;��H;��H;d�H;��H;ָH;�H;��H;��H;'�H;w�H;7�H;C�H;�H;@�H;;�H;�H;      �sH;&tH;�uH;WxH;�{H;V�H;��H;7�H;p�H;�H;��H;8�H;��H;��H;޷H;��H;��H;��H;�H;��H;^�H;j�H;�H;P�H;^�H;�H;X�H;��H;��H;L�H;��H;h�H;��H;�H;X�H;a�H;Z�H;b�H;W�H;�H;��H;i�H;��H;I�H;��H;��H;Z�H;�H;X�H;K�H;�H;k�H;Z�H;��H; �H;��H;��H;��H;�H;��H;��H;8�H;��H;�H;p�H;>�H;��H;S�H;�{H;bxH;�uH;'tH;      hOH;%PH;bRH;�UH;�ZH;�`H;�gH;BoH;wH;�H;ÈH;��H;0�H;��H;X�H;��H;��H;ݾH;��H;��H;�H;�H;v�H;i�H;��H;�H;��H;d�H;��H;��H;H�H;��H;b�H;��H;��H;�H;2�H;�H;��H;��H;g�H;��H;H�H;~�H;��H;`�H;��H;�H;��H;d�H;}�H;�H;�H;��H;��H;ܾH;��H;��H;V�H;��H;0�H;��H;ňH;�H;|wH;BoH;�gH;�`H;�ZH;�UH;mRH;PH;      @H;A H;9#H;�'H;j.H;�6H;�?H;JH;1UH;�`H;[lH;xH;\�H;]�H;ԘH;|�H;c�H;��H;��H;��H;��H;��H;��H;��H;��H;��H;��H;��H;3�H;��H;��H;N�H;��H;r�H;��H;��H;��H;��H;��H;s�H;��H;K�H;��H;��H;-�H;��H;��H;��H;��H;��H;��H;��H;��H;��H;��H;��H;d�H;|�H;ӘH;\�H;]�H;xH;]lH;�`H;/UH;!JH;�?H;�6H;z.H;�'H;:#H;? H;      �G;��G;��G;��G;��G;��G;-H;�H;�(H;�7H;vGH;WH; fH;�tH;<�H;�H;��H;q�H;��H;q�H;��H;~�H;(�H;�H;�H;u�H;U�H;��H;��H;a�H;��H;��H;S�H;��H;M�H;��H;��H;��H;O�H;��H;W�H;��H;��H;b�H;��H;��H;V�H;|�H;�H;��H;/�H;~�H;��H;t�H;��H;o�H;��H;�H;:�H;�tH; fH;WH;vGH;�7H;�(H;�H;-H;��G;��G;�G;��G;��G;      JvG;yG; �G;��G;��G;��G;��G;��G;{�G;hH;H;�,H;�@H;�SH;�eH;XvH;��H;|�H;�H;ܪH;l�H;ѼH;�H;A�H;d�H;��H;\�H;Y�H;��H;��H;[�H;��H;��H;@�H;��H; �H;#�H; �H;��H;A�H;��H;��H;^�H;��H;��H;X�H;]�H;��H;d�H;<�H;"�H;ѼH;k�H;�H;�H;x�H;��H;[vH;�eH;�SH;�@H;�,H;H;fH;z�G;��G;��G;��G;ĝG;��G;�G;yG;      9�F;�F;��F;��F;h�F;cG;CGG;�pG;�G;+�G;��G;e�G;�H;�)H;}AH;KWH;)kH;}H;�H;;�H;��H;$�H;D�H;!�H;��H;)�H;��H;|�H;��H;�H;
�H;��H;��H;��H;7�H;��H;��H;��H;7�H;��H;��H;��H;�H;�H;��H;|�H;��H;0�H;��H;�H;I�H;%�H;��H;@�H;�H;}H;-kH;KWH;AH;�)H;�H;e�G;��G;0�G;�G;�pG;CGG;UG;r�F;��F;��F; �F;      �mD;�~D;F�D;��D;Z\E;��E;l0F;��F;��F;�8G;�vG;�G;7�G;H�G;-H;o0H;0JH;baH;�uH;ׇH;��H;2�H;��H;��H;��H;��H;c�H;�H;��H;��H;[�H;>�H;��H;��H;��H;��H;(�H;��H;��H;��H;��H;=�H;_�H;��H;��H;�H;d�H;��H;��H;��H;��H;4�H;��H;ۇH;�uH;^aH;3JH;n0H;.H;I�G;<�G;�G;�vG;�8G;��F;ÔF;k0F;��E;c\E;��D;H�D;�~D;      `?;��?;��?;س@;��A;r�B;��C;�D;>iE;�F; �F;�G;EnG;�G;��G;D H;e!H;?H;cYH;VpH;B�H;q�H;��H;?�H;��H;�H;<�H;�H;��H;l�H;R�H;��H;��H;��H;��H;7�H;M�H;9�H;��H;��H;��H;��H;V�H;p�H;��H;�H;?�H;#�H;��H;A�H;�H;s�H;B�H;ZpH;eYH;?H;f!H;E H;��G;�G;GnG;�G;�F;�F;8iE;�D;��C;i�B;��A;�@;��?;��?;      &�4;��4;�5;�l7;o_9;H�;;��=;�?;U�A;ÚC;e�D;u�E;èF;X)G;��G;��G;��G;?H;�6H;�SH;�lH;m�H;��H;�H;��H;D�H;�H;-�H;��H;x�H;�H;��H;/�H;��H;��H;_�H;��H;^�H;��H;��H;/�H;��H;�H;�H;��H;/�H;�H;L�H;��H;�H;��H;n�H;�lH;�SH;�6H;8H;��G;��G;��G;U)G;ŨF;u�E;f�D;ÚC;Q�A;�?;��=;F�;;o_9;�l7;�5;��4;      e; ;Y";T%;��(;j-;02;��6;��:;�0>;�A;>YC;'�D;F;�F;�XG;��G;E�G;�H;N1H;�PH;�kH;k�H;t�H;1�H;"�H;мH;�H;��H;�H;j�H;��H;r�H;m�H;��H;Z�H;��H;]�H;��H;k�H;s�H;��H;p�H;�H;��H;~�H;ӼH;(�H;/�H;x�H;n�H;�kH;�PH;P1H;�H;@�G;��G;�XG;�F;F;)�D;>YC;�A;�0>;��:;��6;*2;	j-;��(;F%;[";� ;      ���:�B�:ʆ�:ox;|�
;�;-�;�}$;0|,;Y�3;�_9;4>;zA;��C;�E;��F;5G;o�G;Q�G;8H;�/H;�PH;�lH;C�H;��H;��H;e�H;��H;��H;�H;Y�H;��H;��H;��H;g�H;E�H;��H;G�H;g�H;��H;��H;��H;\�H;�H;�H;��H;h�H;��H;��H;E�H;�lH;�PH;�/H;:H;Q�G;m�G;5G;��F;�E;��C;	zA;3>;�_9;[�3;.|,;�}$;/�;�;��
;ix;��:�B�:      �w[:NBd:��}:��:-�:ɳ�:��:
�;�;P ;�+;��3;ҡ:;	�?;��B;�E;?ZF;�G;�G;k�G;>H;Q1H;�SH;ZpH;ׇH;@�H;ݪH;u�H;��H;��H;��H;��H;p�H;!�H;��H;�H;Y�H;�H;��H;�H;n�H;��H;��H;��H;��H;u�H;ߪH;D�H;ԇH;`pH;�SH;M1H;:H;k�G;�G;�G;AZF;�E;��B;
�?;ҡ:;��3;�+;P ;�;�;��:���:3�:��:��}:2Bd:      p�S���D����0��� (7X�9d�R:��:7��:��:�>;�";�P.;m7;��=;QB;԰D;r9F;G;�G;R�G;�H;�6H;bYH;�uH;�H;�H;��H;��H;��H;�H;��H;�H;6�H;^�H;��H;��H;��H;\�H;4�H;�H;��H;�H;��H;��H;��H;�H;�H;�uH;iYH;�6H;�H;N�G;�G;G;p9F;ְD;LB;��=;m7;�P.;�";�>; ��:5��:!��:\�R:8�9 (7@�������D�      E^��/X�rF�8}*�&���P����D��̬�Pi:��::��:/�;��;>�);��4;�<;�A;�D;p9F;�G;k�G;@�G;:H;?H;[aH;}H;t�H;q�H;��H;ܾH;��H;]�H;{�H;�H;��H;#�H;��H;#�H;��H;�H;y�H;\�H;��H;�H;��H;q�H;x�H;}H;UaH;?H;:H;>�G;g�G;�G;m9F;�D;�A;�<;��4;=�);��;.�;@��:��:Pi:@ͬ���D��P��)��?}*�"rF��/X�      ��ﻱ��k�ܻK�ƻj󩻼���FL���ĸ�� ��(�-:��:���:�;�>&;��3;M9<;�A;ְD;>ZF;5G;��G;��G;f!H;/JH;)kH;��H;��H;e�H;��H;��H;��H;��H;��H;��H;a�H;��H;a�H;��H;��H;��H;��H;��H;��H;c�H;��H;��H;(kH;(JH;f!H;��G;��G;5G;?ZF;԰D;	�A;K9<;��3;�>&;�;���:��:(�-: ���������FL����p�O�ƻp�ܻ���      m�V��5S��6H���6�F� �T,��?ػ;G���D^������D�H��9u4�:� �:%�;�%;��3;�<;OB;�E;��F;�XG;��G;B H;i0H;IWH;UvH;�H;{�H;��H;��H;��H;l�H;O�H;��H;��H;4�H;��H;��H;H�H;i�H;��H;��H;��H;x�H;�H;TvH;DWH;b0H;A H;��G;�XG;��F;�E;NB;�<;��3;�%;#�;� �:q4�:8��9��D�����D^�<G���?ػT,�I� ���6��6H��5S�      ��.��MȤ���������<�f�w�=����A�ܻ�*��[o5�r��� t(7P�}:�n�:%�;�>&;��4;��=;��B;�E;�F;��G;��G;+H;}AH;�eH;:�H;ԘH;V�H;ٷH;b�H;�H;��H;h�H;��H;K�H;��H;e�H;��H;�H;_�H;׷H;X�H;ԘH;7�H;�eH;xAH;&H;��G;��G;�F;܍E;��B;��=;��4;�>&; �;�n�:H�}: r(7t���[o5��*��?�ܻ���w�=�=�f� �������MȤ�.��      �c��8���������Ҽ����������r�JE:�H,�Nߵ��/X���º�Ǭ�T�}:� �:�;>�);m7;
�?;��C;F;X)G;�G;H�G;�)H;�SH;�tH;_�H;{�H;�H;��H;��H;��H;�H;��H;I�H;��H;�H;��H;��H;��H;�H;�H;_�H;�tH;�SH;�)H;?�G;�G;V)G;F;��C;�?;m7;=�);�;� �:D�}:�Ǭ���º�/X�Oߵ�G,�JE:���r�����������Ҽ�켷����8�      $'K���G��>��0�]y��c����U��� ��Y�V�+���ƻ�od���º w(7}4�:���:��;�P.;ϡ:;zA;'�D;ɨF;KnG;9�G;�H;�@H; fH;`�H;,�H;��H;ѸH;��H;��H;��H;z�H;5�H;z�H;��H;��H;��H;θH;��H;.�H;]�H;fH;�@H;�H;2�G;GnG;ŨF;&�D;zA;ҡ:;�P.;��;���:w4�: v(7��º�od��ƻ+��Y�V� ��U�����伖c�_y��0��>���G�      ���1Z��ϐ����}��c���D�2/%��8���Ҽ2c��4�f�����ƻ�/X�j���X��9��:/�;�";��3;=>;=YC;u�E;�G;�G;b�G;�,H;�VH;xH;��H;/�H;�H;�H;��H;-�H;A�H;-�H;A�H;*�H;��H;�H;�H;-�H;��H;xH;�VH;�,H;[�G;�G;�G;u�E;;YC;3>;��3;�";0�;��:8��9l����/X��ƻ���5�f�2c����Ҽ�8�3/%���D��c���}�ϐ��1Z��      �Pν�ʽO8���������ΐ��b�f���;�2�����CȤ�5�f�+��Qߵ�\o5���D��-:0��:�>;�+;�_9;�A;c�D;�F;�vG;��G;H;tGH;[lH;��H;��H;�H;)�H;��H;��H;�H;"�H;�H;��H;��H;&�H;�H;��H;��H;ZlH;oGH;H;��G;�vG;�F;c�D;�A;�_9;�+;�>;,��:�-: �D�_o5�Qߵ�,��6�f�CȤ����2����;�b�f�ΐ���������O8���ʽ      ���g9�Z[��s�{�ؽ���t����}���G������1c��Y�V�H,��*�����p��}�:��:M ;_�3;�0>;C;�F;�8G;'�G;eH;�7H;�`H;�H;�H;��H;H�H;��H;D�H;��H;�H;��H;B�H;��H;E�H;��H;�H;�H;�`H;�7H;dH;#�G;�8G;�F;ÚC;�0>;T�3;M ; ��:{�:p������*��H,�Z�V�2c���������G���}�t�����|�ؽ�s�Z[�g9�      ��=�׀:���0��Q"�~������Pν�榽@����G�2����Ҽ ��KE:�A�ܻ�D^�̸��,i:3��:�;2|,;��:;G�A;:iE;��F;�G;z�G;�(H;/UH;vwH;m�H;�H;��H;�H;��H;��H;�H;��H;��H;�H;��H;�H;l�H;{wH;/UH;�(H;{�G;�G;��F;<iE;H�A;��:;,|,;�;/��:4i:ʸ���D^�A�ܻKE:� ����Ҽ2����G�@���榽�Pν����~��Q"���0�ր:�      0Dx�4�s���f�tS�׀:����Z[��7ս�榽��}���;��8�V�����r����?G�����ά���:�;�}$;��6;��?;�D;ÔF;�pG;��G;�H;JH;:oH;9�H;u�H;��H;4�H;��H;��H;"�H;��H;��H;3�H;��H;o�H;6�H;AoH;JH;�H;��G;�pG;��F;�D;��?;��6;�}$;�;��:`ά���@G�������r�V����8���;���}��榽�7սZ[����׀:�tS���f�4�s�      �*���0��ޥ��;����k��H��#%�Z[��Pνt��a�f�3/%���伇���w�=��?ػ�FL���D�@�R:��:-�;.2;��=;��C;a0F;BGG;��G;H;�?H;�gH;��H;)�H;��H;��H;z�H;��H;p�H;��H;}�H;��H;��H;'�H;�H;�gH;�?H;!H;��G;FGG;a0F;��C;��=;*2;&�;��:8�R:��D��FL��?ػw�=��������3/%�a�f�t���PνZ[��#%��H��k�;���ޥ���0��      '�þ��� ����R��|쏾5�s��H�����������ϐ����D��c�����>�f�V,�����P�� �9���:�;j-;E�;;l�B;��E;UG;��G;��G;|6H;�`H;W�H;J�H;ѩH;K�H;��H;L�H;��H;L�H;��H;J�H;ЩH;I�H;S�H;�`H;~6H;��G;��G;[G;��E;n�B;E�;;j-;�;���:��9�P�����V,�>�f������c���D�ΐ�������������H�5�s�|쏾�R�� ������      @��/�待Yؾ(�þĪ�|쏾�k�׀:�~�|�ؽ�����c�^y���Ҽ����F� �o�8�� (73�:��
;��(;v_9;��A;a\E;e�F;��G;��G;�.H;�ZH;�{H;�H;E�H;M�H;�H;��H;r�H;��H;�H;J�H;D�H;�H;�{H;�ZH;�.H;��G;��G;o�F;`\E;��A;v_9;��(;��
;;�: (74��o�F� �������Ҽ^y��c�����{�ؽ~�׀:��k�|쏾Ī�(�þ�Yؾ/��      #��N������>I�(�þ�R��;���tS��Q"��s������}��0��켊�����6�L�ƻD}*�P�����:tx;P%;�l7;ҳ@;��D;��F;��G;}�G;�'H;�UH;[xH;J�H;B�H;��H;��H;��H;w�H;��H;��H;��H;B�H;J�H;XxH;�UH;�'H;}�G;��G;��F;��D;ӳ@;�l7;N%;sx;��:`���@}*�K�ƻ��6��������0���}�����s��Q"�tS�;����R��(�þ>Iᾣ���O��      ���R��8�
������Yؾ���ޥ����f���0�Z[�O8��ϐ���>�����KȤ��6H�f�ܻrF�����}:��:[";%�5;��?;R�D;��F;�G;��G;*#H;]RH;�uH;C�H;��H;q�H;��H;�H;��H;�H;��H;q�H;��H;B�H;�uH;dRH;*#H;��G;	�G;��F;M�D;��?;!�5;X";���:�}:��rF�g�ܻ�6H�KȤ������>�ϐ��N8��Z[���0���f�ޥ������Yؾ����8�
�R��      �� ����R��N��/������0��4�s�׀:�g9��ʽ1Z����G��8�.���5S����
0X���D�JBd:�B�:� ;��4;��?;�~D;�F;	yG;��G;I H;'PH;tH;�H;ʢH;ðH;)�H;m�H;2�H;j�H;)�H;ðH;ȢH;�H;tH;.PH;J H;��G;yG;�F;�~D;��?;��4;� ;�B�:^Bd:��D�0X���껰5S�.���8���G�1Z���ʽg9�׀:�4�s��0�����/��N��R�����      GF�Wh����VVھ8�������~���S��#��o��8S��p₽2�6�q���jy��YFB��Eֻ�A?��	�[Y�:���:_�";_46;T@;[�D;��F;�nG;��G;�H;@H;�fH;>�H;+�H;��H;̳H;ʹH;��H;ƹH;˳H;��H;(�H;;�H;�fH;@H;�H;��G;�nG;��F;X�D;T@;Y46;]�";���:aY�:�	��A?��EֻYFB�jy��q���3�6�p₽8S���o���#��S��~������7��VVھ��Wh��      Vh���b���쾧*־�v��(���*��(�O�V� �s��r���؀�H�3���@ݜ�?�>�X�ѻ�9� ���o�:5% ;jM#;;�6;DA@;��D;��F;qG;F�G;H;�@H;dgH;��H;��H;٩H;�H;��H;ڻH;�H;�H;٩H;��H;��H;^gH;�@H;H;F�G;qG;��F;��D;BA@;5�6;fM#;3% ;o�:����9�X�ѻ?�>�@ݜ���H�3��؀��r��s�V� �'�O�*��)����v���*־���b��      ���쾳�޾/5ʾL;���:��(�v��E�`'����r����u���+��W��A����4���Ļ(9)��j��iW�:Z�;%;�k7;�@;��D;��F;�wG;N�G;.H;:CH;$iH;�H;��H;��H;��H;��H;o�H;��H;��H;��H;��H;�H; iH;@CH;.H;P�G;�wG;��F;��D;�@;�k7;�%;Z�;qW�:�j��&9)���Ļ��4��A���W缄�+���u�q�����`'��E�(�v��:��L;��/5ʾ��޾��      VVھ�*־/5ʾr��������M���9b��5�����ս����Xc���̖ռ�I��X�$�rT���Z��]����:��;c�';�8;RA;�9E;��F;��G;��G;=H;GH;lH;?�H;8�H;ޫH;��H;��H;M�H;��H;��H;ޫH;4�H;>�H;lH;GH;?H;��G;��G;��F;�9E;RA;�8;a�';��;�:�]���Z�qT��X�$��I��̖ռ���Xc������ս���5��9b��M������r���05ʾ�*־      7���v��M;������RP��E�r�z�H�U� ���6@��ѓ����K�b��վ���s�u���񕻲ܺP4u9�%�:�;%�+;v�:;�"B;h�E;��F;ΐG;��G;*H;3LH;�oH;9�H;q�H;��H;2�H;ּH;�H;мH;3�H;��H;n�H;4�H;�oH;8LH;*H;��G;АG;��F;h�E;�"B;r�:;%�+;�;&�:@4u9�ܺ��u����s��վ�b���K�ѓ��6@����U� �z�H�E�r�RP������M;���v��      ����(����:���M��E�r�&�O�#,�X�
��gٽqĥ���u�y1�j���+Ϥ���P�[��.o��p��:O��:�P;6�/;0�<;�
C;�E;f!G;0�G;��G;�%H;�RH;�tH;�H;C�H;ӯH;��H;X�H;�H;R�H;��H;ЯH;@�H;�H;�tH;�RH;�%H;��G;0�G;n!G;�E;�
C;/�<;4�/;�P;W��::�p���.o�[򻭎P�+Ϥ�j���x1���u�qĥ��gٽX�
�#,�&�O�E�r��M���:��(���      �~��*��(�v��9b�z�H�#,�MZ����7S��x^����N������μ�I���%+�����.������j~:9��:%m;��3;�>;6�C;6PF;yFG;L�G;��G;r/H;�YH;qzH;B�H;��H;Y�H;�H;&�H;��H;#�H;�H;Y�H;�H;@�H;nzH;ZH;u/H;��G;L�G;~FG;7PF;4�C;�>;��3;"m;C��:�j~:�����.�����%+��I����μ�����N�x^��7S�����MZ�#,�z�H��9b�(�v�*��      �S�'�O��E��5�U� �X�
���罥9��(l���Xc���(��������[�����ݎ�Xܺ�:9��:&�	;=d';] 8;6�@;x�D;ߩF;jG;��G;HH;j:H;=bH;��H;�H;.�H;?�H;z�H;3�H;��H;2�H;}�H;@�H;+�H;��H;��H;DbH;m:H;KH;��G;jG;�F;t�D;6�@;_ 8;<d';,�	;��:�:9Wܺ�ݎ������[��������(��Xc�'l���9�����X�
�U� ��5��E�'�O�      �#�U� �`'������gٽ7S��'l��O�j�D�3��i��վ�{���
(���ĻjA?���B���@:�[�:Q;��.;��;;ttB;�E;y�F;�G;��G;�H;NFH;!kH;��H;�H;�H;d�H;�H;p�H;��H;n�H;
�H;d�H;�H;�H;��H;&kH;RFH;�H;��G;"�G;}�F;�E;wtB;��;;��.;
Q;�[�:��@:��B�jA?���Ļ	(�{����վ��i�D�3�N�j�'l��7S���gٽ����`'�U� �      �o��s��罫�ս5@��qĥ�x^���Xc�D�3���	�ˌ˼�]��UFB�[򻲜���Ӻ���8��:ԛ;�M#;n=5;?;E�C;w@F; :G;�G;�G;*'H;�RH;vtH;��H;x�H;(�H;��H;��H;��H;>�H;��H;��H;��H;&�H;t�H;��H;|tH;�RH;-'H;�G;�G;:G;u@F;H�C;?;n=5;�M#;՛;��:@��8Ӻ���� [�UFB��]��ˌ˼��	�D�3��Xc�x^��pĥ�6@����ս���s�      8S���r��r�����ѓ����u���N���(��i�̌˼�A����P�js��D|�����x\:!�:i�;pn-;ܞ:;�A;t,E;d�F;#oG;��G;�H;�7H;6_H;~H;�H; �H;q�H;	�H;w�H;9�H;�H;9�H;w�H;�H;p�H;��H;�H;~H;;_H;�7H;�H;��G;)oG;f�F;y,E;�A;ޞ:;{n-;k�;!�:�\:����B|��js���P��A��̌˼�i���(���N���u�ѓ�����r���r��      p₽�؀���u��Xc���K�y1�������վ��]����P����FT����9�,�o�h3�9f&�:Y�	;T%;?�5;��>;��C;�F;�!G;��G;��G;@H;[HH;�kH;��H;F�H;��H;��H;q�H;I�H;��H;��H;��H;H�H;u�H;��H;��H;I�H;��H;�kH;^HH;AH;��G;��G;�!G;�F;��C;��>;K�5;W%;V�	;p&�:p3�9(�o���9�ET�������P��]���վ�����x1���K��Xc���u��؀�      3�6�G�3���+���a�k�����μ���{���TFB�is�FT��3�D��{���9u9�q�:k��:xY;�t0;��;;�B;�9E;߻F;�gG;ԿG;��G;v0H;�XH;#xH;�H;r�H;��H;��H;��H;�H;,�H;0�H;,�H;�H;��H;�H;��H;u�H;&�H;)xH;�XH;w0H;��G;ٿG;�gG;�F;�9E;�B;��;;�t0;sY;w��:�q�: :u9�{��2�D�DT��is�TFB�z��������μj���b�����+�G�3�      n�����W�͖ռ�վ�,Ϥ��I����[�
(��Z����9��{�� ;9=X�:JX�:3Q;8,;��8;�A@;BD;�@F;�,G;��G;��G;bH;�DH;hH;)�H;O�H;a�H;[�H; �H;�H;��H;��H;b�H;��H;��H;�H;�H;X�H;e�H;X�H;3�H;hH;�DH;^H;��G;��G;�,G;�@F;BD;�A@;��8;6,;9Q;HX�:EX�:0;9�{����9���Z�(���[��I��+Ϥ��վ�͖ռ�W���      hy��Aݜ��A���I����s���P��%+������Ļ����@|�@�o��9u9CX�:�+�:P;�);̈́6;p�>;zPC;^�E;��F;�xG;&�G;vH;a1H;XH;�vH;��H;�H;��H;z�H;�H;>�H;~�H;��H;��H;��H;}�H;?�H;�H;w�H;��H;�H;��H;wH;XH;\1H;xH;)�G;�xG;��F;b�E;�PC;t�>;Ǆ6;�);P;�+�:IX�: :u9,�o�<|�������Ļ����%+���P���s��I���A��@ݜ�      SFB�>�>���4�W�$�u��[�����ݎ�oA?�|Ӻ����X3�9�q�:JX�:P;��';|=5;y�=;��B;GE;E�F;UG;�G;��G;PH;�HH;jH;�H;q�H;D�H;-�H;F�H;��H;>�H;�H;�H;��H;�H;	�H;=�H;��H;C�H;3�H;I�H;x�H;�H;jH;�HH;SH;��G;�G;�UG;I�F;GE;�B;t�=;�=5;��';R;HX�:�q�:h3�9x���yӺhA?��ݎ����[�x��X�$���4�;�>�      �EֻV�ѻ��ĻuT�����.o���.�Pܺ��B����8�\:f&�:s��:7Q;�);�=5;�:=;%#B;~�D;�uF;�6G;��G;Y�G;oH;�:H;^H;�zH;��H;]�H;��H;�H;��H;Z�H;�H;j�H;/�H;��H;*�H;h�H;�H;U�H;��H;�H;ŲH;a�H;��H;�zH;	^H;�:H;rH;V�G;��G;�6G;�uF;��D; #B;�:=;=5;�);9Q;s��:l&�:�\:���8��B�Mܺ�.��.o���xT����ĻQ�ѻ      }A?��9�,9)��Z��ܺ�p������ ;9��@:��:'�:R�	;oY;6,;Ƅ6;o�=;#B;��D;ZXF;�!G;v�G;�G;�H;�.H;uSH;_qH;ۉH;��H;_�H;��H;m�H;��H;��H;��H;�H;�H;��H;�H;|�H;��H;��H;��H;o�H;��H;c�H;��H;ىH;ZqH;ySH;�.H;�H;�G;z�G;�!G;^XF;��D;#B;m�=;Ʉ6;4,;oY;R�	;1�:��:��@:0;9����|p���ܺ�Z�$9)��9�      ��	������j��@]��@4u9@:�j~:��:�[�:؛;r�;Q%;�t0;��8;s�>;�B;�D;cXF;1G;[�G;��G;��G;�%H; KH;�iH;��H;��H;4�H;s�H;�H;Z�H;��H;��H;0�H;~�H;��H;P�H;��H;z�H;/�H;��H;��H;[�H;�H;q�H;4�H;��H;݂H;�iH;KH;�%H;��G;��G;_�G;4G;]XF;��D;��B;t�>;��8;�t0;U%;r�;՛;�[�:��:�j~:(:P4u9�^���j������      KY�:o�:sW�:�:�%�:W��:U��:&�	;Q;�M#;xn-;G�5;��;;�A@;�PC;GE;�uF;�!G;\�G;��G;�G;C H;	EH;�cH;4}H;q�H;��H;��H;��H;��H;��H;(�H;Q�H;P�H;K�H;y�H;��H;r�H;H�H;P�H;O�H;%�H;��H;��H;��H;��H;��H;n�H;8}H;�cH;EH;E H;�G;��G;_�G;�!G;�uF;GE;�PC;�A@;��;;H�5;{n-;�M#;Q;-�	;O��:c��:�%�:��:[W�:�n�:      ���:#% ;<�;��;�;�P;$m;9d';��.;n=5;ޞ:;��>;�B;BD;_�E;I�F;�6G;��G;��G;�G;pH;�AH;`H;GyH;z�H;�H;M�H;߹H;H�H;��H;��H;/�H;��H;@�H;��H;��H;C�H;��H;��H;>�H;��H;*�H;��H;��H;G�H;޹H;H�H;�H;|�H;FyH;`H;�AH;rH;�G;��G;|�G;�6G;H�F;_�E;BD;�B;��>;�:;m=5;��.;6d';(m;�P;�;��;F�;% ;      R�";lM#;%;m�';#�+;6�/;��3;Z 8;��;;?;��A;��C;�9E;�@F;��F;�UG;��G; �G;��G;E H;�AH;�^H;BwH;�H;~�H;۫H;��H;+�H;��H;"�H;�H;��H;��H;��H;k�H;I�H;y�H;B�H;i�H;��H;��H;��H;�H;%�H;��H;(�H;��H;٫H;��H;�H;=wH;�^H;�AH;E H;��G;�G;��G;UG;��F;�@F;�9E;��C;��A;?;��;;d 8;��3;/�/;6�+;a�';�%;`M#;      t46;8�6;�k7;"�8;n�:;7�<;#�>;@�@;tB;M�C;�,E;�F;�F;�,G;�xG;"�G;\�G;�H;�%H;EH;`H;@wH;-�H;1�H;C�H;�H;��H;k�H;��H;��H;%�H;=�H;��H;\�H;��H;o�H;��H;i�H;��H;]�H;��H;9�H;(�H;��H;��H;j�H;��H;�H;G�H;.�H;&�H;AwH;`H;EH;�%H;�H;Z�G; �G;�xG;�,G;�F;�F;�,E;H�C;~tB;@�@;!�>;4�<;|�:;�8;�k7;�6;      U@;LA@;�@;RA;�"B;�
C;8�C;x�D;�E;{@F;j�F;�!G;�gG;��G;)�G;��G;rH;�.H;KH;�cH;DyH;�H;.�H;��H;�H;z�H;t�H;��H;�H;K�H;��H;I�H;7�H;��H;��H;^�H;��H;X�H;��H;��H;7�H;F�H;��H;J�H;�H;��H;n�H;{�H;�H;��H;*�H;�H;CyH;�cH;�JH;�.H;qH;��G;(�G;��G;�gG;�!G;m�F;y@F;�E;~�D;7�C;�
C;�"B;RA;�@;EA@;      {�D;��D;��D;�9E;a�E;"�E;APF;�F;}�F;:G;3oG;��G;ٿG;��G;{H;YH;�:H;�SH;�iH;=}H;��H;��H;F�H;�H;9�H;��H;,�H;j�H;��H;'�H;��H;�H;��H;��H;��H;$�H;b�H;�H;��H;��H;��H;�H;��H;(�H;��H;i�H;#�H;��H;:�H;�H;F�H;��H;�H;8}H;�iH;|SH;�:H;WH;zH;��G;ٿG;��G;1oG;:G;��F;�F;APF;�E;j�E;}9E;��D;��D;      ��F;��F;��F;�F;��F;q!G;�FG;jG;%�G;�G;��G;��G;�G;kH;a1H;�HH;^H;aqH;݂H;k�H;�H;֫H;ߵH;x�H;��H;�H;�H;X�H;��H;��H;��H;��H;��H;��H;w�H;��H;�H;��H;u�H;��H;��H;|�H;��H;��H;��H;U�H;�H;�H;��H;u�H;ߵH;׫H;�H;j�H;܂H;ZqH;^H;�HH;_1H;dH;��G;��G;��G;�G;#�G;jG;�FG;f!G;��F;��F;��F;��F;      �nG;qG;�wG;��G;ŐG;+�G;Z�G;��G;��G;�G;�H;>H;u0H;�DH;XH;jH;�zH;߉H;��H;��H;Q�H;��H;��H;t�H;)�H;�H;;�H;��H;Z�H;z�H;H�H;��H;��H;��H;4�H;��H;��H;��H;0�H;��H;��H;��H;H�H;w�H;Y�H;��H;2�H;�H;)�H;p�H;��H;��H;O�H;��H;��H;ىH;�zH;jH;XH;�DH;u0H;@H;�H;�G;��G;��G;T�G;)�G;ܐG;��G;�wG;�pG;      ��G;C�G;I�G;��G;��G;��G;��G;HH;�H;3'H;�7H;bHH;�XH;hH;�vH;�H;��H;��H;4�H;��H;߹H;&�H;e�H;��H;h�H;U�H;��H;7�H;t�H;>�H;��H;��H;��H;`�H;��H;�H;�H;��H;��H;a�H;��H;��H;��H;=�H;t�H;6�H;��H;W�H;j�H;��H;h�H;'�H;޹H;��H;4�H;��H;��H;�H;�vH;hH;�XH;dHH;�7H;3'H;�H;HH;��G;��G;��G;��G;I�G;8�G;      �H;�H;+H;JH;H;�%H;y/H;i:H;HFH;�RH;=_H;�kH;)xH;.�H;��H;u�H;b�H;f�H;v�H;��H;I�H;��H;��H;	�H;��H;��H;U�H;t�H;�H;��H;��H;��H;R�H;��H;B�H;u�H;��H;p�H;B�H;��H;V�H;��H;��H;��H;�H;s�H;O�H;��H;��H;�H;��H;��H;G�H;��H;t�H;c�H;b�H;w�H;��H;-�H;&xH;�kH;@_H;�RH;KFH;i:H;y/H;�%H;&H;GH;+H;H;      @H;�@H;DCH;GH;:LH;�RH;ZH;<bH;%kH;|tH;~H;��H;$�H;Y�H;�H;D�H;ŲH;��H;�H;��H;��H;�H;��H;D�H;'�H;��H;v�H;=�H;��H;��H;��H;g�H;��H;L�H;��H;��H;��H;��H;��H;L�H;��H;a�H;��H;��H;��H;;�H;q�H;��H;'�H;C�H;��H;�H;��H;��H;�H;��H;ŲH;E�H;�H;V�H;#�H;��H;~H;~tH;#kH;AbH;ZH;�RH;:LH;GH;ECH;�@H;      �fH;vgH;*iH;lH;�oH;�tH;xzH;��H;��H;��H;�H;P�H;z�H;m�H;�H;5�H;�H;r�H;^�H;��H;��H;�H;"�H;��H;��H;��H;H�H;��H;��H;��H;e�H;�H;]�H;��H;��H;�H;&�H;�H;��H;��H;^�H;��H;e�H;��H;��H;��H;E�H;��H;��H;��H;(�H;�H;��H;��H;]�H;q�H;�H;4�H;�H;k�H;}�H;Q�H;�H;��H;��H;��H;�zH;�tH;�oH;lH;+iH;ygH;      <�H;��H;	�H;7�H;6�H;�H;H�H;�H; �H;z�H;�H;��H;�H;e�H;}�H;H�H;��H;��H;��H;,�H;2�H;��H;9�H;C�H;�H;{�H;��H;��H;��H;g�H;��H;s�H;��H;��H;$�H;?�H;?�H;?�H;#�H;��H;��H;n�H;��H;e�H;��H;��H;��H;|�H;	�H;>�H;=�H;��H;.�H;(�H;��H;��H;��H;K�H;~�H;b�H;�H;��H;�H;{�H;�H;�H;P�H;�H;A�H;8�H;�H;��H;      .�H;��H;��H;6�H;x�H;@�H;��H;*�H;�H;-�H;w�H;��H;��H;'�H;�H;��H;\�H;��H;��H;T�H;��H;��H;��H;2�H;��H;��H;��H;��H;W�H;��H;[�H;��H;�H;5�H;S�H;t�H;{�H;t�H;P�H;5�H;�H;��H;X�H;��H;V�H;��H;��H;��H;��H;2�H;��H;��H;��H;Q�H;��H;��H;^�H;��H;�H;'�H;��H;��H;x�H;.�H;�H;+�H;��H;:�H;|�H;1�H;��H;��H;      ��H;ԩH;��H;ԫH;��H;ɯH;c�H;B�H;i�H;��H;�H;|�H;��H;$�H;E�H;D�H;�H;��H;3�H;S�H;B�H;��H;U�H;��H;��H;��H;��H;c�H;��H;O�H;��H;��H;2�H;o�H;~�H;��H;��H;��H;}�H;p�H;4�H;��H;��H;J�H;��H;^�H;��H;��H;��H;��H;\�H;��H;=�H;M�H;2�H;��H;"�H;D�H;E�H;#�H;��H;|�H;�H;��H;l�H;I�H;g�H;ȯH;��H;׫H;��H;�H;      ɳH; �H;��H;õH;B�H;��H;&�H;z�H;�H;��H;��H;Q�H;�H;��H;��H;�H;m�H;}�H;}�H;L�H;��H;g�H;��H;��H;��H;m�H;,�H;��H;B�H;��H;��H;&�H;Q�H;�H;��H;��H;��H;��H;��H;��H;U�H;&�H;��H;��H;>�H;��H;,�H;n�H;��H;��H;��H;f�H;��H;E�H;z�H;�H;q�H;�H;��H;��H;�H;T�H;��H;��H;�H;��H;*�H;��H;B�H;ĵH;´H;%�H;      ʹH;��H;��H;��H;ԼH;M�H;5�H;6�H;r�H;��H;B�H;��H;0�H;��H;��H;�H;/�H;�H;��H;u�H;��H;D�H;d�H;L�H;�H;��H;��H; �H;w�H;��H;�H;C�H;z�H;��H;��H;��H;��H;��H;��H;��H;}�H;C�H;�H;��H;u�H;��H;��H;��H;�H;M�H;k�H;B�H;��H;p�H;��H;�H;2�H;�H;��H;��H;0�H;��H;D�H;��H;v�H;<�H;:�H;O�H;ּH;��H;��H;�H;      ŻH;ٻH;��H;L�H;|�H;�H;��H;��H;��H;C�H;��H;��H;>�H;o�H;��H;��H;��H;��H;S�H;��H;K�H;|�H;��H;��H;b�H; �H;��H;�H;��H;��H;#�H;C�H;}�H;��H;��H;��H;��H;��H;��H;��H;��H;B�H;$�H;��H;��H;�H;��H;�H;b�H;��H;��H;|�H;F�H;��H;S�H;��H;��H;��H;��H;o�H;=�H;��H;��H;H�H;��H;��H;��H;�H;~�H;J�H;��H;�H;      ˹H;��H;��H;��H;ԼH;R�H;4�H;7�H;r�H;��H;@�H;��H;2�H;��H;��H;�H;-�H;�H;��H;u�H;��H;E�H;d�H;L�H;�H;��H;��H; �H;y�H;��H;�H;D�H;{�H;��H;��H;��H;��H;��H;��H;��H;}�H;C�H;�H;��H;u�H;��H;��H;��H;�H;M�H;k�H;A�H;��H;p�H;��H;�H;0�H; �H;��H;��H;0�H;��H;D�H;��H;v�H;=�H;7�H;O�H;ؼH;��H;��H;��H;      ��H;#�H;��H;��H;D�H;��H;)�H;~�H;�H;��H;��H;Q�H;�H;��H;��H;�H;m�H;�H;}�H;L�H;��H;i�H;��H;��H;��H;k�H;,�H;��H;C�H;��H;��H;&�H;S�H;�H;��H;��H;��H;��H;��H;��H;W�H;&�H;��H;��H;>�H;��H;,�H;p�H;��H;��H;��H;g�H;��H;E�H;z�H;�H;q�H;�H;��H;��H;�H;V�H;��H;��H;�H;��H;/�H;��H;G�H;��H;��H;&�H;      ��H;שH;��H;ګH;��H;ͯH;b�H;G�H;k�H;��H;�H;{�H;��H;$�H;F�H;B�H; �H;��H;3�H;S�H;B�H;��H;U�H;��H;��H;��H;��H;c�H;��H;P�H;��H;��H;1�H;o�H;~�H;��H;��H;��H;}�H;p�H;5�H;��H;��H;J�H;��H;^�H;��H;��H;��H;��H;\�H;��H;;�H;N�H;2�H;��H;!�H;E�H;F�H;#�H;��H;|�H;�H;��H;l�H;L�H;i�H;̯H;��H;׫H;��H;ةH;      .�H;��H;��H;5�H;u�H;C�H;��H;-�H;�H;-�H;w�H;��H;��H;'�H;�H;��H;\�H;��H;��H;U�H;��H;��H;��H;2�H;��H;��H;��H;��H;Z�H;��H;Z�H;��H; �H;4�H;Q�H;w�H;{�H;t�H;S�H;5�H;�H;��H;Z�H;��H;R�H;��H;��H;��H;��H;/�H;��H;��H;��H;R�H;��H;��H;^�H;��H;�H;'�H;��H;��H;w�H;.�H;�H;1�H;��H;@�H;y�H;;�H;��H;��H;      .�H;��H;��H;5�H;2�H;��H;L�H;�H;�H;z�H;�H;��H;�H;b�H;�H;J�H;��H;��H;��H;+�H;5�H;��H;:�H;B�H;�H;|�H;��H;��H;��H;e�H;��H;o�H;��H;��H;'�H;=�H;?�H;?�H;#�H;��H;��H;o�H;��H;e�H;��H;��H;��H;}�H;�H;;�H;@�H;��H;+�H;(�H;��H;��H;��H;J�H;}�H;b�H;�H;��H;�H;{�H;#�H;�H;O�H;�H;3�H;5�H;�H;��H;      �fH;ugH;-iH;lH;�oH;�tH;xzH;��H;��H;��H;�H;Q�H;z�H;k�H;�H;5�H;�H;r�H;]�H;��H;��H;�H;#�H;��H;��H;��H;D�H;��H;��H;��H;e�H;�H;^�H;��H;��H;�H;&�H;�H;��H;��H;`�H;�H;d�H;��H;��H;��H;D�H;��H;��H;��H;)�H;�H;��H;��H;^�H;o�H;�H;4�H;�H;m�H;|�H;S�H;�H;��H;��H;��H;zH;�tH;pH;lH;2iH;vgH;      @H;�@H;>CH;GH;1LH;�RH;ZH;DbH;&kH;~tH;~H;��H;$�H;V�H;�H;E�H;ŲH;��H;�H;��H;��H;!�H;��H;D�H;(�H;��H;t�H;=�H;��H;��H;��H;e�H;��H;M�H;��H;��H;��H;��H;��H;M�H;��H;e�H;��H;��H;��H;:�H;s�H;��H;&�H;?�H;��H;�H;��H;��H;�H;��H;ŲH;G�H;�H;X�H;&�H;��H;~H;�tH;%kH;DbH;ZH;�RH;:LH;GH;KCH;�@H;      �H;H;<H;GH;H;�%H;v/H;i:H;QFH;�RH;=_H;�kH;)xH;0�H;��H;x�H;a�H;f�H;q�H;��H;I�H;��H;��H;	�H;��H;��H;P�H;t�H;!�H;��H;��H;��H;S�H;��H;C�H;s�H;��H;s�H;C�H;��H;V�H;��H;��H;��H;�H;p�H;R�H;��H;��H;�H;��H;��H;G�H;��H;v�H;b�H;`�H;x�H;��H;.�H;'xH;�kH;>_H;�RH;OFH;m:H;{/H;�%H;#H;DH;=H;�H;      ��G;7�G;<�G;��G;��G;�G;��G;NH;�H;3'H;�7H;bHH;�XH;hH; wH;�H;��H;��H;1�H;��H;߹H;(�H;d�H;��H;j�H;P�H;��H;6�H;w�H;;�H;��H;��H;��H;a�H;��H;��H;�H;��H;��H;c�H;��H;��H;��H;;�H;s�H;3�H;��H;X�H;h�H;��H;k�H;'�H;ܹH;��H;4�H;��H;��H;�H; wH;hH;�XH;bHH;�7H;2'H;�H;IH;��G;��G;��G;��G;J�G;7�G;      �nG;qG;�wG;ǂG;ԐG;4�G;X�G;��G;��G;�G;�H;@H;r0H;�DH;XH;jH;�zH;߉H;��H;��H;Q�H;��H;��H;w�H;'�H;�H;5�H;��H;\�H;v�H;G�H;��H;��H;��H;4�H;��H;��H;��H;2�H;��H;��H;��H;I�H;w�H;W�H;��H;6�H;�H;)�H;q�H;��H;��H;O�H;��H;��H;܉H;�zH;jH;XH;�DH;s0H;BH;�H;�G;��G;��G;Z�G;1�G;ڐG;łG;�wG;qG;      x�F;��F;��F;}�F;��F;v!G;zFG; jG;&�G;�G;��G;��G;�G;eH;b1H;�HH;^H;aqH;܂H;j�H;�H;֫H;ܵH;x�H;��H;�H;�H;U�H;��H;��H;��H;��H;��H;��H;x�H;��H;
�H;��H;u�H;��H;��H;��H;��H;��H;��H;U�H;�H;�H;��H;w�H;�H;׫H;�H;m�H;߂H;^qH;^H;�HH;f1H;gH;�G;��G;��G;�G;!�G;jG;|FG;g!G;��F;|�F;��F;y�F;      z�D;��D;��D;�9E;a�E;$�E;BPF;�F;��F;:G;0oG;��G;׿G;��G;}H;YH;�:H;�SH;�iH;;}H;�H;��H;C�H;�H;:�H;��H;%�H;i�H;��H;$�H;��H;�H;��H;��H;��H;"�H;c�H;!�H;��H;��H;��H;�H;��H;(�H;��H;h�H;)�H;��H;9�H;�H;H�H;��H;�H;?}H;�iH;|SH;�:H;ZH;H;��G;ۿG;��G;0oG;:G;}�F;�F;APF;�E;h�E;9E;��D;��D;      5@;7A@;
�@;RA;�"B;C;:�C;z�D;�E;w@F;k�F;�!G;�gG;��G;(�G;��G;qH;�.H; KH;�cH;DyH;�H;*�H;��H;�H;t�H;q�H;��H;�H;G�H;��H;J�H;9�H;��H;��H;Z�H;��H;[�H;��H;��H;:�H;I�H;��H;K�H;�H;��H;q�H;{�H;�H;��H;.�H;�H;FyH;�cH;KH;�.H;rH;��G;)�G;��G;�gG;�!G;k�F;x@F;�E;t�D;8�C;�
C;�"B;,RA;�@;A@;      h46;7�6;�k7;*�8;l�:;3�<;�>;>�@;�tB;I�C;|,E;�F;�F;�,G;�xG;"�G;Z�G;�H;�%H;EH;`H;AwH;(�H;0�H;F�H;ߵH;��H;h�H;��H;��H;&�H;?�H;��H;\�H;��H;o�H;��H;l�H;��H;[�H;��H;?�H;*�H;��H;��H;h�H;��H;�H;D�H;1�H;*�H;AwH;`H;EH;�%H;�H;\�G;!�G;�xG;�,G;�F;�F;},E;K�C;tB;D�@;�>;3�<;j�:;&�8;�k7; �6;      X�";nM#;�%;f�';#�+;:�/;��3;^ 8;��;;?;��A;��C;�9E;�@F;��F;�UG;��G;�G;��G;E H;�AH;�^H;>wH;�H;��H;ҫH;��H;(�H;��H;�H;�H;��H;��H;��H;i�H;E�H;y�H;G�H;g�H;��H;��H;��H; �H;%�H;��H;'�H;��H;ګH;�H;�H;AwH;�^H;�AH;F H;��G;�G;��G;UG;��F;�@F;�9E;��C;��A;?;��;;a 8;��3;%�/;:�+;X�';�%;`M#;      ���:<% ;N�;��;�;�P;&m;9d';��.;k=5;�:;��>;�B;BD;b�E;I�F;�6G;�G;��G;�G;qH;�AH;`H;FyH;{�H;�H;H�H;ܹH;G�H;��H;��H;/�H;��H;B�H;��H;��H;D�H;��H;��H;=�H;��H;-�H;��H;��H;G�H;ܹH;M�H;�H;{�H;IyH;`H;�AH;qH;�G;��G;|�G;�6G;I�F;d�E;BD;�B;��>;�:;n=5;��.;=d';+m;�P;�;��;\�;(% ;      {Y�:o�:iW�:�:�%�:c��:W��:0�	;Q;�M#;{n-;G�5;��;;�A@;�PC;GE;�uF;�!G;^�G;��G;�G;E H;EH;�cH;8}H;m�H;��H;��H;��H;��H;��H;(�H;Q�H;S�H;K�H;u�H;��H;u�H;H�H;M�H;O�H;'�H;��H;��H;��H;��H;��H;q�H;5}H;�cH;EH;C H;�G;��G;^�G;�!G;�uF;GE;�PC;�A@;��;;G�5;|n-;�M#;Q;)�	;Q��:Q��:�%�:��:kW�:o�:      ��	������j�� ]�� 4u9@:�j~:��:�[�:՛;p�;R%;�t0;��8;u�>;�B;�D;`XF;1G;\�G;��G;��G;�%H; KH;�iH;݂H;��H;3�H;s�H;�H;Z�H;��H;��H;0�H;}�H;��H;P�H;��H;{�H;/�H;��H;��H;[�H;�H;q�H;3�H;��H;߂H;�iH;KH;�%H;��G;��G;^�G;2G;]XF;�D;��B;u�>;��8;�t0;R%;r�;כ;�[�:��:�j~:<:�3u9`]���j��X���      �A?�ڡ9�09)��Z��ܺnp������p;9��@:��:+�:R�	;oY;4,;ʄ6;r�=;#B;��D;\XF;�!G;z�G;�G;�H;�.H;ySH;[qH;؉H;��H;c�H;��H;n�H;��H;��H;��H;|�H;�H;��H;�H;y�H;��H;��H;��H;o�H;��H;b�H;��H;ۉH;[qH;tSH;�.H;�H;�G;v�G;�!G;\XF;��D;#B;n�=;ʄ6;4,;nY;R�	;/�:��:��@:P;9����zp���ܺ�Z�89)�١9�      �EֻV�ѻ��ĻrT�����.o��.�Mܺ��B����8�\:n&�:s��:6Q;�);�=5;�:=;"#B;�D;�uF;�6G;��G;\�G;qH;�:H;^H;�zH;��H;b�H;��H;�H;��H;X�H;�H;i�H;,�H;��H;,�H;f�H;�H;T�H;��H;�H;òH;`�H;��H;�zH;^H;�:H;rH;\�G;��G;�6G;�uF;~�D;#B;�:=;=5;�);7Q;s��:j&�:�\:���8��B�Mܺ�.��.o���vT����ĻR�ѻ      SFB�>�>���4�V�$�u��[�����ݎ�lA?�|Ӻp���x3�9�q�:HX�:T;��';|=5;u�=;��B;GE;L�F;�UG;!�G;��G;VH;�HH;jH;�H;x�H;D�H;0�H;D�H;��H;@�H;�H;�H;��H;�H;�H;:�H;��H;A�H;0�H;G�H;u�H;�H;jH;�HH;PH;��G; �G;UG;B�F;GE;��B;q�=;~=5;��';R;JX�:�q�:X3�9x���|ӺlA?��ݎ����[�x��W�$���4�=�>�      iy��@ݜ��A���I����s���P��%+������Ļ����>|�0�o��9u9IX�:�+�:T;�);Ʉ6;s�>;�PC;d�E;��F;�xG;(�G;zH;b1H;XH;�vH;��H;�H;��H;z�H;�H;?�H;~�H;��H;��H;��H;}�H;>�H;�H;v�H;��H;�H;��H;�vH;XH;^1H;tH;)�G;�xG;��F;[�E;�PC;p�>;Ƅ6;�);N;�+�:CX�:�9u98�o�@|�������Ļ����%+���P���s��I���A��@ݜ�      n�����W�͖ռ�վ�+Ϥ��I����[�	(��Z����9��{��0;9IX�:RX�:7Q;4,;��8;�A@;BD;�@F;�,G;��G;��G;dH;�DH;hH;0�H;R�H;e�H;[�H;�H;�H;��H;��H;a�H;��H;��H;�H;�H;W�H;c�H;U�H;.�H;hH;�DH;^H;��G;��G;�,G;�@F;BD;�A@;��8;4,;7Q;FX�:CX�: ;9�{����9���Z�
(���[��I��+Ϥ��վ�͖ռ�W���      3�6�G�3���+���a�j�����μ���{���TFB�is�ET��0�D��{��@:u9�q�:o��:sY;�t0;��;;�B;�9E;�F;�gG;ٿG;��G;u0H;�XH;*xH; �H;u�H;��H;��H;��H;�H;+�H;0�H;+�H;�H;��H;�H;��H;s�H;#�H;)xH;�XH;s0H;��G;ҿG;�gG;�F;�9E;�B;��;;�t0;oY;o��:�q�: :u9�{��4�D�FT��is�UFB�z��������μj���c�����+�G�3�      p₽�؀���u��Xc���K�x1�������վ��]����P����ET����9��o�p3�9j&�:S�	;U%;F�5;��>;��C;�F;�!G;��G;��G;@H;[HH;�kH;��H;J�H;��H;��H;t�H;H�H;��H;��H;��H;E�H;r�H;��H;��H;G�H;��H;�kH;XHH;=H;��G;��G;�!G;�F;��C;��>;F�5;R%;S�	;h&�:X3�9(�o���9�FT�������P��]���վ�����x1���K��Xc���u��؀�      8S���r��r�����ѓ����u���N���(��i�ˌ˼�A����P�is��@|������\:�:i�;un-;�:;�A;z,E;f�F;(oG;��G;�H;�7H;:_H;~H;�H;��H;q�H;�H;v�H;8�H;�H;9�H;t�H;
�H;o�H;��H;�H;	~H;:_H;�7H;�H;��G;#oG;g�F;y,E;�A;؞:;un-;f�;�:�\:����C|��js���P��A��̌˼�i���(���N���u�ғ�����r���r��      �o��s��罬�ս5@��qĥ�x^���Xc�D�3���	�ˌ˼�]��UFB� [򻲜��|Ӻ ��8��:՛;�M#;q=5;?;I�C;x@F;:G;�G;�G;*'H;�RH;wtH;��H;w�H;(�H;��H;��H;��H;<�H;��H;��H;��H;&�H;t�H;��H;wtH;�RH;*'H;�G;�G; :G;w@F;K�C;?;g=5;�M#;қ;��: ��8�Ӻ����[�UFB��]��ˌ˼��	�D�3��Xc�x^��qĥ�6@����ս���s�      �#�U� �`'������gٽ7S��'l��N�j�D�3��i��վ�{���
(���ĻhA?���B���@:�[�:Q;�.;��;;xtB;�E;}�F;!�G;��G;�H;QFH;"kH;��H;�H;�H;e�H;�H;n�H;��H;l�H;�H;d�H;�H;�H;��H;#kH;OFH;�H;��G;"�G;{�F;�E;xtB;��;;��.;	Q;�[�:��@:��B�jA?���Ļ
(�{����վ��i�D�3�N�j�'l��8S���gٽ����`'�U� �      �S�'�O��E��5�U� �X�
���罥9��(l���Xc���(��������[�����ݎ�Wܺ�:9��:)�	;@d';_ 8;8�@;z�D;�F;jG;��G;GH;k:H;=bH;��H;�H;/�H;@�H;x�H;3�H;��H;2�H;z�H;@�H;+�H;��H;��H;CbH;k:H;HH;��G;jG;�F;x�D;6�@;] 8;:d';,�	;��:�:9Tܺ�ݎ������[��������(��Xc�(l���9�����X�
�U� ��5��E�'�O�      �~��*��(�v��9b�z�H�#,�MZ����7S��x^����N������μ�I���%+�����.������j~:;��:&m;��3;�>;7�C;6PF;yFG;J�G;��G;t/H;�YH;rzH;B�H;��H;[�H;�H;&�H;��H;#�H;�H;[�H;�H;A�H;pzH;ZH;u/H;��G;M�G;~FG;6PF;8�C;�>;��3;!m;E��:�j~:�����.�����%+��I����μ�����N�x^��7S�����MZ�#,�z�H��9b�)�v�*��      ����(����:���M��E�r�'�O�#,�X�
��gٽqĥ���u�y1�j���+Ϥ���P�[��.o��p��:U��:�P;4�/;2�<;�
C;�E;g!G;.�G;��G;�%H;�RH;�tH;�H;A�H;ӯH;��H;U�H; �H;U�H;��H;ӯH;@�H;�H;�tH;�RH;�%H;��G;0�G;n!G;�E;�
C;0�<;1�/;�P;Y��::�p���.o�[򻭎P�+Ϥ�j���y1���u�qĥ��gٽX�
�#,�'�O�E�r��M���:��(���      8���v��M;������RP��E�r�z�H�U� ���6@��ѓ����K�b��վ���s�u���񕻹ܺP4u9 &�:�;&�+;t�:;�"B;h�E;��F;͐G;��G;*H;0LH;�oH;6�H;n�H;��H;-�H;ԼH;�H;мH;0�H;��H;n�H;4�H;�oH;8LH;*H;��G;ӐG;��F;g�E;�"B;r�:;%�+;�;&�:@4u9�ܺ��u����s��վ�b���K�ѓ��6@����U� �z�H�E�r�RP������M;���v��      VVھ�*־/5ʾr��������M���9b��5�����ս����Xc���̖ռ�I��X�$�qT���Z��]���:��;a�';�8;RA;�9E;}�F;��G;��G;<H;GH;lH;?�H;5�H;ޫH;��H;��H;M�H;��H;��H;۫H;5�H;?�H;
lH;GH;=H;��G;��G;��F;�9E;RA;�8;`�';��;�:�]���Z�qT��X�$��I��̖ռ���Xc������ս���5��9b��M������r���05ʾ�*־      ���쾳�޾/5ʾM;���:��)�v��E�`'����r����u���+��W��A����4���Ļ(9)��j��kW�:Z�;�%;�k7;�@;��D;��F;�wG;N�G;.H;:CH;&iH;	�H;��H;��H;��H;��H;o�H;��H;��H;��H;��H;�H;!iH;@CH;/H;P�G;�wG;��F;��D;�@;�k7;�%;X�;sW�:�j��&9)���Ļ��4��A���W缄�+���u�r�����`'��E�)�v��:��M;��/5ʾ��޾��      Vh���b���쾧*־�v��(���*��(�O�U� �s��r���؀�H�3���@ݜ�?�>�X�ѻ�9����o�:7% ;jM#;;�6;DA@;��D;��F;qG;F�G;H;�@H;dgH;��H;��H;٩H;�H;��H;ۻH;�H;�H;۩H;��H;��H;^gH;�@H;H;F�G;qG;��F;��D;DA@;5�6;fM#;3% ;o�: ����9�Y�ѻ?�>�@ݜ���H�3��؀��r��s�V� �(�O�*��(����v���*־���b��      ���^�T_ݾ��ɾj*��쫖�{x�&G�P,�����b��^@{���/�����䙼�J;�S�ͻ��4�XW����:.;��#;�6;[@;,�D;��F;�lG;��G;3H;�:H;�bH;ۀH;(�H;*�H;ձH;�H;عH;�H;ԱH;*�H;&�H;׀H;�bH;�:H;2H;��G;�lG;��F;,�D;	[@;�6;��#;,;���:XW���4�R�ͻ�J;��䙼����/�^@{��b�����P,�&G�{x�쫖�j*����ɾT_ݾ^�      ^�3���:پ|�žg�����9t�p�C� �����䪫�X`w�F-����+`����7�:Sɻ�K/�yƹ���:�/;�f$;�7;�~@;D�D;U�F;�nG;��G;H;;H;ecH;l�H;}�H;m�H;�H;*�H;�H;&�H;�H;k�H;|�H;i�H;`cH;�;H;H;��G;�nG;`�F;D�D;�~@;�7;�f$;�/;���:yƹ�K/�:Sɻ��7�+`�����F-�X`w�䪫���� ��p�C�9t���g���|�ž�:پ3��      U_ݾ�:پ�V;+���Ƥ�La����g��$:��Z�pݽ�ƣ�{l�f.%��߼i���9.�д��VV� 2p��@�:x;F(&;+�7;3�@;�
E;��F;duG;�G;KH;�=H;IeH;��H;p�H;I�H;��H;��H;��H;��H;��H;I�H;n�H;��H;CeH;�=H;KH;!�G;euG;��F;�
E;/�@;'�7;D(&;
x;�@�:02p�VV�ϴ���9.�h���߼f.%�{l��ƣ�pݽ�Z��$:���g�La���Ƥ�+���V;�:پ      ��ɾ|�ž+��qת�쫖�!�����T��J+�;��2̽�s���yZ����Oμgy����aϨ�X,� 
�6��:��
;W�(;ON9;��A;wNE;+�F;�G;��G;wH;�AH;-hH;�H;=�H;ѩH;ɳH;��H;t�H;��H;˳H;ЩH;9�H;߄H;)hH;�AH;wH;��G;�G;3�F;wNE;��A;IN9;U�(;��
;��: �6V,�aϨ���gy��Oμ����yZ��s���2̽;��J+���T�!���쫖�qת�+��|�ž      j*��h����Ƥ�쫖��/��>�c��G=�����zｑж��ɇ�R�C���$"��t;k��&��-����˺�X�9d��:9;�h,;�	;;�PB;]�E;� G;،G;��G;dH;	GH;JlH;��H;��H;��H;6�H;�H;ѼH;��H;8�H;��H;��H;��H;FlH;GH;dH;��G;ڌG;� G;^�E;�PB;�	;;�h,;9;n��:�X�9��˺�-���&�s;k�$"����R�C��ɇ��ж��z�����G=�>�c��/��쫖��Ƥ�h���      쫖���La��!���>�c�p�C�z#���SvϽ����{l�eg*����
���I�����\c�퀺�t,:���:�;�_0;_�<;�1C;��E;p#G;O�G;�G; H;�MH;2qH;��H;y�H;٭H;(�H;��H;[�H;��H;(�H;׭H;v�H;��H;1qH;�MH; H;�G;O�G;w#G;��E;�1C;\�<;�_0;�;���:�t,:퀺�\c�����I��
�����eg*�{l�����RvϽ��z#�p�C�>�c�!���La����      {x�9t���g���T��G=�z#�6�oݽ�b������BG������Ǽiy��M�$�i���(�$�vƹ?��:�&�:�� ;E4;o�>;HD;�[F;�FG;|�G;��G;�)H;ZUH;�vH;��H;�H;~�H;h�H;��H;'�H;~�H;h�H;~�H;�H;�H;�vH;bUH;�)H; �G;z�G;�FG;�[F;HD;l�>;F4;�� ;�&�:?��: vƹ$�$�j���L�$�iy����Ǽ���BG������b��oݽ6�z#��G=���T���g�9t�      &G�p�C��$:��J+� ����oݽ^���.I���yZ��"����ԫ��fT��� � M����˺�m9)ٶ:^�;`(;�8;_�@;��D;رF;:hG;{�G;~H;+5H;�]H;a}H;�H;��H;P�H;ĻH;��H;2�H;��H;ȻH;R�H;��H;�H;_}H;�]H;-5H;�H;|�G;@hG;ܱF;��D;_�@;	�8;`(;e�;)ٶ: m9��˺ M���� �eT�ԫ������"��yZ�.I��]���pݽ�� ���J+��$:�p�C�      P,�����Z�;��z�SvϽ�b��.I��g]a�G-�h� �""��y�{�H�!�������4��P(��nQ:�L�:��;Ί/;�'<;՟B;��E;��F;��G;��G;.H;8AH;gH;I�H;0�H;̪H;��H;{�H;��H;O�H;��H;�H;��H;ȪH;/�H;J�H;gH;<AH;2H;��G;��G;��F;��E;؟B;�'<;ϊ/;��;�L�:�nQ:�P(���4�����G�!�y�{�""��i� �G-�f]a�-I���b��RvϽ�z�:��Z����      ������pݽ�2̽�ж����������yZ�G-�ַ�/aļZO���J;���軅�|���º�M@9���:6�;�f$;��5;�N?;3D;�LF;�:G;��G;��G;�!H;�MH;�pH;��H;͟H;,�H;�H;<�H;p�H;��H;p�H;?�H;�H;)�H;ɟH;��H;�pH;�MH;�!H;��G;��G;�:G;�LF;7D;�N?;��5;�f$;7�;���: N@9��º��|�����J;�ZO��/aļַ�G-��yZ����������ж��2̽pݽ���      �b��䪫��ƣ��s���ɇ�{l�BG��"�i� �0aļc���I��C��ۙ�L�puƹ*�k:���:�;6>.;
;;��A;�AE;X�F;mG;��G;��G;Q2H;�ZH;�zH;ҒH;��H;��H;U�H;)�H;��H;�H;��H;*�H;X�H;��H;��H;ӒH;�zH;�ZH;T2H;��G;��G;mG;X�F;�AE;��A;
;;B>.;�;���:B�k:`uƹI��ۙ��C��I�c��/aļh� ��"�BG�{l��ɇ��s���ƣ�䪫�      ]@{�X`w�zl��yZ�R�C�eg*�������#"��ZO���I�@|�>Ϩ�vK/��$T�Q:B��:��;�(&;�#6;�%?;|�C;l#F;�#G;�G;��G;�H;%CH;�gH;y�H;T�H;h�H;�H;��H;�H;�H;��H;�H;�H;��H;�H;c�H;V�H;��H;�gH;&CH;�H;��G;�G;�#G;s#F;��C;�%?;�#6;�(&;��;P��:Q:�$T�rK/�=Ϩ�?|��I�ZO��""����鼮��dg*�S�C��yZ�zl�X`w�      ��/�F-�f.%����
�������Ǽӫ��y�{��J;��C�>Ϩ�RO:� �[�9���:h;|�;3.1;�'<;�5B;�NE;�F;,fG;޹G;*�G;�*H;�SH;�tH;�H;��H;�H;I�H;u�H;��H;��H;�H;��H;��H;v�H;H�H;�H;��H;$�H;�tH;�SH;�*H;&�G;�G;-fG;�F;�NE;�5B;(<;:.1;x�;n;���: [�9����PO:�<Ϩ��C��J;�x�{�ҫ����Ǽ��������f.%�F-�      ������߼Pμ""���
��iy��eT�H�!�����ۙ�yK/�
�Pm9�A�:���:(�;<�,;�N9;9@;�^D;�LF;P.G;ޗG;��G;�H;�?H;dH;�H;j�H;�H;��H;��H;��H;��H;��H;u�H;��H;��H;��H;��H;��H;�H;t�H;�H;dH;�?H;�H;��G;ߗG;V.G;�LF;�^D;B@;�N9;9�,;/�;���:�A�:�m9�tK/��ۙ����F�!�cT�iy���
��$"��Qμ�߼���      �䙼,`��j��hy��r;k��I�L�$��� �������|�H��$T��Z�9�A�:V��:�;�);#7;��>;�tC;�E;��F;�uG;�G;��G;�+H;�SH;�sH;|�H;]�H;�H;ȻH;��H;3�H;m�H;��H;��H;��H;k�H;4�H;��H;ŻH;
�H;b�H;��H;�sH;�SH;�+H;��G;�G;�uG;��F;�E;�tC;��>;7;�);�;V��:�A�:[�9�$T�D���|������� �L�$��I�v;k�hy��j��+`��      �J;���7��9.����&����d���M����4���ºXuƹQ:���:���:�;��(;��5;��=;��B;�[E;=�F;�TG;��G;��G;�H;�CH;fH;āH;q�H;�H;��H;��H;��H;R�H;��H;;�H;�H;:�H;��H;Q�H;��H;��H;��H;��H;v�H;ǁH;fH;�CH;�H;��G;��G;�TG;C�F;�[E;��B;��=;��5;��(;�;���:���:Q:Huƹ��º��4�M��f�����軭&����9.���7�      N�ͻ8Sɻմ��dϨ��-���\c�"�$���˺�P(�`N@9F�k:D��:l;,�;�);��5;C�=;#QB;dE;�F; 8G;=�G;>�G;�	H;Q5H;�YH;=wH;ӎH;��H;ΰH;��H;��H;Q�H;�H;~�H;r�H;�H;n�H;|�H; �H;M�H;��H;��H;ѰH;��H;ՎH;>wH;�YH;W5H;�	H;>�G;A�G;"8G;�F;hE;QB;E�=;��5;�);.�;l;J��:N�k:PN@9�P(���˺&�$��\c��-��hϨ�ڴ��3Sɻ      ��4��K/�\V�N,�h�˺퀺�uƹ0m9�nQ:���:���:��;t�;9�,;7;��=;QB;��D;~cF;$G;ƇG;��G;��G;t)H;�NH;�mH;؆H;��H;!�H;�H;�H;��H;��H;��H;��H;u�H;�H;r�H;��H;��H;��H;��H;�H;�H;#�H;��H;؆H;�mH;�NH;s)H;��G;��G;ʇG;$G;�cF;��D;QB;��=;7;7�,;u�;��;���:���:�nQ:�m9�uƹ퀺c�˺V,�TV��K/�      �VṐyƹ@2p� �6�X�9�t,:Q��:3ٶ:�L�:9�;�;�(&;7.1;�N9;��>;��B;eE;�cF;�G;%�G;��G;��G;Q H;�EH;�eH;�H;��H;ΥH;��H;��H;	�H;��H;��H;O�H;��H;G�H;��H;D�H;��H;N�H;��H;��H;�H;��H;��H;ХH;��H;�H;�eH;�EH;M H;��G;��G;)�G;�G;�cF;hE;��B;��>;�N9;7.1;�(&;�;9�;�L�:5ٶ:M��:�t,:�X�9 ��6P2p��yƹ      笊:���:�@�:��:^��:���:�&�:^�;��;�f$;@>.;�#6;�'<;@@;�tC;�[E;�F;!$G;'�G;��G;�G;�H;�?H;�_H;�yH;Z�H;�H;��H;-�H;s�H;��H;L�H;o�H;��H;��H;��H;d�H;��H;��H;��H;m�H;G�H;��H;s�H;-�H;��H;�H;V�H;�yH;�_H;�?H;�H;�G;��G;*�G;$G;�F;�[E;�tC;<@;�'<;�#6;@>.;�f$;��;e�;�&�:���:f��::�@�:{��:      P;�/;�w;�
;�8;�;�� ;�_(;̊/;��5;
;;�%?;�5B;�^D;�E;B�F; 8G;ӇG;��G;�G;�H;�<H;�[H;�uH;�H;Q�H;5�H;;�H;��H;��H;��H;g�H;�H;��H;y�H;}�H;��H;v�H;y�H;��H;�H;a�H;��H;��H;��H;:�H;3�H;P�H;��H;�uH;�[H;�<H;�H;�G;��G;͇G;!8G;@�F;�E;�^D;�5B;�%?;
;;��5;ʊ/;�_(;�� ;�;9;�
;�w;�/;      ��#;�f$;R(&;_�(;�h,;�_0;B4;�8;�'<;�N?;��A;|�C;�NE;�LF;��F;�TG;>�G;��G;��G;�H;�<H;jZH;�sH;��H;��H;��H;еH;ƿH;��H;�H;9�H;2�H;Q�H;u�H;��H;��H;�H;��H;��H;u�H;N�H;,�H;;�H;�H;��H;ƿH;˵H;��H;��H;�H;�sH;jZH;�<H;�H;��G;��G;@�G;�TG;��F;�LF;�NE;}�C;��A;�N?;�'<;�8;F4;�_0;�h,;T�(;D(&;{f$;      %�6;�7;&�7;\N9;�	;;d�<;�>;i�@;ߟB;;D;�AE;s#F;�F;^.G;�uG;��G;C�G;��G;Q H;�?H;�[H;�sH;3�H;T�H;�H;&�H;��H;"�H;��H;!�H;M�H;��H;A�H;,�H;;�H;��H;.�H;��H;9�H;.�H;>�H;��H;O�H;!�H;��H;$�H;��H;&�H;�H;Q�H;.�H;�sH;�[H;�?H;Q H;��G;A�G;��G;�uG;W.G;�F;t#F;�AE;4D;ݟB;i�@;}�>;a�<;�	;;YN9;#�7;y7;      [@;�~@;$�@;�A;�PB;�1C;KD;��D;�E;�LF;\�F;�#G;-fG;�G;�G;��G;�	H;{)H;�EH;�_H;�uH;��H;Q�H;`�H;7�H;�H;&�H;��H;P�H;��H;�H;��H;��H;h�H;h�H;��H;@�H;��H;e�H;h�H;��H;��H;�H;��H;N�H;��H; �H;�H;:�H;]�H;M�H;�H;�uH;�_H;�EH;s)H;�	H;��G;�G;ޗG;*fG;�#G;\�F;�LF;�E;��D;KD;�1C;�PB;�A;'�@;�~@;      N�D;@�D;�
E;mNE;W�E;��E;�[F;رF;��F;�:G;mG;!�G;�G;��G;��G;�H;[5H;�NH;�eH;�yH;��H;��H;�H;>�H;��H;��H;&�H;��H;��H;w�H;O�H;��H;P�H;y�H;x�H;��H;�H;��H;w�H;z�H;N�H;��H;R�H;w�H;��H;��H;�H;��H;��H;;�H;�H;��H;��H;�yH;�eH;�NH;[5H;�H;��G;��G;�G;$�G;mG;�:G;��F;رF;�[F;��E;`�E;gNE;�
E;@�D;      ��F;Y�F;��F;(�F;� G;x#G;�FG;HhG;��G;��G;��G;��G;-�G;�H;�+H;�CH;�YH;�mH;�H;U�H;P�H;��H; �H;�H;��H;��H;1�H;��H;�H;�H;Z�H;�H;��H;}�H;\�H;��H;��H;��H;Y�H;}�H;��H; �H;Z�H;�H;�H;��H;*�H;��H;��H;�H; �H;��H;P�H;R�H;�H;�mH;�YH;�CH;�+H;�H;,�G;��G;��G;��G;��G;IhG;�FG;m#G;� G;2�F;��F;\�F;      �lG;�nG;cuG;�G;ΌG;K�G;��G;x�G;��G;��G;��G;�H;�*H;�?H;�SH;fH;AwH;݆H;��H;�H;:�H;͵H;��H;(�H;%�H;1�H;Q�H;��H;��H;'�H;�H;g�H;��H;m�H;��H;\�H;x�H;U�H;��H;n�H;��H;b�H;�H;&�H;��H;��H;I�H;3�H;&�H;!�H;��H;εH;:�H;�H;��H;ֆH;AwH;fH;�SH;�?H;�*H;�H;��G;��G;��G;z�G;��G;E�G;�G;�G;duG;�nG;      ��G;��G;�G;��G;��G;�G;�G;~H;4H;�!H;V2H;,CH;�SH;dH;�sH;ƁH;ӎH;��H;ХH;��H;<�H;ſH;�H;��H;��H;��H;��H;��H;�H;��H;b�H;��H;r�H;6�H;|�H;��H;�H;��H;|�H;7�H;r�H;��H;b�H;��H;�H;��H;��H;��H;��H;��H;�H;ĿH;:�H;��H;ͥH;��H;ӎH;ǁH;�sH;dH;�SH;*CH;Y2H;�!H;2H;~H;�G;��G;��G;��G;�G;��G;      -H;H;GH;�H;UH;
 H;�)H;'5H;2AH;�MH;�ZH;�gH;�tH;�H;��H;t�H;��H;(�H;��H;,�H;��H;��H;��H;M�H;��H;�H;��H;�H;��H;J�H;p�H;��H;3�H;��H;�H;L�H;V�H;F�H;�H;��H;4�H;��H;q�H;I�H;��H;�H;��H;�H;��H;G�H;��H;��H;��H;)�H;��H;#�H;��H;u�H;��H;�H;�tH;�gH;�ZH;�MH;4AH;&5H;�)H; H;^H;�H;GH;H;      �:H;x;H;�=H;�AH;GH;�MH;_UH;�]H;gH;�pH;�zH;��H;"�H;t�H;`�H;�H;ӰH;�H;��H;o�H;��H;�H;�H;��H;v�H;�H;$�H;��H;I�H;��H;i�H;(�H;��H;1�H;��H;��H;��H;��H;��H;0�H;��H;#�H;i�H;��H;I�H;��H;�H;�H;w�H;��H;�H;�H;��H;l�H;��H;�H;ӰH;�H;`�H;q�H;"�H;��H;�zH;�pH;gH;�]H;_UH;�MH;GH;�AH;�=H;v;H;      �bH;vcH;MeH;.hH;IlH;5qH;�vH;b}H;L�H;��H;ܒH;]�H;áH;�H;�H;��H;��H;�H;�H;��H;��H;:�H;M�H;�H;P�H;X�H;�H;g�H;s�H;n�H;;�H;��H;&�H;��H;��H;��H;�H;��H;��H;��H;)�H;��H;:�H;k�H;q�H;b�H;�H;[�H;S�H;�H;O�H;:�H;��H;��H;�H;�H;��H;��H;�H;�H;ġH;`�H;ܒH;��H;O�H;e}H;wH;+qH;SlH;-hH;NeH;ycH;      ڀH;p�H;��H;ۄH;��H;��H;��H;�H;5�H;ϟH;��H;n�H;!�H;��H;˻H;��H;��H;��H;��H;N�H;k�H;0�H;��H;��H;��H; �H;b�H;��H;��H;)�H;��H;;�H;��H;��H;�H;8�H;+�H;8�H;�H;��H;��H;8�H;��H;(�H;��H;��H;a�H;�H;��H;��H;��H;2�H;e�H;J�H;��H;��H;��H;��H;ͻH;��H;!�H;n�H;��H;ϟH;5�H;�H;�H;��H;�H;݄H;ȂH;w�H;      )�H;��H;|�H;=�H;��H;v�H;�H;��H;ǪH;-�H;��H;�H;Q�H;��H;��H;��H;T�H;��H;��H;s�H;�H;Q�H;<�H;��H;P�H;��H;��H;x�H;7�H;��H;%�H;��H;��H;�H;P�H;a�H;.�H;a�H;M�H;�H;��H;��H;#�H;��H;6�H;u�H;��H;��H;S�H;��H;A�H;O�H;�H;o�H;��H;��H;V�H;��H;��H;��H;Q�H;�H;��H;/�H;ʪH;��H;�H;r�H;��H;7�H;��H;��H;      *�H;h�H;L�H;ʩH;��H;ЭH;��H;U�H;��H;�H;c�H;��H;��H;��H;:�H;X�H;$�H;��H;R�H;��H;��H;u�H;'�H;^�H;u�H;x�H;g�H;7�H;��H;3�H;��H;��H;�H;G�H;f�H;m�H;��H;l�H;c�H;G�H;�H;��H;��H;.�H;��H;3�H;f�H;z�H;w�H;]�H;,�H;s�H;��H;��H;Q�H;��H;(�H;X�H;:�H;��H;~�H;��H;e�H;��H;��H;Y�H;��H;ЭH;��H;ʩH;V�H;u�H;      ұH;�H;��H;ͳH;I�H;"�H;t�H;ȻH;��H;I�H;3�H;%�H;��H;��H;t�H;��H;��H;��H;��H;��H;|�H;��H;2�H;X�H;q�H;R�H;��H;y�H;�H;��H;��H;�H;P�H;h�H;o�H;�H;��H;��H;l�H;h�H;Q�H;�H;��H;��H;�H;u�H;��H;T�H;s�H;X�H;9�H;��H;v�H;��H;��H;��H;��H;��H;r�H;��H;��H;&�H;8�H;J�H;��H;̻H;w�H;%�H;G�H;гH;��H;�H;      �H;)�H;��H;��H;�H;��H;��H;��H;��H;{�H;�H;��H;�H;��H;��H;:�H;r�H;r�H;G�H;��H;~�H;��H;��H;��H;��H;��H;V�H;��H;M�H;��H;��H;=�H;f�H;q�H;��H;��H;��H;��H;��H;v�H;i�H;<�H;��H;��H;J�H;��H;W�H;��H;��H;��H;��H;��H;x�H;��H;F�H;u�H;w�H;<�H;��H;��H;�H;��H;�H;~�H; �H;��H;��H;��H;�H;��H;��H;7�H;      ߹H;�H;̺H;r�H;μH;]�H;0�H;6�H;W�H;��H;�H;��H;(�H;��H;��H;!�H;%�H;�H;��H;h�H;��H;�H;*�H;5�H;�H;��H;t�H;�H;X�H;��H;�H;/�H;/�H;��H;��H;��H;��H;��H;��H;��H;4�H;.�H;�H;��H;T�H;�H;t�H;��H;�H;5�H;0�H;�H;��H;d�H;��H;�H;%�H;#�H;��H;��H;(�H;��H;�H;��H;[�H;:�H;4�H;]�H;мH;q�H;κH;'�H;      �H;,�H;��H;��H;�H;��H;��H;��H;��H;}�H;�H;��H;�H;��H;��H;:�H;r�H;r�H;G�H;��H;�H;��H;��H;��H;��H;��H;V�H;��H;O�H;��H;��H;=�H;h�H;s�H;��H;��H;��H;��H;��H;t�H;i�H;<�H;��H;��H;J�H;��H;V�H;��H;��H;��H;��H;��H;x�H;��H;F�H;u�H;u�H;<�H;��H;��H;�H;��H;�H;}�H; �H;��H;��H;��H;�H;��H;��H;4�H;      ʱH;�H;��H;ųH;I�H;!�H;v�H;˻H;��H;J�H;5�H;%�H;��H;��H;u�H;��H;��H;��H;��H;��H;}�H;��H;2�H;X�H;s�H;Q�H;��H;y�H;�H;��H;��H;�H;N�H;h�H;o�H;��H;��H;��H;m�H;i�H;T�H;�H;��H;��H;�H;t�H;��H;V�H;q�H;W�H;9�H;��H;u�H;��H;��H;��H;��H;��H;r�H;��H;��H;(�H;5�H;J�H;��H;һH;{�H;�H;J�H;ƳH;��H;�H;      *�H;h�H;L�H;ΩH;��H;ԭH;��H;W�H;��H;�H;e�H;��H;~�H;��H;;�H;V�H;'�H;��H;R�H;��H;��H;w�H;'�H;`�H;y�H;x�H;i�H;7�H;��H;3�H;��H;��H;�H;G�H;e�H;l�H;��H;m�H;e�H;G�H;�H;��H;��H;0�H;��H;3�H;f�H;{�H;v�H;Z�H;.�H;v�H;��H;��H;R�H;��H;'�H;Y�H;;�H;��H;~�H;��H;c�H;�H;��H;\�H;��H;ѭH;��H;ʩH;V�H;j�H;      *�H;��H;|�H;:�H;��H;y�H;�H;��H;ȪH;/�H;��H;�H;Q�H;��H;��H;��H;S�H;��H;��H;s�H;�H;R�H;:�H;��H;U�H;��H;��H;x�H;:�H;��H;#�H;��H;��H;�H;N�H;b�H;/�H;b�H;N�H;�H;��H;��H;#�H;��H;2�H;t�H;��H;��H;P�H;��H;C�H;O�H;�H;p�H;��H;��H;V�H;��H;��H;��H;S�H;�H;��H;/�H;̪H;��H;�H;v�H;��H;A�H;��H;��H;      ̀H;w�H;��H;ڄH;��H;��H;�H;�H;2�H;͟H;��H;m�H; �H;��H;ͻH;��H;��H;��H;��H;M�H;l�H;3�H;��H;��H;��H; �H;a�H;��H;��H;(�H;��H;:�H;��H;��H;�H;6�H;-�H;8�H;�H;��H;��H;:�H;��H;&�H;��H;��H;^�H;�H;��H;��H;��H;3�H;d�H;J�H;��H;��H;��H;��H;̻H;��H;!�H;n�H;��H;ПH;7�H;�H;�H;��H;��H;ۄH;��H;o�H;      �bH;vcH;PeH;*hH;OlH;5qH;�vH;a}H;M�H;��H;ڒH;`�H;áH;�H;�H;��H;��H;�H;�H;��H;��H;=�H;K�H;�H;S�H;U�H;�H;d�H;v�H;m�H;:�H;��H;&�H;��H;��H;��H;�H;��H;��H;��H;*�H;��H;:�H;j�H;o�H;a�H;�H;[�H;P�H;�H;R�H;=�H;��H;��H;�H;�H;��H;��H;�H;�H;áH;b�H;ڒH;��H;M�H;h}H; wH;2qH;XlH;8hH;XeH;xcH;      �:H;};H;�=H;�AH;GH;�MH;^UH;�]H;gH;�pH;�zH;��H;"�H;r�H;b�H;�H;ѰH;�H;��H;o�H;��H;�H;�H;��H;y�H;�H;!�H;��H;L�H;��H;i�H;(�H;��H;1�H;��H;��H;��H;��H;��H;1�H;��H;&�H;i�H;��H;F�H;��H; �H;�H;v�H;��H;"�H;�H;��H;l�H;��H;�H;ӰH;�H;b�H;r�H;"�H;��H;�zH;�pH;gH;�]H;bUH;�MH;GH;�AH;�=H;v;H;      :H;H;YH;�H;LH; H;�)H;'5H;;AH;�MH;�ZH;�gH;�tH;�H;��H;u�H;��H;)�H;��H;*�H;��H;��H;��H;L�H;��H;
�H;��H;�H;��H;H�H;p�H;��H;4�H;��H;�H;J�H;V�H;I�H;�H;��H;6�H;��H;q�H;I�H;��H;�H;��H;�H;��H;F�H;��H;��H;��H;*�H;��H;#�H;��H;u�H;��H;�H;�tH;�gH;�ZH;�MH;9AH;-5H;*H; H;^H;~H;YH;H;      ��G;��G;�G;��G;��G;�G;�G;�H;2H;�!H;V2H;(CH;�SH;dH;�sH;ǁH;ӎH;ÚH;ͥH;��H;>�H;ƿH;�H;��H;��H;��H;��H;��H;�H;��H;d�H;��H;q�H;7�H;{�H;��H;�H;��H;{�H;7�H;u�H;��H;d�H;��H;�H;��H;��H;��H;��H;��H;$�H;ĿH;8�H;��H;ΥH;��H;ՎH;ǁH;�sH;dH;�SH;*CH;X2H;�!H;4H;H;�G;�G;��G;��G;�G;��G;      �lG;�nG;`uG;�G;܌G;S�G;��G;{�G;��G;��G;��G;�H;�*H;�?H;�SH;fH;AwH;݆H;��H;�H;:�H;εH;��H;(�H;%�H;-�H;M�H;��H;��H;$�H;�H;h�H;��H;m�H;��H;W�H;x�H;W�H;��H;n�H;��H;e�H;�H;&�H;��H;��H;M�H;5�H;&�H;$�H;��H;еH;8�H;�H;��H;؆H;AwH;fH;�SH;�?H;�*H;�H;��G;��G;��G;�G;��G;N�G;�G;�G;euG;�nG;      ~�F;\�F;��F;(�F;� G;#G;�FG;KhG;��G;��G;��G;��G;-�G;�H;�+H;�CH;�YH;�mH;�H;P�H;Q�H;��H;�H;�H;��H;��H;-�H;��H;�H;�H;X�H;�H;��H;~�H;\�H;��H;��H;��H;[�H;~�H;��H;�H;\�H;�H;�H;��H;.�H;��H;��H;�H;#�H;��H;P�H;U�H;�H;�mH;�YH;�CH;�+H;�H;.�G;��G;��G;��G;��G;GhG;�FG;p#G;� G;&�F;��F;K�F;      L�D;=�D;�
E;nNE;W�E;��E;�[F;رF;��F;�:G;mG;"�G;�G;��G;��G;�H;Z5H;�NH;�eH;�yH;��H;��H;�H;>�H;��H;��H;!�H;��H;��H;s�H;P�H;��H;N�H;y�H;z�H;��H;�H;��H;x�H;|�H;P�H;��H;U�H;w�H;��H;��H;#�H;��H;��H;;�H;�H;��H;��H;�yH;�eH;�NH;\5H;�H;��G;��G;�G;$�G;mG;�:G;��F;ڱF;�[F;��E;`�E;jNE;�
E;=�D;      �Z@;�~@;!�@;��A;�PB;�1C;LD;��D;��E;�LF;^�F;�#G;)fG;��G;�G;��G;�	H;x)H;�EH;�_H;�uH;��H;L�H;`�H;;�H;�H;!�H;��H;P�H;��H;�H;��H;��H;h�H;g�H;��H;@�H;��H;e�H;g�H;��H;��H;�H;��H;P�H;��H;$�H;�H;9�H;a�H;Q�H;�H;�uH;�_H;�EH;v)H;�	H;��G;�G;��G;*fG;�#G;^�F;�LF;��E;��D;KD;�1C;�PB;�A; �@;�~@;      �6;�7;�7;cN9;�	;;a�<;w�>;f�@;��B;7D;�AE;s#F;�F;Z.G;�uG;��G;A�G;��G;P H;�?H;�[H;�sH;.�H;T�H;�H;�H;��H;!�H;��H;�H;N�H;��H;?�H;,�H;;�H;��H;1�H;��H;9�H;+�H;?�H;��H;R�H;"�H;��H;!�H;��H;&�H;�H;S�H;1�H;�sH;�[H;�?H;T H;��G;C�G;��G;�uG;W.G;�F;s#F;�AE;8D;��B;j�@;x�>;`�<;�	;;^N9;�7;7;      ��#;�f$;H(&;W�(;�h,;�_0;H4;�8;�'<;�N?;��A;��C;�NE;�LF;��F;�TG;>�G;��G;��G;�H;�<H;jZH;�sH;��H;��H;��H;͵H;ƿH;��H;�H;;�H;2�H;O�H;u�H;��H;��H;�H;��H;��H;s�H;Q�H;0�H;>�H;�H;��H;ƿH;εH;��H;��H;��H;�sH;kZH;�<H;�H;��G;��G;=�G;�TG;��F;�LF;�NE;�C;��A;�N?;�'<;�8;A4;�_0;�h,;K�(;H(&;{f$;      F;�/;x;�
;�8;�;�� ;�_(;ϊ/;��5;
;;�%?;�5B;�^D;�E;C�F;!8G;ЇG;��G;�G;�H;�<H;�[H;�uH;��H;N�H;1�H;8�H;��H;��H;��H;g�H;�H;��H;y�H;x�H;��H;z�H;w�H;��H;�H;e�H;��H;��H;��H;8�H;5�H;Q�H;��H;�uH;�[H;�<H;�H;�G;��G;̇G; 8G;B�F;�E;�^D;�5B;�%?;
;;��5;Ί/;`(;�� ;�;9;�
;x;�/;      ��:���:�@�:��:b��:���:�&�:h�;��;�f$;D>.;�#6;�'<;>@;�tC;�[E;�F;$G;'�G;��G;�G;�H;�?H;�_H;�yH;U�H;�H;��H;-�H;n�H;��H;L�H;q�H;��H;��H;��H;e�H;��H;��H;��H;o�H;J�H;��H;r�H;,�H;��H;�H;W�H;�yH;�_H;�?H;�H;�G;��G;)�G;$G;�F;�[E;�tC;>@;�'<;�#6;B>.;�f$;��;a�;�&�:���:n��:��:�@�:���:      �V�xyƹ02p� �6�X�9�t,:M��:3ٶ:�L�:9�;�;�(&;7.1;�N9;��>;��B;dE;�cF;�G;'�G;��G;��G;S H;�EH;�eH;�H;��H;ͥH;��H;��H;	�H;��H;��H;Q�H;��H;F�H;��H;F�H;��H;N�H;��H;��H;�H;��H;��H;ͥH;��H;�H;�eH;�EH;Q H;��G;��G;)�G;�G;�cF;eE;��B;��>;�N9;6.1;�(&;�;7�;�L�:7ٶ:Q��:�t,:�X�9 �6�2p�`yƹ      ��4��K/�`V�P,�`�˺퀺�uƹ�m9�nQ:���:���:��;v�;9�,; 7;��=;QB;��D;cF;$G;ɇG;��G;��G;t)H;�NH;�mH;ӆH;��H;%�H;�H;�H;��H;��H;��H;��H;s�H;�H;u�H;��H;��H;��H;��H;�H;�H;#�H;��H;؆H;�mH;�NH;t)H;��G;��G;ƇG;$G;~cF;��D;QB;��=; 7;6�,;t�;��;���:���:�nQ:�m9�uƹ퀺h�˺U,�hV��K/�      M�ͻ8SɻԴ��bϨ��-���\c�$�$���˺�P(�`N@9J�k:L��:l;,�;�);��5;F�=;QB;dE;�F;%8G;@�G;A�G;�	H;X5H;�YH;=wH;юH;��H;ͰH;��H;��H;P�H;!�H;~�H;r�H;�H;r�H;|�H;�H;M�H;��H;��H;аH;��H;юH;>wH;�YH;S5H;�	H;A�G;>�G;8G;�F;dE;QB;C�=;��5;�);,�;l;H��:J�k:@N@9�P(���˺'�$��\c��-��fϨ�ٴ��4Sɻ      �J;���7��9.����&����d���M����4���º@uƹ Q:���:���:�;��(;��5;��=;��B;�[E;D�F;�TG;��G;��G;�H;�CH;fH;āH;u�H;�H;��H;��H;��H;T�H;��H;:�H;�H;8�H;��H;O�H;��H;��H;��H;�H;t�H;āH;fH;�CH;�H;��G;��G;�TG;;�F;�[E;��B;��=;��5;��(;�;���:���:Q:Puƹ��º��4�M��h�����軭&����9.���7�      �䙼+`��k��gy��r;k��I�L�$��� �������|�F��$T�[�9�A�:^��:�;�); 7;��>;�tC;�E;��F;�uG;�G;��G;�+H;�SH;�sH;��H;^�H;�H;ȻH;��H;6�H;m�H;��H;��H;��H;h�H;3�H;��H;ĻH;
�H;^�H;��H;�sH;�SH;�+H;��G;�G;�uG;��F;�E;�tC;��>;7;�);�;V��:�A�:�Z�9�$T�H���|������� �L�$��I�v;k�iy��j��+`��      ������߼Pμ""���
��iy��cT�F�!���軿ۙ�tK/���m9�A�:���:,�;7�,;�N9;<@;�^D;�LF;V.G;�G;��G;�H;�?H;dH;�H;m�H;�H;��H;��H;��H;��H;��H;u�H;��H;��H;��H;��H;��H;�H;q�H;�H;dH;�?H;�H;��G;��G;X.G;�LF;�^D;?@;�N9;7�,;+�;��:�A�:`m9�uK/��ۙ����G�!�cT�iy���
��$"��Pμ�߼���      ��/�F-�f.%����
�������Ǽӫ��y�{��J;��C�=Ϩ�PO:�����0[�9���:j;y�;6.1;�'<;�5B;�NE;�F;0fG;�G;*�G;�*H;�SH;�tH;�H;��H;�H;I�H;y�H;��H;��H;�H;��H;��H;u�H;F�H;�H;��H;!�H;�tH;�SH;�*H;&�G;ܹG;,fG;�F;�NE;�5B;�'<;3.1;u�;j;���: [�9����RO:�>Ϩ��C��J;�x�{�ӫ����Ǽ��������g.%�F-�      ^@{�X`w�zl��yZ�R�C�eg*�������""��ZO���I�?|�=Ϩ�tK/��$T�Q:H��:��;�(&;�#6;�%?;�C;s#F;�#G;�G;��G;�H;%CH;�gH;z�H;X�H;e�H;�H;��H;�H;|�H;��H;~�H;�H;��H;�H;d�H;U�H;}�H;�gH;"CH;�H;��G;�G;�#G;s#F;}�C;�%?;�#6;�(&;��;H��:Q:�$T�vK/�>Ϩ�@|��I�ZO��""����鼯��dg*�T�C��yZ�{l�W`w�      �b��䪫��ƣ��s���ɇ�{l�BG��"�i� �/aļc���I��C��ۙ�H�huƹ2�k:���:�;<>.;
;;��A;�AE;[�F;mG;��G;��G;U2H;�ZH;�zH;ՒH;��H;��H;X�H;'�H;��H;�H;��H;'�H;W�H;��H;��H;ҒH;�zH;�ZH;R2H;��G;��G;mG;Y�F;�AE;��A;
;;<>.;�;���::�k:xuƹJ��ۙ��C��I�c��/aļi� ��"�CG�zl��ɇ��s���ƣ�䪫�      ������pݽ�2̽�ж����������yZ�G-�ַ�/aļZO���J;���軂�|���º N@9���:7�;�f$;��5;�N?;6D;�LF;�:G;��G;��G;�!H;�MH;�pH;��H;˟H;,�H;�H;<�H;p�H;��H;p�H;<�H;�H;)�H;ɟH;��H;�pH;�MH;�!H;��G;��G;�:G;�LF;8D;�N?;��5;�f$;4�;���: N@9��º��|�����J;�ZO��/aļַ�G-��yZ����������ж��2̽pݽ���      P,�����Z�:��z�RvϽ�b��.I��g]a�G-�i� �""��y�{�G�!�������4��P(��nQ:�L�:��;Ҋ/;�'<;ٟB;��E;��F;��G;��G;1H;;AH;gH;L�H;0�H;̪H;��H;{�H;��H;P�H;��H;|�H;��H;ȪH;/�H;J�H;gH;;AH;/H;��G;��G;��F;��E;ٟB;�'<;ˊ/;��;�L�:�nQ:�P(���4�����G�!�y�{�""��i� �G-�g]a�.I���b��RvϽ�z�:��Z����      &G�p�C��$:��J+������pݽ^���.I���yZ��"����ԫ��fT��� � M����˺�m9-ٶ:a�;`(;
�8;b�@;��D;۱F;;hG;z�G;H;+5H;�]H;b}H;�H;��H;R�H;ĻH;��H;2�H;��H;ƻH;P�H;��H;�H;a}H;�]H;+5H;H;z�G;=hG;رF;��D;`�@;�8;�_(;d�;'ٶ:m9��˺ M���� �fT�ԫ������"��yZ�.I��]���pݽ�� ���J+��$:�p�C�      {x�9t���g���T��G=�z#�6�oݽ�b������BG������Ǽiy��M�$�j���$�$�8vƹ?��:�&�:�� ;F4;o�>;ID;�[F;�FG;y�G;��G;�)H;[UH;�vH;��H;�H;��H;f�H;�H;'�H;~�H;h�H;~�H;�H;��H;�vH;aUH;�)H; �G;z�G;�FG;�[F;KD;p�>;C4;�� ;�&�:;��:(vƹ$�$�j���L�$�iy����Ǽ���BG������b��oݽ6�z#��G=���T���g�9t�      쫖���La��!���>�c�p�C�z#���SvϽ����{l�eg*����
���I�����\c�!퀺�t,:���:�;�_0;a�<;�1C;��E;n#G;N�G;�G; H;�MH;6qH;��H;x�H;٭H;(�H;��H;[�H;��H;(�H;حH;v�H;��H;2qH;�MH; H;�G;N�G;w#G;��E;�1C;]�<;�_0;�;���:�t,:!퀺�\c�����I��
�����eg*�{l�����SvϽ��z#�p�C�>�c�!���La����      j*��g����Ƥ�쫖��/��>�c��G=�����zｑж��ɇ�R�C���$"��t;k��&��-����˺�X�9j��:
9;�h,;�	;;�PB;`�E;� G;׌G;��G;dH;GH;JlH;��H;��H;��H;4�H;�H;ѼH;��H;6�H;��H;��H;��H;HlH;GH;eH;��G;یG;� G;^�E;�PB;�	;;�h,;9;n��:�X�9�˺�-���&�s;k�$"����R�C��ɇ��ж��z�����G=�>�c��/��쫖��Ƥ�g���      ��ɾ|�ž+��qת�쫖�!�����T��J+�;��2̽�s���yZ����Oμhy����aϨ�Z,� �6��:��
;U�(;NN9;��A;xNE;(�F;�G;��G;wH;�AH;.hH;�H;:�H;ЩH;ɳH;��H;u�H;��H;ɳH;ΩH;:�H;�H;,hH;�AH;wH;��G;�G;2�F;wNE;��A;IN9;T�(;��
;��: 
�6U,�`Ϩ���gy��Oμ����yZ��s���2̽;��J+���T�!���쫖�qת�+��|�ž      U_ݾ�:پ�V;+���Ƥ�La����g��$:��Z�pݽ�ƣ�{l�f.%��߼i���9.�ϴ��VV� 2p��@�:x;D(&;+�7;3�@;�
E;��F;duG;�G;KH;�=H;JeH;��H;o�H;H�H;��H;��H;��H;��H;��H;H�H;n�H;��H;DeH;�=H;KH;!�G;guG;��F;�
E;2�@;&�7;D(&;
x;�@�:2p�VV�ϴ���9.�h���߼f.%�{l��ƣ�pݽ�Z��$:���g�La���Ƥ�+���V;�:پ      ^�3���:پ{�žh�����9t�p�C� �����䪫�X`w�F-����+`����7�:Sɻ�K/�yƹ���:�/;�f$;�7;�~@;D�D;S�F;�nG;��G;H;;H;ecH;j�H;|�H;m�H;�H;)�H; �H;&�H;�H;m�H;|�H;j�H;`cH;�;H;H;��G;�nG;a�F;C�D;�~@;�7;�f$;�/;���: yƹ�K/�;Sɻ��7�+`�����F-�X`w�䪫���� ��p�C�9t���h���{�ž�:پ4��      GF�Wh����UVھ8�������~���S��#��o��8S��p₽2�6�p���jy��YFB��Eֻ�A?���	�^Y�:���:a�";b46;X@;Y�D;��F;�nG;��G;�H;@H;�fH;<�H;)�H;��H;̳H;˹H;��H;ƹH;̳H;��H;+�H;>�H;�fH;@H;�H;��G;�nG;��F;Y�D;T@;Y46;a�";���:bY�:��	��A?��EֻXFB�iy��p���2�6�p₽8S���o���#��S��~������7��UVھ��Wh��      Vh���b���쾧*־�v��)���*��(�O�V� �s��r���؀�F�3���@ݜ�?�>�V�ѻ�9� ���o�:6% ;lM#;<�6;HA@;��D;��F;qG;H�G;H;�@H;dgH;��H;��H;٩H;�H;��H;ٻH;�H;�H;٩H;��H;��H;`gH;�@H;H;H�G;qG;��F;��D;DA@;7�6;jM#;6% ;o�:����9�V�ѻ?�>�@ݜ���F�3��؀��r��s�V� �'�O�*��)����v���*־���b��      ���쾳�޾05ʾM;���:��(�v��E�`'����r����u���+��W��A����4���Ļ&9)��j��kW�:Z�;%;�k7;�@;��D;��F;�wG;Q�G;.H;9CH;&iH;	�H;��H;��H;��H;��H;n�H;��H;��H;��H;��H;	�H; iH;ACH;1H;Q�G;�wG;��F;��D;�@;�k7;�%;Z�;sW�:�j��&9)���Ļ��4��A���W缄�+���u�q�����`'��E�(�v��:��L;��05ʾ��޾��      UVھ�*־/5ʾr��������M���9b��5�����ս����Xc���̖ռ�I��X�$�qT���Z��]����:��;f�';�8;RA;�9E;��F;��G;��G;=H;GH;lH;?�H;6�H;ݫH;��H;��H;L�H;��H;��H;ޫH;5�H;>�H;lH;GH;@H;��G;��G;��F;�9E;RA;�8;c�';��;�:�]���Z�pT��X�$��I��̖ռ���Xc������ս���5��9b��M������r���/5ʾ�*־      7���v��L;������SP��E�r�z�H�U� ���6@��ѓ����K�b��վ���s�t���񕻰ܺP4u9�%�:�;'�+;x�:;�"B;g�E;��F;ΐG;��G;*H;1LH;�oH;7�H;q�H;��H;0�H;ԼH;�H;мH;4�H;��H;n�H;6�H;�oH;:LH;+H;��G;АG;��F;h�E;�"B;t�:;&�+;�;&�:P4u9�ܺ��u����s��վ�b���K�ѓ��6@����U� �z�H�E�r�SP������M;���v��      ����)����:���M��E�r�'�O�#,�X�
��gٽqĥ���u�x1�j���+Ϥ���P�[��.o��p��:Q��:�P;7�/;4�<;�
C;�E;g!G;0�G;��G;�%H;�RH;�tH;�H;C�H;ӯH;��H;V�H; �H;R�H;��H;үH;@�H;�H;�tH;�RH;�%H;��G;0�G;n!G;�E;�
C;0�<;6�/;�P;[��: :�p���.o�[򻬎P�*Ϥ�j���w1���u�qĥ��gٽX�
�#,�'�O�E�r��M���:��)���      �~��*��(�v��9b�z�H�#,�MZ����7S��x^����N������μ�I���%+�����.������j~:9��:&m;��3;�>;7�C;6PF;yFG;L�G;��G;r/H;�YH;qzH;A�H;��H;Y�H;�H;&�H;��H;#�H;�H;[�H;��H;@�H;pzH;ZH;u/H;��G;J�G;�FG;8PF;6�C;�>;��3;%m;C��:�j~:�����.�����%+��I����μ�����N�x^��6S�����MZ�#,�z�H��9b�(�v�*��      �S�'�O��E��5�V� �X�
���罥9��(l���Xc���(��������[�����ݎ�Wܺ�:9��:&�	;@d';^ 8;6�@;z�D;�F;jG;��G;HH;k:H;<bH;��H;�H;.�H;=�H;x�H;3�H;��H;2�H;{�H;?�H;-�H;��H;��H;FbH;p:H;KH;��G;jG;�F;t�D;8�@;_ 8;=d';-�	;��:�:9Rܺ�ݎ������[��������(��Xc�(l���9�����X�
�V� ��5��E�'�O�      �#�U� �`'������gٽ6S��(l��P�j�C�3��i��վ�{���	(���ĻhA?���B���@:�[�:Q; �.;��;;xtB;�E;y�F;�G;��G;�H;NFH;kH;��H;�H;�H;b�H;�H;o�H;��H;l�H;�H;e�H;�H;�H;��H;(kH;TFH;�H;��G;"�G;}�F;�E;ztB;��;;��.;
Q;�[�:��@:��B�gA?���Ļ	(�{����վ��i�C�3�O�j�(l��6S���gٽ����`'�V� �      �o��s��罬�ս5@��qĥ�y^���Xc�D�3���	�ˌ˼�]��UFB��Z򻲜��}Ӻ���8��:ԛ;�M#;p=5;?;F�C;w@F; :G;�G;�G;*'H;�RH;stH;��H;x�H;(�H;��H;��H;��H;<�H;��H;��H;��H;&�H;u�H;��H;}tH;�RH;/'H;�G;�G;:G;u@F;K�C;?;n=5;�M#;՛;��:���8|Ӻ�����Z�TFB��]��ˌ˼��	�C�3��Xc�x^��qĥ�6@����ս���s�      8S���r��r�����ѓ����u���N���(��i�ˌ˼�A����P�is��D|�����|\:"�:h�;pn-;ܞ:;�A;v,E;d�F;&oG;��G;�H;�7H;4_H;~H;�H;��H;p�H;	�H;t�H;6�H;|�H;8�H;v�H;�H;p�H;��H;�H;~H;=_H;�7H;�H;��G;,oG;f�F;z,E;�A;ޞ:;|n-;l�;"�:�\:����B|��is���P��A��ˌ˼�i���(���N���u�ғ�����r���r��      p₽�؀���u��Xc���K�w1�������վ��]����P����FT����9�(�o�p3�9d&�:W�	;T%;@�5;��>;��C;�F;�!G;��G;��G;@H;ZHH;�kH;��H;F�H;��H;��H;q�H;F�H;��H;��H;��H;F�H;u�H;��H;��H;J�H;��H;�kH;`HH;BH;��G;��G;�!G;�F;��C;��>;K�5;W%;V�	;r&�:�3�9 �o���9�DT�������P��]���վ�����w1���K��Xc���u��؀�      3�6�F�3���+���a�j�����μ���{���TFB�is�FT��6�D��{�� :u9�q�:k��:xY;�t0;��;;�B;�9E;߻F;�gG;ӿG;��G;u0H;�XH;"xH;�H;r�H;��H;��H;��H;�H;+�H;/�H;+�H;�H;��H;��H;��H;w�H;&�H;,xH;�XH;y0H;��G;ۿG;�gG;�F;�9E;�B;��;;�t0;sY;y��:�q�:0:u9�{��4�D�CT��hs�TFB�z��������μj���b�����+�F�3�      n�����W�͖ռ�վ�,Ϥ��I����[�
(��Z����9��{�� ;9?X�:HX�:3Q;8,;��8;�A@;
BD;�@F;�,G;��G;��G;aH;�DH;hH;)�H;N�H;a�H;Z�H; �H;�H;��H;��H;a�H;��H;��H;�H;�H;X�H;g�H;Y�H;3�H;hH;�DH;`H;��G;��G;�,G;�@F;BD;�A@;��8;6,;;Q;HX�:EX�:@;9�{����9���Z�(���[��I��+Ϥ��վ�͖ռ�W���      hy��@ݜ��A���I����s���P��%+������Ļ����@|�<�o��9u9CX�:�+�:P;�);̈́6;n�>;zPC;^�E;��F;�xG;%�G;tH;_1H;XH;�vH;��H;�H;��H;z�H;�H;<�H;}�H;��H;��H;��H;}�H;?�H;�H;w�H;��H;�H;��H;wH;XH;^1H;{H;)�G;�xG;��F;b�E;�PC;t�>;Ǆ6;�);P;�+�:GX�::u9,�o�=|�������Ļ����%+���P���s��I���A��@ݜ�      SFB�=�>���4�V�$�u��[�����ݎ�nA?�yӺ����X3�9�q�:HX�:P;��';~=5;x�=;��B;GE;E�F;}UG;�G;��G;NH;�HH;jH;�H;q�H;D�H;,�H;D�H;��H;;�H;�H;�H;��H;�H;
�H;;�H;��H;A�H;3�H;I�H;x�H;��H;jH;�HH;VH;��G;�G;�UG;I�F;GE; �B;t�=;�=5;��';T;HX�:�q�:p3�9x���vӺgA?��ݎ����[�w��X�$���4�:�>�      �EֻT�ѻ��ĻsT�����.o���.�Qܺ��B����8�\:h&�:q��:9Q;�);�=5;�:=;$#B;~�D;�uF;�6G;��G;V�G;oH;�:H;^H;�zH;��H;[�H;��H;�H;��H;Z�H;�H;j�H;/�H;��H;*�H;h�H;�H;U�H;��H;�H;ĲH;b�H;��H;�zH;^H;�:H;rH;X�G;��G;�6G;�uF;��D;#B;�:=;�=5;�);:Q;s��:l&�:�\:���8��B�Kܺ�.��.o���vT����ĻO�ѻ      }A?��9�,9)��Z��ܺ�p������ ;9��@:��:(�:P�	;qY;4,;Ƅ6;o�=;#B;��D;\XF;�!G;v�G;�G;�H;�.H;uSH;_qH;ۉH;��H;_�H;��H;m�H;��H;��H;��H;�H;�H;��H;�H;|�H;��H;��H;��H;q�H;��H;c�H;��H;܉H;[qH;{SH;�.H;�H;�G;z�G;�!G;^XF;��D;#B;m�=;Ʉ6;4,;qY;S�	;2�:��:��@:P;9����zp���ܺ�Z�$9)��9�      ��	������j���\��@4u9H:�j~:��:�[�:כ;r�;T%;�t0;��8;s�>;�B;~�D;dXF;1G;[�G;��G;��G;�%H;�JH;�iH;��H;��H;5�H;s�H;�H;X�H;��H;��H;0�H;}�H;��H;P�H;��H;{�H;/�H;��H;��H;[�H;�H;s�H;5�H;��H;߂H;�iH;KH;�%H;��G;��G;_�G;4G;\XF;��D;��B;u�>;��8;�t0;T%;r�;՛;�[�:��:�j~:0:`4u9`^���j��p���      NY�:o�:uW�:�:�%�:Y��:U��:&�	;Q;�M#;yn-;G�5;��;;�A@;�PC;GE;�uF;�!G;^�G;��G;�G;B H;EH;�cH;5}H;q�H;��H;��H;��H;��H;��H;)�H;Q�H;P�H;K�H;w�H;��H;r�H;H�H;N�H;O�H;'�H;��H;��H;��H;��H;��H;p�H;;}H;�cH;EH;E H;�G;��G;b�G;�!G;�uF;GE;�PC;�A@;��;;H�5;|n-;�M#;Q;-�	;O��:c��:�%�:��:aW�:�n�:      ���:$% ;>�;��;�;�P;$m;7d';��.;n=5;ޞ:;��>;�B;BD;a�E;I�F;�6G;��G;��G;�G;qH;�AH;`H;IyH;x�H;�H;N�H;޹H;H�H;��H;��H;.�H;��H;@�H;��H;��H;A�H;��H;��H;>�H;��H;(�H;��H;��H;H�H;߹H;K�H;�H;|�H;FyH;`H;�AH;tH;�G;��G;z�G;�6G;E�F;_�E;BD;�B;��>;�:;m=5;��.;6d';(m;�P;�;��;H�;"% ;      U�";nM#;%;n�';#�+;4�/;��3;X 8;��;;?;��A;��C;�9E;�@F;��F;�UG;��G;�G;��G;E H;�AH;�^H;BwH;�H;~�H;ݫH;��H;+�H;��H;"�H;�H;��H;��H;��H;k�H;I�H;y�H;D�H;j�H;��H;��H;��H;�H;#�H;��H;*�H;��H;۫H;��H;�H;=wH;�^H;�AH;F H;��G;�G;��G;~UG;��F;�@F;�9E;��C;��A;?;��;;a 8;��3;/�/;7�+;c�';�%;bM#;      t46;:�6;�k7;"�8;p�:;7�<;$�>;@�@;tB;M�C;�,E;�F;�F;�,G;�xG;!�G;Z�G;�H;�%H;EH;`H;AwH;/�H;3�H;D�H;�H;��H;k�H;��H;��H;%�H;?�H;��H;]�H;��H;o�H;��H;i�H;��H;_�H;��H;<�H;(�H;��H;��H;k�H;��H;�H;H�H;.�H;(�H;BwH;`H;	EH;�%H;�H;\�G;�G;�xG;�,G;�F;�F;~,E;F�C;~tB;@�@; �>;6�<;~�:;!�8;�k7;�6;      W@;NA@;�@;RA;�"B;�
C;7�C;w�D;�E;y@F;h�F;�!G;�gG;��G;)�G;��G;tH;�.H;KH;�cH;GyH;�H;0�H;��H;�H;{�H;u�H;��H;�H;K�H;��H;J�H;:�H;��H;��H;^�H;��H;X�H;��H;��H;7�H;H�H;��H;J�H;�H;��H;p�H;|�H;�H;��H;*�H;�H;DyH;�cH; KH;�.H;qH;��G;(�G;��G;�gG;�!G;h�F;w@F;�E;~�D;7�C;�
C;�"B;RA;�@;GA@;      {�D;��D;��D;�9E;`�E;!�E;APF;�F;|�F;:G;0oG;��G;ڿG;��G;{H;ZH;�:H;�SH;�iH;?}H;��H;��H;H�H;�H;:�H;��H;*�H;j�H;��H;*�H;��H;	�H;��H;��H;��H;%�H;c�H;�H;��H;��H;��H;�H;��H;(�H;��H;j�H;#�H;��H;=�H;�H;F�H;��H;�H;;}H;�iH;|SH;�:H;VH;zH;��G;ٿG;��G;0oG;:G;�F;ߩF;?PF;�E;j�E;}9E;��D;��D;      ~�F;��F;��F;|�F;��F;n!G;�FG;jG;#�G;�G;��G;��G;�G;lH;b1H;�HH;^H;cqH;��H;n�H;�H;׫H;�H;{�H;��H;�H;�H;X�H;��H;��H;��H;��H;��H;��H;x�H;��H;�H;��H;u�H;��H;��H;}�H;��H;��H;��H;W�H;�H;
�H;��H;x�H;�H;׫H;�H;k�H;܂H;[qH;^H;�HH;_1H;dH;��G;��G;��G;�G;#�G;jG;�FG;a!G;��F;��F;��F;��F;      �nG;qG;�wG;��G;ƐG;+�G;X�G;��G;��G;�G;�H;>H;u0H;�DH;XH;jH;�zH;�H;��H;��H;T�H;��H;��H;x�H;)�H;�H;;�H;��H;Z�H;x�H;I�H;��H;��H;��H;4�H;��H;��H;��H;2�H;��H;��H;��H;I�H;x�H;W�H;��H;5�H;�H;,�H;r�H;��H;��H;Q�H;��H;��H;؉H;�zH;jH;XH;�DH;r0H;@H;�H;�G;��G;��G;Q�G;&�G;ڐG;��G;�wG;�pG;      ��G;B�G;J�G;��G;��G;��G;��G;GH;�H;2'H;�7H;dHH;�XH; hH;�vH;��H;��H;��H;7�H;��H;�H;'�H;h�H;��H;i�H;W�H;��H;9�H;t�H;>�H;��H;��H;��H;a�H;��H; �H;�H;��H;��H;c�H;��H;��H;��H;>�H;s�H;6�H;��H;X�H;l�H;��H;j�H;(�H;߹H;��H;5�H;��H;��H;�H;�vH;hH;�XH;aHH;�7H;0'H;�H;HH;��G;��G;��G;��G;I�G;:�G;      �H;H;+H;JH;H;�%H;v/H;d:H;HFH;�RH;=_H;�kH;*xH;.�H;��H;w�H;b�H;i�H;x�H;��H;K�H;��H;��H;�H;��H;��H;V�H;t�H;!�H;��H;��H;��H;U�H;��H;C�H;u�H;��H;p�H;C�H;��H;V�H;��H;��H;��H;�H;s�H;P�H;��H;��H;�H;��H;��H;H�H;��H;v�H;e�H;d�H;w�H;��H;,�H;%xH;�kH;=_H;�RH;JFH;g:H;v/H;�%H;&H;FH;*H;H;      @H;�@H;DCH;GH;:LH;�RH;�YH;:bH;#kH;|tH;~H;��H;#�H;Y�H;�H;G�H;ǲH;��H;�H;��H;��H;�H;��H;G�H;'�H;��H;w�H;>�H;��H;��H;��H;g�H;��H;M�H;��H;��H;��H;��H;��H;M�H;��H;d�H;��H;��H;��H;;�H;q�H;��H;*�H;D�H;��H;!�H;��H;��H;�H;��H;ŲH;H�H;�H;V�H;#�H;��H;~H;}tH;"kH;@bH;ZH;�RH;8LH;GH;ECH;�@H;      �fH;tgH;+iH;lH;�oH;�tH;{zH;��H;��H;��H;�H;P�H;z�H;m�H;�H;5�H;�H;u�H;`�H;��H;��H;�H;%�H;��H;��H;��H;H�H;��H;��H;��H;g�H;�H;^�H;��H;��H;�H;'�H;�H;��H;��H;`�H;�H;g�H;��H;��H;��H;E�H;��H;��H;��H;)�H;�H;��H;��H;^�H;r�H;�H;5�H;�H;k�H;}�H;Q�H;�H;��H;��H;��H;�zH;�tH;�oH;lH;-iH;vgH;      A�H;��H;�H;;�H;7�H;�H;K�H;�H;!�H;{�H;�H;��H;�H;d�H;{�H;J�H;��H;��H;��H;,�H;5�H;��H;<�H;E�H;�H;|�H;��H;��H;��H;h�H;��H;u�H;��H;��H;&�H;@�H;@�H;@�H;#�H;��H;��H;o�H;��H;g�H;��H;��H;��H;}�H;	�H;?�H;?�H;��H;/�H;)�H;��H;��H;��H;K�H;~�H;b�H;�H;��H;�H;z�H; �H;�H;P�H;�H;B�H;;�H;�H;��H;      .�H;��H;��H;8�H;{�H;@�H;��H;+�H;	�H;-�H;w�H;��H;��H;'�H;�H;��H;^�H;��H;��H;V�H;��H;��H;��H;3�H;��H;��H;��H;��H;Z�H;��H;[�H;��H;�H;5�H;T�H;w�H;}�H;w�H;Q�H;6�H;�H;��H;Z�H;��H;U�H;��H;��H;��H;��H;3�H;��H;��H;��H;R�H;��H;��H;_�H;��H;�H;'�H;��H;��H;x�H;.�H;�H;-�H;��H;:�H;}�H;2�H;��H;��H;      ��H;שH;��H;׫H;��H;ɯH;d�H;C�H;k�H;��H;�H;~�H;��H;$�H;E�H;D�H;�H;��H;4�H;T�H;D�H;��H;X�H;��H;��H;��H;��H;c�H;��H;P�H;��H;��H;2�H;p�H;�H;��H;��H;��H;~�H;q�H;5�H;��H;��H;M�H;��H;]�H;��H;��H;��H;��H;]�H;��H;=�H;N�H;3�H;��H;$�H;E�H;E�H;$�H;��H;{�H;�H;��H;o�H;I�H;i�H;ɯH;��H;֫H;��H;�H;      ɳH;"�H;��H;ĵH;B�H;��H;(�H;{�H;�H;��H;��H;S�H;�H;��H;��H;�H;o�H;�H;}�H;L�H;��H;i�H;��H;��H;��H;m�H;,�H;��H;E�H;��H;��H;'�H;T�H;��H;��H;��H;��H;��H;��H;��H;U�H;'�H;��H;��H;?�H;��H;,�H;p�H;��H;��H;��H;f�H;��H;G�H;{�H;��H;s�H;�H;��H;��H;�H;T�H;��H;��H;�H;�H;)�H;��H;B�H;ƵH;ôH;#�H;      ʹH;�H;��H;��H;ԼH;N�H;5�H;7�H;r�H;��H;C�H;��H;2�H;��H;��H;�H;/�H;�H;��H;w�H;��H;E�H;e�H;N�H;�H;��H;��H;�H;y�H;��H;�H;D�H;}�H;��H;��H;��H;��H;��H;��H;��H;�H;D�H;�H;��H;u�H;��H;��H;��H;�H;N�H;k�H;D�H;��H;r�H;��H;�H;3�H; �H;��H;��H;0�H;��H;D�H;��H;v�H;<�H;:�H;O�H;׼H;��H;��H;�H;      ŻH;ٻH;��H;M�H;|�H;�H;��H;��H;��H;E�H;��H;��H;>�H;o�H;��H;��H;��H;��H;U�H;��H;M�H;�H;��H;��H;b�H; �H;��H;�H;��H;��H;$�H;D�H;~�H;��H;��H;��H;��H;��H;��H;��H;��H;D�H;$�H;��H;��H;�H;��H;�H;b�H;��H;��H;|�H;F�H;��H;U�H;��H;��H;��H;��H;p�H;=�H;��H;��H;F�H;��H;��H;��H;�H;~�H;L�H;��H;�H;      ʹH;��H;��H;��H;ּH;R�H;3�H;6�H;r�H;��H;B�H;��H;3�H;��H;��H;�H;/�H;�H;��H;w�H;��H;G�H;e�H;N�H;�H;��H;��H; �H;y�H;��H;�H;D�H;}�H;��H;��H;��H;��H;��H;��H;��H;�H;D�H;�H;��H;u�H;��H;��H;��H;�H;M�H;k�H;B�H;��H;r�H;��H;�H;0�H; �H;��H;��H;0�H;��H;D�H;��H;v�H;<�H;7�H;O�H;ڼH;��H;��H;��H;      ��H;&�H;��H;��H;D�H;��H;)�H;~�H;�H;��H;��H;S�H;�H;��H;��H;�H;o�H;��H;}�H;L�H;��H;j�H;��H;��H;��H;k�H;-�H;��H;C�H;��H;��H;(�H;T�H;��H;��H;��H;��H;��H;��H;��H;W�H;'�H;��H;��H;?�H;��H;,�H;r�H;��H;��H;��H;g�H;��H;G�H;{�H;�H;q�H;�H;��H;��H;�H;V�H;��H;��H;�H;��H;/�H;��H;E�H;��H;��H;%�H;      ��H;թH;��H;ګH;��H;ͯH;b�H;G�H;l�H;��H;�H;|�H;��H;$�H;H�H;D�H;!�H;��H;4�H;T�H;E�H;��H;X�H;��H;��H;��H;��H;c�H;��H;O�H;��H;��H;4�H;p�H;�H;��H;��H;��H;~�H;o�H;4�H;��H;��H;L�H;��H;^�H;��H;��H;��H;��H;]�H;��H;;�H;P�H;3�H;��H;!�H;D�H;F�H;#�H;��H;{�H;�H;��H;o�H;J�H;i�H;˯H;��H;֫H;��H;ةH;      /�H;��H;��H;5�H;u�H;A�H;��H;.�H;	�H;.�H;w�H;��H;��H;(�H;�H;��H;^�H;��H;��H;V�H;��H;��H;��H;3�H;��H;��H;��H;��H;Z�H;��H;[�H;��H;�H;5�H;T�H;x�H;}�H;v�H;S�H;4�H;�H;��H;Z�H;��H;S�H;��H;��H;��H;��H;2�H;��H;��H;��H;T�H;��H;��H;\�H;��H;�H;'�H;��H;��H;w�H;+�H;�H;1�H;��H;=�H;y�H;;�H;��H;��H;      0�H;��H;��H;7�H;3�H;��H;N�H;�H;�H;z�H;�H;��H;�H;d�H;�H;K�H;��H;��H;��H;,�H;6�H;��H;:�H;C�H;	�H;|�H;��H;��H;��H;e�H;��H;r�H;��H;��H;'�H;?�H;@�H;@�H;$�H;��H;��H;p�H;��H;e�H;��H;��H;��H;��H;�H;>�H;A�H;��H;-�H;)�H;��H;��H;��H;J�H;}�H;b�H;�H;��H;�H;{�H;#�H;�H;P�H;�H;7�H;8�H;�H;��H;      �fH;ugH;-iH;lH;�oH;�tH;zzH;��H;��H;��H;�H;S�H;|�H;m�H;�H;5�H;�H;u�H;`�H;��H;��H;�H;%�H;��H;��H;��H;E�H;��H;��H;��H;g�H;�H;^�H;��H;��H;�H;'�H;�H;��H;��H;`�H;�H;e�H;��H;��H;��H;E�H;��H;��H;��H;*�H;�H;��H;��H;^�H;q�H;�H;4�H;�H;k�H;z�H;S�H;�H;��H;��H;��H;zH;�tH;pH;lH;4iH;vgH;      @H;�@H;@CH;GH;0LH;�RH;�YH;CbH;&kH;~tH;~H;��H;$�H;X�H;�H;G�H;ǲH;��H;�H;��H;��H;"�H;��H;F�H;(�H;��H;t�H;>�H;��H;��H;��H;g�H;��H;M�H;��H;��H;��H;��H;��H;M�H;��H;e�H;��H;��H;��H;;�H;s�H;��H;(�H;A�H;��H;!�H;��H;��H;�H;��H;ŲH;E�H;�H;X�H;$�H;��H;~H;~tH;%kH;DbH;ZH;�RH;;LH;GH;PCH;�@H;      �H;H;=H;DH;H;�%H;u/H;i:H;QFH;�RH;;_H;�kH;)xH;.�H;��H;w�H;`�H;j�H;t�H;��H;K�H;��H;��H;�H;��H;��H;R�H;t�H;!�H;��H;��H;��H;V�H;��H;C�H;s�H;��H;s�H;C�H;��H;W�H;��H;��H;��H;�H;q�H;R�H;��H;��H;�H;��H;��H;H�H;��H;v�H;b�H;`�H;x�H;��H;.�H;)xH;�kH;@_H;�RH;QFH;m:H;{/H;�%H;#H;CH;?H;�H;      ��G;8�G;<�G;��G;��G;�G;��G;KH;�H;3'H;�7H;aHH;�XH;hH;�vH;�H;��H;��H;3�H;��H;�H;(�H;d�H;��H;l�H;Q�H;��H;6�H;w�H;;�H;��H;��H;��H;a�H;��H;��H;�H;��H;��H;c�H;��H;��H;��H;>�H;t�H;4�H;��H;U�H;i�H;��H;m�H;(�H;۹H;��H;5�H;��H;��H;�H; wH;hH;�XH;aHH;�7H;2'H;�H;IH;��G;��G;��G;��G;J�G;8�G;      �nG;qG;�wG;ʂG;ӐG;4�G;W�G;��G;��G;�G;�H;@H;r0H;�DH;XH;jH;�zH;��H;��H;��H;T�H;��H;��H;x�H;*�H;�H;6�H;��H;\�H;w�H;H�H;��H;��H;��H;4�H;��H;��H;��H;2�H;��H;��H;��H;K�H;z�H;Y�H;��H;6�H;�H;*�H;t�H;��H;��H;Q�H;��H;��H;ۉH;�zH;jH;XH;�DH;s0H;AH;�H;�G;��G;��G;[�G;0�G;ڐG;ǂG;�wG;qG;      {�F;��F;��F;|�F;��F;v!G;|FG;"jG;(�G;�G;��G;��G;�G;gH;a1H;�HH;^H;aqH;݂H;k�H;�H;׫H;޵H;x�H;��H;�H;�H;W�H;��H;��H;��H;��H;��H;��H;x�H;��H;
�H;��H;u�H;��H;��H;��H;��H;��H;��H;U�H;�H;�H;��H;x�H;�H;׫H;�H;m�H;߂H;\qH;^H;�HH;f1H;gH;�G;��G;��G;�G;!�G;jG;}FG;g!G;��F;}�F;��F;y�F;      z�D;��D;��D;�9E;`�E;$�E;APF;ߩF;}�F;:G;/oG;��G;׿G;��G;{H;YH;�:H;�SH;�iH;;}H;��H;��H;D�H;�H;<�H;��H;&�H;j�H;��H;$�H;��H;	�H;��H;��H;��H;"�H;c�H;"�H;��H;��H;��H;�H;��H;(�H;��H;f�H;'�H;��H;:�H;�H;K�H;��H;�H;?}H;�iH;}SH;�:H;YH;~H;��G;ڿG;��G;/oG;:G;}�F;�F;BPF;�E;j�E;�9E;��D;��D;      8@;6A@;�@;RA;�"B;C;8�C;x�D;�E;u@F;h�F;�!G;�gG;��G;)�G;��G;qH;�.H; KH;�cH;GyH;�H;,�H;��H;�H;t�H;r�H;��H;�H;G�H;��H;L�H;9�H;��H;��H;\�H;��H;^�H;��H;��H;<�H;J�H;��H;K�H;�H;��H;t�H;{�H;�H;éH;.�H;�H;FyH;�cH;KH;�.H;rH;��G;+�G;��G;�gG;�!G;k�F;w@F;�E;t�D;8�C;�
C;�"B;,RA;�@;A@;      h46;5�6;�k7;,�8;n�:;3�<;�>;>�@;�tB;I�C;z,E;�F;�F;�,G;�xG;"�G;Z�G;�H;�%H;EH;`H;BwH;)�H;3�H;G�H;ߵH;��H;k�H;��H;��H;(�H;@�H;��H;]�H;��H;p�H;��H;n�H;��H;[�H;��H;@�H;-�H;��H;��H;j�H;��H;�H;F�H;1�H;,�H;AwH;`H;EH;�%H;�H;\�G;!�G;�xG;�,G;�F;�F;},E;L�C;�tB;B�@;�>;3�<;l�:;&�8;�k7; �6;      Z�";pM#;%;d�';#�+;;�/;��3;] 8;��;;?;��A;��C;�9E;�@F;��F;�UG;��G; �G;��G;F H;�AH;�^H;>wH;�H;��H;֫H;��H;*�H;��H;!�H;�H;��H;��H;��H;i�H;E�H;{�H;H�H;j�H;��H;��H;��H; �H;#�H;��H;'�H;��H;ګH;~�H;�H;BwH;�^H;�AH;F H;��G;�G;��G;UG;��F;�@F;�9E;��C;��A;?;��;;a 8;��3;&�/;:�+;Y�';%;`M#;      ���:<% ;N�;��;�;�P;&m;9d'; �.;k=5;��:;��>;�B;BD;b�E;I�F;�6G;��G;��G;�G;qH;�AH;`H;IyH;{�H;�H;J�H;ܹH;H�H;��H;��H;/�H;��H;B�H;��H;��H;C�H;��H;��H;@�H;��H;-�H;��H;��H;E�H;۹H;M�H;�H;z�H;JyH;`H;�AH;pH;�G;��G;|�G;�6G;H�F;d�E;BD;�B;��>;�:;m=5;��.;=d';+m;�P;�;��;\�;(% ;      �Y�:o�:oW�:�:�%�:c��:W��:0�	;	Q;�M#;~n-;G�5;��;;�A@;�PC;GE;�uF;�!G;^�G;��G;�G;F H;EH;�cH;9}H;m�H;��H;��H;��H;��H;��H;(�H;R�H;S�H;K�H;s�H;��H;u�H;H�H;M�H;Q�H;(�H;��H;��H;��H;��H;��H;p�H;5}H;�cH;	EH;C H;�G;��G;^�G;�!G;�uF;GE;�PC;�A@;��;;G�5;|n-;�M#;Q;)�	;Q��:Q��: &�:��:oW�:o�:      ��	�p����j���\�� 4u9H:�j~:��:�[�:כ;p�;U%;�t0;��8;w�>;�B;�D;`XF;1G;_�G;��G;��G;�%H;KH;�iH;݂H;��H;3�H;t�H;�H;[�H;��H;��H;0�H;~�H;��H;P�H;��H;{�H;/�H;��H;��H;[�H;�H;q�H;1�H;��H;��H;�iH;KH;�%H;��G;��G;^�G;1G;]XF;�D;��B;u�>;��8;�t0;T%;r�;՛;�[�: ��:�j~:@: 4u9 ]���j��H���      �A?�ܡ9�.9)��Z��ܺlp�������;9��@:��:,�:U�	;qY;4,;ʄ6;r�=;#B;��D;ZXF;�!G;|�G;�G;�H;�.H;ySH;\qH;׉H;��H;e�H;��H;o�H;��H;��H;��H;}�H;�H;��H;�H;{�H;��H;��H;��H;o�H;��H;b�H;��H;ۉH;[qH;uSH;�.H;�H;�G;v�G;�!G;\XF;��D;#B;n�=;ʄ6;4,;oY;R�	;0�:��:��@:p;9����vp���ܺ�Z�89)�ܡ9�      �EֻT�ѻ��ĻqT�����.o��.�Mܺ��B����8�\:p&�:s��:9Q;�);�=5;�:=; #B;|�D;�uF;�6G;��G;Z�G;rH;�:H;^H;�zH;��H;b�H;��H;�H;��H;Z�H;�H;j�H;-�H;��H;-�H;h�H;�H;T�H;��H;�H;òH;`�H;�H;�zH;^H;�:H;qH;Z�G;��G;�6G;�uF;|�D;#B;�:=;�=5;�);9Q;s��:j&�:�\:���8��B�Mܺ�.��.o���uT����ĻP�ѻ      SFB�=�>���4�V�$�u��[�����ݎ�jA?�yӺh����3�9�q�:LX�:V;��';~=5;u�=;��B;GE;K�F;�UG;"�G;��G;VH;�HH;jH;�H;x�H;G�H;1�H;G�H;��H;@�H;�H;�H;��H;�H;	�H;:�H;��H;A�H;.�H;E�H;u�H;�H;jH;�HH;NH;��G;!�G;UG;B�F;GE;��B;r�=;~=5;��';R;HX�:�q�:X3�9p���{ӺjA?��ݎ����[�x��W�$���4�=�>�      hy��@ݜ��A���I����s���P��%+������Ļ����>|�0�o�:u9IX�:�+�:R;�);ʄ6;q�>;�PC;e�E;��F;�xG;)�G;zH;c1H;XH;�vH;��H;�H;��H;z�H;�H;A�H;~�H;��H;��H;��H;}�H;>�H;�H;w�H;��H;�H;��H;�vH;XH;\1H;tH;)�G;�xG;��F;\�E;�PC;n�>;Ƅ6;�);N;�+�:CX�:�9u94�o�@|�������Ļ����%+���P���s��I���A��@ݜ�      n�����W�̖ռ�վ�+Ϥ��I����[�(��Z����9��{��@;9KX�:RX�:7Q;4,;��8;�A@;BD;�@F;�,G;��G;��G;eH;�DH;hH;0�H;T�H;g�H;]�H; �H;�H;��H;��H;a�H;��H;��H;�H;�H;W�H;c�H;V�H;.�H;hH;�DH;^H;��G;��G;�,G;�@F;BD;�A@;��8;4,;7Q;HX�:CX�: ;9�{����9���Z�	(���[��I��+Ϥ��վ�̖ռ�W���      2�6�F�3���+���a�j�����μ���{���TFB�hs�DT��3�D��{��P:u9�q�:q��:uY;�t0;��;;�B;�9E;�F;�gG;ٿG;��G;v0H;�XH;*xH;!�H;v�H;��H;��H;��H;�H;+�H;/�H;+�H;�H;��H;�H;��H;s�H;!�H;'xH;�XH;r0H;��G;ӿG;�gG;�F;�9E;�B;��;;�t0;qY;q��:�q�:0:u9�{��5�D�ET��is�TFB�{��������μj���b�����+�F�3�      p₽�؀���u��Xc���K�w1�������վ��]����P����DT����9��o��3�9l&�:R�	;U%;D�5;��>;��C;�F;�!G;��G;��G;@H;]HH;�kH;��H;J�H;��H;��H;t�H;F�H;��H;��H;��H;F�H;r�H;��H;��H;G�H;��H;�kH;ZHH;;H;��G;��G;�!G;�F;��C;��>;F�5;R%;U�	;j&�:X3�9 �o���9�ET�������P��]���վ�����w1���K��Xc���u��؀�      8S���r��r�����ѓ����u���N���(��i�ˌ˼�A����P�is��@|������\:�:i�;un-;�:;�A;|,E;g�F;)oG;��G;�H;�7H;;_H;~H;�H;��H;p�H;�H;t�H;9�H;~�H;8�H;t�H;
�H;m�H;��H;�H;	~H;;_H;�7H;�H;��G;#oG;g�F;z,E;�A;؞:;wn-;h�;�:�\:����C|��is���P��A��ˌ˼�i���(���N���u�ғ�����r���r��      �o��s��罬�ս5@��qĥ�x^���Xc�C�3���	�ʌ˼�]��UFB��Z򻰜��{Ӻ���8��:ԛ;�M#;r=5;?;K�C;x@F;:G;�G;�G;,'H;�RH;ztH;��H;u�H;(�H;��H;��H;��H;<�H;��H;��H;��H;&�H;t�H;��H;ytH;�RH;)'H;�G;�G; :G;x@F;K�C;?;j=5;�M#;ћ;��:`��8}Ӻ�����Z�UFB��]��ˌ˼��	�C�3��Xc�y^��qĥ�6@����ս���s�      �#�U� �`'������gٽ6S��(l��P�j�C�3��i��վ�{���	(���ĻfA?���B���@:�[�:Q;�.;��;;ztB;�E;}�F;"�G;��G;�H;QFH;!kH;��H;�H;�H;e�H;�H;o�H;��H;n�H;�H;d�H;�H;�H;�H;"kH;QFH;�H;��G;"�G;{�F;�E;ztB;��;;��.;
Q;�[�:��@:��B�hA?���Ļ	(�{����վ��i�C�3�O�j�(l��7S���gٽ����`'�U� �      �S�'�O��E��5�U� �X�
���罥9��(l���Xc���(��������[�����ݎ�Uܺ�:9��:)�	;Ad';_ 8;:�@;{�D;�F;jG;��G;GH;j:H;<bH;��H;�H;.�H;@�H;x�H;3�H;��H;3�H;z�H;@�H;*�H;��H;��H;@bH;m:H;HH;��G;jG;�F;z�D;8�@;^ 8;:d';-�	;��:�:9Qܺ�ݎ������[��������(��Xc�(l���9�����X�
�U� ��5��E�'�O�      �~��*��(�v��9b�z�H�#,�MZ����7S��x^����N������μ�I���%+�����.������j~:?��:)m;��3;�>;7�C;7PF;zFG;I�G;��G;t/H;�YH;rzH;A�H;��H;[�H;�H;&�H;��H;#�H;�H;Y�H;��H;@�H;pzH;ZH;u/H;��G;J�G;~FG;6PF;7�C;�>;��3;"m;E��:�j~:�����.�����%+��I����μ�����N�x^��6S�����MZ�#,�z�H��9b�)�v�*��      ����)����:���M��E�r�'�O�#,�X�
��gٽqĥ���u�x1�j���+Ϥ���P�[��.o��p�� :Y��:�P;7�/;4�<; C;�E;f!G;.�G;��G;�%H;�RH;�tH;�H;A�H;ӯH;��H;V�H; �H;V�H;��H;ӯH;@�H;�H;�tH;�RH;�%H;��G;.�G;n!G;�E; C;3�<;4�/;�P;]��::�p���.o�[򻬎P�+Ϥ�i���w1���u�qĥ��gٽX�
�#,�'�O�E�r��M���:��)���      8���v��L;������SP��E�r�z�H�U� ���6@��ѓ����K�b��վ���s�t���񕻵ܺ`4u9 &�:�;&�+;x�:;�"B;h�E;��F;͐G;��G;(H;0LH;�oH;6�H;o�H;��H;/�H;ּH;�H;мH;2�H;��H;n�H;7�H;�oH;:LH;+H;��G;ѐG;��F;g�E;�"B;t�:;&�+;�;&�:P4u9�ܺ��t����s��վ�b���K�ѓ��6@����U� �z�H�E�r�SP������M;���v��      UVھ�*־/5ʾr��������M���9b��5�����ս����Xc���̖ռ�I��X�$�pT���Z�`]���:��;d�';�8;RA;�9E;}�F;��G;��G;=H;GH;lH;?�H;4�H;ݫH;��H;��H;N�H;��H;��H;۫H;6�H;?�H;lH;GH;?H;��G;��G;��F;�9E;RA;�8;c�';��;�:�]���Z�oT��W�$��I��̖ռ���Xc������ս���5��9b��M������r���/5ʾ�*־      ���쾴�޾05ʾM;���:��)�v��E�`'����r����u���+��W��A����4���Ļ(9)��j��mW�:Z�;%;�k7; �@;��D;��F;�wG;P�G;.H;9CH;$iH;	�H;��H;��H;��H;��H;o�H;��H;��H;��H;��H;	�H;!iH;ACH;1H;Q�G;�wG;��F;��D;�@;�k7;�%;Z�;uW�:�j��&9)���Ļ��4��A���W缄�+���u�r�����`'��E�)�v��:��M;��05ʾ��޾��      Vh���b���쾧*־�v��)���*��(�O�U� �s��r���؀�G�3���@ݜ�?�>�V�ѻ�9����o�:8% ;lM#;<�6;HA@;��D;��F;qG;H�G;H;�@H;cgH;��H;��H;٩H;�H;��H;ڻH;�H;�H;۩H;��H;��H;`gH;�@H;H;H�G;qG;��F;��D;EA@;7�6;jM#;6% ;o�:����9�W�ѻ?�>�@ݜ���F�3��؀��r��s�V� �'�O�*��)����v���*־���b��      1�$��� ����#��@��(�þ�*��1Dx���=�����Pν���#'K��c���r�V����E^���S�jw[:���:e;%�4;A`?;�mD;M�F;FvG;�G;:H;]OH;�sH;��H;w�H;|�H;�H;P�H;#�H;L�H;�H;}�H;u�H;��H;�sH;hOH;:H;�G;JvG;X�F;�mD;=`?;�4;e;���:vw[:��S�E^����q�V����c�"'K�����Pν�����=�1Dx��*��(�þ@��#������� �      �� ����R��O��/������0��5�s�׀:�g9��ʽ2Z����G��8�.���5S����0X���D�NBd:�B�: ;��4;Ĉ?;�~D;	�F;	yG;��G;L H;&PH;tH;�H;ȢH;°H;'�H;m�H;1�H;j�H;)�H;ðH;ȢH;�H;tH;0PH;O H;��G;yG;�F;�~D;��?;��4;� ;�B�:^Bd:��D�0X���껰5S�.���8���G�2Z���ʽg9�׀:�4�s��0�����/��O��R�����      ���R��8�
������Yؾ ���ޥ����f���0�[[�N8��ϐ���>�����KȤ��6H�f�ܻrF�����}:��:]";+�5;��?;M�D;��F;�G;��G;-#H;]RH;�uH;B�H;��H;s�H;��H;�H;��H;�H;��H;s�H;��H;B�H;�uH;dRH;/#H;��G;�G;��F;O�D;��?;$�5;[";��:�}:��rF�f�ܻ�6H�JȤ������>�ϐ��N8��Z[���0���f�ޥ�� ����Yؾ����8�
�R��      #��N������=I�(�þ�R��;���tS��Q"��s������}��0��켉�����6�L�ƻ@}*�X�����:vx;T%;�l7;ֳ@;��D;��F;��G;��G;�'H;�UH;ZxH;H�H;B�H;��H;��H;��H;t�H;��H;��H;��H;@�H;H�H;WxH;�UH;�'H;�G;��G;��F;��D;ҳ@;�l7;R%;tx;��:X���>}*�K�ƻ��6��������0���}�����s��Q"�tS�;����R��(�þ=Iᾤ���O��      @��0�待Yؾ(�þ
Ī�|쏾�k�׀:�~�{�ؽ�����c�]y���Ҽ����F� �n�2�� (75�:��
;��(;}_9;��A;a\E;h�F;��G;��G;�.H;�ZH;�{H;�H;E�H;M�H;�H;��H;t�H;��H;	�H;M�H;D�H;�H;�{H;�ZH;�.H;��G;��G;p�F;c\E;��A;v_9;��(;��
;?�: (71��m�F� �������Ҽ]y��c�����|�ؽ~�׀:��k�|쏾
Ī�(�þ�Yؾ0��      '�þ�������R��|쏾5�s��H�����������ΐ����D��c�����?�f�V,�����P�� �9���:�;j-;K�;;n�B;��E;VG;��G;��G;~6H;�`H;T�H;H�H;ЩH;J�H;��H;O�H;��H;L�H;��H;H�H;ΩH;H�H;S�H;�`H;�6H;��G;��G;]G;��E;k�B;E�;;j-;�;ų�: �9�P�����V,�>�f������c���D�ΐ�������������H�5�s�|쏾�R�� ������      �*���0��ޥ��;����k��H��#%�Z[��Pνt��a�f�3/%���伆���w�=��?ػ�FL���D�D�R:��:-�;.2;��=;��C;a0F;@GG;��G;!H;�?H;�gH;��H;&�H;��H;��H;|�H;��H;p�H;��H;}�H;��H;��H;%�H;�H;�gH;�?H;!H;��G;GGG;d0F;��C;��=;.2;+�;��:H�R:��D��FL��?ػv�=��������2/%�a�f�t���PνZ[��#%��H��k�;���ޥ���0��      1Dx�4�s���f�tS�׀:����Z[��7ս�榽��}���;��8�V�����r����?G���� ά���:�;�}$;��6;��?;�D;��F;�pG;��G;�H;JH;;oH;6�H;r�H;��H;3�H;��H;��H;#�H;��H;��H;6�H;��H;p�H;7�H;DoH;!JH;�H;��G;�pG;ĔF;�D;��?;��6;�}$;
�;��: ά���>G�������r�V����8���;���}��榽�7սZ[����׀:�tS���f�4�s�      ��=�׀:���0��Q"�~������Pν�榽@����G�2����Ҽ ��KE:�B�ܻ�D^�ʸ��<i:/��:�;2|,;��:;G�A;;iE;��F;�G;}�G;�(H;.UH;vwH;l�H;�H;��H;�H;��H;��H;�H;��H;��H;�H;��H;�H;l�H;}wH;2UH;�(H;{�G;�G;��F;:iE;K�A;��:;2|,;�;3��:<i:¸���D^�@�ܻJE:� ����Ҽ2����G�@���榽�Pν����~��Q"���0�׀:�      ���g9�Z[��s�{�ؽ���t����}���G������2c��Y�V�H,��*����������:��:J ;^�3;�0>;��C;�F;�8G;&�G;eH;�7H;�`H;�H;�H;��H;G�H;��H;B�H;��H;�H;��H;G�H;��H;E�H;��H;�H;�H;�`H;�7H;fH;'�G;�8G;�F;ÚC;�0>;\�3;Q ;��:��:@������*��G,�X�V�1c���������G���}�t�����|�ؽ�s�Z[�g9�      �Pν�ʽO8���������ΐ��a�f���;�2�����CȤ�6�f�,��Rߵ�^o5���D��-:6��:�>;�+;�_9;�A;a�D;�F;�vG;��G;H;nGH;TlH;��H;��H;�H;)�H;��H;��H;�H;!�H;�H;��H;��H;(�H;�H;��H;ňH;^lH;tGH;H;��G;�vG;�F;e�D;�A;�_9;�+;�>;6��:(�-:��D�Zo5�Pߵ�+��5�f�CȤ����2����;�a�f�ΐ���������O8���ʽ      ���2Z��ϐ����}��c���D�2/%��8���Ҽ1c��5�f�����ƻ�/X�j���P��9��:5�;�";��3;7>;;YC;n�E;�G;�G;^�G;�,H;�VH;xH;��H;+�H;�H;�H;��H;-�H;A�H;,�H;B�H;.�H;��H;�H;�H;/�H;��H;xH;WH;�,H;_�G;�G;�G;u�E;DYC;8>;��3;�";5�;�:P��9f����/X��ƻ���4�f�1c����Ҽ�8�2/%���D��c���}�ϐ��2Z��      #'K���G��>��0�\y��c����U��� ��X�V�+���ƻ�od���º s(7y4�:���:��;�P.;ˡ:;zA;&�D;¨F;GnG;2�G;�H;�@H;fH;Y�H;(�H;��H;иH;��H;��H;��H;w�H;5�H;x�H;��H;��H;��H;θH;��H;0�H;a�H;!fH;�@H;�H;;�G;JnG;ƨF;,�D;zA;֡:;�P.;��;���:�4�: v(7��º�od��ƻ*��X�V� ��T�����伖c�]y��0��>���G�      �c��8���������Ҽ����������r�KE:�G,�Pߵ��/X���º@Ȭ�@�}:� �:�;A�);m7;�?;��C;F;O)G;	�G;?�G;�)H;�SH;�tH;X�H;w�H;�H;��H;��H;��H;�H;��H;I�H;��H;�H;��H;��H;��H;�H;��H;c�H;�tH;�SH;�)H;H�G;�G;Y)G;F;��C;�?;!m7;?�);�;� �:L�}:�Ǭ���º�/X�Nߵ�G,�HE:���r�����������Ҽ�켸����8�      ��.��KȤ���������>�f�v�=����B�ܻ�*��Zo5�v��� r(7H�}:�n�:#�;�>&;��4;��=;��B;�E;�F;��G;��G;$H;}AH;�eH;7�H;͘H;T�H;׷H;d�H;�H;��H;h�H;��H;N�H;��H;g�H;��H;�H;b�H;ڷH;[�H;֘H;=�H;�eH;zAH;.H;��G;��G;�F;�E;��B;��=;��4;�>&;#�;�n�:T�}: u(7l���Vo5��*��=�ܻ���v�=�<�f���������LȤ�.��      l�V��5S��6H���6�F� �W,��?ػ<G���D^������D�8��9s4�:� �:#�;�%;��3;�<;NB;�E;��F;�XG;��G;? H;d0H;HWH;UvH;�H;u�H;��H;��H;��H;m�H;K�H;��H;��H;5�H;��H;��H;K�H;j�H;��H;��H;��H;|�H;�H;YvH;DWH;i0H;B H;��G;�XG;��F;�E;RB;�<;��3;�%;'�;� �:u4�:H��9��D�����D^�:G���?ػT,�H� ���6��6H��5S�      ��ﻰ��k�ܻN�ƻj󩻽���FL���¸�� �� �-:��:���:�;�>&;��3;J9<;�A;԰D;;ZF;5G;��G;��G;c!H;'JH;*kH;��H;��H;^�H;��H;��H;��H;��H;��H;��H;a�H;��H;^�H;��H;��H;��H;��H;��H;��H;d�H;��H;��H;(kH;/JH;h!H;��G;��G;5G;BZF;װD;	�A;M9<;��3;�>&;�;���:��:4�-: ���������FL����n�P�ƻp�ܻ���      �D^� 0X�rF�6}*�$���P����D��ͬ�@i:��::��:/�;��;>�);��4;�<;�A; �D;o9F;�G;h�G;>�G;7H;?H;UaH;}H;x�H;q�H;��H;߾H;��H;_�H;|�H;�H;��H;%�H;��H;#�H;��H;�H;x�H;\�H;��H;�H;��H;s�H;y�H;}H;[aH;?H;7H;B�G;k�G;�G;r9F;�D;�A;�<;��4;>�);��;0�;D��:��:Pi: ͬ���D��P��"��<}*�rF��/X�      h�S���D���� ��� (7`�9l�R:��:3��:��:�>;�";�P.; m7;��=;QB;ְD;y9F;G;�G;M�G;�H;�6H;eYH;�uH;�H;�H;��H;��H;��H;�H;��H;�H;5�H;^�H;��H;��H;��H;]�H;4�H;�H;��H;�H;��H;��H;��H;�H;�H;�uH;iYH;�6H;�H;Q�G;�G;G;p9F;װD;LB;��=; m7;�P.;�";�>;��:9��:��:\�R:0�9 (7���������D�      >w[:>Bd:�}:��:1�:���:��:�;�;P ;�+;��3;ҡ:;�?;��B;�E;AZF;�G;�G;k�G;8H;N1H;�SH;[pH;ԇH;D�H;�H;u�H;��H;��H;��H;��H;o�H;!�H;��H;�H;X�H;�H;��H;�H;o�H;��H;��H;��H;��H;y�H;�H;B�H;هH;^pH;�SH;P1H;>H;k�G;�G;�G;AZF;�E;��B;	�?;ѡ:;��3;�+;O ;�;	�;��:ϳ�:5�:��:��}:Bd:      ��:�B�:���:hx;��
;�;)�;�}$;.|,;^�3;�_9;3>;zA;��C;�E;��F;5G;q�G;P�G;8H;�/H;�PH;�lH;C�H;��H;��H;k�H;��H;�H;�H;Z�H;��H;��H;��H;i�H;K�H;��H;D�H;j�H;��H;��H;��H;\�H;�H;��H;��H;h�H;��H;��H;C�H;�lH;�PH;�/H;8H;Q�G;m�G;5G;��F;�E;��C;zA;3>;�_9;[�3;,|,;�}$;/�;�;��
;hx;Ć�:�B�:      e; ;j";`%;��(;j-;*2;��6;��:;�0>;�A;;YC;)�D;F;�F;�XG;��G;C�G;�H;P1H;�PH;�kH;r�H;x�H;.�H;+�H;ӼH;��H;��H;�H;j�H;��H;u�H;n�H;��H;`�H;��H;Z�H;��H;m�H;s�H;��H;m�H;�H;��H;��H;μH;)�H;2�H;w�H;k�H;�kH;�PH;P1H;�H;@�G;��G;�XG;�F;�F;&�D;;YC;�A;�0>;��:;��6;.2;j-;��(;R%;]";� ;      7�4;��4;!�5;�l7;t_9;M�;;��=;�?;O�A;ĚC;j�D;u�E;ƨF;[)G;��G; �G;��G;AH;�6H;�SH;�lH;p�H;��H;�H;��H;N�H;�H;/�H;��H;�H;�H;��H;2�H;��H;��H;a�H;��H;[�H;��H;��H;.�H;��H;�H;~�H;��H;2�H;�H;N�H;��H;�H;��H;p�H;�lH;�SH;�6H;7H;��G;��G;��G;U)G;èF;u�E;h�D;��C;N�A;�?;��=;K�;;�_9;�l7;�5;��4;      @`?;ˈ?;��?;ѳ@;��A;n�B;��C;�D;0iE;�F;�F;�G;JnG;�G;��G;E H;f!H;?H;iYH;[pH;E�H;s�H;�H;B�H;��H;#�H;?�H;�H;��H;r�H;R�H;��H;��H;��H;��H;<�H;M�H;6�H;��H;��H;��H;��H;S�H;p�H;��H;�H;:�H;%�H;��H;?�H; �H;v�H;A�H;WpH;cYH;?H;f!H;B H;��G;�G;EnG;�G;�F;�F;5iE;�D;��C;[�B;��A;˳@;��?;È?;      �mD;�~D;I�D;��D;\\E;��E;m0F;��F;��F;�8G;�vG;�G;9�G;L�G;-H;p0H;3JH;eaH;�uH;��H;��H;4�H;��H;��H;��H;��H;g�H;�H;��H;��H;\�H;@�H;��H;��H;��H;��H;)�H;��H;��H;��H;��H;:�H;^�H;��H;��H;�H;c�H;��H;��H;��H;��H;2�H;��H;ڇH;�uH;^aH;0JH;l0H;+H;F�G;8�G;�G;�vG;�8G;��F;��F;k0F;��E;d\E;��D;H�D;�~D;      B�F;�F;��F;��F;b�F;[G;JGG;�pG;�G;-�G;��G;c�G;�H;*H;}AH;LWH;-kH;}H;�H;B�H;��H;%�H;K�H;%�H;��H;-�H;��H;}�H;��H;�H;�H;��H;��H;��H;:�H;��H;��H;��H;7�H;��H;��H;��H;�H;�H;��H;}�H;��H;0�H;��H;"�H;I�H;'�H;��H;@�H;�H;}H;,kH;HWH;zAH;�)H;�H;b�G;��G;+�G;�G;�pG;FGG;OG;u�F;��F;��F;�F;      [vG;yG;��G;��G;��G;��G;��G;��G;x�G;fH;H;�,H;�@H;�SH;�eH;YvH;��H;}�H;�H;�H;o�H;ѼH;"�H;D�H;e�H;��H;`�H;[�H;��H;��H;^�H;��H;��H;@�H;��H;%�H;#�H;�H;��H;A�H;��H;��H;^�H;��H;��H;Y�H;\�H;��H;h�H;?�H; �H;ӼH;n�H;ߪH;�H;v�H;��H;UvH;�eH;�SH;�@H;�,H;H;dH;w�G;��G;��G;�G;��G;}�G; �G;�xG;      �G;��G;��G;��G;��G;��G;,H;�H;�(H;�7H;tGH;WH; fH;�tH;9�H;�H;��H;s�H;��H;u�H;��H;~�H;-�H;�H;�H;|�H;[�H;��H;��H;e�H;��H;��H;V�H;��H;O�H;��H;��H;��H;M�H;��H;V�H;��H;��H;d�H;��H;��H;U�H;}�H;�H;�H;-�H;�H;��H;t�H;��H;o�H;��H;�H;6�H;�tH;fH;WH;vGH;�7H;�(H;�H;*H;{�G;��G;��G;��G;��G;      4H;A H;*#H;�'H;p.H;~6H;�?H;JH;'UH;�`H;[lH;xH;]�H;]�H;јH;|�H;g�H;��H; �H;��H;��H;��H;��H;��H;��H;��H;��H;��H;1�H;��H;��H;O�H;��H;r�H;��H;��H;��H;��H;��H;s�H;��H;I�H;��H;��H;.�H;��H;��H;��H;��H;��H;��H;��H;��H;��H;��H;��H;d�H;|�H;јH;\�H;Y�H;xH;]lH;�`H;(UH;JH;�?H;z6H;|.H;�'H;(#H;C H;      \OH;PH;iRH;�UH;�ZH;�`H;�gH;:oH;{wH;�H;H;��H;/�H;��H;U�H;��H;��H;߾H;��H;��H;�H;�H;z�H;n�H;��H;�H;��H;d�H;��H;��H;H�H;��H;g�H;��H;��H;�H;4�H;�H;��H;��H;g�H;��H;H�H;�H;��H;a�H;��H;�H;��H;i�H;{�H;�H;�H;��H;��H;ݾH;��H;��H;U�H;�H;/�H;��H;ÈH;�H;ywH;@oH;�gH;�`H;�ZH;�UH;gRH;PH;      �sH;&tH;�uH;]xH;�{H;V�H;��H;:�H;p�H;�H;��H;4�H;��H;��H;ݷH;��H;��H;��H; �H;��H;a�H;m�H;�H;R�H;\�H;
�H;]�H;��H;��H;O�H;��H;k�H;��H;�H;X�H;c�H;[�H;a�H;W�H;�H;��H;h�H;��H;N�H;��H;��H;Z�H;�H;a�H;P�H;�H;k�H;]�H;��H; �H;��H;��H;��H;ݷH;��H;��H;6�H;��H;�H;p�H;=�H;��H;J�H;�{H;[xH;�uH;)tH;      ��H;�H;C�H;G�H;�H;?�H;0�H;s�H;&�H;��H;��H;�H;׸H;��H;c�H;��H;��H;c�H;��H;��H;��H;��H;��H;��H;=�H;��H;��H;��H;L�H;��H;d�H;��H;�H;Z�H;��H;�H;��H;��H;��H;[�H;�H;��H;b�H;��H;I�H;��H;��H;��H;@�H;��H;��H;��H;��H;��H;��H;d�H;��H;��H;d�H;��H;ָH;�H;��H;��H;$�H;u�H;5�H;A�H;�H;G�H;M�H;
�H;      ~�H;֢H;̣H;C�H;N�H;ΩH;��H;��H;��H;K�H;/�H;�H;��H;��H; �H;p�H;��H;��H;�H;s�H;��H;v�H;.�H;��H;��H;��H;��H;Z�H;��H;k�H;��H;�H;P�H;��H;��H;��H;��H;��H;��H;��H;S�H;�H;��H;g�H;��H;U�H;��H;��H;��H;��H;2�H;u�H;��H;r�H;�H;��H;��H;s�H; �H;��H;��H;�H;0�H;K�H;��H;��H;��H;ɩH;S�H;=�H;֣H;֢H;      z�H;��H;t�H;��H;Q�H;A�H;��H;9�H;�H;��H;��H;��H;��H;��H;��H;R�H;��H;�H;9�H;#�H;��H;n�H;��H;��H;��H;��H;:�H;��H;r�H;��H;�H;[�H;��H;��H;��H;��H;��H;��H;��H;��H;��H;Z�H;�H;��H;n�H;��H;9�H;��H;��H;��H;��H;m�H;��H;�H;8�H;�H;��H;T�H;��H;��H;��H;��H;��H;��H;��H;;�H;��H;@�H;X�H;��H;~�H;ʰH;      �H;=�H;κH;��H;�H;��H;��H;��H;��H;O�H;��H;:�H;��H;�H;o�H;��H;��H;��H;^�H;��H;m�H;��H;��H;��H;��H;0�H;��H;O�H;��H;�H;Q�H;��H;��H;��H;��H;��H;��H;��H;��H;��H;��H;��H;P�H;��H;��H;J�H;��H;0�H;��H;��H;��H;��H;f�H;��H;\�H;��H;��H;��H;n�H;�H;��H;:�H;��H;P�H;��H;��H;��H;��H;�H;��H;ϺH;<�H;      L�H;j�H;�H;��H;��H;D�H;��H;��H;��H;��H;�H;I�H;~�H;��H;��H;��H;b�H;!�H;��H;�H;L�H;[�H;X�H;+�H;��H;��H;"�H;��H;��H;$�H;a�H;��H;��H;��H;��H;��H;��H;��H;��H;��H;��H;��H;_�H;�H;��H;��H; �H;��H;��H;,�H;\�H;X�H;E�H;�H;��H;&�H;c�H;��H;��H;��H;}�H;H�H;�H;��H;��H;��H;�H;G�H;��H;��H;�H;y�H;      +�H;/�H;��H;w�H;r�H;��H;z�H;&�H;�H;�H;0�H;:�H;A�H;W�H;X�H;<�H;��H;��H;��H;_�H;��H;��H;��H;C�H;)�H;��H;�H;��H;��H;<�H;X�H;��H;��H;��H;��H;��H;��H;��H;��H;��H;��H;��H;W�H;8�H;��H;��H; �H;��H;(�H;D�H;��H;��H;��H;[�H;��H;��H;��H;<�H;V�H;W�H;@�H;:�H;0�H;�H;�H;*�H;|�H;��H;t�H;w�H;��H;8�H;      N�H;n�H;�H;��H;��H;I�H;��H;��H;��H;��H;	�H;H�H;�H;��H;��H;��H;b�H;#�H;��H;�H;N�H;]�H;X�H;+�H;��H;��H;"�H;��H;��H;#�H;a�H;��H;��H;��H;��H;��H;��H;��H;��H;��H;��H;��H;_�H;�H;��H;��H;�H;��H;��H;,�H;^�H;X�H;E�H;�H;��H;%�H;b�H;��H;��H;��H;~�H;H�H;�H;��H;��H;��H; �H;E�H;��H;��H;�H;v�H;      ܹH;A�H;ȺH;��H;�H;��H;��H;��H;��H;O�H;��H;:�H;��H;�H;q�H;��H;��H;��H;]�H;��H;n�H;��H;��H;��H;��H;/�H;��H;M�H;��H; �H;Q�H;��H;��H;��H;��H;��H;��H;��H;��H;��H;��H;��H;Q�H;��H;��H;I�H;��H;4�H;��H;��H;��H;��H;d�H;��H;\�H;��H;��H;��H;m�H;�H;��H;;�H;��H;N�H;��H;��H;��H;��H;�H;��H;κH;?�H;      z�H;��H;t�H;��H;Q�H;F�H;��H;;�H;��H;��H;��H;��H;��H;��H;��H;R�H;��H;!�H;9�H;"�H;��H;p�H;��H;��H;��H;��H;=�H;��H;r�H;��H;�H;[�H;��H;��H;��H;��H;��H;��H;��H;��H;��H;X�H;�H;��H;l�H;��H;:�H;��H;��H;��H;��H;m�H;��H;�H;6�H;�H;��H;T�H;��H;��H;��H;��H;��H;��H;��H;=�H;��H;C�H;Z�H;��H;}�H;��H;      |�H;ܢH;ˣH;@�H;I�H;ѩH;��H;��H;��H;K�H;0�H;�H;��H;��H;"�H;q�H;��H;��H;�H;v�H;��H;v�H;,�H;��H;��H;��H;��H;Z�H;��H;l�H;��H;�H;N�H;��H;��H;��H;��H;��H;��H;��H;Q�H;�H;��H;g�H;��H;U�H;��H;��H;��H;��H;5�H;u�H;��H;r�H;�H;�H;��H;q�H; �H;��H;��H;�H;/�H;I�H;��H;��H;��H;˩H;O�H;G�H;ףH;բH;      ��H;�H;4�H;C�H;�H;P�H;1�H;v�H;#�H;��H;��H;�H;ָH;��H;g�H;��H;��H;d�H;��H;��H;��H;��H;��H;��H;@�H;��H;��H;��H;O�H;��H;d�H;��H;�H;X�H;��H;�H;��H;��H;��H;Z�H;�H;��H;`�H;��H;H�H;��H;��H;��H;>�H;��H;��H;��H;��H;��H;��H;c�H;��H;��H;d�H;��H;ָH;�H;��H;��H;&�H;w�H;7�H;C�H;�H;D�H;:�H;�H;      �sH;&tH;�uH;WxH;�{H;V�H;��H;9�H;p�H;�H;��H;8�H;��H;��H;޷H;��H;��H;��H; �H;��H;c�H;n�H;�H;R�H;^�H;�H;Z�H;��H;��H;N�H;��H;l�H;��H;�H;Z�H;b�H;[�H;c�H;W�H;�H;��H;i�H;��H;I�H;��H;��H;[�H;�H;^�H;O�H;�H;n�H;]�H;��H;"�H;��H;��H;��H;�H;��H;��H;6�H;��H;�H;p�H;@�H;��H;Q�H;�{H;bxH;�uH;'tH;      kOH;&PH;bRH;�UH;�ZH;�`H;�gH;DoH;wH;�H;ňH;��H;0�H;�H;Y�H;��H;��H;�H;��H;��H;�H;	�H;v�H;k�H;��H;�H;��H;b�H;��H;��H;I�H;��H;e�H;��H;��H;�H;4�H;�H;��H;��H;h�H;��H;H�H;|�H;��H;^�H;��H;�H;��H;h�H;��H;�H;�H;��H;��H;ھH;��H;��H;V�H;��H;/�H;��H;ÈH;
�H;{wH;BoH;�gH;�`H;�ZH;�UH;tRH;PH;      DH;A H;;#H;�'H;g.H;�6H;�?H;JH;/UH;�`H;ZlH;xH;\�H;_�H;ԘH;~�H;e�H;��H;��H;��H;��H;��H;��H;��H;��H;��H;��H;��H;3�H;��H;��H;P�H;��H;s�H;��H;��H;��H;��H;��H;r�H;��H;N�H;��H;��H;-�H;��H;��H;��H;��H;��H;��H;��H;��H;��H;��H;��H;e�H;|�H;ӘH;]�H;]�H;xH;^lH;�`H;1UH;JH;�?H;6H;z.H;�'H;:#H;; H;      �G;��G;��G;��G;��G;��G;*H;�H;�(H;�7H;tGH;WH;fH;�tH;:�H;�H;��H;t�H;��H;u�H;��H;��H;*�H;�H;�H;u�H;V�H;��H;��H;a�H;��H;��H;U�H;��H;P�H;��H;��H;��H;O�H;��H;W�H;��H;��H;a�H;��H;��H;X�H;{�H;�H; �H;3�H;�H;��H;t�H;��H;m�H;��H;�H;<�H;�tH; fH;WH;vGH;�7H;�(H;�H;*H;��G;��G;��G;��G;��G;      IvG;yG; �G;��G;��G;��G;��G;��G;x�G;dH;H;�,H;�@H;�SH;�eH;XvH;��H;}�H;�H;ݪH;p�H;ԼH;�H;D�H;g�H;��H;]�H;[�H;��H;��H;]�H;��H;��H;A�H;��H; �H;#�H; �H;��H;B�H;��H;��H;`�H;��H;��H;Y�H;]�H;��H;h�H;?�H;&�H;ӼH;n�H;�H;�H;x�H;��H;YvH;�eH;�SH;�@H;�,H;H;eH;z�G;��G;��G;��G;��G;��G;�G;yG;      <�F;�F;��F;��F;h�F;cG;CGG;�pG;�G;*�G;��G;e�G;�H;�)H;{AH;IWH;)kH;}H;�H;@�H;��H;%�H;G�H;%�H;��H;*�H;��H;�H;��H;�H;�H;��H;��H;��H;:�H;��H;��H;��H;7�H;��H;��H;��H;�H;�H;��H;y�H;��H;/�H;��H;"�H;N�H;%�H;��H;A�H;�H;}H;-kH;KWH;�AH;�)H;�H;c�G;��G;.�G;�G;�pG;DGG;UG;p�F;��F;��F;��F;      �mD;�~D;H�D;��D;Z\E;��E;k0F;��F;��F;�8G;�vG;�G;7�G;H�G;.H;n0H;0JH;baH;�uH;ۇH;��H;5�H;��H;��H;��H;��H;c�H;�H;��H;��H;\�H;A�H;��H;��H;��H;��H;(�H;��H;��H;��H;��H;A�H;b�H;��H;��H;�H;d�H;��H;��H;��H;��H;5�H;��H;݇H;�uH;^aH;2JH;n0H;1H;I�G;9�G;�G;�vG;�8G;��F;��F;l0F;��E;d\E;��D;I�D;�~D;      "`?;��?;��?;ڳ@;��A;w�B;��C;�D;>iE;�F;�F;�G;EnG;�G;��G;D H;e!H;?H;bYH;XpH;C�H;s�H;��H;B�H;��H;�H;<�H;�H;��H;n�H;S�H;��H;��H;��H;��H;7�H;O�H;9�H;��H;��H;��H;��H;W�H;p�H;��H;�H;?�H;#�H;��H;B�H;�H;s�H;C�H;[pH;fYH;?H;h!H;E H;��G;�G;GnG;�G; �F;�F;8iE;�D;��C;k�B;��A;�@;��?;��?;      )�4;��4;�5;�l7;r_9;H�;;��=;�?;R�A;��C;e�D;u�E;èF;Y)G;��G;��G;��G;>H;�6H;�SH;�lH;p�H;��H;�H;��H;H�H;�H;0�H;��H;z�H;�H;��H;0�H;��H;��H;a�H;��H;_�H;��H;��H;0�H;��H;�H;��H;��H;/�H;�H;L�H;��H;�H;��H;p�H;�lH;�SH;�6H;:H;��G;��G;��G;X)G;ƨF;t�E;e�D;C;O�A;�?;��=;K�;;r_9;�l7;�5;��4;      e; ;]";T%;��(;j-;02;��6;��:;�0>;�A;>YC;)�D;F;�F;�XG;��G;C�G;�H;Q1H;�PH;�kH;m�H;w�H;4�H;$�H;мH;��H;��H;�H;m�H;��H;s�H;n�H;��H;[�H;��H;]�H;��H;k�H;u�H;��H;p�H;�H;��H;~�H;ѼH;)�H;.�H;z�H;q�H;�kH;�PH;T1H;�H;@�G;��G;�XG;�F;F;)�D;;YC;�A;�0>;��:;6;*2;	j-;��(;F%;]";� ;       ��:�B�:҆�:px;~�
;�;,�;�}$;2|,;Y�3;�_9;4>;zA;��C;�E;��F;5G;q�G;P�G;:H;�/H;�PH;�lH;E�H;��H;��H;e�H;��H;��H;�H;Z�H;��H;��H;��H;j�H;G�H;��H;H�H;i�H;��H;��H;��H;^�H;�H;�H;��H;i�H;��H;��H;E�H;�lH;�PH;�/H;:H;Q�G;n�G;5G;��F;�E;��C;	zA;3>;�_9;^�3;2|,;�}$;0�;�;��
;ox;��:�B�:      �w[:bBd:��}:��:1�:ϳ�:�:�;�;P ;�+;��3;ӡ:;�?;��B;�E;AZF;�G;�G;k�G;>H;S1H;�SH;]pH;ڇH;B�H;ܪH;u�H;��H;��H;��H;��H;p�H;!�H;��H;�H;[�H;�H;��H;�H;p�H;��H;��H;��H;��H;t�H;�H;D�H;ԇH;`pH;�SH;P1H;;H;k�G;�G;�G;?ZF;�E;��B;
�?;ӡ:;��3;�+;O ;�;�;��:���:;�:��:�}:>Bd:      `�S���D���(��� (7X�9d�R:��:=��:��:�>;�";�P.; m7;��=;QB;԰D;t9F;G;�G;R�G;�H;�6H;fYH;�uH;�H;�H;��H;��H;��H;�H;��H;�H;6�H;^�H;��H;��H;��H;]�H;5�H;�H;��H;�H;��H;��H;��H;�H;�H;�uH;iYH;�6H;�H;P�G;�G;G;p9F;ְD;NB;��=; m7;�P.;�";�>;��:9��:!��:d�R:P�9 (7(�������D�      
E^��/X�rF�9}*� ���P����D��̬�Xi:��:B��:2�;��;?�);��4;�<;�A;�D;p9F;�G;m�G;@�G;;H;?H;[aH;}H;u�H;q�H;��H;ݾH;��H;]�H;|�H;�H;��H;#�H;��H;&�H;��H;�H;|�H;\�H;��H;�H;��H;p�H;x�H;}H;UaH;?H;8H;>�G;g�G;�G;o9F;�D;�A;�<;��4;;�);��;/�;D��:��:Ti: ͬ���D��P��"��=}*�rF��/X�      ��ﻱ��k�ܻK�ƻi󩻻���FL�	������ ��0�-:��:���:�;�>&;��3;M9<;�A;԰D;?ZF;5G;��G;��G;i!H;/JH;*kH;��H;��H;e�H;��H;��H;��H;��H;��H;��H;a�H;��H;a�H;��H;��H;��H;��H;��H;��H;d�H;��H;��H;(kH;)JH;i!H;��G;��G;5G;AZF;԰D;	�A;K9<;��3;�>&;�;���:��:(�-: ������
���FL����o�O�ƻp�ܻ���      l�V��5S��6H���6�F� �T,��?ػ9G���D^������D�P��9w4�:� �:)�;�%;��3;�<;NB;�E;��F;�XG; �G;D H;i0H;IWH;UvH;�H;{�H;��H;��H;��H;m�H;Q�H;��H;��H;5�H;��H;��H;J�H;j�H;��H;��H;��H;z�H;�H;TvH;GWH;d0H;? H;��G;�XG;��F;�E;KB;�<;��3;�%;&�;� �:y4�:@��9��D�����D^�;G���?ػT,�H� ���6��6H��5S�      ��.��LȤ���������=�f�v�=����@�ܻ�*��Vo5�p��� u(7T�}:�n�:&�;�>&;��4;��=;��B;�E;�F;��G;��G;-H;~AH;�eH;:�H;ԘH;V�H;۷H;d�H;�H;��H;g�H;��H;N�H;��H;g�H;��H;�H;_�H;ٷH;U�H;ԘH;7�H;�eH;zAH;'H;��G;��G;�F;ލE;��B;��=;��4;�>&;"�;�n�:L�}: r(7p���Yo5��*��?�ܻ���v�=�<�f���������LȤ�.��      �c��8���������Ҽ����������r�IE:�G,�Nߵ��/X���º�Ǭ�X�}:� �:�;>�);m7;
�?;��C;F;V)G;�G;I�G;�)H;�SH;�tH;_�H;|�H;�H;��H;��H;��H;�H;��H;J�H;��H;�H;��H;��H;��H;�H;~�H;_�H;�tH;�SH;�)H;?�G;�G;V)G;F;��C;�?;m7;>�);�;� �:H�}: Ȭ���º�/X�Oߵ�G,�JE:���r�����������Ҽ�켷����8�      #'K���G��>��0�\y��c����T��� ��X�V�*���ƻ�od���º z(74�:���:��;�P.;ϡ:;zA;'�D;ƨF;NnG;;�G;�H;�@H; fH;`�H;,�H;��H;ӸH;��H;��H;��H;z�H;3�H;x�H;��H;��H;��H;͸H;��H;+�H;]�H;fH;�@H;�H;2�G;HnG;ƨF;'�D;zA;ҡ:;�P.;��;���:y4�: x(7��º�od��ƻ+��X�V� ��T�����伕c�^y��0��>���G�      ���2Z��ϐ����}��c���D�2/%��8���Ҽ1c��4�f�����ƻ�/X�f���h��9��:0�;�";��3;;>;=YC;w�E;�G;�G;b�G;�,H;�VH;xH;��H;1�H;�H;�H;��H;-�H;@�H;,�H;A�H;,�H;��H;�H;�H;+�H;��H;xH;�VH;�,H;^�G;�G;�G;u�E;=YC;3>;��3;�";2�;��:H��9f����/X��ƻ���5�f�1c����Ҽ�8�2/%���D��c���}�ϐ��2Z��      �Pν�ʽO8���������ΐ��a�f���;�2�����CȤ�5�f�+��Pߵ�Yo5���D��-:0��:�>;�+;�_9;�A;f�D;�F;�vG;��G;H;tGH;[lH;��H;��H;�H;*�H;��H;��H;�H;!�H;�H;��H;��H;&�H;�H;��H;��H;ZlH;oGH;H;��G;�vG;�F;e�D;�A;�_9;�+;�>;0��:�-:��D�[o5�Rߵ�+��6�f�CȤ����2����;�a�f�ΐ���������O8���ʽ      ���g9�Z[��s�{�ؽ���t����}���G������1c��X�V�G,��*�����P��~�:��:O ;b�3;�0>;ÚC;�F;�8G;'�G;eH;�7H;�`H;�H;�H;��H;G�H;��H;B�H;��H;�H;��H;B�H;��H;D�H;�H;�H;�H;�`H;�7H;aH;&�G;�8G;�F;ÚC;�0>;X�3;P ; ��:~�:`������*��H,�Y�V�1c���������G���}�t�����|�ؽ�s�[[�g9�      ��=�׀:���0��Q"�~������Pν�榽@����G�2����Ҽ ��JE:�@�ܻ�D^�ȸ��4i:7��:�;4|,;��:;J�A;<iE;��F;�G;{�G;�(H;/UH;xwH;m�H;�H;��H;�H;��H;��H;�H;��H;��H;�H;��H;�H;l�H;ywH;/UH;�(H;x�G;�G;��F;>iE;H�A;��:;,|,;�;1��:<i:ȸ���D^�@�ܻJE:� ����Ҽ2����G�@���榽�Pν����~��Q"���0�׀:�      1Dx�4�s���f�tS�׀:����Z[��7ս�榽��}���;��8�V�����r����>G�����ά���:�;�}$;��6;��?;�D;ƔF;�pG;��G;�H;JH;;oH;7�H;r�H;��H;4�H;��H;��H;"�H;��H;��H;4�H;��H;p�H;7�H;BoH; JH;�H;��G;�pG;��F;�D;��?;��6;�}$;	�;��: ά���?G�������r�V����8���;���}��榽�7սZ[����׀:�tS���f�4�s�      �*���0��ޥ��;����k��H��#%�Z[��Pνt��a�f�2/%���伆���w�=��?ػ�FL���D�H�R:��:-�;.2;��=;��C;b0F;@GG;��G;H;�?H;�gH;��H;&�H;��H;��H;z�H;��H;p�H;��H;~�H;��H;��H;'�H;��H;�gH;�?H;H;��G;GGG;_0F;��C;��=;,2;)�;��:@�R:��D��FL��?ػw�=��������3/%�a�f�t���PνZ[��#%��H��k�;���ޥ���0��      '�þ��� ����R��|쏾5�s��H�����������ΐ����D��c�����?�f�V,�����P�� �9ó�:�;j-;K�;;o�B;��E;TG;��G;��G;~6H;�`H;W�H;I�H;ЩH;K�H;��H;N�H;��H;O�H;��H;K�H;ЩH;I�H;T�H;�`H;�6H;��G;��G;]G;��E;p�B;H�;;j-;�;ǳ�:��9�P�����U,�>�f������c���D�ΐ�������������H�5�s�|쏾�R�� ������      A��/�待Yؾ(�þ
Ī�|쏾�k�׀:�~�{�ؽ�����c�]y���Ҽ����E� �m�4�� (7;�:��
;��(;{_9;��A;c\E;e�F;��G;��G;�.H;�ZH;�{H;�H;D�H;O�H;�H;��H;t�H;��H;	�H;L�H;D�H;�H;�{H;�ZH;�.H;��G;��G;o�F;a\E;��A;w_9;��(;��
;?�: (70��m�F� �������Ҽ]y��c�����{�ؽ~�׀:��k�|쏾
Ī�(�þ�Yؾ/��      #��O������=I�(�þ�R��;���tS��Q"��s������}��0��켉�����6�K�ƻ@}*�H�����:vx;T%;�l7;ճ@;��D;��F;��G;�G;�'H;�UH;[xH;H�H;@�H;��H;��H;��H;u�H;��H;��H;��H;B�H;J�H;ZxH;�UH;�'H;��G;��G;��F;��D;ճ@;�l7;R%;tx;��:X���<}*�J�ƻ��6��������0���}�����s��Q"�tS�;����R��(�þ=Iᾤ���O��      ���R��8�
������Yؾ ���ޥ����f���0�Z[�N8��ϐ���>�����KȤ��6H�f�ܻrF�����}:��:\";)�5;��?;O�D;��F;�G;��G;,#H;\RH;�uH;B�H;��H;q�H;��H;�H;��H;�H;��H;s�H;��H;B�H;�uH;dRH;/#H;��G;�G;��F;O�D;��?;$�5;[";��:�}:��rF�f�ܻ�6H�JȤ������>�ϐ��N8��Z[���0���f�ޥ�� ����Yؾ����8�
�R��      �� ����R��N��0������0��4�s�׀:�h9��ʽ2Z����G��8�.���5S����0X���D�RBd:�B�: ;��4;Ĉ?;�~D;�F;yG;��G;J H;&PH;tH; �H;ȢH;°H;(�H;k�H;2�H;k�H;)�H;ŰH;ȢH;�H;tH;0PH;M H;��G;yG;�F;�~D;��?;��4;� ;�B�:bBd:��D�0X���껰5S�.���8���G�2Z���ʽh9�׀:�4�s��0�����/��N��R�����      FEb�`]��N��7����s� ���˾��(�j��!,�p���L��Cm�,��9,˼��x�]���1�� ���8�:`�:�;�1;3,>;^�C;OwF;�G;j H;�>H;�hH;'�H;>�H;�H;�H;��H;�H;i�H;�H;��H;�H;�H;>�H;&�H;�hH;�>H;m H;�G;\wF;`�C;0,>;�1;�;b�:H�: ����1��]����x�8,˼,��Cm�L��p����!,�(�j�����˾s� �����7��N�`]�      `]�d�W��TI�v3��D�������Ǿv����f�8)�$��s;���Fi��k���Ǽ�[t�P�	�.Ȅ�.X����:���:��;(J2;OZ>; 	D;7F;4�G;�H;�?H;siH;��H;��H;M�H;�H;��H;3�H;��H;.�H;��H;�H;M�H;��H;��H;ziH;�?H;�H;6�G;DF;#	D;LZ>;"J2;��;���:Ƞ:*X��,Ȅ�O�	��[t���Ǽ�k��Fi�r;��%��8)��f�v�����Ǿ�����D�v3��TI�d�W�      �N��TI���;�/�'�l��쾀���y󐾴Z��K ��s�A����&^���"����g����بu�!���2<:��:�
;7g3;��>;QBD;s�F;ڔG;gH;BH;WkH;)�H;��H;�H;��H;<�H;��H;�H;��H;>�H;��H;�H;��H;'�H;`kH;BH;iH;ܔG;~�F;SBD;��>;1g3;�
;��:�2<:!��֨u������g��"����&^�A����s潥K ��Z�y󐾀�����l�/�'���;��TI�      �7�v3�/�'����s� ��{Ծ���H���y�F�����ӽ���_�L�Jv��뮼ST����PV���=�>)i:h��:�z ;{$5;��?;�D;��F;�G;oH;_FH;nnH;^�H;G�H;F�H;��H;�H;-�H;��H;(�H;�H;��H;F�H;G�H;[�H;unH;dFH;oH;�G;��F;�D;��?;v$5;�z ;h��:V)i:��=��PV���ST��뮼Jv�_�L�����ӽ���y�F�H�������{Ծs� ����/�'�v3�      ����D�l�s� �V�ݾk���V͓��f��>/�����'���섽P�6�t�w��`�:�+Tʻ�.�p۷�2t�:�;��$;�Y7;M�@;�	E;��F;&�G;�H;LH;�rH;��H;��H;��H;�H;�H; �H;��H;�H;�H;�H;��H;��H;��H;�rH;LH;�H;&�G;��F;�	E;I�@;~Y7;��$;�;>t�:p۷��.�*Tʻ`�:�w��t�P�6��섽�'������>/��f�V͓�k���V�ݾs� �l��D�      s� ��������{Ծk���v���Z�x��SC��^��޽@���x�e�(��D�Ѽ%G������R������ܤ8���:�Y;@�);��9;��A;��E;|G;	�G;<!H;SH;�wH;E�H;U�H;�H;��H;G�H;S�H;��H;O�H;H�H;��H;�H;V�H;D�H;�wH;SH;>!H;�G;�G;��E;��A;��9;@�);�Y;���:�ܤ8����R�����%G��D�Ѽ(��x�e�@����޽�^��SC�Z�x�v���k����{Ծ�쾠���      ��˾��Ǿ�������V͓�Z�x���J��K �m���������?����뮼+�[�!���3|��W��h�:3�:�';[/;<g<;C;@F;�NG;��G;-H;6[H;�}H;��H;��H;��H;|�H;��H;��H;��H;��H;��H;|�H;��H;��H;��H;�}H;:[H;-H;��G;�NG;AF;C;;g<;]/;�';;�:d�:�W��3|�"���+�[��뮼���?������m����K ���J�Z�x�V͓����������Ǿ      ��v���y�H����f��SC��K �nn�� �Ž����Z��k�}ռ.X��cy-�0���x.����P�:�+�:w�;	4;�>;�D;�wF;��G;��G;�9H;#dH;P�H;|�H;.�H;E�H;��H;{�H;(�H;B�H;'�H;~�H;��H;B�H;,�H;|�H;W�H;'dH;�9H;��G;��G;�wF;�D;�>;
4;t�;�+�:�P�:���u.�/���ay-�.X��}ռ�k��Z������Žnn���K ��SC��f�H���y�v���      (�j��f��Z�y�F��>/��^�m�����ŽF ���Fi��Q+�|t�oT��p�W�����1��<Ⱥ�W�9gP�:{Y;}�(;��8;�A;�E;��F;6�G;mH;�FH;�mH;e�H;��H;�H;D�H;��H;]�H;��H;��H;��H;^�H;��H;A�H;�H;��H;m�H;�mH;�FH;mH;4�G;��F;�E;�A;��8;{�(;�Y;kP�:�W�92Ⱥ�1�����o�W�nT��|t�Q+��Fi�F ����Žm����^��>/�y�F��Z��f�      �!,�8)��K ��������޽������Fi��0����鷼��x�����.��[�(� ���*i:f��: �;��0;2�<;mC;�E;�<G;��G;�$H;5TH;�wH;ÒH;�H;�H;U�H;�H;`�H;p�H;M�H;o�H;c�H;�H;S�H;�H;�H;˒H;�wH;8TH;�$H;��G;�<G;|�E;qC;6�<;��0;'�;p��:�*i:��Y�(��.�������x�鷼����0��Fi�������޽�������K �8)�      o���%��s��ӽ�'��@�������Z��Q+�����"��G��»0���׻ԕb�NW���X�9ġ�:`;x*';�Y7;�#@; �D;ۖF;�G;��G;8H;�aH;ɁH;0�H;w�H;D�H;i�H;u�H;T�H;"�H;
�H;#�H;W�H;v�H;g�H;C�H;y�H;9�H;ЁH;�aH;8H;��G;�G;ܖF;�D;�#@;�Y7;�*';`;ơ�:�X�9HW��ҕb���׻»0�G���"������Q+��Z����?����'���ӽ�s�$��      K��r;��@�������섽x�e��?��k�|t�鷼G���e7����Ȅ��0�@�t�
u�:�+�:f;f1;=�<;E�B;��E;�G;��G;/H;MJH;/oH;͋H;��H;�H;j�H;��H;��H;g�H;��H;��H;��H;g�H;��H;��H;i�H;�H;��H;ًH;2oH;NJH;-H;��G;�G;�E;K�B;>�<;q1;j;�+�:u�:��t�~0�Ȅ���껅e7�G��鷼{t��k��?�x�e��섽���A���r;��      Cm��Fi��&^�`�L�O�6�(����}ռoT����x���0�������!���ط��n`:p�:�;�*;�8;��@;�D;>�F;�}G;v�G;h1H;�[H;?|H;��H;��H;V�H;��H;��H;[�H;e�H;��H;B�H;��H;d�H;[�H;��H;��H;Z�H;��H;��H;C|H;�[H;e1H;|�G;�}G;D�F;�D;��@;!�8;�*;�;~�:�n`:�ط���
��������0���x�nT��}ռ��(��P�6�`�L��&^��Fi�      *���k��Kv�}t�E�Ѽ�뮼-X��p�W������׻Ȅ�%��`���4<:F��:�Y;�t%;�$5;�Z>;�`C;��E;*G;=�G;�H;�GH;AlH;ÈH;ϞH;��H;��H;k�H;��H;��H;H�H;C�H;��H;C�H;G�H;��H;��H;j�H;��H;��H;ٞH;ǈH;ClH;�GH;�H;>�G;*G;��E;�`C;�Z>;�$5;�t%;�Y;H��:�4<:8�� ��Ȅ���׻���n�W�-X���뮼D�Ѽt�Kv���k�      7,˼��Ǽ�"���뮼w��%G��*�[�`y-�����.��ҕb��0��ط��4<:�L�:�\;h�!;�J2;zg<;(0B;CE;�F; �G;��G;Z4H;r\H;�{H;z�H;t�H;,�H;��H;�H;g�H;!�H;#�H;��H;~�H;��H;"�H;#�H;e�H;�H;��H;2�H;y�H;��H;�{H;o\H;_4H;��G;$�G;�F;CE;10B;�g<;�J2;p�!;�\;�L�:�4<:�ط��0�Εb��.�����`y-�*�[�#G��w���뮼�"����Ǽ      ��x��[t���g�PT�`�:�������,����1��W�(�HW����t��n`:F��:�\;�z ;|�0;J;;�<A;�D;�wF;�cG;&�G;�!H;|MH;UoH;F�H;V�H;��H;b�H;6�H;��H;,�H;A�H;��H;j�H;��H;j�H;��H;A�H;)�H;��H;:�H;g�H;��H;Z�H;J�H;OoH;�MH;�!H;-�G;�cG;�wF;��D;�<A;G;;��0;�z ;�\;H��:�n`:��t�BW��V�(��1��+���������b�:�RT���g��[t�      Z��M�	������'Tʻ�R��3|�q.�4Ⱥ����X�9u�:z�:�Y;l�!;��0;͕:;��@;�BD;_2F;S8G;��G;�H;<@H;�cH;��H;E�H;�H;�H;�H;b�H;��H;��H;=�H;��H;��H;W�H;��H;�H;@�H;��H;��H;f�H;!�H;�H;�H;H�H;��H;�cH;?@H;�H;��G;W8G;e2F;�BD;��@;Е:;��0;p�!;�Y;~�:u�:�X�9���(Ⱥp.�3|��R��*Tʻ�����K�	�      �1��*Ȅ�ڨu��PV�w.�����W������W�9�*i:ơ�:�+�:
�;~t%;�J2;C;;��@;VD;�F;�G;Q�G;aH;S5H;RZH; xH;�H;��H;�H;�H;*�H;<�H;��H;��H;��H;�H;0�H;��H;.�H;�H;��H;��H;��H;@�H;0�H;�H;�H;��H;�H;xH;RZH;S5H;eH;U�G;G;�F;SD;��@;@;;�J2;|t%;�;�+�:ԡ�:�*i:X�9p��W�����s.��PV�Шu�*Ȅ�      򥥺FX��!����=��۷�@ޤ8��:�P�:oP�:p��:`;f;�*;�$5;~g<;�<A;�BD;�F;�G;Q�G;:�G;r-H;�RH;(qH;��H;��H;M�H;�H;�H;��H;��H;��H;%�H;��H;r�H;j�H;��H;g�H;p�H;��H;"�H;��H;��H;��H;�H;�H;N�H;��H;��H;-qH;�RH;w-H;=�G;U�G;�G;�F;�BD;�<A;g<;�$5;�*;f; `;p��:uP�:�P�:|�:�ݤ8h۷���=�!��FX��      �:��:�2<:�)i:.t�:���:I�:�+�:{Y;%�;�*';o1;�8;�Z>;10B;��D;c2F;G;S�G;��G;Q)H;WNH;FlH;�H;4�H;T�H;m�H;��H;W�H;��H;�H;��H;�H;/�H;��H;��H;��H;��H;��H;.�H;�H;��H;	�H;��H;X�H;�H;m�H;S�H;9�H;�H;ElH;ZNH;W)H;��G;V�G;G;c2F;��D;10B;�Z>;�8;o1;�*';$�;�Y;�+�:C�:ɇ�:4t�:.)i:�2<:��:      ��:���:���:R��:�;�Y;�';q�;y�(;��0;�Y7;9�<;�@;�`C;CE;�wF;S8G;[�G;=�G;P)H;�LH;�iH;�H;+�H;u�H;��H;��H;4�H;��H;��H;��H;,�H;��H;o�H;��H;}�H;��H;v�H;��H;n�H;��H;(�H;��H;��H;��H;7�H;��H;��H;z�H;+�H;�H;�iH;�LH;Q)H;=�G;W�G;T8G;�wF;CE;�`C;�@;9�<;�Y7;��0;v�(;n�;�';�Y;�;R��:���:���:      �;��;;�z ;��$;>�);Y/;4;��8;6�<;�#@;D�B;�D;��E;
�F;�cG;��G;gH;w-H;ZNH;�iH;�H;��H;��H;��H;��H;v�H;s�H;�H;��H;G�H;�H;�H;��H;��H;F�H;��H;@�H;��H;��H;�H;�H;J�H;��H;�H;v�H;t�H;��H;��H;��H;��H;�H;�iH;ZNH;v-H;dH;��G;�cG;
�F;��E;�D;D�B;�#@;2�<;��8;4;[/;:�);��$;�z ;�
;��;      #�1;$J2;-g3;�$5;yY7;��9;Kg<;�>;�A;rC;�D;�E;D�F;*G;$�G;.�G;�H;[5H;�RH;ClH;�H;��H;��H;��H;\�H;<�H;0�H;�H;��H;�H;`�H;��H;]�H;��H;��H;�H;I�H;��H;��H;��H;Z�H;��H;b�H;�H;��H;�H;/�H;<�H;^�H;��H;��H;��H;	�H;ClH;�RH;S5H;�H;*�G;#�G;*G;A�F;�E;	�D;kC;�A;�>;Dg<;��9;�Y7;�$5;*g3;
J2;      0,>;VZ>;��>;��?;B�@;��A;�C;�D;�E;��E;ݖF;�G;�}G;A�G;��G;�!H;?@H;YZH;-qH;�H;+�H;}�H;��H;�H;��H;��H;�H;��H;��H;��H;:�H;�H;�H;x�H;>�H;��H;��H;��H;;�H;x�H;~�H;�H;<�H;��H;��H;��H;�H;��H;��H;�H;��H;��H;+�H;�H;'qH;RZH;>@H;�!H;��G;:�G;�}G;�G;ݖF;~�E;�E;�D;}C;��A;K�@;��?;��>;MZ>;      �C;	D;JBD;ښD;�	E;��E;KF;�wF;��F;�<G;�G;��G;z�G;�H;a4H;�MH;�cH;xH;��H;@�H;�H;��H;a�H;��H;!�H;��H;��H;M�H;V�H;��H;��H;X�H;x�H;0�H;��H;<�H;>�H;7�H;��H;2�H;t�H;S�H;��H;��H;R�H;M�H;��H;��H;"�H;��H;^�H;��H;�H;<�H;��H;xH;�cH;�MH;_4H;�H;z�G;��G;�G;�<G;��F;�wF;JF;��E;�	E;ښD;IBD;	D;      DwF;;F;u�F;��F;��F;�G;�NG;�G;5�G;��G;��G;2H;i1H;�GH;p\H;YoH;��H;�H;��H;S�H;��H;��H;;�H;��H;��H;>�H;�H;�H;��H;y�H;�H;G�H;(�H;��H;e�H;��H;��H;��H;b�H;��H;&�H;C�H;�H;x�H;��H;�H;�H;B�H;��H;��H;8�H;��H;��H;P�H;��H;�H;��H;SoH;o\H;�GH;g1H;0H;��G;��G;5�G;�G;�NG;vG;��F;��F;s�F;>F;      ��G;:�G;ԔG;�G;�G;�G;��G;��G;iH;�$H;8H;JJH;�[H;ClH;�{H;K�H;N�H; �H;S�H;p�H;��H;v�H;3�H;"�H;��H;�H;��H;W�H;>�H;��H;'�H;�H;��H;}�H;��H;��H;	�H;��H;��H;}�H;��H;�H;'�H;��H;;�H;U�H;��H;�H;��H;�H;2�H;w�H;��H;m�H;P�H;��H;I�H;H�H;�{H;<lH;�[H;JJH;8H;�$H;hH;��G;��G;��G;0�G;ݣG;ՔG;%�G;      k H;�H;aH;uH;�H;<!H;-H;�9H;�FH;>TH;�aH;6oH;A|H;ɈH;y�H;Z�H;�H;�H;�H; �H;9�H;s�H;�H;��H;I�H;	�H;U�H;N�H;��H;��H;��H;��H;o�H;��H;�H;W�H;[�H;S�H;�H;��H;l�H;��H;��H;��H;��H;K�H;Q�H;�H;M�H;��H;�H;s�H;6�H;��H;�H;�H;�H;Y�H;z�H;ǈH;?|H;3oH;�aH;:TH;�FH;�9H;-H;/!H;�H;rH;aH;�H;      �>H;x?H;BH;pFH;�KH;SH;=[H;dH;�mH;�wH;΁H;ԋH;��H;՞H;v�H;��H;�H;�H;�H;Z�H;��H;�H;��H;��H;P�H;~�H;7�H;��H;�H;��H;��H;d�H;��H;.�H;h�H;��H;��H;��H;f�H;/�H;��H;^�H;��H;��H;�H;��H;3�H;�H;S�H;��H;��H;�H;��H;U�H;�H;�H;�H;��H;u�H;ӞH;��H;ӋH;ЁH;�wH;�mH; dH;9[H;SH;LH;lFH;BH;y?H;      �hH;fiH;ckH;jnH;�rH;�wH;�}H;P�H;h�H;ȒH;6�H;��H;��H;��H;,�H;d�H;"�H;-�H;��H;��H;��H;��H;{�H;��H;��H;o�H;��H;��H;��H;��H;h�H;��H;�H;t�H;��H;��H;��H;��H;��H;t�H;�H;��H;h�H;��H;��H;��H;��H;u�H;��H;��H;}�H;��H;��H;��H;��H;,�H;"�H;d�H;.�H;��H;��H;��H;7�H;˒H;h�H;S�H;�}H;�wH;�rH;mnH;ckH;iiH;      .�H;шH;0�H;a�H;��H;H�H;��H;��H;��H;�H;}�H;�H;^�H;��H;��H;=�H;k�H;D�H;��H;�H;��H;J�H;`�H;<�H;��H;�H;'�H;��H;��H;n�H;��H;(�H;�H;��H;��H;��H;��H;��H;��H;��H;��H;&�H;��H;n�H;��H;��H;"�H;�H;��H;9�H;b�H;J�H;��H;�H;��H;C�H;m�H;?�H;��H;��H;`�H;�H;}�H;�H;��H;��H;��H;=�H;��H;a�H;2�H;ӈH;      G�H;��H;��H;G�H;��H;N�H;��H;/�H;�H;�H;H�H;n�H;��H;t�H;�H;��H;��H;��H;��H;�H;2�H;�H;��H;�H;U�H;@�H; �H;��H;`�H;��H; �H;v�H;��H;��H;��H;��H;�H;��H;��H;��H;��H;t�H; �H;��H;[�H;��H;��H;D�H;X�H;�H;��H;�H;,�H;��H;��H;��H;��H;��H;�H;q�H;��H;p�H;M�H;�H;�H;0�H;��H;N�H;��H;G�H;��H;��H;      �H;Z�H;�H;J�H;�H;�H;��H;A�H;?�H;W�H;l�H;��H;��H;��H;h�H;0�H;��H;�H;)�H;�H;��H;�H;[�H;}�H;w�H;#�H;��H;r�H;��H;�H;{�H;��H;��H;��H;�H;�H;��H;�H;�H;��H;��H;��H;{�H;�H;��H;l�H;��H;&�H;z�H;}�H;^�H;�H;��H;�H;)�H;�H;��H;3�H;i�H;��H;��H;��H;o�H;W�H;A�H;A�H;��H;�H;�H;C�H;�H;[�H;      �H;
�H;��H;��H;��H;��H;��H;��H;��H;�H;��H;��H;e�H;��H;'�H;G�H;D�H; �H;��H;3�H;u�H;��H;��H;p�H;/�H;��H;w�H;��H;-�H;v�H;��H;��H;��H;��H;%�H;/�H;�H;/�H;%�H;��H;��H;��H;��H;t�H;(�H;��H;v�H;��H;2�H;n�H;��H;��H;o�H;,�H;��H;�H;I�H;H�H;(�H;��H;b�H;��H;��H;�H;��H;��H;��H;��H;��H;��H;��H;�H;      ��H;��H;L�H;�H;�H;B�H;��H;~�H;a�H;j�H;`�H;q�H;r�H;Q�H;*�H;��H;��H;�H;q�H;��H;��H;��H;|�H;2�H;��H;[�H;��H;�H;h�H;��H;��H;��H;�H;'�H;	�H;$�H;A�H;%�H;	�H;)�H;�H;��H;��H;��H;c�H;	�H;��H;`�H;��H;2�H;��H;��H;��H;��H;q�H;�H;��H;��H;)�H;O�H;p�H;q�H;a�H;k�H;e�H;��H;��H;B�H;�H;�H;M�H;��H;      �H;0�H;��H;.�H;�H;K�H;��H;,�H;��H;w�H;*�H;��H;��H;H�H;��H;j�H;��H;.�H;h�H;��H;�H;A�H;��H;��H;7�H;��H;��H;W�H;��H;��H;��H;��H;�H;0�H;'�H;�H;.�H;�H;%�H;6�H;�H;��H;��H;��H;��H;S�H;��H;��H;5�H;��H;�H;A�H;z�H;~�H;g�H;2�H;��H;m�H;��H;I�H;��H;��H;,�H;x�H;��H;,�H;��H;L�H;!�H;+�H;��H;?�H;      q�H;��H;9�H;��H;��H;��H;��H;G�H;��H;O�H;�H;��H;N�H;	�H;��H;��H;_�H;��H;��H;��H;��H;��H;I�H;��H;A�H;��H;�H;a�H;��H;��H;��H;�H;��H;�H;C�H;+�H;�H;.�H;C�H;�H;�H;�H;��H;��H;��H;\�H;�H;��H;>�H;��H;N�H;��H;��H;��H;��H;��H;_�H;��H;��H;	�H;L�H;��H;�H;Q�H;��H;G�H;��H;��H;��H;��H;:�H;��H;      �H;5�H;��H;.�H; �H;P�H;��H;+�H;��H;w�H;)�H;��H;��H;J�H;��H;j�H;��H;.�H;h�H;��H;��H;C�H;��H;��H;7�H;��H;��H;W�H;��H;��H;��H;��H;�H;2�H;)�H;�H;.�H;�H;%�H;5�H;�H;��H;��H;��H;��H;Q�H;��H;��H;5�H;��H;�H;?�H;z�H;��H;g�H;2�H;��H;k�H;��H;H�H;��H;��H;,�H;t�H;��H;.�H;��H;L�H;$�H;/�H;��H;<�H;      ��H;��H;E�H;�H;�H;>�H;��H;��H;d�H;k�H;`�H;q�H;p�H;Q�H;,�H;��H;��H;�H;q�H;��H;��H;��H;|�H;0�H;��H;Z�H;��H;�H;h�H;��H;��H;��H;�H;'�H;�H;%�H;D�H;(�H;�H;)�H;�H;��H;��H;��H;c�H;�H;��H;`�H;��H;0�H;��H;��H;��H;��H;p�H;�H;��H;��H;'�H;O�H;p�H;r�H;^�H;j�H;b�H;��H;��H;;�H;�H;	�H;L�H;��H;      �H;�H;��H;��H;��H;��H;��H;��H;��H;�H;��H;��H;d�H;��H;*�H;G�H;G�H;�H;��H;2�H;u�H;��H;��H;q�H;2�H;��H;y�H;��H;.�H;w�H;��H;��H;��H;��H;(�H;.�H;�H;/�H;%�H;��H;��H;��H;��H;q�H;&�H;��H;w�H;��H;/�H;m�H;��H;��H;k�H;/�H;��H; �H;G�H;H�H;(�H;��H;b�H;��H;��H;�H;��H;��H;��H;��H; �H;��H;��H;
�H;      �H;a�H;�H;F�H;��H;�H;��H;E�H;@�H;W�H;n�H;��H;��H;��H;l�H;2�H;��H;�H;)�H;�H;��H;�H;X�H;}�H;z�H;�H;��H;r�H;��H;�H;{�H;��H;��H;��H;�H;�H;��H;�H;�H;��H;��H;��H;z�H;�H;��H;l�H;��H;&�H;x�H;{�H;a�H;�H;��H;�H;(�H;�H;��H;2�H;i�H;��H;��H;��H;n�H;T�H;A�H;E�H;��H;�H;�H;K�H;�H;Z�H;      6�H;��H;��H;@�H;��H;]�H;��H;3�H;�H;�H;H�H;p�H;��H;r�H;�H;��H;��H;��H;��H;�H;3�H;�H;��H;
�H;X�H;?�H;��H;��H;d�H;��H; �H;v�H;��H;��H;��H;��H;�H;��H;��H;��H;��H;t�H;�H;��H;[�H;��H;��H;D�H;W�H;�H;��H;�H;,�H;��H;��H;��H;��H;��H;�H;q�H;��H;p�H;J�H;�H;�H;2�H;��H;P�H;��H;C�H;��H;��H;      "�H;шH;0�H;[�H;��H;G�H;��H;~�H;��H;�H;~�H;�H;^�H;��H;��H;?�H;m�H;D�H;��H;�H;��H;K�H;^�H;:�H;��H;�H;"�H;��H;��H;n�H;��H;(�H;��H;��H;��H;��H;��H;��H;��H;��H;��H;'�H;��H;i�H;��H;��H;"�H;	�H;��H;7�H;e�H;K�H;��H;�H;��H;C�H;n�H;=�H;��H;��H;^�H;�H;}�H;�H;��H;��H;��H;B�H;��H;h�H;7�H;шH;      �hH;piH;^kH;wnH;�rH;�wH;�}H;X�H;m�H;˒H;6�H;��H;��H;��H;0�H;e�H;"�H;/�H;��H;��H;��H;��H;x�H;��H;��H;n�H;��H;��H;��H;��H;i�H;��H;�H;t�H;��H;��H;��H;��H;��H;t�H;�H;��H;g�H;��H;��H;��H;��H;t�H;��H;��H;��H;��H;��H;��H;��H;,�H;"�H;g�H;0�H;��H;��H;��H;7�H;˒H;j�H;W�H;�}H;�wH;�rH;znH;okH;iiH;      �>H;x?H; BH;lFH;�KH;SH;9[H;"dH;�mH;�wH;΁H;ԋH;��H;՞H;y�H;��H;�H;�H;�H;W�H;��H;�H;��H;��H;R�H;x�H;4�H;��H;�H;��H;��H;d�H;��H;.�H;h�H;��H;��H;��H;f�H;.�H;��H;a�H;��H;��H;�H;��H;4�H;�H;R�H;��H;��H;�H;��H;Z�H;�H;�H;�H;��H;y�H;֞H;��H;ӋH;ЁH;�wH;�mH;%dH;>[H;SH;�KH;kFH;BH;q?H;      u H;�H;WH;uH;|H;G!H;-H;�9H;�FH;<TH;�aH;4oH;A|H;ʈH;|�H;Y�H;�H;�H;�H;��H;9�H;u�H;�H;��H;L�H;�H;S�H;L�H;��H;��H;��H;��H;l�H;��H;�H;T�H;\�H;U�H;�H;��H;o�H;��H;��H;��H;��H;H�H;S�H;
�H;I�H;��H;	�H;s�H;6�H; �H;�H;�H;�H;Z�H;~�H;ʈH;A|H;4oH;�aH;;TH;�FH;�9H;-H;6!H;�H;uH;bH;�H;      �G;?�G;הG;�G;)�G;�G;��G;��G;iH;�$H;8H;MJH;�[H;AlH;�{H;J�H;I�H;�H;P�H;m�H;��H;w�H;-�H;"�H;��H;�H;��H;W�H;@�H;��H;%�H;�H;��H;}�H;��H;��H;	�H;��H;��H;~�H;��H;�H;'�H;��H;:�H;T�H;��H;�H;��H;�H;6�H;w�H;��H;p�H;Q�H;��H;K�H;K�H;�{H;AlH;�[H;KJH;8H;�$H;iH;��G;��G;�G;1�G;�G;۔G;0�G;      ;wF;;F;�F;��F;��F;�G;�NG;	�G;9�G;��G;��G;3H;i1H;�GH;r\H;VoH;��H;�H;��H;Q�H;��H;��H;7�H;��H;��H;;�H;�H;�H;��H;u�H;�H;G�H;&�H;��H;e�H;��H;��H;��H;b�H;��H;(�H;G�H;	�H;u�H;�H;
�H;
�H;A�H;��H;��H;<�H;��H;��H;S�H;��H;�H;��H;WoH;u\H;�GH;i1H;2H;��G;��G;2�G;�G;�NG;{G;��F;��F;g�F;,F;      ~�C;	D;IBD;ߚD;�	E;��E;KF;�wF;��F;�<G;�G;��G;y�G;�H;b4H;�MH;�cH;xH;��H;=�H;�H;��H;]�H;��H;"�H;��H;��H;M�H;V�H;��H;��H;X�H;u�H;2�H;��H;:�H;?�H;:�H;��H;3�H;x�H;X�H;��H;��H;P�H;H�H;��H;��H;!�H;��H;c�H;��H;�H;<�H;��H;
xH;�cH;�MH;e4H;�H;|�G;��G;�G;�<G;��F;�wF;MF;��E;�	E;ܚD;JBD;	D;      ,>;<Z>;��>;��?;=�@;��A;�C;�D;�E;�E;ߖF;�G;�}G;>�G;��G;�!H;<@H;XZH;(qH;�H;,�H;~�H;��H;�H;��H;��H;�H;��H;��H;��H;<�H;�H;�H;z�H;=�H;��H;��H;��H;;�H;x�H;��H;�H;?�H;��H;��H;��H;�H;��H;��H;�H;��H;}�H;+�H;�H;+qH;UZH;?@H;�!H;��G;@�G;�}G;�G;��F;�E;�E;�D;�C;��A;T�@;��?;��>;'Z>;      �1;J2;!g3;�$5;wY7;��9;Cg<;�>;�A;oC;�D;�E;A�F;*G;'�G;.�G;�H;X5H;�RH;ElH;�H;��H;��H;��H;^�H;5�H;,�H;	�H;��H;{�H;a�H;��H;[�H;��H;��H;�H;L�H;�H;��H;��H;^�H;��H;e�H;�H;��H;�H;0�H;:�H;Z�H;��H;��H;��H;�H;ElH;�RH;T5H;�H;-�G;(�G;*G;D�F;�E;�D;qC;�A;�>;Dg<;��9;wY7;�$5;!g3;J2;      �;��;�
;�z ;��$;E�);^/;
4;��8;4�<;�#@;I�B;�D;��E;�F;�cG;��G;gH;t-H;ZNH;�iH;�H;��H;��H;��H;��H;s�H;v�H;�H;��H;H�H;�H;�H;��H;��H;A�H;��H;D�H;��H;��H;�H;�H;K�H;��H;�H;s�H;v�H;��H;��H;��H;��H;�H;�iH;\NH;v-H;eH;��G;�cG;�F;��E;�D;G�B;�#@;4�<;��8;4;W/;/�);��$;�z ;�
;��;      ��:��:���:`��:�;�Y;�';t�;~�(;��0;�Y7;;�<;��@;�`C;CE;�wF;T8G;Z�G;<�G;Q)H;�LH;�iH;�H;,�H;z�H;��H;��H;6�H;��H;��H;��H;-�H;��H;o�H;��H;x�H;��H;z�H;��H;k�H;��H;,�H;��H;��H;��H;4�H;��H;��H;u�H;,�H;�H;�iH;�LH;T)H;>�G;X�G;T8G;�wF;CE;�`C;��@;7�<;�Y7;��0;{�(;w�;�';�Y;�;`��:��:���:      ��:��:�2<:~)i:2t�:ɇ�:O�:�+�:�Y;%�;�*';o1;�8;�Z>;40B;��D;c2F;G;S�G;��G;W)H;\NH;FlH;�H;9�H;Q�H;i�H;�H;Z�H;��H;�H;��H;�H;0�H;��H;��H;��H;��H;��H;,�H;�H;��H;�H;��H;W�H;��H;m�H;S�H;5�H; �H;FlH;YNH;U)H;��G;S�G;G;c2F;��D;30B;�Z>;�8;m1;�*';$�;�Y;�+�:C�:���::t�:N)i:�2<:��:      �DX��!����=��۷�`ޤ8��:�P�:uP�:p��: `;h;�*;�$5;�g<;�<A;�BD;�F;�G;S�G;=�G;w-H;�RH;*qH;��H;��H;L�H;�H;�H;��H;��H;��H;%�H;��H;r�H;h�H;��H;h�H;p�H;��H;%�H;��H;��H;��H;�H;�H;M�H;��H;��H;-qH;�RH;t-H;=�G;U�G;�G;�F;�BD;�<A;�g<;�$5;�*;d;`;p��:qP�:�P�:��: ޤ8�۷���=�!��<X��      �1��%Ȅ�ܨu��PV�p.�����W��H�� X�9�*i:Ρ�:�+�:�;�t%;�J2;F;;��@;UD;�F; G;U�G;eH;W5H;UZH;xH;�H;��H;�H;�H;)�H;?�H;��H; �H;��H;�H;0�H;��H;2�H;�H;��H;��H;��H;@�H;/�H;�H;�H;��H;�H; xH;TZH;U5H;cH;Q�G;G;�F;SD;��@;C;;�J2;|t%;
�;�+�:Ρ�:�*i:X�9`��W�����q.��PV��u�'Ȅ�      Z��N�	������&Tʻ�R��3|�n.�.Ⱥ����X�9u�:|�:�Y;r�!;��0;ѕ:;��@;�BD;b2F;W8G;��G;�H;@@H;�cH;��H;E�H;�H;�H;�H;d�H;��H;��H;B�H;��H;��H;Z�H;��H;��H;=�H;��H;��H;f�H; �H;�H;�H;E�H;��H;�cH;>@H;�H;��G;Q8G;e2F;�BD;��@;Ε:;��0;p�!;�Y;|�:u�:�X�9 ��,Ⱥo.�3|��R��+Tʻ�����L�	�      ��x��[t���g�QT�`�:�������*����1��V�(�>W��@�t��n`:H��:�\;�z ;�0;H;;�<A;��D;�wF;�cG;.�G;�!H;�MH;VoH;F�H;V�H;��H;b�H;9�H;��H;,�H;D�H;��H;j�H;��H;h�H;��H;@�H;)�H;��H;9�H;b�H;��H;V�H;D�H;RoH;}MH;�!H;+�G;�cG;�wF;��D;�<A;D;;}�0;�z ;�\;D��:�n`:��t�DW��W�(��1��+��� ������c�:�QT���g��[t�      7,˼��Ǽ�"���뮼w��$G��*�[�_y-�����.��Εb��0��ط��4<:�L�:�\;n�!;�J2;~g<;-0B;CE;
�F;(�G;��G;_4H;s\H;�{H;}�H;x�H;.�H;��H;�H;g�H;$�H;#�H;��H;~�H;��H;"�H;#�H;e�H;�H;��H;.�H;y�H;z�H;�{H;p\H;[4H;��G;%�G;
�F;CE;/0B;zg<;�J2;l�!;�\;�L�:�4<:�ط��0�Еb��.�����`y-�*�[�$G��w���뮼�"����Ǽ      *���k��Jv�}t�D�Ѽ�뮼-X��n�W������׻Ȅ���8���4<:R��:�Y;�t%;�$5;�Z>;�`C;��E;*G;B�G;�H;�GH;AlH;ƈH;՞H;��H;��H;k�H;��H;��H;G�H;B�H;��H;E�H;F�H;��H;��H;i�H;��H;��H;֞H;ňH;>lH;�GH;�H;A�G;*G;��E;�`C;�Z>;�$5;~t%;�Y;D��:�4<:X��"��Ȅ���׻���o�W�,X���뮼D�Ѽt�Jv���k�      Cm��Fi��&^�`�L�O�6�(����}ռnT����x���0����
������ط��n`:z�:�;�*;�8;��@;�D;E�F;�}G;|�G;i1H;�[H;A|H;��H;��H;Y�H;��H;��H;^�H;e�H;��H;B�H;��H;d�H;[�H;��H;��H;W�H;��H;��H;?|H;�[H;g1H;v�G;�}G;B�F;�D;�@;�8;�*;�;z�:�n`:�ط� ����������0���x�nT��}ռ��(��P�6�`�L��&^��Fi�      K��r;��@�������섽x�e��?��k�|t�鷼G���e7����Ȅ�z0�@�t�u�:�+�:f;m1;B�<;H�B;�E;�G;��G;0H;KJH;0oH;ӋH;��H;�H;i�H;��H;��H;f�H;��H;��H;��H;f�H;��H;��H;g�H;�H;��H;֋H;0oH;IJH;-H;��G;�G;�E;E�B;:�<;o1;d;�+�:u�:@�t��0�Ȅ���껆e7�G��鷼|t��k��?�x�e��섽���A���r;��      o���%��s��ӽ�'��@�������Z��Q+�����"��G����0���׻Еb�HW���X�9���:`;|*';�Y7;�#@;�D;ݖF;�G;��G;8H;�aH;́H;3�H;z�H;F�H;i�H;x�H;T�H;#�H;�H;#�H;V�H;v�H;g�H;C�H;w�H;6�H;΁H;�aH;8H;��G;�G;ܖF;�D;�#@;�Y7;~*';`;���:�X�9LW��ӕb���׻»0�G���"������Q+��Z����?����'���ӽ�s�%��      �!,�8)��K ��������޽������Fi��0����鷼��x�����.��W�(����*i:l��:"�;��0;4�<;qC;��E;�<G;��G;�$H;5TH;�wH;ǒH;�H;�H;U�H;�H;`�H;o�H;M�H;o�H;b�H;�H;S�H;�H;�H;ȒH;�wH;7TH;�$H;��G;�<G;�E;oC;2�<;��0;%�;d��:�*i:��Z�(��.�������x�鷼����0��Fi�������޽�������K �8)�      (�j��f��Z�y�F��>/��^�m�����ŽF ���Fi��Q+�|t�nT��p�W�����1��8Ⱥ�W�9kP�:�Y;~�(;��8;�A;�E;��F;4�G;lH;�FH;�mH;j�H;��H;�H;F�H;��H;[�H;��H;��H;��H;]�H;��H;A�H;�H;��H;j�H;�mH;�FH;kH;6�G;��F;�E;�A;��8;y�(;�Y;cP�:�W�98Ⱥ�1�����p�W�nT��|t�Q+��Fi�F ����Žm����^��>/�y�F��Z��f�      ��v���y�H����f��SC��K �nn����Ž����Z��k�}ռ.X��by-�/���u.����P�:�+�:{�;
4;�>;�D;�wF;��G;��G;�9H;"dH;P�H;}�H;/�H;E�H;��H;{�H;(�H;B�H;'�H;|�H;��H;B�H;,�H;}�H;V�H;'dH;�9H;��G; �G;�wF;�D;�>;	4;t�;�+�:�P�:���t.�0���by-�.X��}ռ�k��Z������Žnn���K ��SC��f�H���y�v���      ��˾��Ǿ�������V͓�Z�x���J��K �m���������?����뮼+�[�!���3|��W��d�:5�:�';[/;=g<;�C;AF;�NG;��G;-H;7[H;�}H;��H;��H;��H;~�H;��H;��H;��H;��H;��H;|�H;��H;��H;��H;�}H;;[H;-H;��G;�NG;?F;�C;<g<;Z/;�';=�:\�:�W��3|�"���+�[��뮼���?������m����K ���J�Z�x�V͓����������Ǿ      s� ��������{Ծk���v���Z�x��SC��^��޽@���x�e�(��D�Ѽ%G������R������ܤ8���:�Y;>�);��9;��A;��E;{G;�G;<!H;SH;�wH;I�H;W�H;�H;��H;G�H;S�H;��H;S�H;H�H;��H;�H;W�H;E�H;�wH;	SH;@!H;�G;�G;��E;��A;��9;>�);�Y;Ç�:�ܤ8����R�����%G��D�Ѽ(��x�e�@����޽�^��SC�Z�x�v���k����{Ծ�쾠���      ����D�l�s� �V�ݾk���V͓��f��>/�����'���섽O�6�t�w��`�:�*Tʻ�.�p۷�8t�:�;��$;�Y7;O�@;�	E;��F;#�G;�H;LH;�rH;��H;��H;��H;��H;��H;"�H;��H;�H;�H;�H;��H;��H;��H;�rH;LH;�H;)�G;��F;�	E;M�@;~Y7;��$;�;<t�:x۷�.�*Tʻ`�:�w���t�P�6��섽�'������>/��f�V͓�k���V�ݾs� �l��D�      �7�v3�/�'����s� ��{Ծ���H���y�F�����ӽ���_�L�Jv��뮼ST����PV���=�J)i:l��:�z ;{$5;��?;�D;��F;�G;nH;_FH;mnH;a�H;G�H;D�H;��H;�H;-�H;��H;*�H;�H;��H;G�H;J�H;]�H;wnH;dFH;pH;�G;��F;�D;��?;v$5;�z ;h��:^)i:��=��PV���RT��뮼Jv�_�L�����ӽ���y�F�H�������{Ծs� ����/�'�v3�      �N��TI���;�/�'�l��쾀���y󐾴Z��K ��s�A����&^���"����g����بu�!���2<:��:�
;5g3;��>;QBD;p�F;ؔG;gH;BH;WkH;+�H;��H;�H;��H;;�H;��H;�H;��H;>�H;��H;�H;��H;'�H;`kH;BH;kH;ޔG;~�F;SBD;��>;.g3;�
;��:�2<:!��Ԩu������g��"����&^�A����s潥K ��Z�y󐾀�����l�/�'���;��TI�      `]�d�W��TI�v3��D�������Ǿv����f�8)�%��r;���Fi��k���Ǽ�[t�P�	�.Ȅ�,X����:���:��;(J2;OZ>; 	D;6F;4�G;�H;�?H;siH;��H;��H;M�H;�H;��H;1�H;��H;.�H;��H;�H;M�H;��H;��H;ziH;�?H;�H;7�G;EF;!	D;MZ>; J2;��;���:̠:.X��,Ȅ�O�	��[t���Ǽ�k��Fi�s;��%��8)��f�v�����Ǿ�����D�v3��TI�d�W�      �?��}h��=v��� ��6�X��O/�0y�A�;ఖ��+X����ѽ����_n;�[�������B(�ݚ��d���e9�:�;�Y.;O�<;_WC;�ZF;�G;�/H;/jH;5�H;C�H;}�H;$�H;��H;T�H;��H;��H;��H;S�H;��H;"�H;}�H;A�H;<�H;1jH;�/H;��G;�ZF;aWC;M�<;�Y.;�;�:`�e9f��ܚ���B(�����[��_n;������ѽ���+X�ఖ�A�;0y��O/�6�X�� ��=v��}h��      |h��/���b�����y�VvS�pM+��v�9ɾ�����T� ]�\ν����y\8�����x��%�Q������0�9b-�:c�;��.;�<;�nC;�dF;�G;�1H;�jH;��H;��H;ƵH;d�H;��H;`�H;��H;��H;��H;a�H;��H;c�H;ƵH;��H;��H;�jH;�1H;�G;�dF;�nC;�<;��.;a�;f-�:X�9���O���%��x�����y\8�����\ν ]��T�����9ɾ�v�pM+�VvS���y�b���/���      =v��b���W ��a�h�6E�X��j���|㼾}���nH�ӈ�y�ý�Ȅ��s/��o��#�����'J��6к(	�9Ig�:�l; 0;]=;ղC;ӀF;k�G;6H;mH;$�H;��H;z�H;��H;=�H;��H;�H;��H;��H;��H;:�H;��H;z�H;��H;)�H;mH;6H;m�G;��F;زC;]=;0;�l;Mg�:X	�9:к&J������#���o��s/��Ȅ�y�ýӈ��nH�}��|㼾j���W��6E�a�h�W ��b���      � ����y�a�h��N��O/����B�߾B���*|��6�p}�䳽jSt�<�!�prμCF{��_��X��ړ��4: ��:�Z;�2;�O>;iD;&�F;v�G;=H;�pH;��H;E�H;ƷH;��H;��H;X�H;w�H;Z�H;s�H;X�H;��H;��H;ƷH;A�H;��H;�pH;=H;v�G;/�F;jD;�O>;�2;�Z;"��:P:ړ���X���_�CF{�orμ<�!�jSt�䳽p}��6��*|�B��B�߾����O/���N�a�h���y�      6�X�VvS�6E��O/��S�HW����������LS\��� ���:����Y�{��Ѓ����]�����)�b���Y�0�Y:��:^`;5�4;�?;5�D;��F;�G; FH;CuH;��H;��H;~�H;�H;��H;�H;�H;��H;�H;�H;��H;�H;}�H;��H;ēH;CuH;FH;	�G;��F;8�D;�?;1�4;``;��:@�Y:��Y�'�b�������]�Ѓ��{���Y�9����彑� �LS\���������HW���S��O/�6E�VvS�      �O/�pM+�X�����HW��9ɾ@���Mw�� :�i��w�ý�L��\n;�^���tv���E<��˻��-�X��`y�:�^;�%;}�7;r�@;5E;�"G;�G;3PH;�zH;��H;V�H;u�H;��H;��H;�H;��H;��H;��H;�H;��H;��H;u�H;Q�H;��H;�zH;6PH;�G;�"G;5E;o�@;|�7;�%;�^;dy�:P����-��˻�E<�sv��^���\n;��L��w�ýi��� :��Mw�@��9ɾHW�����X��pM+�      0y��v�j���B�߾����@��?����nH���CὝu����d�0O�jrμJ"�����	������q89S;�:Z�;�+;Q|:;u7B;��E;�aG;mH;�ZH;_�H;'�H;��H;�H;C�H;@�H; �H;��H;q�H;��H;�H;@�H;B�H;�H;��H;-�H;c�H;�ZH;iH;�aG;��E;t7B;N|:;�+;Z�;[;�: r89���	�����J"��irμ0O���d��u��C����nH�?���@������B�߾j����v�      @�;9ɾ{㼾B�������Mw��nH�����Z�䳽ʕ��r\8�o#������^N�P���b�Ix� 5:ծ�:*�;��0;]=;<�C;�[F;ҞG;�)H;�eH;n�H;�H;9�H;~�H;�H;��H;$�H;��H;i�H;��H;(�H;��H;�H;}�H;7�H;&�H;p�H;�eH;�)H;՞G;�[F;8�C;]=;��0;)�;��:(5:Ix��b�O��^N�����n#��q\8�ʕ��䳽�Z񽰯��nH��Mw�����B��{㼾9ɾ      ఖ�����}���*|�LS\�� :����Z�l$�������K�v���Oļ����������F&�p��5/�:�^;��#;�G6;7�?;��D;D�F;��G;�?H;�pH;ڏH;q�H;�H;G�H;,�H;g�H;k�H;��H;v�H;��H;n�H;i�H;)�H;H�H;�H;t�H;ۏH;�pH;�?H;��G;E�F;��D;;�?;�G6;��#;�^;;/�:P��B&������������Oļv���K�����k$���Z���� :�LS\��*|�}������      �+X��T��nH��6��� �i��C�䳽�����mR����ټ�����E<��?ݻ<d\������ :�d�:��;"�,;s�:;V7B;��E;kLG;+H;VSH;�{H;y�H;�H;�H;9�H;O�H;�H;��H;��H;��H;��H;��H;�H;N�H;7�H;�H;�H;}�H;�{H;USH;)H;nLG;��E;Y7B;v�:;"�,;��;�d�:� :����9d\��?ݻ�E<�����ټ����mR�����䳽C�i���� ��6��nH��T�      �� ]�ӈ�p}���w�ý�u��ʕ���K�����o�jv���&R�!��Z^����� �>����:UB;3";`�4;��>;=D;��F;�G;�)H;adH;m�H;�H;\�H;#�H;'�H;|�H;��H;�H;�H;��H;
�H;�H;��H;|�H;'�H;%�H;a�H;	�H;p�H;cdH;�)H;�G;��F;AD;��>;c�4;>";[B;���: �>����X^�����&R�iv���o�����K�ʕ���u��w�ý��p}�ӈ� ]�       �ѽ\νy�ý䳽9����L����d�q\8�v��ټiv����Y��_����D���[�t�Y:G��:Am;�r-;�:;j�A;(oE;�"G;F�G;UGH;�sH;ߐH;��H;�H;�H;�H;��H;r�H;z�H;%�H;��H;%�H;{�H;x�H;��H;�H;#�H;�H;��H;�H;�sH;UGH;J�G;�"G;0oE;l�A;�:;�r-;Hm;Q��:��Y:�[�@������_���Y�iv��ټu��q\8���d��L��:���䳽y�ý\ν      ���������Ȅ�jSt��Y�\n;�/O�n#���Oļ�����&R��_������N3���Y��3:��:̯;�?&;�G6;xX?;�D;"xF;��G;'!H;�^H;��H;�H;��H;8�H;��H;��H;��H;�H;��H;M�H;�H;M�H;��H;�H;��H;��H;��H;B�H;ƭH;�H;��H;^H;.!H;��G;&xF;�D;}X?;�G6;�?&;ί;��:�3:�Y��N3������_��&R������Oļm#��/O�[n;��Y�jSt��Ȅ�����      ]n;�x\8��s/�=�!�y��_���irμ��������E<�������N3�lHx�x�9��:�^;J ;"2;[�<;�B;��E;!5G;��G;$FH;vqH;��H;;�H;��H;C�H;��H;��H;��H;��H;�H;k�H; �H;k�H;�H;��H;��H;��H;��H;M�H;��H;A�H;��H;sqH;*FH;��G;(5G;��E;�B;f�<;)2;M ;�^;��:��9XHx��N3�������E<��������irμ^���z��=�!��s/�w\8�      Y������o�orμσ��sv��I"��^N�����?ݻX^��H�� �Y�x�9��:ʦ�:��;G�.;t|:;�>A;��D; �F;��G;�)H;aH;�H;r�H;جH;)�H;�H;,�H;T�H;��H;�H;M�H;��H;��H;��H;K�H;�H;��H;S�H;/�H;�H;/�H;ݬH;r�H;�H;aH;�)H;��G;#�F;��D;�>A;{|:;F�.;��;̦�:��:��9�Y�C��V^���?ݻ���^N�I"��rv��у��prμ�o����      �����x���#��@F{���]��E<����L�뻬���7d\�����[��3:��:̦�:r[;X�,;��8;!@;�0D;l[F;{G;�
H;8PH;vH;אH;4�H;�H;�H;[�H;o�H;��H;��H;q�H;m�H;��H;��H;��H;j�H;s�H;��H;��H;q�H;`�H; �H;�H;5�H;ѐH;vH;:PH;�
H;{G;p[F;�0D;!@;��8;a�,;s[;Ԧ�:��:�3:�[����5d\�����K�뻢���E<���]�AF{��#���x��      �B(�%�����_������˻	���b�@&����� �>���Y:��:�^;��;^�,;`8;[�?;��C;gF;�FG;<�G;�?H;kH;�H;��H;�H;I�H;��H;_�H;h�H;�H;r�H;��H;��H;}�H;��H;x�H;~�H;��H;p�H;�H;l�H;`�H;��H;L�H;�H;�H;�H;kH;�?H;@�G;�FG;qF;��C;W�?;`8;_�,;��;�^;��:��Y: �>�����;&��b�	���˻�����_����%�      Ϛ��K���(J���X���b���-���� Ix�@��� :���:A��:ǯ;I ;D�.;��8;P�?;�C;��E;&#G;��G;�1H;�aH;=�H;g�H;l�H;��H;��H;P�H;�H;%�H;-�H;��H;�H;��H;3�H;��H;0�H;~�H;�H;��H;-�H;)�H;�H;R�H;��H;��H;f�H;n�H;=�H;�aH;�1H;��G;+#G;��E;�C;T�?;��8;F�.;I ;ȯ;C��:���:� :����Hx������-��b��X��"J��L���      4�����<кʓ��ćY����pr8985:?/�:�d�:_B;Cm;�?&;'2;z|:;!@;��C;��E;kG;��G;H(H;�ZH;]zH;,�H;ŤH;��H;Y�H;��H;��H;S�H;��H;��H;B�H;$�H;C�H;��H;u�H;��H;@�H;!�H;@�H;��H;��H;W�H;��H;��H;W�H;��H;̤H;/�H;\zH;�ZH;L(H;��G;nG;��E;��C;!@;z|:;&2;�?&;Cm;aB;�d�:A/�:85:Pr89 ����Y�䓤�<к���      ��e9�9p	�9|: �Y:`y�:g;�:ծ�:�^;��;=";�r-;�G6;a�<;�>A;�0D;mF;1#G;��G;�$H;OWH;�vH;f�H;1�H;4�H;l�H;�H;�H;n�H;-�H;��H;u�H;��H;!�H;�H;��H;��H;��H;�H; �H;��H;u�H;��H;-�H;m�H;��H;��H;k�H;:�H;4�H;d�H;�vH;UWH;�$H;��G;-#G;nF;�0D;�>A;]�<;�G6;�r-;>";��;�^;ۮ�:a;�:jy�:0�Y:4: 	�9��9      A�:D-�:g�:��:��:�^;Y�;%�;��#; �,;_�4; �:;zX?;�B;��D;r[F;�FG;��G;K(H;MWH;YuH;|�H;
�H;�H;�H;��H;��H;��H;��H;��H;��H;��H;��H;��H;��H;Q�H;L�H;J�H;��H;��H;��H;��H;��H;��H;��H;��H;��H;��H;�H;�H;�H;��H;_uH;OWH;L(H;��G;�FG;o[F;��D;�B;xX?;��:;c�4;�,;��#;"�;]�;�^;��:
��:+g�:@-�:      �;m�;�l;�Z;\`;�%;�+;��0;�G6;y�:;��>;j�A;�D;��E;#�F;{G;B�G;�1H;�ZH;�vH;��H;=�H;��H;¸H;{�H;J�H;��H;��H;��H;��H;0�H;1�H;��H;��H;d�H;��H;��H;��H;a�H;��H;��H;.�H;4�H;��H;��H;��H;��H;H�H;~�H;��H;��H;?�H;��H;�vH;�ZH;�1H;C�G;{G;#�F;��E;�D;g�A;��>;s�:;�G6;��0;�+;�%;p`;�Z;�l;a�;      �Y.;��.;0;�2;*�4;��7;_|:;"]=;<�?;Z7B;BD;,oE;$xF;/5G;��G;�
H;�?H;�aH;`zH;f�H;	�H;��H;A�H;��H;Z�H;��H;��H;��H;�H;��H;��H;U�H;O�H;?�H;��H;�H;?�H;�H;��H;A�H;N�H;U�H;��H;��H;�H;��H;��H;��H;^�H;��H;;�H;��H;
�H;d�H;`zH;�aH;�?H;�
H;��G;)5G;$xF;,oE;AD;R7B;>�?;"]=;X|:;}�7;9�4;�2;0;��.;      M�<; �<;]=;�O>;ہ?;u�@;x7B;:�C;�D;��E;��F;�"G;��G; �G;�)H;?PH;kH;E�H;/�H;2�H;�H;��H;��H;/�H;(�H;*�H;<�H;��H;�H;3�H;��H;�H;�H;��H;?�H;{�H;��H;t�H;<�H;��H;�H;�H;��H;3�H;�H;��H;8�H;-�H;*�H;+�H;��H;��H;�H;/�H;.�H;=�H;kH;;PH;�)H;��G;��G;�"G;��F;��E;�D;=�C;q7B;`�@;�?;�O>;]=;�<;      ~WC;�nC;βC;aD;1�D;5E;��E;�[F;E�F;oLG;��G;M�G;.!H;1FH;aH;vH;��H;v�H;֤H;A�H;�H;~�H;a�H;3�H;��H;��H;9�H;��H;��H;��H;��H;��H;��H;.�H;��H;��H;��H;��H;��H;/�H;��H;��H;��H;��H;��H;��H;6�H;��H;��H;/�H;^�H;��H;�H;;�H;ԤH;q�H;��H;vH;aH;+FH;-!H;P�G;��G;nLG;E�F;�[F;��E;5E;9�D;cD;˲C;�nC;      �ZF;�dF;ڀF;"�F;��F;�"G;�aG;۞G;��G;/H;�)H;YGH;�^H;}qH;�H;ېH;��H;m�H;��H;k�H;��H;D�H;��H;0�H;��H;�H;��H;��H;e�H;��H;��H;��H;�H;q�H;��H;�H;�H;�H;��H;q�H;�H;��H;��H;��H;c�H;��H;��H;!�H;��H;-�H;��H;G�H;��H;i�H;��H;i�H;��H;ڐH;�H;xqH;�^H;XGH;�)H;.H;��G;۞G;�aG;�"G;��F;-�F;׀F;�dF;      �G;�G;d�G;w�G;��G;�G;tH;�)H;�?H;WSH;ddH;�sH;��H;��H;q�H;6�H;�H;��H;]�H;�H;��H;��H;��H;B�H;6�H;��H;��H;;�H;{�H;��H;[�H;��H;m�H;��H;��H;3�H;N�H;,�H;��H;��H;l�H;��H;[�H;��H;x�H;8�H;�H;��H;;�H;>�H;��H;��H;��H;��H;Z�H;��H;�H;6�H;n�H;��H;�H;�sH;cdH;SSH;�?H;�)H;nH;��G;�G;o�G;f�G;֪G;      �/H;�1H;6H;=H;�EH;4PH;�ZH;�eH;�pH;�{H;n�H;�H;�H;B�H;׬H;�H;J�H;��H;��H;��H;��H;��H;��H;��H;��H;��H;6�H;r�H;Y�H;H�H;��H;_�H;��H;�H;?�H;T�H;?�H;O�H;=�H;�H;��H;[�H;��H;F�H;W�H;q�H;5�H;��H;��H;��H;��H;��H;��H;~�H;��H;��H;I�H;�H;֬H;>�H;�H;�H;r�H;�{H;�pH;�eH;�ZH;(PH;FH;=H;6H;�1H;      'jH;�jH;mH;�pH;2uH;�zH;h�H;l�H;ӏH;{�H;�H;��H;ƭH;��H;*�H;!�H;��H;Y�H;��H;r�H;��H;��H;�H;�H;��H;b�H;u�H;Z�H;P�H;��H;J�H;��H;��H;.�H;]�H;d�H;U�H;`�H;[�H;/�H;��H;��H;L�H;��H;M�H;Y�H;q�H;c�H;��H;�H;�H;��H;��H;m�H;��H;U�H;��H;#�H;*�H;��H;ĭH;��H;
�H;|�H;ԏH;n�H;b�H;�zH;>uH;�pH;mH;�jH;      4�H;��H;.�H;��H;��H;��H;*�H; �H;r�H;�H;_�H;�H;?�H;M�H;�H;]�H;f�H;�H;S�H;.�H;��H;��H;��H;3�H;��H;��H;��H;F�H;��H;@�H;��H;��H;.�H;V�H;b�H;w�H;��H;u�H;_�H;U�H;)�H;��H;��H;=�H;��H;F�H;}�H;��H;��H;.�H;��H;��H;��H;*�H;Q�H;�H;c�H;`�H;�H;I�H;>�H;�H;a�H;�H;q�H;!�H;,�H;��H;��H;��H;.�H;��H;      H�H;��H;��H;G�H;��H;T�H;��H;;�H;�H;�H;,�H;*�H;�H;��H;2�H;v�H;s�H;/�H;��H;��H;��H;6�H;��H;��H;��H;��H;[�H;��H;P�H;��H;��H;!�H;X�H;f�H;�H;~�H;x�H;{�H;|�H;g�H;V�H; �H;��H;��H;J�H;��H;W�H;��H;��H;��H;��H;6�H;��H;��H;��H;-�H;s�H;w�H;3�H;��H;�H;*�H;*�H;�H;�H;>�H;��H;J�H;��H;G�H;��H;��H;      ��H;εH;{�H;ŷH;z�H;m�H;�H;��H;N�H;9�H;+�H;�H;��H;��H;V�H;��H;�H;3�H;��H;{�H;��H;2�H;V�H;	�H;��H;��H;��H;a�H;��H;��H;�H;9�H;b�H;~�H;��H;��H;��H;��H;��H;�H;b�H;7�H;�H;��H;��H;^�H;��H;��H;��H; �H;Y�H;4�H;��H;x�H;��H;4�H;�H;��H;V�H;��H;��H;�H;.�H;9�H;N�H;��H;��H;n�H;��H;ƷH;��H;˵H;      ,�H;p�H;�H;��H;�H;��H;E�H;�H;&�H;Q�H;��H;��H;��H;��H;��H;��H;w�H;��H;H�H;��H;��H;��H;O�H;�H;��H;�H;o�H;��H;��H;0�H;T�H;c�H;w�H;��H;��H;��H;��H;��H;��H;��H;t�H;c�H;R�H;,�H;��H;��H;j�H;�H;��H;�H;R�H;��H;��H;��H;H�H;��H;z�H;��H;��H;��H;��H;��H;��H;R�H;*�H;�H;E�H;{�H;�H;��H;�H;p�H;      ��H;��H;>�H;��H;��H;��H;G�H;��H;k�H;�H;��H;|�H;�H;��H;�H;v�H;��H;�H;'�H;'�H;��H;��H;<�H;��H;*�H;o�H;��H;	�H;.�H;X�H;`�H;�H;��H;�H;��H;��H;��H;��H;��H;�H;��H;�H;`�H;U�H;)�H;�H;��H;p�H;-�H;��H;B�H;��H;��H; �H;&�H;�H;��H;w�H;�H;��H;�H;|�H;��H;�H;n�H;��H;K�H;��H;��H;��H;E�H;��H;      P�H;u�H;��H;b�H;+�H;�H;�H;*�H;r�H;��H;!�H;��H;��H;�H;T�H;o�H;��H;�H;A�H;�H;��H;a�H;��H;2�H;��H;��H;��H;=�H;_�H;d�H;x�H;��H;��H;��H;��H;��H;��H;��H;��H;��H;��H;��H;w�H;_�H;X�H;9�H;��H;��H;��H;2�H;��H;`�H;��H;�H;A�H;��H;��H;t�H;U�H;�H;��H;��H;$�H;��H;w�H;-�H;�H; �H;)�H;c�H;��H;v�H;      ��H;��H;�H;w�H;�H;��H;��H;��H;��H;��H;�H;)�H;N�H;p�H;��H;��H;{�H;/�H;��H;��H;S�H;��H;�H;l�H;��H;�H;.�H;R�H;i�H;|�H;{�H;��H;��H;��H;��H;��H;��H;��H;��H;��H;��H;��H;z�H;w�H;c�H;N�H;,�H;�H;��H;l�H;�H;��H;M�H;��H;��H;5�H;�H;��H;��H;q�H;P�H;'�H;�H;��H;��H;��H;��H;��H;�H;v�H;�H;��H;      ��H;��H;��H;^�H;��H;��H;y�H;l�H;z�H;��H;��H;��H;�H;
�H;��H;��H;��H;��H;x�H;��H;T�H;��H;B�H;��H;��H;�H;M�H;F�H;\�H;��H;t�H;��H;��H;��H;��H;��H;��H;��H;��H;��H;��H;��H;t�H;��H;U�H;@�H;J�H;	�H;��H;��H;C�H;��H;M�H;��H;x�H;��H;��H;��H;��H;�H;�H;��H;��H;��H;}�H;o�H;}�H;��H;��H;_�H;��H;��H;      ��H;��H;��H;y�H;�H;��H;��H;��H;��H;��H;�H;)�H;Q�H;r�H;��H;��H;}�H;0�H;��H;��H;T�H;��H;�H;l�H;��H;�H;.�H;R�H;j�H;{�H;{�H;��H;��H;��H;��H;��H;��H;��H;��H;��H;��H;��H;z�H;u�H;c�H;M�H;+�H;�H;��H;j�H;�H;��H;M�H;��H;��H;5�H;~�H;��H;��H;p�H;Q�H;'�H;�H;��H;��H;��H;��H;��H;�H;z�H;�H;��H;      F�H;w�H;��H;[�H;)�H;��H;�H;-�H;r�H;��H;!�H;��H;��H;�H;U�H;q�H;��H;��H;A�H;�H;��H;d�H;��H;4�H;��H;��H;��H;=�H;]�H;c�H;w�H;��H;��H;��H;��H;��H;��H;��H;��H;��H;��H;��H;w�H;]�H;X�H;6�H;��H;��H;��H;1�H;��H;a�H;��H;�H;A�H;��H;��H;t�H;T�H;�H;��H;��H;!�H;��H;t�H;1�H;�H;��H;.�H;\�H;��H;y�H;      ��H;��H;;�H;��H;��H;��H;D�H;��H;m�H;�H;��H;|�H;�H;��H;�H;w�H;��H;�H;'�H;%�H;��H;��H;>�H;��H;.�H;o�H;��H;	�H;.�H;X�H;`�H;�H;��H;�H;��H;��H;��H;��H;��H;�H;��H;�H;_�H;U�H;'�H;�H;��H;p�H;+�H;��H;B�H;��H;��H;!�H;'�H;�H;��H;z�H;�H;��H;�H;|�H;��H;�H;p�H;��H;L�H;��H;��H;��H;D�H;��H;      ,�H;x�H;�H;��H;�H;��H;B�H;�H;'�H;Q�H;��H;��H;��H;��H;��H;��H;z�H;��H;G�H;��H;��H;��H;N�H;�H;��H;�H;m�H;��H;��H;0�H;R�H;`�H;u�H;��H;��H;��H;��H;��H;��H;��H;t�H;c�H;R�H;+�H;��H;��H;j�H;�H;��H;��H;S�H;��H;��H;��H;E�H;��H;y�H;��H;��H;��H;��H;��H;��H;O�H;)�H;�H;J�H;|�H;�H;��H;�H;p�H;      s�H;ѵH;n�H;��H;x�H;|�H;��H;��H;L�H;9�H;-�H;�H;��H;��H;X�H;��H;�H;4�H;��H;|�H;��H;6�H;U�H;�H;��H;��H;��H;a�H;��H;��H;�H;7�H;c�H;|�H;��H;��H;��H;��H;��H;~�H;b�H;7�H;�H;��H;��H;[�H;��H;��H;��H;��H;Y�H;4�H;��H;w�H;��H;2�H;�H;��H;W�H;��H;��H;�H;-�H;<�H;O�H;��H;��H;o�H;}�H;·H;t�H;˵H;      <�H;��H;��H;A�H;��H;T�H;��H;=�H;�H;�H;*�H;-�H;�H;��H;3�H;w�H;u�H;-�H;��H;��H;��H;7�H;��H;��H;��H;��H;X�H;��H;P�H;��H;��H;!�H;X�H;f�H;��H;|�H;x�H;~�H;|�H;g�H;Y�H;!�H;��H;��H;I�H;��H;V�H;��H;��H;��H;��H;6�H;��H;��H;��H;-�H;u�H;w�H;5�H;��H;�H;,�H;*�H;�H;�H;A�H;��H;Q�H;��H;N�H;��H;��H;      E�H;��H;)�H;��H;��H;ėH;)�H;(�H;u�H;�H;_�H;�H;A�H;L�H;�H;_�H;d�H;�H;S�H;.�H;��H;��H;��H;0�H;��H;��H;��H;I�H;��H;B�H;��H;��H;(�H;V�H;b�H;u�H;��H;w�H;_�H;V�H;,�H;��H;��H;=�H;��H;C�H;|�H;��H;��H;-�H;��H;��H;��H;*�H;S�H;�H;c�H;_�H;�H;L�H;?�H;�H;_�H;�H;r�H;'�H;-�H;��H;ƓH;��H;:�H;��H;      8jH;�jH;)mH;�pH;+uH;�zH;c�H;o�H;ۏH;x�H;�H;��H;ǭH;��H;/�H;#�H;��H;Y�H;��H;o�H;��H;��H;�H;�H;��H;^�H;r�H;Z�H;Q�H;��H;L�H;��H;��H;.�H;\�H;c�H;U�H;c�H;[�H;.�H;��H;��H;L�H;��H;J�H;S�H;q�H;b�H;��H;�H;�H;��H;��H;n�H;��H;U�H;��H;$�H;/�H;��H;ƭH;��H;�H;y�H;ݏH;r�H;h�H;�zH;<uH;�pH;)mH;�jH;      
0H;�1H;6H;=H;�EH;APH;�ZH;�eH;�pH;�{H;q�H;�H;�H;B�H;ڬH;��H;J�H;��H;��H;~�H;��H;��H;��H;��H;��H;��H;5�H;r�H;\�H;E�H;��H;a�H;��H;�H;?�H;Q�H;@�H;R�H;<�H;�H;��H;^�H;��H;E�H;U�H;m�H;2�H;��H;��H;��H;��H;��H;��H;~�H;��H;��H;L�H;��H;ڬH;?�H;�H;�H;r�H;�{H;�pH;�eH;�ZH;/PH;FH;=H;6H;�1H;      ��G;�G;g�G;��G;�G;
�G;uH;�)H;�?H;USH;ddH;�sH;�H;��H;r�H;8�H;�H;��H;Z�H;��H;��H;��H;��H;C�H;9�H;��H;�H;9�H;|�H;��H;Z�H;��H;m�H;��H;��H;/�H;O�H;/�H;��H;��H;o�H;��H;[�H;��H;w�H;5�H;|�H;��H;7�H;>�H;��H;��H;��H;�H;\�H;��H;�H;9�H;t�H;��H;~�H;�sH;cdH;SSH;�?H;�)H;zH;�G;�G;��G;k�G;�G;      �ZF;�dF;�F;�F;��F;�"G;�aG;ݞG;��G;0H;�)H;\GH;�^H;yqH;�H;ݐH;��H;o�H;��H;k�H;��H;G�H;��H;0�H;��H;�H;��H;��H;h�H;��H;��H;��H;�H;s�H;��H;�H;�H;�H;��H;q�H;�H;��H;��H;��H;a�H;��H;��H;�H;��H;-�H;��H;F�H;��H;i�H;��H;i�H;��H;ݐH;	�H;xqH;�^H;WGH;�)H;/H;��G;ٞG;�aG;�"G;��F;"�F;ˀF;zdF;      }WC;�nC;˲C;bD;-�D;!5E;��E;�[F;K�F;oLG;��G;P�G;-!H;-FH;aH;vH;��H;v�H;ԤH;<�H;�H;��H;\�H;3�H;��H;��H;6�H;��H;��H;��H;��H;��H;��H;/�H;��H;��H;��H;��H;��H;/�H;��H;��H;��H;��H;��H;��H;7�H;��H;��H;0�H;b�H;��H;�H;>�H;֤H;r�H;��H;vH;aH;-FH;.!H;M�G;��G;nLG;G�F;�[F;��E;5E;;�D;bD;̲C;�nC;      0�<;�<;]=;�O>;ׁ?;|�@;v7B;<�C;��D;��E;��F;�"G;��G;��G;�)H;>PH;kH;D�H;.�H;/�H;�H;��H;��H;/�H;*�H;'�H;:�H;��H;�H;1�H;��H;
�H;�H;��H;=�H;x�H;��H;z�H;<�H;��H;�H;	�H;��H;3�H;�H;��H;<�H;,�H;)�H;/�H;��H;��H;�H;2�H;0�H;>�H;kH;=PH;�)H;��G;��G;�"G;��F;��E;�D;6�C;u7B;r�@;��?;�O>;]=;��<;      �Y.;��.;
0;�2;(�4;|�7;W|:;"]=;?�?;V7B;=D;/oE;$xF;,5G;��G;�
H;�?H;�aH;^zH;d�H;	�H;��H;;�H;��H;^�H;��H;��H;��H;�H;��H;��H;V�H;N�H;?�H;��H;�H;B�H;�H;��H;>�H;O�H;V�H;��H;��H;�H;��H;��H;��H;[�H;��H;?�H;��H;
�H;f�H;`zH;�aH;�?H;�
H;��G;)5G;$xF;,oE;@D;X7B;?�?;%]=;X|:;~�7;(�4;�2;	0;~�.;      �;m�;�l;�Z;\`;�%;�+;��0;�G6;u�:;��>;n�A;�D;��E;&�F;{G;B�G;�1H;�ZH;�vH;��H;?�H;��H;��H;�H;D�H;��H;��H;��H;��H;3�H;2�H;��H;��H;a�H;��H;��H;��H;a�H;��H;��H;1�H;6�H;��H;��H;��H;��H;H�H;|�H;øH;��H;?�H;��H;�vH;�ZH;�1H;B�G;{G;%�F;��E;�D;i�A;��>;v�:;�G6;��0;�+;�%;t`;�Z;�l;`�;      7�:t-�:5g�:��:��:�^;Z�;'�;��#;�,;c�4;�:;zX?;�B;��D;r[F;�FG;��G;K(H;MWH;\uH;��H;�H;�H;�H;��H;��H;��H;��H;��H;��H;��H;��H;��H;��H;M�H;M�H;O�H;��H;��H;��H;��H;��H;��H;��H;��H;��H;��H;�H;�H;	�H;|�H;\uH;PWH;L(H;��G;�FG;o[F;��D;�B;zX?;��:;c�4; �,;��#;*�;^�;�^;��:��:Ig�:F-�:      `�e9X�9X	�9x:$�Y:ny�:o;�:��:�^;��;A";�r-;�G6;a�<;�>A;�0D;nF;0#G;��G;�$H;UWH;�vH;f�H;2�H;:�H;i�H;��H;��H;n�H;*�H;��H;w�H;��H;"�H;�H;��H;��H;��H;�H;�H;��H;u�H;��H;*�H;n�H;~�H;�H;l�H;5�H;5�H;g�H;�vH;RWH;�$H;��G;+#G;lF;�0D;�>A;]�<;�G6;�r-;@";��;�^;ۮ�:c;�:\y�:<�Y:D:X	�9 �9      0�����8кΓ��ЇY����Pr89<5:G/�:�d�:aB;Em;�?&;'2;~|:;!@;��C;��E;lG;��G;N(H;�ZH;`zH;.�H;̤H;��H;U�H;��H;��H;S�H;��H;��H;A�H;$�H;D�H;��H;u�H;��H;C�H;#�H;A�H;��H;��H;U�H;��H;��H;Y�H;��H;ǤH;/�H;^zH;�ZH;K(H;��G;kG;��E;��C;!@;||:;%2;�?&;Cm;_B;�d�:C/�:<5:Pr89 ��ЇY�Г��Fк���      ֚��F���(J���X���b���-�����Hx����� :���:I��:˯;J ;J�.;��8;S�?;�C;��E;*#G;��G;�1H;�aH;>�H;n�H;j�H;��H;��H;U�H;�H;(�H;-�H;��H;�H;�H;2�H;��H;3�H;}�H;�H;��H;,�H;)�H;�H;R�H;��H;��H;i�H;g�H;=�H;�aH;�1H;��G;*#G;��E;��C;Q�?;��8;J�.;G ;ʯ;C��:���:� :����Hx������-��b��X��,J��H���      �B(�%�����_������˻	���b�<&����� �>���Y:��:�^;��;d�,;`8;Z�?;��C;mF;�FG;@�G;�?H;kH;��H;��H;�H;H�H;��H;]�H;l�H;�H;s�H;��H;��H;{�H;��H;{�H;~�H;��H;o�H;�H;l�H;`�H;��H;H�H;�H;��H;�H;kH;�?H;=�G;�FG;nF;��C;U�?;`8;_�,;��;�^;��:��Y: �>�����;&��b�	���˻�����_����%�      �����x���#��@F{���]��E<����J�뻪���5d\�~�뺼[��3:��:ڦ�:w[;]�,;��8;!@;�0D;r[F;{G;�
H;=PH;vH;ؐH;4�H;�H; �H;[�H;q�H;��H;��H;t�H;o�H;��H;��H;��H;j�H;p�H;��H;��H;p�H;]�H;�H;�H;1�H;ԐH;	vH;8PH;�
H;{G;i[F;�0D;!@;��8;[�,;r[;Ҧ�:��:�3:�[����7d\�����K�뻤���E<���]�AF{��#���x��      Z������o�orμσ��rv��I"��^N�����?ݻV^��D���Y���9��:Ԧ�:��;G�.;z|:;�>A;��D;#�F;��G;�)H;aH;�H;p�H;۬H;/�H;�H;/�H;V�H;��H;�H;M�H;��H;��H;��H;M�H;�H;��H;Q�H;.�H;�H;/�H;ڬH;n�H;�H;aH;�)H;��G;#�F;��D;�>A;u|:;C�.;��;Ʀ�:��:��9��Y�F��X^���?ݻ���^N�J"��rv��у��prμ�o����      ]n;�x\8��s/�<�!�y��^���irμ��������E<�������N3�XHx���9��:�^;K ;%2;_�<;�B;��E;'5G;�G;+FH;yqH;��H;>�H;��H;F�H;��H;��H;��H;��H;�H;j�H; �H;m�H;�H;��H;��H;��H;��H;J�H;��H;>�H;��H;uqH;&FH; �G;)5G;��E;�B;b�<; 2;I ;�^;��:��9`Hx��N3�������E<��������jrμ^���z��<�!��s/�w\8�      ���������Ȅ�jSt��Y�\n;�/O�n#���Oļ�����&R��_������N3�܅Y��3:��:̯;�?&;�G6;�X?;�D;'xF;��G;.!H;�^H;�H;�H;ĭH;<�H;��H;��H;��H;	�H;��H;M�H;�H;M�H;��H;�H;��H;��H;��H;>�H;ƭH;�H;~�H;�^H;)!H;��G;&xF;�D;vX?;�G6;�?&;ȯ;��:�3:�Y��N3������_��&R������Oļm#��/O�[n;��Y�jSt��Ȅ�����       �ѽ\νy�ý䳽9����L����d�q\8�u��ټiv����Y��_����@���[���Y:C��:Em;�r-;�:;j�A;/oE;�"G;K�G;WGH;�sH;ߐH;��H;�H;%�H;�H;��H;v�H;{�H;#�H;��H;%�H;z�H;t�H;��H;�H;!�H;�H;��H;ߐH;sH;UGH;D�G;�"G;-oE;j�A;�:;�r-;Am;C��:��Y:�[�@������_���Y�iv��ټv��q\8���d��L��:���䳽y�ý\ν      �� ]�ӈ�p}���w�ý�u��ʕ���K�����o�jv���&R� ��V^����� �>����:WB;9";g�4;��>;BD;��F;�G;�)H;`dH;n�H;�H;^�H;&�H;*�H;}�H;��H;�H;
�H;��H;	�H;�H;��H;z�H;&�H;"�H;^�H;
�H;n�H;^dH;�)H;�G;��F;AD;��>;\�4;7";UB;���: �>����X^�� ���&R�jv���o�����K�ʕ���u��w�ý��p}�ӈ� ]�      �+X��T��nH��6��� �i��C�䳽�����mR����ټ�����E<��?ݻ8d\������ :�d�:��;'�,;u�:;Z7B;��E;nLG;,H;USH;�{H;|�H;�H;�H;7�H;O�H;
�H;��H;��H;��H;��H;��H;�H;M�H;6�H;�H;�H;�H;�{H;SSH;,H;hLG;��E;Y7B;u�:;�,;��;�d�:� :����<d\��?ݻ�E<�����ټ����mR�����䳽C�i���� ��6��nH��T�      ఖ�����}���*|�LS\�� :����Z�l$�������K�v���Oļ����������C&����9/�:�^;��#;�G6;8�?;��D;H�F;��G;�?H;�pH;ݏH;r�H;�H;G�H;-�H;j�H;m�H;��H;w�H;��H;m�H;g�H;)�H;G�H;�H;r�H;ޏH;�pH;�?H;��G;D�F;��D;9�?;�G6;��#;�^;//�:`��D&������������Oļv���K�����k$���Z���� :�LS\��*|�}������      @�;9ɾ{㼾B�������Mw��nH�����Z�䳽ʕ��q\8�o#������^N�O���b�$Ix�,5:ٮ�:-�;��0;]=;=�C;�[F;ҞG;�)H;�eH;o�H; �H;:�H;��H;�H;��H;&�H;��H;i�H;��H;'�H;��H;�H;|�H;9�H;$�H;r�H;�eH;�)H;֞G;�[F;<�C;]=;��0;&�;��:5:Ix��b�P��^N�����o#��q\8�ʕ��䳽�Z񽰯��nH��Mw�����B��{㼾9ɾ      0y��v�j���B�߾����@��?����nH���CὝu����d�0O�jrμJ"�����	������q89Y;�:[�;�+;Q|:;v7B;��E;�aG;jH;�ZH;b�H;)�H;��H;�H;E�H;B�H; �H;��H;q�H;��H;�H;A�H;B�H;�H;��H;,�H;c�H;�ZH;kH; bG;��E;u7B;R|:;�+;W�;];�:�q89���	�����J"��jrμ0O���d��u��C����nH�?���@������B�߾j����v�      �O/�pM+�X�����HW��9ɾ@���Mw�� :�i��w�ý�L��\n;�^���sv���E<��˻��-�P��by�:�^;�%;~�7;t�@;5E;�"G;�G;4PH;�zH;��H;W�H;v�H;��H;��H;�H;��H;��H;��H;�H;��H;��H;v�H;S�H;��H;�zH;7PH;�G;�"G;5E;t�@;}�7;�%;�^;hy�:h����-��˻�E<�sv��^���\n;��L��w�ýj��� :��Mw�@��9ɾHW�����X��pM+�      7�X�VvS�6E��O/��S�HW����������LS\��� ���:����Y�{��Ѓ����]�����*�b���Y�<�Y:��:``;6�4;�?;7�D;��F;�G;�EH;@uH;��H;��H;}�H;�H;��H;�H;�H;��H;�H;�H;��H;�H;}�H;��H;ēH;DuH;FH;�G;��F;7�D;�?;2�4;``;��:@�Y:��Y�%�b�������]�Ѓ��{���Y�9����彑� �LS\���������HW���S��O/�6E�VvS�      � ����y�a�h��N��O/����B�߾B���*|��6�p}�䳽jSt�<�!�prμCF{��_��X��֓��@:"��:�Z;�2;�O>;iD;"�F;p�G;=H;�pH;��H;G�H;ƷH;��H;��H;X�H;w�H;[�H;u�H;X�H;��H;��H;ȷH;D�H;��H;�pH;=H;w�G;/�F;jD;�O>;�2;�Z; ��:X:ړ���X���_�BF{�orμ<�!�jSt�䳽p}��6��*|�B��B�߾����O/��N�a�h���y�      =v��b���W ��a�h�6E�X��j���|㼾}���nH�ӈ�y�ý�Ȅ��s/��o��#�����(J��8к0	�9Mg�:�l;0;]=;ֲC;ҀF;g�G;6H;mH;$�H;��H;{�H;��H;;�H;��H;�H;��H;��H;��H;;�H;��H;z�H;��H;)�H;mH;6H;n�G;��F;ֲC;]=;0;�l;Mg�:X	�96к%J������#���o��s/��Ȅ�y�ýӈ��nH�}��|㼾j���X��6E�a�h�W ��b���      |h��/���b�����y�VvS�pM+��v�9ɾ�����T� ]�\ν����x\8�����x��%�Q������@�9f-�:c�;��.;�<;�nC;�dF;�G;�1H;�jH;��H;��H;ǵH;d�H;��H;a�H;��H;��H;��H;b�H;��H;c�H;ǵH;��H;��H;�jH;�1H;�G;�dF;�nC;�<;��.;a�;f-�:`�9���O���%��x�����x\8�����\ν ]��T�����9ɾ�v�pM+�VvS���y�b���/���      dܿ3�ֿ�aǿ=^��/���Xo���7����iþ�(���-=��` �A���_�1]�/p����I�U�ѻ��)���R���:*�
;�*;�:;��B;�HF;!�G;�lH;�H;q�H;:�H;��H;{�H;J�H;y�H;	�H;��H;�H;y�H;L�H;{�H;��H;9�H;y�H;�H;�lH;'�G; IF;��B;�:;�*;*�
;��:`�R���)�R�ѻ��I�/p��1]��_�A���` ��-=��(���iþ����7�Xo�/���>^���aǿ3�ֿ      2�ֿCpѿ�¿������_Xi�ϕ3��
�VD��Fl��A�9��.���R�� \� �ex��2�E��ͻ#�$�� �э�:8�;H�*;1�:;�B;�TF;��G;%nH;��H;��H;i�H;��H;��H;X�H;|�H;�H;��H;�H;�H;W�H;��H;��H;d�H;·H;��H;&nH;��G;�TF;�B;.�:;B�*;8�;Ս�:@ �"�$��ͻ2�E�ex�� �!\��R���.��A�9�Fl��VD���
�ϕ3�_Xi��������¿Cpѿ      �aǿ�¿����������"Y��f'�����7o���.}��k/����$ڟ�!<Q�-#�ע��(;�0���?�� l7���:�;q,;��;;�C;�vF;�G;�rH;�H;��H;�H;��H;��H;��H;��H;J�H;��H;C�H;��H;��H;��H;��H;
�H;��H;�H;�rH;�G;wF;�C;�;;j,;�;��: e7�@��.����(;�ע�-#�"<Q�$ڟ�����k/��.}�7o�������f'��"Y�����������¿      =^������k���Yo���@�(�$�޾����:ce�0����ڽ���� g@������R���O*�LG�� ���PC^9$��: ;Zd.;��<;��C;�F;��G;�yH;��H;�H;�H;��H;g�H;��H;��H;~�H;�H;x�H;��H;��H;e�H;��H;�H;�H;��H;�yH;��G;��F;��C;��<;Sd.;�;&��:�C^9 ���IG���O*��R������ g@�������ڽ0��:ce�����$�޾(���@�Yo�k�������      /����������Yo��!J�K�#��\��VD������zPH�����b�� C��� +���ټ)��������T�:��:>�;�Y1;>;�0D;y�F;[H;A�H;��H;�H;X�H;��H;�H;_�H;E�H;��H;\�H;��H;F�H;^�H;�H;��H;T�H;�H;¨H;B�H;^H;��F;�0D;>;�Y1;A�;��:p�:�������)����ټ� +� C���b�����zPH�����VD���\��K�#��!J�Yo��������      Xo�_Xi��"Y���@�K�#��
��о�A���i���(�~��ur���_��5��ɺ�r�`��<��k�d�|�\�D�X:�P�:�`;ȱ4;��?;��D;r8G;g0H;��H;g�H;p�H; �H;��H;��H;��H;��H;�H;��H;�H;��H;��H;��H;��H;��H;t�H;j�H;��H;g0H;y8G;��D;��?;ű4;�`;�P�:L�X:x�\�f�d��<��r�`��ɺ��5��_�ur��~����(��i��A���о�
�K�#���@��"Y�_Xi�      ��7�ϕ3��f'�(��\���о�����.}��-=�{
���Ľ[��,:����������7�&GĻʃ$�@O�����:�{;D&;�+8;JA;�E;��G;wLH;�H;r�H;/�H;��H;��H;��H;��H;�H;~�H;�H;{�H;�H;��H;��H;��H;��H;4�H;u�H;�H;tLH;��G;�E;JA;�+8;�D&;�{;���:@O��ǃ$�$GĻ�7���������+:�[����Ľ{
��-=��.}������о�\��(��f'�ϕ3�      ���
�����#�޾VD���A���.}�(�D�ht���ڽ�!��\����\�ļ�
v�?��̿���Iɺ�R�9���:(;�-;��;;��B;cIF;��G;fH;��H;�H;)�H;��H;`�H;��H;W�H;��H;��H;d�H;��H;��H;Y�H;��H;`�H;��H;.�H;�H;��H;fH;��G;fIF;��B;��;;�-;(;���:�R�9�Iɺʿ��>���
v�[�ļ���\��!����ڽht�(�D��.}��A��VD��#�޾�����
�      �iþUD��7o�����������i��-=�ht�����R��hys�z +����y񗼕(;�.�ѻ�s@���!��3j:�P�:��;�D3;0�>;FD;��F;�	H;8|H;��H;o�H;2�H;��H;��H;��H;�H;+�H;k�H;��H;j�H;,�H;�H;��H;��H;��H;4�H;q�H;��H;7|H;�	H;��F;FD;3�>;�D3;��;�P�:�3j:�!��s@�,�ѻ�(;�x����z +�hys��R�����ht��-=��i���������7o��UD��      �(��Fl���.}�:ce�zPH���(�{
���ڽ�R�� �{�C�6�� �-p��`�`�Ψ��,��TIҺ�K^9���:գ;�~(;)�8;�IA;|E;	jG;�=H;?�H;ҬH;�H;[�H;"�H;e�H;��H;��H;��H;��H;H�H;��H;��H;��H;��H;f�H;#�H;_�H;�H;ԬH;?�H;�=H;jG;�{E;�IA;/�8;�~(;ޣ;���: L^9BIҺ�,��ͨ�^�`�-p��� �C�6���{��R����ڽ{
���(�zPH�:ce��.}�Fl��      �-=�A�9��k/�0�����~��Ľ�!��iys�C�6�%#��ɺ��vz����D^��p�$��$�r:���:��;�Y1;�H=;&xC;$wF;�G;�eH;E�H;�H;��H;�H;M�H;��H;��H;��H;`�H;u�H;��H;v�H;c�H;��H;��H;��H;N�H;��H;��H;��H;H�H;�eH;�G;"wF;)xC;�H=;�Y1;��;���:8�r:�~�k�$�A^������vz��ɺ�$#�C�6�hys��!����Ľ~���0���k/�A�9�      �` �.�����ڽ�b��ur��[��\�z +�� ��ɺ�@��O*�Hͻ�5R� ǅ���:��:|�;�);�t8;`�@;T*E;i8G;:$H;>�H;>�H;�H;�H;��H;h�H;]�H;��H;J�H;��H;��H;�H;��H;��H;N�H;��H;^�H;n�H;��H;&�H;�H;>�H;;�H;>$H;i8G;\*E;d�@;�t8;�);��;$��:М:ǅ��5R�Dͻ�O*�?��ɺ�� �y +�\�[��ur���b����ڽ���.��      A���R��$ڟ�����C���_�+:�������-p���vz��O*��4ֻk�:�����09�:1;H� ;�D3;B�=;��C;�kF;��G;�\H;��H;K�H;��H;4�H;��H;s�H;��H;��H;�H;��H;T�H;��H;T�H;��H;�H;��H;��H;z�H;��H;>�H; �H;L�H;��H;�\H;��G;�kF;��C;E�=;�D3;Q� ;1;4�:�09,���k��4ֻ�O*��vz�-p����輤��+:��_� C������$ڟ��R��      �_� \�!<Q�g@�� +��5�����[�ļx�_�`����Hͻk�Iɺ �6�/�:�P�:!�;�d.;@�:;�A;#|E;tNG;?'H;��H;ĥH;X�H;��H;!�H;F�H;U�H;0�H;��H;��H;	�H;��H;��H;��H;	�H;��H;��H;3�H;\�H;O�H;*�H;��H;[�H;��H;��H;@'H;}NG;)|E; �A;L�:;�d.;%�;�P�:7�: �6�Iɺk�Eͻ���^�`�w�Z�ļ�����5�� +�g@�!<Q�\�      0]� �-#�������ټ�ɺ������
v��(;�Ψ�B^���5R�>��� �6����:���:�;"�*;�+8;|!@;Q�D;]�F;��G;�eH;{�H;��H;��H;��H;��H;��H;�H;o�H;��H;b�H;z�H;+�H;V�H;+�H;z�H;e�H;��H;p�H;!�H;��H;��H;��H;��H;��H;�H;�eH;��G;a�F;U�D;�!@;�+8;�*;��;���:���: �6�0����5R�>^��Ψ��(;��
v������ɺ���ټ����.#� �      ,p��dx��ע��R��)��r�`���7�<��.�ѻ�,��k�$�ǅ���095�:���:|;�~(;�Z6;|�>;ǨC;�HF;נG;�DH;D�H;��H;��H;�H;&�H;�H;��H;��H;��H;��H;�H;��H;��H;��H;��H;��H;�H;��H;��H;��H;��H;�H;)�H;�H;��H;��H;D�H;�DH;۠G;�HF;ϨC;��>;�Z6;�~(;~;���:5�:��09ǅ�g�$��,��*�ѻ<�� �7�o�`�*���R��ע�cx��      ��I�/�E��(;��O*����<��"GĻƿ���s@�<IҺ�~�:.�:�P�:��;�~(;�5;�>;1C;+�E;tcG;6$H;�{H;5�H;�H;��H;��H;7�H;��H;�H;T�H;��H;O�H;��H;A�H;��H;��H;��H;=�H;��H;J�H;��H;Z�H; �H;��H;:�H;��H;��H;�H;7�H;�{H;8$H;wcG;4�E;6C;�>;
�5;�~(;��;�P�:.�:Ȝ:�~�>IҺ�s@�ƿ��$GĻ�<�����O*��(;�.�E�      F�ѻ�ͻ/���CG��꿐�f�d���$��Iɺ��!�PL^90�r:��:�0;!�;�*;�Z6;�>;7�B;��E;�8G;�	H;�mH;�H;F�H;��H;a�H;��H;��H;E�H;��H;�H;t�H;��H;��H;��H;�H;!�H;�H;��H;��H;��H;t�H;��H;�H;G�H;��H;��H;^�H;��H;C�H;�H;�mH;�	H;�8G;��E;5�B;�>;�Z6; �*;"�;1;��:L�r:@L^9ԅ!��IɺÃ$�d�d�濐�FG��*����ͻ      s�)�/�$�A�����,���H�\��N��S�94j:���:��:~�;O� ;�d.;�+8;�>;1C;��E;�)G;��G;dH;|�H;��H;Y�H;��H;5�H;��H;��H;��H;��H;��H;H�H;{�H;`�H; �H;7�H;I�H;4�H;��H;]�H;x�H;F�H;��H;��H;��H;��H;��H;/�H;��H;\�H;��H;�H;dH;��G;�)G;��E;7C;|�>;�+8;�d.;Q� ;�;	��:���:4j:S�9O��`�\�"���*���@��1�$�      ��R�� � a7��D^9X�:D�X:Ϳ�:���:�P�:ޣ;��;�);�D3;G�:;�!@;ΨC;/�E;�8G;��G;�`H;l�H;�H;�H;u�H;7�H;0�H;J�H;[�H;��H;��H;��H;�H;��H;��H;0�H;n�H;c�H;h�H;,�H;��H;��H;	�H;��H;��H;��H;]�H;H�H;-�H;<�H;x�H;�H;�H;r�H;�`H;��G;�8G;1�E;˨C;�!@;E�:;�D3;�);��;ޣ;�P�:���:ǿ�:`�X:d�:`C^9 k7�` �      ��:���:��:��:��:�P�:�{;(;��;�~(;�Y1;�t8;A�=;�A;T�D;�HF;tcG;�	H;dH;j�H;D�H;ѶH;.�H;��H;��H;:�H;G�H;��H; �H;��H;|�H;��H;U�H;��H;H�H;��H;��H;��H;H�H;��H;R�H;��H;~�H;��H;�H;��H;B�H;7�H;��H;��H;,�H;նH;I�H;k�H;dH;�	H;wcG;�HF;T�D;�A;A�=;�t8;�Y1;�~(;��;(;�{;�P�:��:��:��:���:      (�
;C�;��;;<�;�`;D&;�-;�D3;/�8;I=;_�@;��C;)|E;`�F;ܠG;:$H; nH;��H;�H;ضH;��H;6�H;�H;d�H;��H;��H;r�H;i�H;�H;�H;��H;��H;�H;e�H;��H;��H;��H;c�H;�H;��H;��H; �H;�H;f�H;r�H;��H;��H;i�H;�H;2�H;��H;ٶH;�H;��H;�mH;;$H;۠G;a�F;$|E;��C;b�@;I=;,�8;�D3;�-;�D&;�`;Q�;;�;8�;      �*;D�*;e,;bd.;�Y1;α4;�+8;��;;7�>;�IA;-xC;Z*E;�kF;�NG;��G;�DH;�{H;�H;��H;�H;.�H;5�H;��H;��H;��H;\�H;�H;��H;��H;��H;��H;m�H;��H;;�H;��H;��H;��H;��H;��H;;�H;��H;k�H;��H;��H;��H;��H;�H;^�H;��H;��H;��H;6�H;0�H;�H;��H;�H;�{H;�DH;��G;}NG;�kF;[*E;-xC;�IA;8�>;��;;�+8;Ǳ4;�Y1;dd.;c,;-�*;      �:;8�:;y�;;��<;�>;��?;JA;��B;FD;|E;"wF;i8G;��G;C'H;�eH;K�H;8�H;M�H;]�H;u�H;��H;�H;��H;��H;�H;��H;��H;3�H;v�H;o�H;�H;��H;�H;]�H;�H;��H;��H;��H;|�H;]�H;�H;��H;�H;o�H;p�H;3�H;��H;��H;�H;��H;��H;�H;��H;t�H;\�H;E�H;7�H;H�H;�eH;>'H;��G;g8G;%wF;�{E;FD;��B;JA;��?;>;��<;y�;;-�:;      ɣB;�B;�C;��C;�0D;��D;��E;cIF;��F;jG;�G;B$H;�\H;�H;��H;��H;"�H;��H;��H;E�H;��H;j�H;��H; �H;��H;p�H;��H;C�H;*�H;��H;��H;��H;,�H;q�H;��H;��H;��H;��H;��H;t�H;)�H;��H;��H;��H;&�H;B�H;��H;q�H;��H;�H;��H;m�H;��H;?�H;��H;��H;$�H;��H;��H;��H;�\H;D$H;!�G;jG;��F;eIF;��E;��D;�0D;��C;�C;�B;      �HF;�TF;�vF;�F;n�F;x8G;��G;��G;�	H;�=H;�eH;?�H;��H;˥H;��H;��H;��H;e�H;3�H;-�H;;�H;��H;^�H;��H;m�H;��H;"�H;�H;��H;D�H;��H;!�H;4�H;o�H;��H;��H;��H;��H;��H;n�H;3�H;�H;��H;C�H;��H;�H;�H;��H;q�H;��H;Z�H;��H;;�H;,�H;2�H;a�H;��H;��H;��H;ƥH;��H;>�H;�eH;�=H;�	H;��G;��G;k8G;��F;��F;�vF;�TF;      5�G;��G;
�G;��G;SH;g0H;~LH;fH;4|H;A�H;H�H;=�H;G�H;Z�H;��H;�H;��H;��H;��H;M�H;N�H;��H;�H;��H;��H; �H;��H;��H;O�H;��H;��H;0�H;O�H;r�H;��H;��H;��H;}�H;��H;t�H;N�H;-�H;��H;��H;J�H;��H;��H;'�H;��H;��H;�H;��H;K�H;I�H;��H;��H;��H;�H;��H;S�H;E�H;=�H;H�H;>�H;5|H;fH;wLH;_0H;hH;��G;�G;��G;      �lH;%nH;�rH;�yH;:�H;��H;�H;��H;��H;۬H;��H;��H;��H;��H;��H;*�H;:�H;��H;��H;]�H;��H;r�H;��H;7�H;?�H;�H;��H;3�H;��H;��H;�H;:�H;^�H;c�H;|�H;��H;}�H;��H;{�H;c�H;\�H;4�H;�H;��H;��H;3�H;��H;�H;B�H;3�H;��H;p�H;��H;Z�H;��H;��H;:�H;*�H;��H;��H;��H;��H;��H;֬H;��H;��H;�H;��H;C�H;�yH;�rH;nH;      �H;��H;�H;��H;��H;f�H;x�H;�H;f�H;�H;��H;#�H;;�H;&�H;��H;�H;��H;N�H;��H;��H;*�H;g�H;��H;w�H;&�H;��H;H�H;��H;��H;�H;&�H;I�H;^�H;c�H;a�H;m�H;j�H;h�H;`�H;d�H;^�H;E�H;)�H;�H;��H;��H;D�H;��H;'�H;r�H;��H;f�H;&�H;��H;��H;I�H;��H;�H;��H;#�H;9�H;!�H;��H;�H;j�H;�H;u�H;b�H;��H;��H;�H;��H;      q�H;��H;��H;�H;
�H;n�H;1�H;*�H;2�H;_�H;��H;��H;��H;Q�H;��H;��H;!�H;�H;��H;��H;��H;�H;��H;p�H;��H;<�H;��H;��H;�H;"�H;>�H;A�H;O�H;a�H;K�H;Y�H;n�H;W�H;G�H;a�H;K�H;>�H;=�H;�H;	�H;��H;��H;A�H;��H;l�H;��H;�H;��H;��H;��H;��H;!�H;��H;��H;N�H;��H;��H;��H;`�H;2�H;*�H;2�H;j�H;
�H;�H;��H;��H;      ?�H;|�H;�H;"�H;W�H; �H;��H;��H;��H;(�H;S�H;r�H;}�H;^�H;#�H;��H;^�H;��H;��H;��H;��H;#�H;��H;�H;��H;��H;��H;
�H;-�H;D�H;S�H;L�H;>�H;=�H;^�H;L�H;,�H;I�H;Z�H;@�H;=�H;L�H;S�H;B�H;(�H;�H;��H;��H;��H;�H;��H;!�H;��H;��H;��H;��H;`�H;��H;#�H;^�H;{�H;r�H;Q�H;(�H;��H;��H;��H;��H;e�H; �H;�H;|�H;      ��H;��H;��H;��H;��H;��H;�H;b�H;��H;f�H;��H;d�H;��H;7�H;r�H;��H;��H;y�H;M�H;�H;��H;��H;n�H;��H;��H;�H;,�H;:�H;I�H;B�H;G�H;S�H;;�H;4�H;H�H;)�H;"�H;,�H;E�H;6�H;=�H;S�H;E�H;A�H;D�H;6�H;)�H;!�H;��H;��H;r�H;��H;��H;�H;L�H;{�H;��H;��H;r�H;7�H;��H;b�H;��H;f�H;��H;c�H;�H;��H;��H;��H;��H;��H;      ��H;��H;�H;l�H;�H;��H;��H;��H;��H;��H;��H;�H;��H;��H;��H;��H;S�H; �H;�H;��H;_�H;��H;��H;�H;,�H;0�H;O�H;d�H;e�H;R�H;9�H;=�H;D�H;;�H;�H;�H;K�H;�H;�H;>�H;A�H;@�H;7�H;N�H;^�H;^�H;L�H;2�H;0�H;�H;��H;��H;Y�H;��H;�H;�H;T�H;��H;��H;��H;��H;�H;��H;��H;��H;��H;��H;��H;�H;d�H;�H;��H;      F�H;X�H;��H;��H;c�H;��H;��H;Y�H;�H;��H;��H;T�H;�H;��H;h�H;�H;��H;��H;b�H;��H;��H;!�H;:�H;W�H;o�H;k�H;n�H;d�H;d�H;d�H;7�H;7�H;=�H;%�H;�H;�H;%�H;�H;�H;&�H;=�H;7�H;7�H;a�H;^�H;`�H;m�H;m�H;t�H;V�H;>�H;�H;��H;��H;b�H;�H;��H;�H;h�H;��H;�H;T�H;��H;��H;�H;Z�H;��H;��H;j�H;��H;��H;b�H;      u�H;��H;��H;��H;V�H;��H;!�H;��H;0�H;��H;k�H;��H;��H;�H;��H;��H;F�H;��H;��H;2�H;K�H;d�H;��H;r�H;��H;��H;��H;|�H;d�H;N�H;V�H;I�H;�H;�H;!�H;�H;��H;�H;�H;�H;�H;L�H;U�H;H�H;]�H;v�H;��H;��H;��H;r�H;��H;^�H;E�H;*�H;��H;��H;G�H;��H;��H;�H;��H;��H;n�H;��H;5�H;��H;#�H;��H;W�H;��H;��H;��H;      �H;�H;J�H;~�H;��H;�H;��H;��H;k�H;��H;|�H;��H;U�H;��H;,�H;��H;��H;�H;6�H;k�H;��H;��H;��H;��H;��H;��H;�H;��H;n�H;]�H;H�H;-�H;!�H;�H;�H;�H;�H;�H;�H;�H;!�H;0�H;G�H;Y�H;j�H;��H;}�H;��H;��H;��H;��H;��H;��H;g�H;6�H;�H;��H;��H;+�H;��H;U�H;��H;~�H;��H;n�H;��H;��H;�H;��H;~�H;I�H;+�H;      ��H;��H;��H;�H;\�H;��H;�H;h�H;��H;I�H;��H;'�H;��H;�H;_�H;��H;��H;(�H;N�H;k�H;��H;��H;��H;��H;��H;��H;��H;��H;o�H;u�H;)�H;&�H;N�H;"�H;��H;�H;��H;�H;��H;#�H;P�H;)�H;)�H;q�H;h�H;��H;��H;��H;��H;��H;��H;��H;��H;e�H;L�H;)�H;��H;��H;]�H;�H;��H;'�H;��H;J�H;��H;j�H;!�H;��H;_�H;�H;��H;��H;      �H;!�H;D�H;�H;��H;�H;��H;��H;k�H;��H;z�H;��H;W�H;��H;,�H;��H;��H;�H;6�H;k�H;��H;��H;��H;��H;��H;��H;�H;��H;o�H;\�H;H�H;/�H;"�H;�H;�H;�H;�H;�H;�H;�H;!�H;0�H;G�H;W�H;j�H;��H;}�H;��H;��H;��H;��H;��H;��H;g�H;6�H;�H;��H;��H;+�H;��H;W�H;��H;~�H;��H;n�H;��H;��H;�H;��H;��H;L�H;'�H;      m�H;��H;��H;��H;V�H;��H;!�H;��H;0�H;��H;k�H;��H;��H;�H;��H;��H;D�H;��H; �H;2�H;N�H;d�H;��H;r�H;��H;��H;��H;{�H;d�H;K�H;U�H;I�H;�H;�H;#�H;�H;��H;�H;#�H;�H;!�H;I�H;U�H;G�H;]�H;u�H;��H;��H;��H;q�H;��H;`�H;D�H;,�H;��H;��H;G�H;��H;�H;�H;��H;��H;k�H;��H;3�H;��H;'�H;��H;Z�H;��H;��H;��H;      F�H;W�H;��H;��H;e�H;��H;��H;\�H;�H;��H;��H;R�H;�H;��H;i�H;�H;��H;�H;c�H;��H;��H;#�H;:�H;Y�H;t�H;k�H;o�H;d�H;e�H;d�H;7�H;7�H;=�H;%�H;�H;�H;%�H;�H;�H;%�H;>�H;7�H;6�H;`�H;\�H;`�H;m�H;n�H;q�H;S�H;>�H;!�H;��H;��H;c�H;�H;��H;�H;i�H;��H;�H;R�H;��H;��H;�H;]�H;��H;��H;l�H;��H;��H;W�H;      ��H;��H;�H;g�H;�H;��H;��H;��H;��H;��H;��H;�H;��H;��H;��H;��H;S�H;�H;�H;��H;_�H;��H;��H;�H;0�H;-�H;O�H;d�H;e�H;R�H;7�H;:�H;B�H;:�H;�H;�H;K�H;�H;�H;=�H;@�H;>�H;7�H;L�H;\�H;]�H;K�H;2�H;-�H;�H;��H;��H;V�H;��H;�H; �H;S�H;��H;��H;��H;��H;�H;��H;��H;��H;��H;��H;��H;�H;o�H;�H;��H;      z�H;��H;��H;��H;��H;��H;�H;d�H;��H;f�H;��H;d�H;��H;9�H;u�H;��H;��H;|�H;M�H;�H;��H;��H;n�H;��H;��H;�H;*�H;:�H;L�H;A�H;E�H;R�H;;�H;3�H;H�H;(�H;"�H;,�H;E�H;6�H;;�H;S�H;D�H;@�H;D�H;4�H;(�H;�H;��H;��H;t�H;��H;��H;�H;L�H;y�H;��H;��H;r�H;7�H;��H;b�H;��H;h�H;��H;d�H;�H;��H;��H;��H;��H;��H;      5�H;�H;�H;�H;^�H; �H;��H;��H;��H;(�H;S�H;u�H;{�H;`�H;&�H;��H;`�H;��H;��H;��H;��H;#�H;��H;�H;��H;��H;��H;
�H;/�H;B�H;R�H;L�H;=�H;=�H;^�H;K�H;,�H;K�H;Z�H;@�H;=�H;L�H;R�H;@�H;&�H;�H;��H;��H;��H;�H;��H;#�H;��H;��H;��H;��H;a�H;��H;$�H;^�H;z�H;r�H;Q�H;&�H;��H;��H;��H;��H;j�H;&�H;�H;~�H;      ��H;��H;��H;�H;��H;z�H;2�H;1�H;6�H;`�H;��H;��H;��H;O�H;��H;��H;!�H;�H;��H;��H;��H;�H;��H;m�H;��H;:�H;��H;��H;�H;!�H;=�H;@�H;K�H;a�H;I�H;W�H;n�H;W�H;H�H;a�H;L�H;@�H;=�H;�H;�H;��H;��H;@�H;��H;i�H;��H;�H;��H;��H;��H;��H;!�H;��H;��H;N�H;��H;��H;��H;`�H;3�H;0�H;4�H;j�H;�H; �H;��H;��H;      ��H;��H;'�H;��H;��H;m�H;u�H;�H;p�H;�H;��H;%�H;;�H;(�H;��H;�H;��H;N�H;��H;��H;+�H;i�H;��H;w�H;(�H;��H;F�H;��H;��H;
�H;(�H;I�H;]�H;c�H;`�H;j�H;j�H;j�H;`�H;c�H;^�H;I�H;)�H;
�H;��H;��H;C�H;��H;$�H;o�H;��H;i�H;&�H;��H;��H;I�H;��H;�H;��H;&�H;:�H;�H;��H;�H;m�H;�H;{�H;g�H;��H;��H;'�H;|�H;      �lH;nH;�rH;�yH;3�H;��H;�H;��H;��H;٬H;��H;��H;��H;��H;��H;*�H;:�H;��H;��H;]�H;��H;s�H;��H;6�H;B�H;�H;��H;3�H;��H;��H;�H;:�H;]�H;a�H;{�H;��H;�H;��H;{�H;d�H;`�H;7�H;�H;��H;��H;/�H;��H;�H;<�H;2�H;��H;p�H;��H;Z�H;��H;��H;:�H;*�H;��H;��H;��H;�H;��H;֬H;��H;��H;�H;��H;F�H;�yH;�rH;nH;      '�G;��G;�G;��G;aH;n0H;~LH;fH;5|H;>�H;F�H;@�H;E�H;X�H;��H;�H;��H;��H;��H;I�H;O�H;��H;�H;��H;��H;�H;��H;��H;O�H;��H;��H;0�H;N�H;t�H;��H;��H;��H;��H;��H;u�H;O�H;0�H;��H;��H;H�H;��H;��H;%�H;��H;��H;�H;��H;I�H;L�H;��H;��H;��H;�H;��H;T�H;D�H;;�H;F�H;<�H;4|H;fH;�LH;i0H;iH;��G;�G;��G;      �HF;�TF;wF;�F;u�F;�8G;��G;��G;�	H;�=H;�eH;B�H;��H;ȥH;��H;��H;��H;g�H;3�H;-�H;@�H;��H;Z�H;��H;q�H;��H; �H;�H;��H;A�H;��H;!�H;3�H;q�H;��H;��H;��H;��H;��H;o�H;3�H;!�H;��H;A�H;��H;�H; �H;��H;o�H;��H;^�H;��H;;�H;-�H;3�H;`�H;��H;��H;��H;ƥH;��H;<�H; fH;�=H;�	H;��G;��G;p8G;��F;�F;�vF;�TF;      ȣB;�B;�C;��C;�0D;��D;��E;eIF;��F;jG;!�G;D$H;�\H;�H;��H;��H;"�H;��H;��H;A�H;��H;m�H;��H;�H;��H;l�H;��H;C�H;*�H;��H;��H;��H;*�H;r�H;��H;��H;��H;��H;��H;t�H;,�H;��H;��H;��H;$�H;?�H;��H;q�H;��H;�H;��H;m�H;��H;A�H;��H;��H;$�H;��H;��H; �H;�\H;A$H;�G;jG;��F;eIF;��E;��D;�0D;��C;�C;�B;      ��:;�:;v�;;��<;�>;§?;JA;��B;FD; |E;%wF;j8G;��G;@'H;�eH;K�H;8�H;M�H;\�H;t�H;��H;�H;��H;��H;�H;��H;��H;4�H;v�H;m�H;�H;��H;�H;]�H;|�H;��H;��H;��H;|�H;\�H;�H;��H;�H;o�H;r�H;0�H;��H;��H;�H;��H;��H;�H;��H;v�H;]�H;G�H;8�H;I�H;�eH;?'H;��G;f8G;$wF;�{E;FD;��B;JA;��?;>;�<;x�;;�:;      �*;;�*;^,;ld.;�Y1;Ǳ4;�+8;��;;;�>;�IA;)xC;[*E;�kF;~NG;��G;�DH;�{H;�H;��H;�H;/�H;6�H;��H;��H;��H;W�H;�H;��H;��H;��H;��H;n�H;��H;;�H;��H;��H;��H;��H;��H;:�H;��H;n�H;��H;��H;��H;��H;�H;^�H;��H;��H;��H;6�H;2�H;�H;��H;�H;�{H;�DH;��G;{NG;�kF;W*E;)xC;�IA;:�>;��;;�+8;ȱ4;�Y1;nd.;],;&�*;      &�
;F�;��;;=�;�`;�D&;�-;�D3;,�8;I=;d�@;��C;&|E;d�F;ޠG;:$H; nH;�H;�H;ضH;��H;2�H;�H;j�H;��H;��H;r�H;i�H;�H;�H;��H;��H;�H;c�H;��H;��H;��H;a�H;�H;��H;��H;!�H;�H;g�H;p�H;��H;��H;f�H; �H;6�H;��H;ضH;�H;�H;�mH;:$H;۠G;a�F;&|E;��C;`�@;I=;+�8;�D3;�-;|D&;�`;S�;�;�;9�;      ��:ݍ�:��:��:��:�P�:�{;(;��;�~(;�Y1;�t8;B�=;�A;X�D;�HF;vcG;�	H;dH;k�H;E�H;ֶH;,�H;��H;��H;4�H;A�H;��H; �H;��H;~�H;��H;R�H;��H;G�H;��H;��H;��H;G�H;��H;V�H;��H;��H;��H;�H;��H;E�H;7�H;��H;��H;.�H;ӶH;G�H;l�H;dH;�	H;vcG;�HF;U�D;�A;A�=;�t8;�Y1;�~(;��;(;�{;�P�:&��:$��:��:���:      @�R�@ � d7�pD^9X�:d�X:ѿ�:���:�P�:ޣ;��;�);�D3;F�:;�!@;ϨC;1�E;�8G;��G;�`H;o�H;�H;�H;x�H;<�H;,�H;E�H;]�H;��H;��H;��H;�H;��H;��H;/�H;j�H;d�H;k�H;,�H;��H;��H;�H;��H;��H;��H;[�H;J�H;0�H;8�H;y�H;�H;�H;o�H;�`H;��G;�8G;.�E;̨C;�!@;C�:;�D3;�);��;٣;�P�:���:ÿ�:<�X:d�:�C^9 d7�� �      p�)�.�$�>�����.���D�\�O��S�94j:���:��:�;Q� ;�d.;�+8;��>;4C;��E;�)G;��G;dH;�H;��H;[�H;��H;0�H;��H;��H;��H;��H;��H;H�H;{�H;`�H;��H;6�H;I�H;6�H;��H;]�H;{�H;H�H;��H;��H;��H;��H;��H;2�H;��H;]�H;��H;|�H;dH;��G;�)G;��E;1C;|�>;�+8;�d.;N� ;~�;��:���:4j:S�9 O��P�\�,������E��*�$�      M�ѻ�ͻ/���FG��俐�[�d���$��Iɺ̅!�PL^9H�r:��:1;"�;$�*;�Z6;�>;7�B;��E;�8G;�	H;�mH;�H;G�H;��H;a�H;��H;��H;H�H;��H;��H;u�H;��H;��H;��H;�H;"�H;�H;��H;��H;��H;r�H;��H;�H;G�H;��H;��H;`�H;��H;E�H;�H;�mH;�	H;�8G;��E;4�B;�>;�Z6;"�*;�; 1;��:L�r: L^9؅!��Iɺ��$�`�d�濐�GG��3����ͻ      ��I�0�E��(;��O*����<��!GĻƿ���s@�:IҺ�~�М:.�:�P�:��;�~(;	�5;�>;3C;/�E;ycG;8$H;�{H;8�H;�H;��H;��H;9�H;��H;�H;X�H;��H;O�H;��H;@�H;��H;��H;��H;?�H;��H;J�H;��H;Z�H;�H;��H;7�H;��H;��H;�H;7�H;�{H;7$H;scG;1�E;0C;�>;�5;�~(;��;�P�:.�:��:�~�@IҺ�s@�ƿ��#GĻ�<�����O*��(;�/�E�      ,p��dx��ע��R��(��o�`���7�;��*�ѻ�,��g�$�ǅ���095�:���:�;�~(;�Z6;~�>;˨C;�HF;۠G;�DH;I�H;��H;��H;�H;(�H;�H;��H;��H;��H;��H;�H;��H;��H;��H;��H;��H;�H;��H;��H;��H;��H;�H;(�H;	�H;��H;��H;E�H;�DH;ؠG;�HF;̨C;y�>;�Z6;�~(;|;���:1�:��09ǅ�i�$��,��+�ѻ<���7�p�`�*���R��ע�dx��      0]� �.#�������ټ�ɺ������
v��(;�ͨ�?^���5R�4��� �6����:���:��; �*;�+8;�!@;X�D;a�F;��G;�eH;��H;��H;��H;��H;��H;��H; �H;r�H;��H;g�H;{�H;)�H;X�H;)�H;x�H;d�H;��H;n�H;�H;��H;��H;��H;��H;��H;}�H;�eH;��G;`�F;O�D;�!@;�+8;�*;�;���:���: �6�:����5R�@^��Ψ��(;��
v������ɺ���ټ����.#� �      �_�\�!<Q� g@�� +��5�����Z�ļw�^�`����Dͻk�Iɺ �6�?�:�P�:"�;�d.;F�:;$�A;'|E;}NG;E'H;�H;ȥH;X�H;��H;&�H;K�H;\�H;3�H;��H;��H;�H;��H;��H;��H;�H;��H;��H;0�H;W�H;M�H;(�H;��H;V�H;ĥH;��H;C'H;~NG;$|E;�A;G�:;�d.;!�;�P�:5�: �6�Iɺk�Fͻ���^�`�x�Z�ļ�����5�� +� g@�!<Q�\�      A���R��$ڟ�����C���_�+:�������,p���vz��O*��4ֻk�*����09.�:1;N� ;�D3;I�=;��C;�kF;��G;�\H;��H;H�H;��H;=�H;��H;x�H;��H;��H;
�H;��H;T�H;��H;T�H;��H;�H;��H;��H;v�H;��H;=�H;��H;G�H;��H;�\H;��G;�kF;��C;>�=;�D3;J� ;1;(�:��090���k��4ֻ�O*��vz�-p����輤��+:��_� C������$ڟ��R��      �` �.�����ڽ�b��ur��[��\�y +�� ��ɺ�?��O*�Dͻ�5R�ǅ���:��:��;�);�t8;c�@;\*E;m8G;A$H;>�H;=�H;�H;"�H;��H;o�H;`�H;�H;N�H;��H;��H;�H;��H;��H;M�H;��H;[�H;k�H;��H;%�H;�H;:�H;<�H;;$H;k8G;[*E;b�@;�t8;�);|�;��:��:ǅ��5R�Hͻ�O*�@��ɺ�� �z +�\�[��ur���b����ڽ���.��      �-=�A�9��k/�0�����~��Ľ�!��hys�C�6�$#��ɺ��vz����@^��k�$��~�,�r:���:��;�Y1;�H=;+xC;%wF;�G;�eH;B�H;�H;��H;��H;P�H;��H;��H;��H;a�H;w�H;��H;v�H;a�H;��H;��H;��H;M�H;��H;��H;��H;B�H;�eH;�G;%wF;)xC;�H=;�Y1;��;���:,�r:�~�o�$�B^������vz��ɺ�%#�C�6�hys��!����Ľ~���0���k/�A�9�      �(��Fl���.}�:ce�zPH���(�{
���ڽ�R����{�C�6�� �-p��_�`�ͨ��,��HIҺ L^9���:ۣ;�~(;,�8;�IA;|E;jG;�=H;>�H;ҬH;�H;]�H;%�H;e�H;��H;��H;��H;��H;I�H;��H;��H;��H;��H;c�H;"�H;\�H;�H;ԬH;<�H;�=H;	jG;|E;�IA;+�8;�~(;ۣ;���:�K^9HIҺ�,��Ψ�`�`�-p��� �C�6���{��R����ڽ{
���(�zPH�:ce��.}�Fl��      �iþUD��7o�����������i��-=�ht�����R��hys�z +����x񗼔(;�+�ѻ�s@��!��3j:�P�:��;�D3;4�>;FD;��F;�	H;7|H;��H;q�H;3�H;��H;��H;��H;�H;+�H;k�H;��H;j�H;,�H;�H;��H;��H;��H;3�H;s�H;��H;7|H;�	H;��F;FD;3�>;�D3;��;�P�:�3j:��!��s@�-�ѻ�(;�y����z +�hys��R�����ht��-=��i���������7o��UD��      ���
�����#�޾VD���A���.}�(�D�ht���ڽ�!��\����[�ļ�
v�>��ʿ���Iɺ�R�9���:(;�-;��;;��B;hIF;��G;fH;��H;�H;*�H;��H;b�H;��H;Z�H;��H;��H;e�H;��H;��H;V�H;��H;`�H;��H;.�H;�H;��H;fH;��G;eIF;��B;��;;�-;(;���:�R�9�Iɺʿ��>���
v�\�ļ���\��!����ڽht�(�D��.}��A��VD��$�޾�����
�      ��7�ϕ3��f'�(��\���о�����.}��-=�{
���Ľ[��+:����������7�%GĻ˃$�@O�����:�{;�D&;�+8;JA;�E;��G;tLH;�H;t�H;1�H;��H;��H;��H;��H;�H;�H;�H;~�H;�H;��H;��H;��H;��H;4�H;v�H;�H;yLH;��G;�E;JA;�+8;�D&;�{;���:HO��ȃ$�$GĻ�7���������+:�[����Ľ{
��-=��.}������о�\��(��f'�ϕ3�      Xo�_Xi��"Y���@�K�#��
��о�A���i���(�~��ur���_��5��ɺ�q�`��<��k�d�p�\�H�X:�P�:�`;ȱ4;��?;��D;r8G;g0H;��H;i�H;r�H;�H;��H;��H;��H;��H;�H;��H;�H;��H;��H;��H;��H;��H;t�H;j�H;��H;i0H;{8G;��D;��?;Ǳ4;�`;�P�:L�X:��\�i�d��<��q�`��ɺ��5��_�ur��~����(��i��A���о�
�K�#���@��"Y�_Xi�      /����������Yo��!J�K�#��\��VD������zPH�����b��C��� +���ټ)����￐����`�:��:@�;�Y1;>;�0D;v�F;[H;A�H;��H;�H;X�H;��H;�H;b�H;B�H;��H;\�H;��H;E�H;\�H;�H;��H;U�H;�H;¨H;E�H;aH;��F;�0D;>;�Y1;C�;��:h�: ���쿐���)����ټ� +� C���b�����zPH�����VD���\��K�#��!J�Yo��������      =^������k���Yo���@�(�$�޾����:ce�0����ڽ���� g@������R���O*�KG�����pC^9$��:�;Yd.;��<;��C;�F;��G;�yH;��H;�H;�H;��H;g�H;��H;��H;~�H;�H;{�H;��H;��H;g�H;��H;�H;�H;��H;�yH;��G;��F;��C;��<;Td.;�;$��:�C^9"���HG���O*��R������ g@�������ڽ0��:ce�����$�޾(���@�Yo�k�������      �aǿ�¿����������"Y��f'�����7o���.}��k/����$ڟ�"<Q�-#�ע��(;�0���>�� k7���:�;o,;��;;�C;�vF;�G;�rH;�H;��H;�H;��H;��H;��H;��H;I�H;��H;D�H;��H;��H;��H;��H;�H;��H;�H;�rH;�G;wF;�C;��;;j,;�;��: d7�>��.����(;�ע�-#�"<Q�$ڟ�����k/��.}�7o�������f'��"Y�����������¿      2�ֿCpѿ�¿������_Xi�ϕ3��
�VD��Fl��B�9��.���R�� \� �ex��2�E��ͻ!�$�p �Ս�:8�;H�*;2�:;�B;�TF;��G;#nH;��H;��H;i�H;��H;��H;X�H;}�H;�H;��H;�H;�H;X�H;��H;��H;d�H;·H;��H;&nH;��G;�TF;�B;/�:;B�*;8�;Ս�:@ �#�$��ͻ2�E�ex�� � \��R���.��A�9�Fl��VD���
�ϕ3�_Xi��������¿Cpѿ      �� $������꿯�ſ�ޞ�%3s��2�>����� j���yHͽƸ����'�B<ͼt�n�h���EQ^�..�h��:jW;^S%;co8;��A;DF;�H;y�H;��H;��H;�H;	�H;!�H;��H;��H;��H;�H;��H;��H;��H;"�H;�H;�H;��H;��H;{�H;�H;DF;��A;bo8;WS%;jW;n��:�-.�FQ^�e���s�n�B<ͼ��'�Ƹ��yHͽ�� j���>����2�%3s��ޞ���ſ������ $�       $�������忇�����cm�V�-�����Qh��Vde�"-�תɽ�v��(�$���ɼ{mj�:���X�0���ņ:dx;�%;0�8;BB;RF;�H;�H;�H;��H;B�H;�H;�H;u�H;��H;��H;�H;��H;��H;u�H;�H;�H;A�H;��H;�H;�H;�H;*RF;CB;.�8;�%;dx;�ņ:��X�8���{mj���ɼ(�$��v��תɽ"-�Vde�Qh������V�-�cm��������忝����      ����������ԿLw�����:�\�"����k��Y0X�����;����w����������]�$���F� ���ɒ:��; �';��9;�oB;�zF;�!H;p�H;��H; �H;n�H;�H;�H;}�H;��H;��H;��H;��H;��H;}�H;�H;�H;k�H;�H;��H;s�H;�!H;�zF;�oB;��9;��';��;�ɒ:����F�"�黬�]����������w��;�����Y0X�k�����"�:�\����Lw���Կ��𿝏�      ������Կp���ޞ�`F�h�C�-E�#�;�I��D���"��f�c�|��֯���J��ѻ֢)��K���:�
;�M*;j�:;�C;ȸF;�8H;*�H;F�H;X�H;��H;�H;�H;}�H;��H;��H;��H;��H;��H;|�H;�H;�H;��H;\�H;J�H;*�H;�8H;иF;�C;i�:;�M*;�
;��:�K�Ӣ)��ѻ��J��֯�|�f�c�"����D��I��#�;-E�h�C�`F��ޞ�p���Կ��      ��ſ���Lw���ޞ�����?�W�5�%�����hɰ��|x�f{+�ұ����J��  �϶��[�1�,���%+��
9��:��;߷-;��<;Z�C;�G;�TH;!�H;��H;��H;��H;(�H;�H;c�H;��H;r�H;��H;n�H;��H;c�H;�H;(�H;��H;��H;��H;$�H;�TH;�G;Z�C;��<;ܷ-;��;��:@ 
9$+�+���[�1�϶���  ��J���ұ�f{+��|x�hɰ�����5�%�?�W������ޞ�Lw�����      �ޞ�������`F�?�W�W�-����?Kɾ�G����O����ƽȸ��΄-���ۼㄼ64�ǐ�϶�]:��:z;z�1;�c>;A�D;u\G;)sH;s�H;4�H;A�H;��H;G�H;	�H;G�H;g�H;Z�H;��H;W�H;h�H;D�H;
�H;K�H;��H;G�H;4�H;v�H;)sH;|\G;B�D;�c>;x�1;z;��: ]:
϶�ǐ�64�ㄼ��ۼ΄-�Ǹ��ƽ�����O��G��?Kɾ���W�-�?�W�`F�������      %3s�cm�:�\�h�C�5�%����TҾj��
 j��C(����]P����[�|������Y�=��kX���<���k:*��:�� ;ҟ5;.R@;2uE;βG;�H;�H;��H;��H;�H;C�H;�H;>�H;K�H;6�H;k�H;3�H;L�H;@�H;�H;D�H;�H;��H;��H;�H;�H;ҲG;5uE;-R@;ҟ5;�� ;$��: �k:|�<�hX�;����Y����|���[�]P����콪C(�
 j�j���TҾ��5�%�h�C�:�\�cm�      �2�V�-�"�-E�����?Kɾj����s�9�5���u㻽�v��	z0��;��+���*����;6��CS�;M�:I�	;l�(;��9;�/B;GDF;H;��H;Z�H;��H;��H;J�H;`�H;��H;�H;�H;�H;7�H;�H;�H;�H;��H;`�H;J�H;��H;��H;Z�H;��H; H;HDF;�/B;�9;p�(;F�	;MM�:�CS�56�����*��+���;�	z0��v��u㻽��8�5���s�j��?Kɾ����-E�"�V�-�      >����������#�;hɰ��G��
 j�8�5��	�ΪɽY����J�s���沼��]�����	x�b	���m:|��:�v;��/;c-=;��C;�F;�HH;z�H;��H;��H;��H;z�H;c�H;��H;��H;��H;��H;�H;��H;��H;��H;��H;f�H;{�H;�H;��H;��H;z�H;�HH;�F;��C;g-=;��/;�v;���:n:\	���	x������]��沼s���J�Y���Ϊɽ�	�8�5�
 j��G��hɰ�"�;��徶���      ��Ph��k���I���|x���O��C(���Ϫɽ����RDX�H��'<ͼ	ㄼ�X!��s���W�0vK���:�y;��#;�H6;R@;�PE;e�G;[�H;��H;�H;��H;z�H;��H;Q�H;��H;��H;��H;��H;��H;��H;��H;��H;��H;R�H;��H;��H;��H;�H;��H;Y�H;k�G;�PE;
R@;�H6;��#;�y;��:�uK��W��s���X!�	ㄼ'<ͼG��RDX�����Ϊɽ���C(���O��|x��I��k��Ph��       j�Vde�Z0X�D�e{+�������u㻽Y���RDX������ۼ̾����;�J>ۻ'X���y��>":���:��;��-;~�;;��B;izF;�H;^�H;U�H;��H;��H;��H;��H;K�H;��H;z�H;p�H;��H;Y�H;��H;r�H;|�H;��H;K�H;��H;��H;��H;��H;W�H;]�H;�H;hzF;��B;��;;��-;��;���:�>":`�y�#X�G>ۻ��;�˾����ۼ���RDX�Y���u㻽��콂��f{+�D�Z0X�Vde�      ��"-������ѱ�ƽ]P���v���J�H����ۼ��e�J������+���rѺ�'
9�M�:��;n $;��5;��?;Z�D;=\G;�eH;��H;��H;��H;��H;��H;��H;2�H;Q�H;9�H;2�H;D�H;�H;D�H;3�H;=�H;R�H;2�H;��H;�H;��H;��H;��H;��H;�eH;=\G;b�D;��?;��5;z $;��;�M�:0(
9�rѺ�+������d�J�����ۼG���J��v��]P��ƽұ轃����"-�      yHͽ֪ɽ�;��"����Ǹ����[�	z0�s��&<ͼ˾��d�J�����j���*� �ڨ�:,b�:1�;��/;wL<;�C; mF;l�G;ءH;��H;��H;��H;�H;/�H;��H;�H;�H;��H;��H;��H;��H;��H;��H;��H;�H;�H;��H;8�H;�H;��H;��H;��H;ޡH;l�G;mF;�C;~L<;��/;8�;,b�:ꨂ:��*��j�����d�J�˾��&<ͼr��	z0���[�Ǹ����"���;��֪ɽ      Ÿ���v����w�f�c��J�τ-�|��;缆沼ㄼ��;������j���5�����>Q:$��:Hi;�M*;`�8;a�@;�PE;�uG;iH;��H;��H;��H;��H;��H;Q�H;��H;��H;��H;��H;��H;��H;�H;��H;��H;��H;��H;��H;��H;\�H;��H; �H;��H;��H;��H;iH;�uG;�PE;d�@;j�8;�M*;Ki;8��:�>Q:x�깪5��j��������;�ㄼ�沼�;�|�΄-��J�g�c���w��v��      ��'�(�$����|��  ���ۼ����+����]��X!�H>ۻ�+���*���깴�>:���:��;�%;ʟ5;s�>;(D;��F;Q!H;�H;'�H;��H;��H;��H;��H;I�H;��H;��H;h�H;m�H;J�H;4�H;Q�H;4�H;I�H;p�H;j�H;��H;��H;Q�H;��H;��H;��H;��H;+�H;�H;U!H;��F;�(D;}�>;Ο5;�%;��;���:��>:��깁*��+��D>ۻ�X!���]��+�������ۼ�  �|����(�$�      ?<ͼ�ɼ�����֯�ζ��ㄼ��Y��*�����s��"X��rѺ��>Q:���:��
;.�#;K�3;nc=;�#C;DF;��G;�H;��H;��H;�H;��H;3�H;��H;C�H;l�H;D�H;�H;2�H;��H;��H;��H;��H;��H;2�H;�H;F�H;s�H;I�H;�H;8�H;��H;�H;��H;��H;�H;��G;DF;�#C;sc=;H�3;2�#;��
;���:�>Q: ��rѺX��s������*���Y�ㄼ϶���֯�����~�ɼ      p�n�ymj���]���J�Z�1�54�8������	x��W�`�y��'
9樂:2��:��;2�#;5�2;�<;HpB;��E;��G;�eH;��H;�H;��H;��H;��H;��H;�H;'�H;�H;��H;��H;��H;��H;��H;��H;��H;��H;��H;��H;��H;�H;+�H;�H;��H;��H;��H;��H;�H;��H;�eH;��G;�E;KpB;��<;8�2;2�#;��;8��:樂:(
9P�y��W��	x����:��44�[�1���J���]�wmj�      Z���4���"���ѻ(���ǐ�_X�26�^	���uK��>":�M�:"b�:Ei;�%;E�3;ۆ<;(0B;��E;O\G;�HH;�H;t�H;;�H;��H;�H;�H;��H;��H;��H;��H;��H;��H;C�H;8�H;8�H;�H;5�H;4�H;C�H;��H;��H;��H;��H;��H;��H;�H;�H;��H;9�H;s�H;#�H;�HH;X\G;��E;&0B;��<;D�3;�%;Hi;&b�:�M�:�>":�uK�N	��06�dX�ǐ�$����ѻ��6���      1Q^�X��F�͢)�++��ζ�`�<��AS�n:��:���:��;5�;�M*;Ο5;qc=;HpB;��E;�JG;*8H;G�H;a�H;��H;�H;_�H;��H;r�H;��H;��H;��H;s�H;[�H;7�H;��H;��H;��H;��H;��H;��H;��H;5�H;Z�H;v�H;��H;��H;��H;n�H;��H;f�H;�H;��H;e�H;M�H;08H;�JG;��E;NpB;nc=;Ο5;�M*;6�;��;���:��:n: BS�p�<��ζ�%+�ڢ)��F�X�       ..�@����깰~K��
9]:�k:?M�:���:�y;��;v $;��/;f�8;|�>;�#C;�E;[\G;/8H;��H;��H;��H;j�H;�H;d�H;0�H;��H;��H;��H;b�H;�H;��H;��H;��H;�H;v�H;]�H;q�H;{�H;��H;��H;��H;�H;a�H;��H;��H;��H;-�H;j�H;�H;i�H;��H;��H;��H;08H;V\G;�E;�#C;~�>;d�8;��/;x $;��;�y;���:CM�:�k:,]:  
9�K����h��      ���:�ņ:�ɒ:��:��:��:"��:E�	;�v;��#;��-;��5;vL<;^�@;(D;DF;��G;�HH;J�H;��H;��H;%�H;��H;:�H;��H;k�H;��H;��H;A�H;�H;��H;��H;U�H;H�H;�H;�H;�H;	�H;�H;G�H;R�H;��H;��H;�H;>�H;��H;��H;i�H;��H;9�H;��H;*�H;��H;��H;J�H;�HH;��G;DF;�(D;]�@;yL<;��5;��-;��#;�v;B�	;*��:ޤ�:��:��:�ɒ:�ņ:      hW;nx;��;�
;��;|;�� ;j�(;��/;�H6;��;;��?;�C;�PE;��F;��G;�eH;%�H;g�H;��H;*�H;��H;�H;��H;>�H;b�H;i�H;I�H;��H;��H;��H;-�H;��H;��H;��H;��H;��H;��H;��H;��H;��H;*�H;��H;��H;��H;I�H;e�H;b�H;E�H;��H;
�H;��H;,�H;��H;e�H;#�H;�eH;��G;��F;�PE;�C;��?;��;;�H6;��/;p�(;�� ;x;��;�
;��;bx;      sS%; �%;��';�M*;շ-;��1;��5;��9;k-=;R@;��B;`�D;mF;�uG;U!H;�H;��H;z�H;��H;j�H;��H;�H;��H;H�H;^�H;W�H;�H;��H;��H;y�H;�H;��H;��H;�H;p�H;Y�H;:�H;U�H;k�H;��H;��H;��H;
�H;y�H;��H;��H;�H;Z�H;b�H;E�H;��H;�H;��H;j�H;��H;v�H;��H;�H;T!H;�uG;mF;b�D;��B;R@;k-=;��9;ܟ5;z�1;�-;�M*;�';��%;      ^o8;4�8;��9;j�:;u�<;�c>;0R@;�/B;��C;�PE;fzF;<\G;i�G;iH;�H;��H;�H;B�H;
�H;�H;;�H;��H;F�H;Q�H;I�H;*�H;��H;��H;S�H;��H;��H;��H;D�H;�H;�H;�H;��H;	�H;�H;�H;C�H;��H;��H;��H;N�H;��H;��H;-�H;L�H;O�H;A�H;��H;;�H;�H;�H;<�H;�H;��H;�H;iH;h�G;<\G;hzF;�PE;��C;�/B;*R@;�c>;��<;e�:;��9;*�8;      ��A;>B;�oB;�C;R�C;P�D;=uE;FDF;�F;i�G;�H;�eH;ޡH;��H;.�H;��H;��H;��H;n�H;q�H;�H;E�H;g�H;S�H;�H;��H;��H;Y�H;��H;��H;_�H;0�H;��H;��H;��H;��H;��H;��H;��H;��H;��H;,�H;b�H;��H;��H;W�H;��H;��H;�H;P�H;b�H;F�H;�H;m�H;m�H;��H;��H;��H;.�H;��H;ޡH;�eH;�H;i�G;�F;FDF;;uE;D�D;]�C;�C;�oB;?B;      	DF;'RF;�zF;ƸF;�G;{\G;ѲG;'H;�HH;]�H;]�H;��H;��H;��H;��H;�H;��H;�H;��H;.�H;o�H;a�H;X�H;0�H;��H;u�H;H�H;��H;��H;R�H;�H;��H;��H;��H;e�H;U�H;b�H;P�H;c�H;��H;��H;��H;�H;R�H;��H;��H;D�H;x�H;��H;-�H;V�H;b�H;n�H;-�H;��H;�H;��H;�H;��H;��H;��H;��H;a�H;]�H;�HH;)H;ͲG;p\G;�G;͸F;�zF;%RF;      �H;�H;�!H;�8H;�TH;)sH;�H;��H;w�H;��H;U�H;��H;��H;��H;��H;��H;��H;�H;u�H;��H;��H;i�H;�H;��H;��H;G�H;��H;x�H;=�H;�H;��H;��H;U�H;6�H;!�H;��H;�H;��H;�H;8�H;T�H;��H;��H;�H;6�H;u�H;��H;K�H;��H;��H;�H;i�H;��H;��H;r�H;�H;��H;��H;��H;��H;��H;��H;U�H;��H;x�H;��H;�H;"sH;�TH;�8H;�!H;�H;      ��H;�H;l�H;4�H;�H;w�H;*�H;Z�H;��H;�H;��H;��H;��H;��H;��H;7�H;��H;��H;��H;��H;��H;I�H;��H;��H;S�H;��H;u�H;J�H;��H;��H;f�H;<�H;�H;��H;��H;��H;��H;��H;��H;��H;�H;9�H;f�H;��H;��H;G�H;p�H;��H;W�H;��H;��H;I�H;��H;��H;��H;��H;��H;7�H;��H;��H;��H;��H;�H;
�H;��H;Z�H;'�H;i�H;$�H;1�H;l�H;��H;      ��H;�H;��H;X�H;��H;0�H;��H;��H;��H;��H;��H;��H;�H;��H;��H;�H;�H;��H;��H;��H;H�H;��H;��H;U�H;��H;��H;5�H;��H;��H;a�H;*�H;��H;��H;��H;��H;��H;u�H;��H;��H;��H;��H;��H;*�H;_�H;��H;��H;/�H;��H;��H;O�H;��H;��H;E�H;��H;��H;��H;�H;�H;��H;��H;�H;��H;��H;��H;��H;��H;��H;,�H;��H;V�H;��H;�H;      ��H;��H;�H;P�H;��H;A�H;��H;��H;��H;}�H;��H; �H;4�H;\�H;L�H;F�H;-�H;��H;��H;e�H;
�H;��H;v�H;��H;��H;J�H;�H;��H;b�H;#�H;��H;��H;��H;~�H;^�H;C�H;7�H;B�H;Z�H;~�H;��H;��H;��H; �H;\�H;��H;��H;O�H;��H;��H;y�H;��H;�H;b�H;��H;��H;-�H;I�H;J�H;Z�H;2�H;��H;��H;��H;��H;��H;��H;=�H;��H;U�H;�H;��H;      #�H;X�H;u�H;��H;��H;��H;$�H;Q�H;~�H;��H;��H;��H;��H;��H;��H;v�H; �H;��H;z�H;%�H;��H;��H;	�H;��H;_�H;�H;��H;l�H;/�H;��H;��H;|�H;p�H;7�H;�H;�H;�H;�H;�H;:�H;o�H;z�H;��H;��H;*�H;h�H;��H;�H;c�H;��H;�H;��H;��H;�H;z�H;��H; �H;v�H;��H;��H;��H;��H;��H;��H;~�H;Q�H;-�H;��H;��H;��H;v�H;X�H;      �H;�H;�H;�H;!�H;?�H;G�H;b�H;i�H;Q�H;M�H;6�H;	�H;��H;��H;G�H;��H;��H;`�H;��H;��H;0�H;��H;��H;.�H;��H;��H;=�H;��H;��H;v�H;Z�H;:�H;�H;��H;��H;��H;��H;��H;�H;;�H;X�H;u�H;��H;��H;;�H;~�H;��H;2�H;��H;��H;0�H;��H;��H;^�H;��H;��H;J�H;��H;��H;�H;5�H;N�H;Q�H;g�H;`�H;M�H;A�H;0�H;�H;�H;�H;      /�H;#�H;)�H;�H;�H; �H;�H;��H;��H;��H;��H;U�H;�H;��H;j�H;�H;��H;��H;;�H;��H;`�H;�H;��H;D�H;��H;��H;U�H;�H;��H;��H;k�H;:�H;��H;��H;��H;��H;��H;��H;��H;��H;��H;<�H;i�H;��H;��H;�H;S�H;��H;��H;F�H;��H;�H;Z�H;��H;<�H;��H;��H;�H;l�H;��H;�H;U�H;��H;��H;��H;��H;�H;��H;�H;�H;2�H;#�H;      |�H;v�H;�H;{�H;d�H;;�H;B�H;�H;��H;��H;��H;@�H;�H;��H;t�H;6�H;��H;H�H;��H;��H;O�H;��H;�H;�H;��H;��H;2�H;��H;��H;��H;1�H;�H;��H;��H;��H;��H;��H;��H;��H;��H;��H;�H;3�H;}�H;��H;��H;1�H;��H;��H;�H;��H;��H;K�H;��H;��H;J�H;��H;8�H;s�H;��H;�H;?�H;��H;��H;��H;�H;H�H;;�H;k�H;{�H;��H;��H;      ��H;��H;��H;��H;��H;c�H;U�H;!�H;��H;��H;z�H;=�H;�H;��H;S�H;��H;��H;8�H;��H;��H;�H;��H;m�H;�H;��H;\�H;�H;��H;��H;`�H;�H;��H;��H;��H;��H;��H;��H;��H;��H;��H;��H;��H;�H;[�H;��H;��H;�H;_�H;��H;�H;p�H;��H;�H;|�H;��H;;�H;��H;��H;P�H;��H;�H;?�H;|�H;��H;��H;!�H;V�H;c�H;��H;��H;��H;��H;      ��H;��H;��H;��H;j�H;V�H;@�H;�H;��H;��H;��H;H�H;��H;��H;5�H;��H;��H;5�H;��H;u�H;�H;��H;R�H;�H;��H;G�H;��H;��H;��H;F�H;�H;��H;��H;��H;��H;��H;��H;��H;��H;��H;��H;��H;�H;B�H;��H;��H;��H;J�H;��H;�H;X�H;��H;�H;q�H;��H;:�H;��H;��H;6�H;��H;��H;G�H;��H;��H;��H;�H;G�H;W�H;m�H;��H;��H;��H;      �H;�H;
�H;��H;��H;��H;r�H;;�H;�H;��H;c�H;!�H;��H;��H;Z�H;��H;��H;�H;��H;d�H;�H;��H;<�H;��H;��H;[�H;	�H;��H;z�H;<�H;�H;��H;��H;��H;��H;��H;y�H;��H;��H;��H;��H;��H;�H;8�H;u�H;��H;	�H;^�H;��H;��H;?�H;��H;�H;`�H;��H;�H;��H;��H;Z�H;��H;��H; �H;g�H;��H;	�H;=�H;y�H;��H;��H;��H;
�H;�H;      ��H;��H;��H;��H;k�H;Z�H;@�H;�H;��H;��H;��H;H�H;��H;��H;6�H;��H;��H;5�H;��H;u�H;�H;��H;R�H;�H;��H;G�H;��H;��H;��H;E�H;�H;��H;��H;��H;��H;��H;��H;��H;��H;��H;��H;��H;�H;A�H;��H;��H;��H;L�H;��H;�H;X�H;��H;�H;q�H;��H;:�H;��H;��H;6�H;��H;��H;H�H;��H;��H;��H;�H;D�H;V�H;q�H;��H;��H;��H;      ��H;��H;��H;��H;��H;^�H;S�H;#�H;��H;��H;z�H;=�H;�H;��H;S�H;��H;��H;:�H;��H;��H;!�H;��H;m�H;�H;��H;[�H;�H;��H;��H;^�H;�H;��H;��H;��H;��H;��H;��H;��H;��H;��H;��H;��H;�H;X�H;��H;��H;�H;_�H;��H;�H;p�H;��H;�H;{�H;��H;;�H;��H;��H;N�H;��H;�H;@�H;z�H;��H;��H;&�H;Z�H;]�H;��H;��H;��H;��H;      |�H;u�H;}�H;|�H;e�H;B�H;A�H;�H;��H;��H;��H;@�H;�H;��H;v�H;8�H;��H;J�H;��H;��H;O�H;��H;�H;�H;��H;��H;4�H;��H;��H;��H;1�H;�H;��H;��H;��H;��H;��H;��H;��H;��H;��H;�H;1�H;}�H;��H;��H;1�H;��H;��H;�H;��H;��H;G�H;��H;��H;I�H;��H;9�H;v�H;��H;�H;?�H;��H;��H;��H;�H;I�H;=�H;k�H;}�H;��H;u�H;      -�H;)�H;*�H;�H;�H;�H;�H;��H;��H;��H;��H;X�H;�H;��H;o�H;�H;��H;��H;>�H;��H;^�H;�H;��H;F�H;��H;��H;S�H;�H;��H;��H;i�H;8�H;��H;��H;��H;��H;��H;��H;��H;��H;��H;<�H;k�H;��H;��H;�H;S�H;��H;��H;C�H;��H;�H;W�H;��H;<�H;��H;��H;�H;l�H;��H;�H;T�H;��H;��H;��H;��H;�H;��H;�H;"�H;3�H;#�H;      �H;�H;�H;�H;!�H;N�H;J�H;c�H;g�H;Q�H;O�H;6�H;�H;��H;��H;J�H;��H;��H;`�H;��H;��H;3�H;��H;��H;2�H;��H;�H;=�H;��H;��H;s�H;W�H;:�H;�H;��H;��H;��H;��H;��H;�H;:�H;X�H;s�H;��H;��H;9�H;}�H;��H;0�H;��H;��H;2�H;��H;��H;^�H;��H;��H;J�H;��H;��H;�H;6�H;N�H;R�H;i�H;c�H;M�H;A�H;'�H;�H;�H;�H;      �H;[�H;u�H;��H;��H;��H;#�H;Q�H;�H;��H;��H;��H;��H;��H;��H;w�H;#�H;��H;z�H;"�H;��H;��H;
�H;��H;c�H;�H;��H;j�H;/�H;��H;��H;z�H;o�H;7�H;�H;�H;�H;�H;�H;:�H;o�H;|�H;��H;��H;(�H;f�H;��H;	�H;_�H;��H;�H;��H;��H;"�H;z�H;��H;!�H;w�H;��H;��H;��H;��H;��H;��H;~�H;T�H;(�H;��H;��H;��H;|�H;Z�H;      ��H;��H;�H;\�H;��H;M�H;��H;��H;�H;��H;��H;�H;5�H;[�H;N�H;I�H;/�H;��H;��H;g�H;�H;��H;v�H;��H;��H;H�H;�H;��H;b�H;!�H;��H;��H;��H;}�H;]�H;A�H;5�H;C�H;Z�H;~�H;��H;��H;��H; �H;[�H;��H;��H;N�H;��H;��H;|�H;��H;�H;b�H;��H;��H;-�H;I�H;L�H;[�H;4�H; �H;��H;��H;��H;��H;��H;?�H;��H;b�H;�H;��H;      ��H;�H;�H;V�H;��H;7�H;��H;��H;��H;��H;��H;��H;�H;��H;��H;�H;�H;��H;��H;��H;I�H;��H;��H;U�H;��H;��H;3�H;��H;��H;^�H;(�H;��H;��H;��H;��H;��H;s�H;��H;��H;��H;��H;��H;+�H;_�H;��H;��H;0�H;��H;��H;N�H;��H;��H;E�H;��H;��H;��H;�H;�H;��H;��H;�H;��H;��H;��H;��H;��H;��H;1�H;��H;V�H;�H;�H;      ��H;��H;c�H;2�H;�H;��H;)�H;a�H;��H;�H;��H;��H;��H; �H;��H;8�H;��H;��H;��H;��H;��H;J�H;��H;��H;W�H;��H;t�H;J�H;��H;��H;h�H;;�H;�H;��H;��H;��H;��H;��H;��H;��H;�H;;�H;h�H;��H;��H;D�H;q�H;��H;R�H;��H;��H;I�H;��H;��H;��H;��H;��H;8�H;��H;��H;��H;��H;�H;
�H;��H;Z�H;*�H;p�H;'�H;4�H;p�H;��H;      �H;H;�!H;�8H;�TH;0sH;�H;��H;z�H;��H;U�H;��H;��H;��H;��H;��H;��H;�H;s�H;��H;��H;l�H;�H;��H;��H;E�H;��H;z�H;=�H;�H;��H;��H;T�H;6�H;!�H;��H;�H;��H;�H;8�H;T�H;��H;��H;�H;6�H;t�H;��H;K�H;��H;��H;�H;k�H;��H;��H;s�H;�H;��H;��H;��H;��H;��H;��H;U�H;��H;x�H;��H;�H;,sH;�TH;�8H;�!H;�H;      �CF;&RF;�zF;��F;�G;�\G;ʲG;*H;�HH;]�H;a�H;��H;��H;��H;��H;�H;��H;�H;��H;-�H;r�H;a�H;T�H;1�H;��H;r�H;G�H;��H;��H;Q�H;�H;��H;��H;��H;f�H;P�H;b�H;S�H;b�H;��H;��H;��H;	�H;Q�H;��H;��H;G�H;x�H;��H;.�H;X�H;b�H;o�H;.�H;��H;�H;��H;�H;��H;��H;��H;��H;a�H;]�H;�HH;#H;˲G;t\G;�G;ŸF;yzF;RF;      ��A;<B;�oB;�C;P�C;S�D;<uE;GDF;�F;k�G;�H;�eH;ݡH;��H;2�H;��H;��H;��H;n�H;n�H;�H;F�H;b�H;S�H;�H;��H;��H;Y�H;��H;��H;`�H;0�H;��H;��H;��H;��H;��H;��H;��H;��H;��H;0�H;d�H;��H;��H;U�H;��H;��H;�H;Q�H;g�H;H�H;�H;o�H;p�H;��H;��H;��H;1�H;��H;ޡH;�eH;�H;i�G;�F;GDF;<uE;F�D;]�C;�C;�oB;<B;      >o8;�8;��9;n�:;s�<;�c>;-R@;�/B;��C;�PE;izF;>\G;i�G;iH;�H;��H;�H;B�H;�H;�H;=�H;��H;A�H;Q�H;L�H;%�H;��H;��H;S�H;��H;��H;��H;F�H;�H;�H;�H;��H;�H;�H;�H;G�H;��H;��H;��H;P�H;��H;��H;,�H;I�H;S�H;E�H;��H;=�H;�H;�H;>�H;�H;��H;�H;iH;i�G;<\G;kzF;�PE;��C;�/B;.R@;�c>;��<;��:;��9;�8;      ]S%;��%;�';�M*;ѷ-;z�1;؟5;��9;o-=;R@;��B;b�D;mF;�uG;X!H;��H;��H;{�H;��H;j�H;��H;�H;��H;H�H;b�H;Q�H;�H;��H;��H;v�H;
�H;��H;��H;�H;n�H;Y�H;=�H;X�H;m�H;~�H;��H;��H;�H;{�H;��H;��H;�H;X�H;`�H;F�H;��H;�H;��H;l�H;��H;v�H;��H;��H;X!H;�uG;mF;`�D;��B;
R@;m-=;��9;؟5;z�1;Է-;�M*;�';��%;      fW;px;��;
�
;��;�;�� ;p�(;��/;�H6;��;;��?;�C;�PE;��F;��G;�eH;%�H;e�H;��H;,�H;��H;�H;��H;F�H;^�H;h�H;J�H;��H;��H;��H;-�H;��H;��H;��H;��H;��H;��H;��H;��H;��H;-�H;��H;��H;��H;I�H;i�H;b�H;?�H;��H;�H;��H;,�H;��H;e�H;$�H;�eH;��G;��F;�PE;�C;��?;��;;�H6;��/;p�(;�� ;j;��; �
;��;dx;      ���:�ņ:�ɒ:��:��:���:$��:E�	;�v;��#;��-;��5;zL<;`�@;�(D;DF;��G;�HH;J�H;��H;��H;*�H;��H;=�H;��H;h�H;��H;��H;A�H;�H;��H;��H;S�H;I�H;�H;�H;�H;�H;�H;E�H;U�H;��H;��H;�H;>�H;��H;��H;k�H;��H;;�H;��H;'�H;��H;��H;J�H;�HH;��G;DF;�(D;]�@;wL<;��5;��-;��#;�v;K�	;*��:��:��:��:�ɒ:�ņ:      �-.�$������~K��
90]: �k:UM�:���:�y;��;z $;��/;d�8;��>;�#C;�E;Y\G;/8H;��H;��H;��H;l�H;�H;k�H;,�H;��H;��H;��H;`�H;�H;��H;��H;��H;}�H;r�H;^�H;t�H;|�H;��H;��H;��H;�H;a�H;��H;��H;��H;0�H;e�H;�H;l�H;��H;��H;��H;/8H;V\G;�E;�#C;}�>;b�8;��/;v $;��;�y;���:CM�:�k:]: 
9�K����0��      0Q^�X��F�Т)�,+��ζ�d�<��AS�$n:��:���:��;6�;�M*;ҟ5;tc=;KpB;��E;�JG;-8H;M�H;g�H;��H;�H;g�H;��H;o�H;��H;��H;��H;v�H;[�H;7�H;��H;��H;��H;��H;��H;��H;��H;7�H;Z�H;w�H;��H;��H;��H;p�H;��H;b�H;
�H;��H;c�H;J�H;/8H;�JG;��E;HpB;mc=;П5;�M*;5�;��;���:��:n:�AS�p�<��ζ�,+�Ϣ)��F�X�      _���0���"���ѻ"���ǐ�_X�*6�L	���uK��>":�M�:&b�:Hi;�%;H�3;߆<;(0B;��E;U\G;�HH;$�H;y�H;?�H;��H;�H;�H;��H;��H;��H;��H;��H;��H;E�H;5�H;5�H;�H;7�H;4�H;C�H;��H;��H;��H;��H;��H;��H;�H;�H;��H;;�H;w�H; �H;�HH;U\G;~�E;%0B;܆<;E�3;�%;Di;"b�:�M�:�>":�uK�P	��-6�dX�ǐ�$����ѻ&��1���      o�n�ymj���]���J�Y�1�44�8������	x��W�P�y� (
9樂:6��:��;6�#;8�2;�<;JpB;�E;��G;�eH;��H;�H;��H;��H;��H;��H;�H;'�H;�H;��H;��H;��H;��H;��H;��H;��H;��H;��H;��H;��H;�H;(�H;�H;��H;��H;��H;��H;�H;��H;�eH;��G;�E;GpB;߆<;7�2;2�#;��;0��:樂:�'
9`�y��W��	x����:��44�[�1���J���]�xmj�      ?<ͼ�ɼ�����֯�ζ��ㄼ��Y��*�����s��X��rѺ���>Q:���:��
;.�#;I�3;pc=;�#C;DF;��G;�H;��H;��H;�H;��H;4�H; �H;D�H;q�H;G�H;�H;6�H;��H;��H;��H;��H;��H;1�H;�H;D�H;p�H;F�H;��H;5�H;��H;�H;��H;��H;�H;��G;�CF;�#C;lc=;E�3;.�#;��
;���:�>Q: ��rѺ X��s������*���Y�ㄼ϶���֯������ɼ      ��'�(�$����|��  ���ۼ����+����]��X!�E>ۻ�+���*������>:���:��;�%;Ο5;z�>;�(D;��F;\!H;�H;-�H;��H;��H;��H;��H;M�H;��H;��H;j�H;q�H;J�H;2�H;Q�H;4�H;I�H;p�H;h�H;��H;��H;L�H;��H;��H;��H;��H;'�H;�H;W!H;��F;{(D;z�>;ȟ5;�%;��;���:��>:��깅*��+��G>ۻ�X!���]��+�������ۼ�  �|����(�$�      Ÿ���v����w�f�c��J�΄-�|��;缅沼ㄼ��;������j���5�h���>Q:2��:Hi;�M*;d�8;j�@;�PE;�uG;iH;��H;��H;��H;��H;��H;W�H;��H;��H;��H;��H;��H;��H;��H;��H;��H;��H;��H;��H;��H;Z�H;��H;��H;��H;��H;��H;iH;�uG;�PE;]�@;f�8;�M*;Gi;0��:�>Q:��깭5��j��������;�ㄼ�沼�;�|�΄-��J�f�c���w��v��      yHͽ֪ɽ�;��"����Ǹ����[�	z0�s��&<ͼ˾��d�J�����j��~*���⨂:*b�:5�;��/;�L<;�C;mF;p�G;ߡH;��H;��H;��H;�H;4�H;��H;�H;�H;��H;��H;��H;��H;��H;��H;��H;�H;�H;��H;4�H;�H;��H;��H;��H;ڡH;l�G;mF;�C;vL<;��/;1�;$b�:ਂ:���*��j�����d�J�˾��'<ͼs��	z0���[�Ǹ����"���;��֪ɽ      ��"-������ѱ�ƽ]P���v���J�G����ۼ��d�J������+���rѺ�'
9�M�:��;v $;��5;��?;b�D;@\G;�eH;��H;��H;��H;��H;��H;��H;2�H;U�H;=�H;3�H;D�H;�H;D�H;0�H;:�H;Q�H;/�H;��H; �H;��H;��H;��H;��H;�eH;>\G;b�D;��?;��5;v $;��;�M�:�'
9�rѺ�+������d�J�����ۼG���J��v��]P��ƽұ轃����"-�       j�Vde�Z0X�D�e{+�������u㻽Y���RDX������ۼ˾����;�G>ۻ#X�p�y��>":���:��;��-;��;;��B;lzF;�H;a�H;T�H;��H;��H;��H;��H;M�H;��H;~�H;q�H;��H;[�H;��H;p�H;{�H;��H;J�H;��H;��H;��H;��H;Q�H;]�H;�H;lzF;��B;�;;��-;��;���:�>":p�y�&X�H>ۻ��;�̾����ۼ���RDX�Y���u㻽��콂��f{+�D�Z0X�Vde�      ��Ph��k���I���|x���O��C(���Ϊɽ����RDX�H��'<ͼ	ㄼ�X!��s���W� vK���:�y;��#;�H6;R@;�PE;i�G;]�H;��H;�H;��H;��H;��H;R�H;��H;��H;��H;��H;��H;��H;��H;��H;��H;O�H;��H;~�H;��H;�H;��H;[�H;e�G;�PE;R@;�H6;�#;�y;��: vK��W��s���X!�	ㄼ'<ͼH��RDX�����Ϊɽ���C(���O��|x��I��k��Ph��      >����������"�;hɰ��G��
 j�8�5��	�ΪɽY����J�s���沼��]�����	x�b	��n:���:�v;��/;g-=;��C;�F;�HH;z�H;��H;��H;�H;~�H;f�H;��H;��H;��H;��H;�H;��H;��H;��H;��H;d�H;z�H; �H;��H;��H;z�H;�HH;�F;��C;h-=;��/;�v;���: n:^	���	x������]��沼s���J�Y���Ϊɽ�	�9�5�
 j��G��hɰ�"�;��徶���      �2�U�-�"�-E�����?Kɾj����s�9�5���u㻽�v��	z0��;��+���*����<6� CS�AM�:M�	;l�(;�9;�/B;HDF;H;��H;Y�H;��H;��H;L�H;c�H;��H;�H;�H;�H;7�H;�H;�H;�H;��H;_�H;J�H;��H;��H;Z�H;��H; H;GDF;�/B;�9;n�(;E�	;IM�: DS�76�����*��+���;�	z0��v��u㻽��9�5���s�j��?Kɾ����-E�"�U�-�      %3s�cm�:�\�h�C�5�%����TҾj��
 j��C(����]P����[�|������Y�;��lX�|�<���k:0��:�� ;ԟ5;0R@;5uE;ͲG;�H;�H;��H;��H; �H;D�H;�H;A�H;K�H;6�H;k�H;4�H;L�H;>�H;�H;D�H;�H;��H;��H;�H;�H;ҲG;4uE;1R@;֟5;�� ;"��: �k:��<�iX�;����Y����|���[�]P����콪C(�
 j�j���TҾ���5�%�h�C�:�\�cm�      �ޞ�������`F�?�W�W�-����?Kɾ�G����O����ƽǸ��΄-���ۼㄼ54�ǐ�
϶�]:��:y;|�1;�c>;B�D;u\G;'sH;t�H;3�H;D�H;��H;J�H;	�H;H�H;h�H;Z�H;��H;\�H;h�H;E�H;�H;J�H;��H;F�H;7�H;x�H;,sH;~\G;B�D;�c>;|�1;y;��: ]:϶�ǐ�64�ㄼ��ۼ΄-�Ǹ��ƽ�����O��G��?Kɾ���W�-�?�W�`F�������      ��ſ���Lw���ޞ�����?�W�5�%�����hɰ��|x�f{+�ұ����J��  �϶��Z�1�-���$+� 
9��:��;޷-;��<;[�C;�G;�TH; �H;��H;��H;��H;(�H;�H;e�H;��H;t�H;��H;o�H;��H;`�H;�H;(�H;��H;��H;��H;&�H;�TH;�G;Z�C;��<;޷-;��;��:@ 
9%+�*���[�1�϶���  ��J���ұ�f{+��|x�hɰ�����5�%�?�W������ޞ�Lw�����      ������Կp���ޞ�`F�h�C�-E�#�;�I��D���"��f�c�|��֯���J��ѻԢ)��K���:�
;�M*;i�:;�C;ŸF;�8H;*�H;F�H;W�H;��H;�H;�H;�H;��H;��H;��H;��H;��H;{�H;�H;�H;��H;^�H;J�H;+�H;�8H;иF;�C;l�:;�M*;�
;��:�K�֢)��ѻ��J��֯�|�f�c�"����D��I��#�;-E�h�C�`F��ޞ�p���Կ��      ����������ԿLw�����:�\�"����k��Z0X�����;����w����������]�#���F�����ɒ:��;��';��9;�oB;}zF;�!H;q�H;��H; �H;o�H;�H;�H;}�H;��H;��H;��H;��H;��H;|�H;�H;�H;k�H;�H;��H;t�H;�!H;�zF;�oB;��9;��';��;�ɒ:����F�"�黬�]����������w��;�����Y0X�k�����"�:�\����Lw���Կ��𿝏�       $�������忈�����cm�V�-�����Qh��Vde�"-�תɽ�v��(�$���ɼ{mj�;���X�$���ņ:dx;�%;.�8;BB;RF;�H;�H;�H;��H;B�H;�H;�H;v�H;��H;��H;�H;��H;��H;v�H;�H;�H;A�H;��H;�H;�H;�H;,RF;BB;0�8;�%;bx;�ņ:��X�8���|mj���ɼ(�$��v��תɽ"-�Vde�Qh������V�-�cm��������忝����      �>���8���*�O������˿p��E�b�C\�4m־^��Q�:��J�)��E�B�=��������2/��X���ؑ>:it�:p ;�J6;�DA;ZIF;�NH;��H;�!I;�I;�I;zI;LI;�I;H I;��H;	�H;��H;H I;�I;NI;|I;�I;�I;�!I;��H;�NH;hIF;�DA;�J6;
p ;it�:ؑ>:J���2/���������=��E�B�)���J�Q�:�^��4m־C\�E�b�p���˿����O���*���8�      ��8��4��g&�6��<����<ƿ񲗿�>]����O�Ѿ�p���*7����%W��LR?� }�r8�������څ��|�G:q �:�!;�6;�kA;eYF;�TH;C�H;�!I;�I;�I;dI;&I;�I;: I;��H;��H;��H;< I;�I;)I;gI;�I;�I;�!I;G�H;�TH;rYF;�kA;�6;�!;q �:|�G:Ѕ�������r8�� }�LR?�%W�����*7��p��O�Ѿ����>]�񲗿�<ƿ<���6���g&��4�      ��*��g&��#�t�T[�qL�������M�r5��>ľ����,��D�蒐��5�2�ݼ���q
��x�4uk���b:%l�:�#;7;S�A;��F;�dH;�I;!"I;�I;DI;I;�I;�I;��H;X�H;��H;R�H;��H;�I;�I;I;AI;�I;%"I;�I;�dH;��F;T�A;��7;�#;%l�:��b:uk��x��q
���2�ݼ�5�蒐��DὫ�,����>ľr5���M����qL��T[�t��#��g&�      O�6��t����˿@1��7�y�Î6��z �����2�l�+��ͽ#�����&���˼@�k�%�����X�� �p��:6�;�&;}9;k�B;��F;�}H;�	I;."I;I;�I;xI;RI;$I;��H;�H;_�H;��H;��H;"I;RI;{I;�I;I;3"I;�	I;�}H;��F;j�B;z9;�&;6�;p��:� ���X�"���@�k���˼��&�#����ͽ+�2�l������z �Î6�7�y�@1���˿���t�6��      ����<���T[忶˿�T���{�R�����E۾ӗ����M���	������j��3�d����O�>�׻��/�x��9��:� 
;�*;O;;�jC;�'G;ӛH;�I;�!I;�I;tI;�
I;�I;�I;�H;��H;��H;��H;"�H;�I;�I;�
I;sI;�I;�!I;�I;؛H;�'G;�jC;K;;�*;� 
;9��:0����/�<�׻��O�d���3���j������	���M�ӗ���E۾���{�R���T���˿T[�<���      �˿�<ƿqL��@1����>]���)��$��ֳ���{���,�q��'��Q`I��J���,���3/�,��� ��,69�4�:Є;�o.;.=;=aD;��G;P�H;�I;!I;>I;)I;�	I;�I;� I;�H;��H;B�H;��H;��H;� I;�I;�	I;)I;CI;!I;�I;Q�H;��G;?aD;.=;�o.;Є;�4�:�,69� � ,���3/��,���J��Q`I�'��q�齥�,���{�ֳ��$����)��>]��@1��qL���<ƿ      p��񲗿���7�y�{�R���)�nv��>ľ^���I�Xl����������&�ԮҼ�}�3B�ή��*���d�!:�*�:z;X3;Ij?;r\E;��G;��H;HI;|I;jI;�I;VI;�I;��H;��H;B�H;��H;A�H;��H;��H;�I;WI;�I;pI;I;II;��H;��G;t\E;Fj?;Y3;"z;�*�:��!:���ͮ��2B��}�ԮҼ��&��������Xl��I�^���>ľnv���)�{�R�7�y����񲗿      E�b��>]���M�Î6�����$���>ľ#q��y�Z�+�Q9ݽ!W����L����#F���G��׻;�ho�tȊ:~i;�O$;��7;S�A;�IF;CH;��H;� I;BI;TI;�I;I;~I;��H;��H;r�H;��H;r�H;��H;��H;I;I;�I;ZI;EI;� I;��H;CH;�IF;P�A;��7;P$;zi;�Ȋ:Po�;��׻�G�"F�������L�!W��Q9ݽ+�y�Z�#q���>ľ�$�����Î6���M��>]�      C\����r5��z ��E۾ֳ�^��y�Z�L?#����A����j�%��Fϼ�����ε���lۺ(9�9X4�:=�;@�,;U�;;�C;}G;�H;I;�!I;�I;"I;I;pI;#I;��H;��H;��H;��H;��H;��H;��H;#I;sI;I;'I;�I;�!I;�I; �H;�G;�C;Y�;;F�,;;�;l4�:P9�9�lۺʵ�������Eϼ%����j��A�����K?#�y�Z�^��ֳ��E۾�z �r5����      4m־O�Ѿ�>ľ����җ����{��I�+�����V���{�?�/�&���,��A=�F�һu�@�d� ���k:��:�a;��3;j?;P2E;��G;A�H;I;M I;�I;�I;�I;�I;��H;��H;��H;��H;9�H;��H;��H;��H;��H;�I; 	I;�I;�I;P I;I;?�H;��G;N2E;j?;��3;�a;��:��k:H� �m�@�D�һ?=��,��%��>�/��{��V�����+��I���{�ӗ�������>ľO�Ѿ      ^���p����2�l���M���,�Xl�Q9ݽ�A���{���5��J��
;���T[�$?�����nP���O�9��:��;	*; �9;2kB;��F;TNH;V�H;�I;fI;�I;�I;�I; I;C�H;��H;��H;��H;H�H;��H;��H;��H;D�H;!I;�I;I;�I;kI;�I;T�H;ZNH;��F;7kB;�9;*;��;��: P�9ZP������#?��T[�	;���J����5��{��A��Q9ݽXl���,���M�2�l����p��      Q�:��*7���,�+���	�q�齂��� W����j�>�/��J���I���k�n�.��l��x���Ȋ:!o�:�;?r3;��>;�D;L�G;!�H;�I;!I;�I;bI;_
I;�I;? I;��H;x�H;��H;��H;@�H;��H;��H;|�H;��H;? I;�I;g
I;mI;�I;!I;�I;'�H;M�G;�D;�>;Cr3;�;)o�:�Ȋ:(��f��.��l��k��I���J��>�/���j� W������q�齂�	�+���,��*7�      �J�����D��ͽ���'�������L�%��%��	;���k����nI����/��/��>:��:�B;:�,;��:;�B;ixF;t<H;��H;�I;qI;�I;I;�I;�I;m�H;W�H;�H;N�H;~�H;M�H;�H;N�H;�H;W�H;n�H;�I;�I;I;�I;qI;�I;��H;u<H;mxF;�B;��:;H�,;�B;��:0�>:�/���/�lI������k�;��%��%����L����'������ͽ�D����      (��%W��蒐�#�����j�R`I���&����Eϼ�,���T[�m�pI��k;��nk�d:�4�:�;�&;��6;�!@;2E;��G;~�H;�I;� I;/I;�I;�
I;I;P I;��H;��H;��H;?�H;t�H;&�H;v�H;@�H;��H;��H;��H;V I;I;�
I;�I;/I;� I;�I;~�H;��G;2E;�!@;��6;�&;�;�4�:h:�nk�d;�mI��l��T[��,��Dϼ�����&�Q`I���j�#���蒐�$W��      D�B�LR?��5���&��3��J��ԮҼ"F����@=�#?�.����/��nk����9׳:��;!;63;��=;��C;��F;�cH;��H;kI;�I;�I;�I;�I;�I;!�H;��H;r�H;_�H; �H;e�H;�H;e�H; �H;b�H;u�H;��H;%�H;�I;�I;I;�I;�I;oI;��H;�cH; �F;��C;��=;=3;!;��; ׳:���9�nk���/�.��"?�@=���"F��ԮҼ�J���3���&��5�MR?�      :���|�1�ݼ��˼d���,���}��G����D�һ����l���/�\:׳:�;Lb;��0;j<;~�B;�IF;GH;��H;�I;L I;�I;I;6
I;�I;  I;�H;6�H;��H;�H;�H;\�H;�H;\�H;�H;�H;��H;6�H;�H; I;�I;<
I;I;�I;P I;�I;�H;LH;�IF;��B;p<;��0;Rb;�;"׳:h:�/�h������C�һ����G��}��,��d����˼1�ݼ�|�      ����p8����@�k���O��3/�0B��׻ʵ��j�@�ZP��H�� �>:�4�:��;Ob;|�/;;;�A;d�E;��G;ͭH;�
I;D I;�I;�I;�I;�I;�I;e�H;�H;��H;{�H;��H;��H;Q�H;�H;M�H;��H;��H;x�H;��H;�H;i�H;�I;�I;�I;�I;�I;E I;�
I;ҭH;��G;m�E;�A;;;��/;Sb;��;�4�:$�>:8��RP��i�@�ǵ��
�׻2B��3/���O�A�k���o8��      ������q
����8�׻ ,��Ȯ��;��lۺ@� ��O�9�Ȋ:��:|;!;��0;	;;��A;�pE;L�G;��H;��H;�I;I;,I;�I;�I;SI;��H;"�H;W�H;��H;��H;��H;��H;G�H;�H;D�H;��H;��H;��H;��H;[�H;(�H;��H;UI;�I;�I;2I;I;�I;��H;��H;T�G;�pE;��A;;;��0;!;�;��:�Ȋ:8P�9H� ��lۺ;�ʮ�� ,��4�׻����q
���      (/��&����x���X���/�� ����(o�p9�9��k:��:'o�:�B;�&;:3;m<;�A;�pE;@tG;�|H;�H;I;OI; I;�I;J
I;�I;0 I;*�H;�H;��H;^�H;��H;��H;��H;X�H;E�H;X�H;��H;��H;��H;]�H;��H;�H;,�H;4 I;�I;H
I;�I;#I;KI;I;�H;�|H;BtG;�pE; �A;k<;=3;�&;�B;)o�:��:��k:x9�90o����� ���/���X��x�&���      T���䅍�uk��� �x���,69��!:zȊ:f4�:��:��;�;@�,;��6;��=;��B;k�E;V�G;�|H;s�H;TI;�I;_I;6I;�I;I;fI;&�H;��H;�H;��H;��H;��H;��H;��H;n�H;U�H;k�H;��H;��H;��H;��H;��H;�H;��H;+�H;eI;I;�I;6I;^I;�I;ZI;u�H;�|H;S�G;k�E;��B;��=;��6;A�,;�;��;��:p4�:�Ȋ:��!:0-69X���� �@uk�����      T�>:,�G:X�b:b��:��:�4�:�*�:zi;9�;�a;*;;r3;��:;�!@;��C;�IF;��G;��H;�H;SI;�I;I;I;�I;�I;:I;��H;k�H;��H;X�H;)�H;��H;}�H;��H;��H;��H;d�H;��H;��H;��H;z�H;��H;/�H;\�H;��H;m�H;��H;7I;�I;�I;I;I;  I;TI;
�H;��H;��G;�IF;��C;�!@;��:;=r3;*;�a;7�;xi;�*�:�4�:1��:^��:��b:,�G:      ]t�:� �:9l�:H�;� 
;҄;z;�O$;H�,;��3;�9;��>;�B;2E;��F;OH;ԭH;��H;	I;�I;"I;ZI;I;�I;�I;��H;�H;.�H;��H;x�H;��H;��H;t�H;��H;�H;��H;��H;��H;�H;��H;q�H;��H;��H;y�H;��H;1�H;��H;��H;�I;�I;I;]I;$I;�I;	I;��H;խH;LH; �F;2E;�B; �>;	�9;��3;G�,;P$;"z;̄;� 
;<�;!l�:q �:      $p ;�!;�#;�&;�*;�o.;g3;��7;\�;;j?;9kB;�D;jxF;��G;�cH;�H;�
I;�I;QI;_I;I;I;�I;9I;�H;o�H;o�H;	�H;��H;��H;��H;d�H;u�H;��H;9�H;�H;��H;��H;6�H;��H;q�H;d�H;��H;��H;��H;�H;l�H;r�H;�H;6I;�I;I;I;aI;QI;�I;�
I;�H;�cH;��G;jxF;�D;>kB;j?;^�;;��7;b3;�o.;�*;�&;�#;�!;      �J6;�6;��7;y9;@;;.=;Hj?;O�A;�C;M2E;��F;L�G;r<H;�H;��H;�I;G I;I;%I;5I;�I;�I;9I;/�H;��H;��H;A�H;�H;�H;��H;h�H;U�H;w�H;�H;��H;V�H;,�H;P�H;��H;�H;t�H;R�H;j�H;��H;�H;�H;<�H;��H;��H;,�H;2I;�I;�I;3I;"I;I;D I;�I;��H;{�H;o<H;J�G;��F;K2E;�C;T�A;Aj?;�-=;K;;v9;��7;�6;      �DA;�kA;I�A;g�B;�jC;KaD;y\E;�IF;G;��G;]NH;+�H;��H;�I;tI;W I;�I;9I;�I;�I;�I;�I;�H;��H;��H;`�H;�H;/�H;��H;y�H;M�H;e�H;��H;A�H;��H;��H;��H;��H;��H;C�H;��H;a�H;O�H;y�H;��H;0�H;�H;`�H;��H;��H;�H;�I;�I;�I;�I;5I;�I;W I;qI;�I;��H;+�H;^NH;��G;�G;�IF;w\E;?aD;�jC;f�B;F�A;�kA;      VIF;oYF;��F;��F;r'G;��G;��G;CH;�H;E�H;W�H;�I;�I;� I;�I;�I;�I; I;J
I;I;<I;��H;q�H;��H;]�H;8�H;D�H;��H;|�H;\�H;F�H;��H;�H;�H;7�H;�H;�H;�H;3�H;�H;�H;��H;G�H;[�H;y�H;��H;@�H;<�H;`�H;��H;n�H;��H;<I;I;J
I;�I;�I;�I;�I;� I;�I;�I;[�H;E�H; �H;CH;��G;��G;�'G;��F;��F;kYF;      �NH;�TH;�dH;�}H;ʛH;P�H;��H;��H;�I;I;�I;!I;mI;/I;�I;I;�I;�I;�I;iI;�H; �H;r�H;F�H;�H;A�H;��H;�H;N�H;M�H;��H;��H;U�H;��H;��H;��H;x�H;��H;��H;��H;U�H;��H;��H;L�H;H�H;�H;��H;F�H;�H;A�H;o�H;�H;�H;fI;�I;�I;�I;I;�I;+I;mI;!I;�I;I;~I;��H;��H;I�H;�H;�}H;�dH;vTH;      ��H;G�H;�I;�	I;�I;�I;RI;� I;�!I;T I;kI;�I;�I;�I;�I;<
I;�I;RI;4 I;(�H;n�H;-�H;�H;�H;)�H;��H;}�H;]�H;D�H;u�H;��H;2�H;��H;q�H;5�H;�H;��H;�H;2�H;r�H;��H;/�H;��H;u�H;@�H;\�H;y�H;��H;/�H;�H;	�H;0�H;m�H;'�H;1 I;PI;�I;<
I;�I;�I;�I;�I;kI;P I;�!I;� I;PI;�I;�I;�	I;�I;<�H;      �!I;�!I;"I;@"I;�!I;
!I;�I;EI;�I;�I;�I;lI;I;�
I;�I;�I;�I;��H;3�H;��H;��H;��H;��H;�H;��H;u�H;F�H;D�H;��H;��H;"�H;��H;A�H;��H;��H;��H;��H;��H;��H;��H;@�H;��H;"�H;��H;��H;C�H;C�H;v�H;��H;�H;��H;��H;��H;��H;1�H;��H;�I;�I;�I;�
I;I;iI;�I;�I;�I;DI;�I;!I;�!I;@"I;"I;�!I;      �I;|I;�I;I;�I;<I;kI;XI;$I;�I;I;i
I;�I;I;�I; I;m�H;"�H;�H;!�H;_�H;v�H;��H;��H;v�H;T�H;I�H;v�H;��H;�H;��H;<�H;��H;��H;b�H;B�H;1�H;B�H;\�H;��H;��H;:�H;��H;�H;��H;u�H;D�H;V�H;y�H;��H;��H;y�H;[�H;�H;�H;!�H;m�H; I;�I;I;�I;f
I;I;�I;!I;TI;nI;:I;�I;I;�I;|I;      �I;�I;II;�I;sI;)I;�I;�I;	I;	I;�I;�I;�I;X I;(�H;�H;%�H;`�H;��H;��H;4�H;��H;��H;k�H;M�H;F�H;��H;��H;(�H;��H;�H;��H;m�H;1�H;�H;��H;��H;��H;�H;4�H;m�H;��H;�H;��H;!�H;��H;��H;G�H;O�H;h�H;��H;��H;0�H;��H;��H;^�H;%�H;�H;%�H;W I;�I;�I;�I;	I;
I;�I;�I; I;�I;�I;KI;�I;      |I;oI;I;uI;�
I;�	I;XI;	I;vI;�I;"I;C I;q�H;��H;��H;;�H;��H;��H;e�H;��H;��H;��H;c�H;R�H;c�H;��H;��H;4�H;��H;=�H;��H;L�H;�H;��H;��H;��H;��H;��H;��H;��H;�H;J�H;��H;<�H;��H;/�H;��H;��H;f�H;M�H;h�H;��H;��H;��H;d�H;��H;��H;=�H;��H;��H;p�H;B I;$I;�I;tI;I;^I;�	I;�
I;vI;I;nI;      YI;6I;�I;VI;�I;�I;�I;|I;I;��H;F�H;��H;Y�H;��H;v�H;��H;��H;�H;��H;��H;��H;u�H;t�H;t�H;��H;�H;U�H;��H;G�H;��H;i�H;�H;��H;��H;��H;g�H;`�H;g�H;��H;��H;��H;�H;h�H;��H;C�H;��H;R�H;�H;��H;t�H;x�H;t�H;��H;��H;��H;�H;��H;��H;w�H;��H;Y�H;��H;G�H;��H;I;{I;�I;�I;�I;QI;�I;4I;      �I;�I;�I;I;�I;� I;��H;��H;��H;��H;��H;��H;�H;��H;f�H;�H;��H;��H;��H;��H;��H;��H;��H;�H;;�H;x�H;��H;t�H;��H;��H;.�H;��H;��H;g�H;Q�H;B�H;4�H;C�H;P�H;h�H;��H;��H;.�H;��H;��H;p�H;��H;y�H;?�H;�H;��H;��H;��H;��H;��H;��H;��H;�H;f�H;��H;�H;~�H;��H;��H;��H;��H;  I;� I;�I; I;�I;�I;      B I;P I; I;��H;0�H;{�H;��H;��H;��H;��H;��H;��H;Y�H;J�H;+�H;�H;��H;��H;��H;��H;��H;�H;4�H;��H;��H;,�H;��H;2�H;��H;a�H;��H;��H;��H;P�H;.�H;�H;#�H; �H;*�H;Q�H;��H;��H;��H;^�H;��H;.�H;��H;-�H;��H;��H;8�H;�H;��H;��H;��H;��H;��H;�H;*�H;J�H;Y�H;��H;��H;��H;��H;��H;��H;{�H;0�H;��H;  I;Q I;      ��H;��H;X�H;�H;��H;��H;L�H;y�H;��H;��H;��H;��H;��H;x�H;i�H;\�H;R�H;C�H;Z�H;m�H;��H;��H;��H;C�H;��H;�H;��H;�H;��H;D�H;��H;��H;l�H;B�H;#�H;�H;
�H;�H; �H;H�H;l�H;��H;��H;@�H;��H;��H;��H;�H;��H;E�H; �H;��H;��H;h�H;Z�H;I�H;U�H;`�H;h�H;{�H;��H;��H;��H;��H;��H;x�H;S�H;��H;��H;�H;T�H;��H;      �H;��H;��H;f�H;��H;>�H;��H;��H;�H;8�H;T�H;K�H;U�H;/�H; �H;�H;�H;�H;I�H;Z�H;k�H;��H;��H;"�H;��H;��H;r�H;��H;��H;5�H;��H;��H;d�H;3�H;%�H;�H;�H;�H;"�H;4�H;g�H;��H;��H;1�H;��H;��H;t�H; �H;��H;"�H;��H;��H;f�H;V�H;H�H;#�H;�H;#�H;�H;2�H;U�H;G�H;T�H;9�H;�H;��H;��H;>�H;��H;j�H;��H;��H;      ��H;��H;R�H;�H;��H;��H;J�H;v�H;��H;��H;��H;��H;��H;{�H;i�H;\�H;T�H;C�H;Z�H;n�H;��H;��H;��H;C�H;��H;�H;��H;�H;��H;D�H;��H;��H;n�H;C�H;#�H;�H;
�H;�H; �H;F�H;l�H;��H;��H;?�H;��H;��H;��H;�H;��H;E�H; �H;��H;��H;h�H;Z�H;J�H;T�H;a�H;h�H;z�H;��H;��H;��H;��H;��H;y�H;S�H;��H;��H;�H;Y�H;��H;      7 I;P I;��H;��H;/�H;w�H;��H;��H;��H;��H;��H;��H;Z�H;J�H;-�H;�H;��H;��H;��H;��H; �H;�H;4�H;��H;��H;*�H;��H;2�H;��H;_�H;��H;��H;��H;P�H;-�H;�H;%�H;"�H;,�H;Q�H;��H;��H;��H;\�H;��H;,�H;��H;/�H;��H;��H;8�H;�H;��H;��H;��H;��H;��H;�H;(�H;H�H;W�H;��H;��H;��H;��H;��H;��H;u�H;4�H;��H; I;V I;      �I;�I;�I; I;�I;� I;��H;��H;��H;��H;��H;��H;�H;��H;g�H;�H;��H;��H;��H;��H;��H;��H;��H;�H;>�H;x�H;��H;t�H;��H;��H;-�H;��H;��H;g�H;Q�H;A�H;4�H;B�H;P�H;g�H;��H;��H;-�H;��H;��H;p�H;��H;{�H;?�H; �H;��H;��H;��H;��H;��H;��H;��H;�H;f�H;��H;�H;~�H;��H;��H;��H;��H; I;� I;�I;"I;�I;�I;      VI;;I;�I;RI;�I;�I;�I;�I; I;��H;F�H;��H;\�H;��H;y�H;��H;��H;�H;��H;��H;��H;v�H;t�H;v�H;��H;�H;S�H;��H;G�H;��H;f�H;�H;��H;��H;��H;g�H;`�H;g�H;��H;��H;��H;�H;h�H;��H;?�H;��H;S�H;�H;��H;q�H;z�H;t�H;}�H;��H;��H;�H;��H;��H;v�H;��H;Z�H;��H;F�H;��H;I;I;�I;�I;�I;\I;�I;6I;      rI;pI;I;qI;�
I;�	I;]I;	I;tI;�I;%I;F I;r�H;��H;��H;<�H;��H;��H;d�H;��H;��H;��H;e�H;R�H;h�H;��H;��H;3�H;��H;<�H;��H;I�H;�H;��H;��H;��H;��H;��H;��H;��H;�H;J�H;��H;:�H;��H;/�H;��H;��H;c�H;J�H;k�H;��H;��H;��H;b�H;��H;��H;=�H;��H;��H;q�H;C I;$I;�I;vI;I;]I;�	I;�
I;vI;I;kI;      �I;�I;II;�I;zI;)I;�I;�I;
I;	I;�I;�I;�I;[ I;+�H;�H;'�H;`�H;��H;��H;6�H;��H;��H;k�H;R�H;C�H;��H;��H;(�H;��H;�H;��H;l�H;2�H;�H;��H;��H;��H;�H;5�H;m�H;��H;�H;��H;!�H;��H;��H;I�H;M�H;g�H;��H;��H;/�H;��H;��H;^�H;%�H;�H;(�H;X I;�I;�I;�I;	I;
I;�I;�I;&I;�I;�I;OI;�I;      �I;�I;�I;I;�I;II;mI;^I;(I;�I;I;i
I;�I;I;�I; I;m�H;#�H;�H;�H;a�H;y�H;��H;��H;{�H;R�H;I�H;w�H;��H;�H;��H;9�H;��H;��H;_�H;@�H;1�H;C�H;\�H;��H;��H;:�H;��H;�H;��H;s�H;F�H;X�H;u�H;��H;��H;x�H;\�H;�H;�H;"�H;l�H; I;�I;I;�I;d
I; I;�I;$I;[I;mI;;I;�I;$I;�I;I;      �!I;�!I;/"I;<"I;�!I;!I;~I;EI;�I;�I;�I;lI;I;�
I;�I;�I;�I;��H;0�H;��H;��H;��H;��H; �H;��H;q�H;D�H;F�H;��H;��H;!�H;��H;@�H;��H;��H;��H;��H;��H;��H;��H;A�H;��H;"�H;��H;��H;@�H;C�H;v�H;��H;�H;��H;��H;��H;��H;3�H;��H;�I;�I;�I;�
I;I;iI;�I;�I;�I;GI;�I;!I;�!I;@"I;/"I;�!I;      ��H;=�H;xI;�	I;�I;�I;RI;� I;�!I;T I;kI;�I;�I;�I;I;=
I;�I;SI;3 I;'�H;p�H;0�H;�H;�H;/�H;��H;{�H;]�H;F�H;s�H;��H;0�H;��H;q�H;2�H;�H;��H;�H;0�H;r�H;��H;0�H;��H;r�H;@�H;Y�H;y�H;��H;)�H;�H;�H;.�H;k�H;'�H;4 I;OI;�I;:
I;�I;�I;�I;�I;kI;R I;�!I;� I;SI;�I;�I;�	I;�I;=�H;      �NH;�TH;�dH;�}H;ڛH;V�H;��H;��H;�I;I;�I;!I;mI;0I;�I;I;�I;�I;�I;hI;�H;�H;n�H;H�H;�H;@�H;��H;��H;N�H;J�H;��H;��H;U�H;��H;��H;��H;x�H;��H;��H;��H;U�H;��H;��H;J�H;H�H;|�H;��H;G�H;�H;C�H;s�H;�H;�H;iI;�I;�I;�I;I;�I;,I;lI;!I;�I;I;�I;��H;��H;Q�H;ߛH;�}H;�dH;�TH;      KIF;oYF;��F;��F;v'G;��G;��G;CH;&�H;C�H;X�H;�I;�I;� I;�I;�I;�I;I;K
I;I;@I;��H;n�H;��H;`�H;7�H;C�H;��H;�H;[�H;G�H;��H;�H;|�H;7�H;�H;�H;�H;3�H;}�H;�H;��H;I�H;[�H;v�H;��H;A�H;>�H;\�H;��H;q�H;��H;<I;I;K
I;�I;�I;�I;�I;� I;�I;�I;[�H;E�H;�H;	CH;��G;��G;�'G;��F;��F;_YF;      �DA;�kA;F�A;`�B;�jC;KaD;y\E;�IF;�G;��G;]NH;.�H;��H;�I;vI;X I;�I;9I;�I;�I;�I;�I;�H;��H;��H;Y�H;�H;0�H;��H;x�H;N�H;e�H;��H;A�H;��H;��H;��H;��H;��H;A�H;��H;c�H;R�H;x�H;��H;,�H;�H;b�H;��H;��H;�H;�I;�I;�I;�I;6I;�I;X I;uI;�I;��H;)�H;[NH;��G;�G;�IF;y\E;@aD;�jC;g�B;H�A;�kA;      �J6;��6;��7;}9;:;;.=;Bj?;Q�A;�C;K2E;��F;M�G;q<H;~�H;��H;�I;G I;I;#I;3I;�I;�I;3I;-�H;��H;��H;?�H;�H;�H;��H;j�H;T�H;v�H;�H;��H;Q�H;-�H;S�H;��H;	�H;x�H;T�H;m�H;��H;�H;�H;@�H;��H;��H;/�H;6I;�I;�I;6I;%I;I;G I;�I;��H;{�H;n<H;I�G;��F;J2E;�C;J�A;Ej?;.=;S;;�9;��7;�6;      p ;�!;�#;�&;�*;�o.;\3;��7;_�;;j?;7kB;�D;jxF;��G;�cH;�H;�
I;�I;QI;aI;I;I;�I;9I;�H;j�H;n�H;�H;��H;��H;��H;g�H;t�H;��H;8�H;�H;��H;�H;5�H;��H;u�H;e�H;��H;��H;��H;	�H;o�H;q�H;�H;9I;�I;I;I;bI;RI;�I;�
I;�H;�cH;��G;jxF;�D;7kB;j?;_�;;��7;^3;�o.;�*;�&;�#;�!;      [t�:� �:%l�:8�;� 
;؄;$z;P$;H�,;��3;�9;�>;�B;2E;�F;RH;խH;��H;I;�I;$I;\I;I;�I;�I;��H; �H;1�H;��H;x�H;��H;��H;q�H;��H;�H;��H;��H;��H;�H;��H;t�H;��H;��H;{�H;��H;.�H;�H;��H;�I;�I;I;]I;$I;�I;	I;��H;ҭH;NH;��F;2E;�B;��>;�9;��3;J�,;P$;z;��;� 
;.�;'l�:y �:       �>:��G:��b:h��:��:�4�:�*�:zi;=�;�a;*;?r3;��:;�!@;��C;�IF;��G;��H;
�H;TI;�I;I;I;�I;�I;5I;��H;k�H;��H;X�H;-�H;��H;|�H;��H;��H;��H;d�H;��H;��H;��H;|�H;��H;/�H;[�H;��H;j�H;��H;9I;�I;�I;I;I;�I;VI;�H;��H;��G;�IF;��C;�!@;��:;<r3;*;�a;:�;|i;�*�:�4�:?��:p��:��b:H�G:      "���օ��uk��� ����@-69��!:�Ȋ:t4�:��:��;�;F�,;��6;��=;��B;m�E;V�G;�|H;u�H;XI;�I;aI;9I;�I;I;cI;(�H;��H;�H;��H;��H;��H;��H;��H;k�H;V�H;m�H;��H;��H;��H;��H;��H;�H;��H;'�H;fI;I;�I;<I;bI;�I;XI;t�H;�|H;S�G;j�E;��B;��=;��6;A�,;�;��;��:n4�:�Ȋ:��!:�,69`��� �uk�؅��      &/��$����x���X���/�� ����0o칈9�9��k:��:)o�:�B;�&;A3;p<;�A;�pE;BtG;�|H;
�H;I;RI;%I;�I;H
I;�I;3 I;-�H;�H;��H;`�H;��H;��H;��H;X�H;E�H;W�H;��H;��H;��H;^�H;��H;�H;*�H;1 I;�I;H
I;�I;&I;QI;I;�H;�|H;?tG;�pE;�A;j<;=3;�&;�B;#o�:��:��k:�9�90o����� ���/���X�!�x�"���      ������q
����4�׻�+��Ȯ���;��lۺ8� � P�9�Ȋ:��:�;!;��0;;;��A;�pE;Q�G;��H;��H;�I;I;5I;�I;�I;UI;��H;"�H;[�H;��H;��H;��H;��H;F�H;�H;G�H;��H;��H;��H;��H;[�H;"�H;��H;SI;�I;�I;.I;I;�I;��H;��H;Q�G;�pE;��A;	;;��0;!;|;��:�Ȋ: P�9L� ��lۺ�;�ʮ���+��6�׻����q
���      ����p8����>�k���O��3/�0B�
�׻ȵ��g�@�NP�� ��$�>:�4�:��;Tb;��/;;;�A;j�E;��G;ҭH;�
I;G I;�I;�I;�I;�I;�I;e�H;�H;��H;z�H;��H;��H;O�H;�H;O�H;��H;��H;x�H;��H;�H;f�H;�I;�I;�I;�I;�I;D I;�
I;ѭH;��G;j�E;�A;;;|�/;Rb;��;�4�: �>:H��VP��j�@�ǵ���׻2B��3/���O�@�k���o8��      :���|�1�ݼ��˼d���,���}��G����D�һ����f���/�h:(׳:��;Mb;��0;m<;��B;�IF;NH;�H;�I;T I;�I;I;7
I;�I; I;�H;6�H;��H;�H;�H;\�H;�H;\�H;�H;�H;��H;2�H;�H;  I;�I;9
I;I;�I;L I;�I;�H;KH;�IF;��B;i<;��0;Mb;�; ׳:\:�/�l������D�һ����G��}��,��d����˼2�ݼ�|�      E�B�LR?��5���&��3��J��ӮҼ!F����?=�"?�.����/��nk�ح�9"׳:��;!;<3;��=;��C; �F;�cH;��H;rI;�I;�I;I;�I;�I;%�H;��H;s�H;c�H;#�H;d�H;�H;e�H;!�H;`�H;r�H;��H;$�H;�I;�I;I;�I;�I;kI;��H;�cH;��F;��C;��=;63;!;��;׳:���9�nk���/�.��"?�@=���!F��ԮҼ�J���3���&��5�MR?�      (��$W��蒐�#�����j�Q`I���&����Dϼ�,���T[�l�lI��d;��nk�x:�4�:�;�&;��6;�!@;2E;��G;��H;�I;� I;/I;�I;�
I;I;V I;��H;��H;��H;A�H;t�H;'�H;w�H;?�H;��H;��H;��H;Q I;I;�
I;�I;,I;� I;�I;��H;��G;2E;�!@;��6;�&;�;�4�:\:�nk�g;�nI��l��T[��,��Dϼ�����&�Q`I���j�#���蒐�$W��      �J�����D��ͽ���'�������L�%��$��;���k����lI����/��/��>:��:�B;C�,;��:;�B;pxF;y<H;��H;�I;oI;�I; I;�I;�I;n�H;Y�H;�H;P�H;�H;N�H;�H;O�H;�H;U�H;k�H;�I;�I; I;�I;mI;�I;��H;t<H;nxF;�B;��:;D�,;�B;��:�>:�/���/�mI������k�	;��%��%����L����'������ͽ�D����      Q�:��*7���,�+���	�q�齂��� W����j�>�/��J���I���k�l�.��f��X���Ȋ:'o�:�;Gr3;�>;	�D;P�G;)�H;�I;!I;�I;iI;b
I;�I;? I;��H;|�H;��H;��H;B�H;��H;��H;z�H;��H;< I;�I;c
I;lI;�I;
!I;�I;!�H;M�G;�D;��>;<r3;�;o�:�Ȋ:X��l��.��m��k��I���J��>�/���j� W������q�齂�	�+���,��*7�      ^���p����2�l���M���,�Xl�Q9ݽ�A���{���5��J��	;���T[�#?�����`P���O�9��:��;*;�9;9kB;��F;[NH;X�H;�I;kI;�I; I;�I;"I;D�H;��H;��H;��H;J�H;��H;��H;��H;C�H;I;�I;I;�I;iI;�I;T�H;TNH;��F;9kB;�9;*;��;��:�O�9bP������$?��T[�	;���J����5��{��A��Q9ݽXl���,���M�2�l����p��      4m־O�Ѿ�>ľ����җ����{��I�+�����V���{�>�/�%���,��@=�D�һn�@�X� ���k:��:�a;��3;j?;R2E;��G;B�H;I;N I;�I;�I;	I;�I;��H;��H;��H;��H;9�H;��H;��H;��H;��H;�I;�I;�I;�I;P I;I;A�H;��G;P2E;j?;��3;�a;��:|�k:\� �n�@�E�һ@=��,��%��>�/��{��V�����+��I���{�ӗ�������>ľO�Ѿ      C\����r5��z ��E۾ֳ�^��y�Z�L?#����A����j�%��Eϼ�����̵���lۺP9�9f4�:B�;D�,;X�;;�C;�G; �H;�I;�!I;�I;%I;	I;sI;$I;��H;��H;��H;�H;��H;��H;��H;!I;qI;I;"I;�I;�!I;I; �H;~G;�C;Y�;;F�,;9�;h4�:(9�9�lۺ̵�������Eϼ%����j��A�����K?#�y�Z�^��ֳ��E۾�z �r5����      E�b��>]���M�Î6�����$���>ľ#q��y�Z�+�Q9ݽ!W����L����#F���G��׻;�Ho�|Ȋ:�i; P$;��7;V�A;�IF;CH;��H;� I;BI;VI;�I;
I;�I;��H;��H;t�H;��H;q�H;��H;��H;~I;I;�I;XI;DI;� I;��H;CH;�IF;S�A;��7; P$;xi;�Ȋ:ho�
;��׻�G�"F�������L�!W��Q9ݽ+�y�Z�#q���>ľ�$�����Î6���M��>]�      p��񲗿���7�y�{�R���)�nv��>ľ^���I�Xl����������&�ԮҼ�}�2B�ή��"���t�!:�*�:"z;Y3;Ij?;s\E;��G;��H;HI;I;mI;�I;WI;�I;��H;��H;C�H;��H;B�H;��H;��H;�I;WI;�I;nI;I;KI;��H;��G;r\E;Ij?;^3; z;�*�:��!:&���ή��2B��}�ԮҼ��&��������Xl��I�^���>ľnv���)�{�R�7�y����񲗿      �˿�<ƿqL��@1����>]���)��$��ֳ���{���,�q��'��Q`I��J���,���3/�,��� ��,69�4�:Є;�o.;.=;?aD;��G;P�H;�I;!I;BI;,I;�	I;�I;� I;��H;��H;C�H;��H;�H;� I;�I;�	I;)I;AI;!I;�I;S�H;��G;=aD;.=;�o.;Є;�4�: -69� �,���3/��,���J��Q`I�'��q�齥�,���{�ֳ��$����)��>]��@1��qL���<ƿ      ����<���T[忶˿�T���{�R�����E۾ӗ����M���	������j��3�d����O�=�׻��/�H��=��:� 
;�*;L;;�jC;}'G;ћH;�I;�!I;�I;vI;�
I;�I;�I;�H;��H;��H;��H;!�H;I;�I;�
I;tI;�I;�!I;�I;ڛH;�'G;�jC;O;;�*;� 
;5��:@����/�<�׻��O�d���3���j������	���M�ӗ���E۾���{�R���T���˿T[�<���      O�6��t����˿@1��7�y�Î6��z �����2�l�+��ͽ#�����&���˼@�k�%�����X��� �v��:6�;�&;|9;k�B;��F;�}H;�	I;."I;I;�I;xI;TI;%I;��H;�H;b�H;��H;��H;!I;RI;{I;�I;I;2"I;�	I;�}H;��F;j�B;}9;�&;8�;n��:�� ���X�"���@�k���˼��&�#����ͽ+�2�l������z �Î6�7�y�A1���˿���t�6��      ��*��g&��#�t�T[�qL�������M�r5��>ľ����,��D�蒐��5�2�ݼ���q
��x�(uk���b:!l�:�#;×7;T�A;��F;�dH;�I;!"I;�I;EI;I;�I;�I;��H;X�H;��H;R�H;��H;�I;�I;I;AI;�I;%"I;�I;�dH;��F;Q�A;7;�#;%l�:��b:uk��x��q
���2�ݼ�5�蒐��DὫ�,����>ľr5���M����qL��T[�t��#��g&�      ��8��4��g&�6��<����<ƿ񲗿�>]����O�Ѿ�p���*7����%W��LR?� }�r8�������؅����G:q �:�!;�6;�kA;dYF;�TH;C�H;�!I;�I;�I;dI;&I;�I;; I;��H;��H;��H;< I;�I;)I;hI;�I;�I;�!I;G�H;�TH;sYF;�kA;�6;�!;q �:|�G:̅�������r8�� }�LR?�%W�����*7��p��O�Ѿ����>]�񲗿�<ƿ<���6���g&��4�      �Aq���i���U�F:�@�����<���u���{A�d5�� ��~^Z�����A���]�����d��L",��5����Ѻ ��9���:�;[Y4;H�@;LVF;~�H;�GI;�bI;OI;:I;�)I;I;{I;�I;~I;�I;zI;�I;}I;I;�)I;:I;OI;�bI;�GI;��H;XVF;E�@;ZY4;�;���: ��9��Ѻ�5��L",��d������]��A�����~^Z�� ��d5�{A�u���<�������@�F:���U���i�      ��i���b�Z�O�.5�1i�������������q<�����e��`
V�GE	�!���IY�j9�D�����(��R���ȺX�:N��:�;?�4;>�@;hF;��H;II;ubI;�NI;�9I;�)I;�I;ZI;�I;[I;YI;WI;�I;XI;�I;�)I;�9I;�NI;zbI;II;��H;*hF;>�@;=�4;ޔ;J��:T�: �Ⱥ�R����(�D���j9��IY�!��GE	�`
V��e������q<������������1i�.5�Z�O���b�      ��U�Z�O�H-?�.�'���M�ῴ欿a�{�ea/���뾝���I����d���ZN�\5������>H�f ��p���|�":��:x�;��5;�`A;��F;J�H;MI;�aI;�MI;�8I;�(I;@I;�I;7I;I;I;�I;7I;�I;BI;�(I;�8I;�MI;�aI;MI;L�H;��F;�`A;��5;w�;��:|�":h���g ��=H�����\5���ZN�d������I�������ea/�a�{��欿M����.�'�H-?�Z�O�      F:�.5�.�'��������jȿ���l$_���W�Ҿܕ���6�����*���`=�=�漮)��JG�)6����� �Q:��:�/";�7;^&B;��F;��H;�RI;�`I;uKI;7I;�'I;;I;I;�I;oI;n
I;jI;�I;I;<I;�'I;7I;zKI;�`I;�RI;��H;��F;^&B;�7;�/";��:�Q:���(6��IG��)��<���`=��*������6�ܕ��W�Ҿ��l$_����jȿ�������.�'�.5�      @�1i�������I�ѿk��� ���q<��:��a����q����Wн罅���'�Ub̼�zl��.��Q�X�l����:��;Ύ&;ū9;#C;9MG;��H;6YI;�^I;�HI;�4I;�%I;�I;I;�I;�
I;�	I;�
I;�I;I;�I;�%I;�4I;�HI;�^I;9YI;��H;BMG;$C;«9;Ύ&;��;��:T��P�X��.���zl�Ub̼��'�罅��Wн����q��a���:��q<� ��k���I�ѿ������1i�      �������L��jȿk���������O���{]׾z����I�����A��>�d�n�~֮�RH��jλT�$� )�l��:CN;��+;�<;�3D;��G;�I;~^I;j[I;�DI; 2I;�#I;BI;�I;[I;�	I;�I;�	I;]I;�I;CI;�#I; 2I;�DI;k[I;�^I;�I;��G;�3D;�<;��+;CN;f��:�(�Q�$��jλRH�~֮�n�>�d��A������I�z���{]׾����O�����k���jȿL�Ῡ��      <��������欿��� ����O��x����� ���l���"��ܽ���`=����v���k"�1R��Jۺ���9�?�:XL;~�0;��>;�ME;H#H;�%I;�aI;�VI;�@I;�.I;;!I;=I;I;	I;LI;�I;JI;
I;I;@I;=!I;�.I;�@I;�VI;�aI;�%I;N#H;�ME;��>;�0;ZL;�?�:Г�9Dۺ/R���k"�v������`=����ܽ��"��l�� ����뾁x���O� ������欿����      u�������a�{�l$_��q<�������}��w��	�6�����!���h����㷾�� d��.���^e�I[���Z:Z��:�, ;��5;�A;�VF;��H;�@I;nbI;�QI;�;I;;+I;jI;I;6I;{	I;�I;+I;�I;	I;7I;I;kI;;+I;�;I;�QI;sbI;�@I;��H;�VF;�A;��5;�, ;X��:��Z:I[��^e��.��� d�ⷾ�����h�!������	�6�w���}��������q<�l$_�a�{�����      {A��q<�ea/����:�{]׾� ��w��>�DE	�����ڽ����3�_�꼚���",��W��f���Q�p��:�M
;�f);��:;$@C;�?G;O�H;ETI;�_I;#KI;�6I;L'I;dI;�I;:I;�I;mI;�I;lI;�I;;I;�I;hI;O'I;�6I;*KI;�_I;GTI;R�H;�?G;$@C;��:;�f);�M
;���: Q�c���W��",�����^�꼘�3�ڽ������DE	�>�w��� ��{]׾�:���ea/��q<�      d5�������W�Ҿ�a��z����l�	�6�DE	���Ƚk���aG����e֮��W����t�k�<���c,:~��:��;��1;<�>;=E;�G;I;#_I;@ZI;2DI;�1I;/#I;CI;�I;
I;I;�I;I;�I;I;
I;�I;BI;2#I;�1I;9DI;GZI;&_I;I;&�G;=E;A�>;��1;��;���:�c,:0��l�k�����W�d֮�����aG�k����ȽDE	�	�6��l�z����a��W�Ҿ������      � ���e�����ە����q��I���"���������k���ZN�[�"¼Q�y��$��Q���� � |X���:0;#�&;�w8;k B;��F;АH;T@I;�aI;iRI;=I;,I;�I;�I;[I;�I;3I;I;eI;I;7I;�I;\I;�I;�I;,I;=I;pRI;�aI;T@I;ؐH;��F;o B;�w8;%�&;"0;��: dX��� ��Q���$�O�y�!¼[��ZN�k������������"��I���q�ە������e��      ~^Z�`
V��I��6�������ܽ!��ڽ���aG�[��ȼ�)��~�(�j��QG5������Z:�:S;'1;��=;��D;,�G;��H;�XI;^I;|II;�5I;�&I;�I;�I;�
I;�I;KI;` I;��H;a I;MI;�I;�
I;�I;�I;�&I;�5I;�II;^I;�XI;��H;.�G;��D;��=;'1;S;�:��Z:���KG5�h��}�(��)��
�ȼZ��aG�ڽ��!���ܽ������6��I�`
V�      ���GE	��������Wн�A�����h���3����!¼�)��3x/��һy�X��#��x�9F��:�>;+f);b`9;Z&B;��F;d}H;�6I;NaI;�UI;^@I;�.I;� I;FI;'I;�I;LI;P I;��H;��H;��H;P I;NI;�I;(I;KI;!I;�.I;d@I;�UI;NaI;�6I;d}H;��F;a&B;e`9;9f);�>;H��:��9r#��s�X��һ1x/��)�� ¼�����3��h��󑽡A���Wн��콺��GE	�      �A��!��c���*��潅�?�d��`=����^��d֮�O�y�~�(��һ�]e�����@�f9���:2�;>1";�4;�m?;�E;��G;d�H;�WI;}^I;
KI;o7I;�'I;�I;"I;�
I;#I;I;k�H;��H;;�H;��H;k�H;I;!I;�
I;(I;�I;�'I;u7I;KI;z^I;�WI;e�H;��G;�E;�m?;�4;G1";2�;���:p�f9��]e��һ}�(�N�y�d֮�]�꼘���`=�>�d�罅��*��c��!��      �]��IY��ZN��`=���'�n����᷾������W��$�j��z�X������9n��:Q��:l�;��0;��<;M�C;G;��H;�?I;#aI;�TI;<@I;/I;T!I;�I;I;xI;�I;��H;|�H;�H;��H;�H;|�H;��H;�I;vI;I;�I;Z!I;/I;<@I;�TI;'aI;�?I;��H;"G;R�C;��<;��0;l�;c��:t��:9�u�X�h���$��W�����ⷾ����m���'��`=��ZN��IY�      ���i9�[5��:��Ub̼~֮�u��� d�",�����Q��OG5��#��@�f9p��:��:�;��-;��:;�KB;8VF;KH;�I;�\I;\I;�HI;6I;'I;I;�I;
I;AI;��H;��H;��H;Z�H;��H;X�H;��H;��H;��H;AI;
I;�I;I;!'I;6I;�HI;\I;�\I;�I;KH;<VF;�KB;��:;��-;�;��:x��:`�f9�#��KG5��Q�����",�� d�u��|֮�Vb̼;��[5��i9�      �d��C��������)���zl�RH��k"�~.���W��i�k��� ������9���:]��:�;�-;ɫ9;AaA;��E;#�G;r�H;�RI;`I;�OI;�<I;�,I;�I;-I;I;xI;SI;��H;��H;��H;��H;a�H;��H;��H;��H;��H;TI;I;I;/I;�I;�,I;�<I;�OI;`I;�RI;v�H;(�G;��E;EaA;ƫ9;�-;�;e��:���:��9����� �g�k��W��|.���k"�RH��zl��)������B���      E",���(�=H�FG��.���jλ*R���^e�c��*�� lX���Z::��:.�;i�;��-;«9;tA;�cE;�G;��H;LGI;�`I;�UI;7BI;�1I;�#I;�I;�I;�I;�I;��H;H�H;��H;�H;�H;��H;�H;	�H;��H;E�H;��H;�I;�I;�I;�I;�#I;�1I;>BI;�UI;�`I;QGI;��H;"�G;�cE;tA;ȫ9;��-;l�;2�;@��:��Z: HX�(��]���^e�-R���jλ�.��GG�;H���(�      �5���R��f ��&6��W�X�F�$�6ۺ�H[� Q��c,:��:�:�>;D1";��0;��:;AaA;�cE;��G;p�H;�=I;*`I;pYI;�FI;�5I;�'I;�I;�I;�
I;�I;��H;�H;�H;��H;�H;��H;<�H;��H;~�H;��H;�H;�H;��H;�I;�
I;�I;�I;�'I;�5I;�FI;jYI;.`I;�=I;v�H;��G;�cE;GaA;��:;��0;D1";�>;�:��:�c,:�
Q��H[�>ۺL�$�T�X�+6��f ���R��      ��Ѻ�Ⱥb������x���(��9��Z:z��:���:!0;S;0f);�4;��<;�KB;��E;$�G;u�H;[:I;N_I;~[I;!JI;9I;�*I;�I;�I;�I;[I;I;��H;��H;�H;/�H;��H;7�H;��H;3�H;��H;/�H;�H;��H;��H;I;[I;I;�I;�I;�*I;9I;JI;�[I;S_I;]:I;w�H; �G;��E;�KB;��<;�4;0f);S;"0;���:���:��Z:Г�9�(�\�����x���*�Ⱥ      0��9�:�":�Q:��:j��:v?�:T��:�M
;��; �&;'1;_`9;�m?;N�C;<VF;%�G;��H;�=I;L_I;\I;�KI;;I;�,I;� I;�I;�I;�I;GI;��H;5�H;x�H;5�H;��H;��H;��H;��H;��H;��H;��H;4�H;t�H;7�H;��H;FI;�I;�I;�I;� I;�,I;;I;�KI;\I;N_I;�=I;��H;&�G;<VF;P�C;�m?;b`9;'1;'�&;��;�M
;P��:�?�:^��:��:��Q:0�":�:      ���:d��:��:��:��;CN;WL;�, ;�f);��1;�w8;��=;^&B;�E;"G;KH;v�H;RGI;1`I;�[I;�KI;�;I;�-I;/"I;,I;I;	I;aI;��H;��H;��H;j�H;y�H;�H;F�H;��H;e�H;��H;C�H;�H;y�H;h�H;��H;��H;��H;dI;	I;I;0I;."I;�-I;�;I;�KI;�[I;/`I;QGI;y�H;KH;#G;�E;]&B;��=;�w8;��1;�f);�, ;[L;>N;��;��:��:H��:      1�;ݔ;p�;�/";��&;��+;��0;��5;��:;B�>;u B;��D;��F;��G;��H;�I;SI;�`I;pYI; JI;;I;�-I;�"I; I;�I;�	I;*I;G�H;o�H;W�H;��H;��H;��H;��H;��H;��H;a�H;��H;��H;��H;��H;��H;��H;W�H;k�H;L�H;&I;�	I;�I;�I;�"I;�-I;;I; JI;pYI;�`I;�RI;�I;��H;��G;��F;��D;x B;>�>;��:;��5;��0;��+;ю&;�/";l�;Ô;      TY4;D�4;��5;�7;��9;�<;��>;�A;@C;<E;��F;,�G;`}H;d�H;�?I;�\I;`I;�UI;�FI;�8I;�,I;)"I;�I;!I;Y
I;�I;��H;��H;��H;��H;��H;��H;��H;��H;��H;��H;g�H;��H;��H;��H;��H;��H;��H;��H;��H;��H;��H;�I;\
I; I;�I;+"I;�,I;�8I;�FI;�UI;`I;�\I;�?I;a�H;b}H;,�G;��F;:E;@C;�A;��>;�<;��9;��7;��5;:�4;      b�@;:�@;�`A;X&B;C;4D;�ME;�VF;�?G;%�G;ڐH;��H;�6I;�WI;*aI;'\I;�OI;CBI;�5I;�*I;� I;3I;�I;b
I;�I; I;0�H;��H;$�H;��H;��H;��H;L�H;{�H;��H;��H;f�H;��H;��H;{�H;H�H;��H;��H;��H;�H;��H;,�H; I;�I;`
I;�I;4I;� I;�*I;�5I;ABI;�OI;*\I;)aI;�WI;�6I;��H;ڐH;#�G;�?G;�VF;�ME;�3D;#C;W&B;�`A;:�@;      JVF;*hF;��F;��F;-MG;��G;K#H;��H;P�H;I;W@I;�XI;PaI;�^I;�TI;�HI;�<I;�1I;�'I;�I;�I;I;�	I;�I; I;>�H;�H;X�H;��H;��H;w�H;H�H;=�H;x�H;�H;��H;}�H;��H;�H;z�H;=�H;E�H;y�H;��H;��H;X�H;�H;A�H; I;�I;�	I;I;�I;�I;�'I;�1I;�<I;�HI;�TI;�^I;PaI;�XI;[@I;I;O�H;��H;M#H;��G;CMG;��F;��F;$hF;      ��H;��H;A�H;��H;��H;�I;�%I;�@I;GTI;&_I;�aI;^I;�UI;
KI;<@I;6I;�,I;�#I;�I;�I;�I;	I;,I;��H;,�H;�H;H�H;�H;.�H;n�H;&�H;�H;8�H;��H;8�H;��H;��H;��H;5�H;��H;8�H;�H;(�H;l�H;(�H;�H;@�H;�H;.�H;��H;*I;	I;�I;�I;�I;�#I;�,I;	6I;:@I;KI;�UI;^I;�aI;#_I;DTI;�@I;�%I;�I;��H;��H;A�H;��H;      �GI;II;MI;�RI;*YI;�^I;�aI;obI;�_I;GZI;oRI;�II;^@I;u7I;/I;!'I;�I;�I;�I;�I;�I;aI;E�H;��H;��H;R�H;�H;�H;|�H;&�H;��H;�H;e�H;��H;t�H;@�H;4�H;>�H;t�H;��H;d�H;�H;��H;#�H;w�H;�H;�H;V�H;��H;��H;E�H;aI;�I;�I;�I;�I;�I;"'I;/I;r7I;]@I;�II;pRI;EZI;�_I;kbI;�aI;u^I;6YI;�RI;MI;II;      �bI;qbI;�aI;�`I;�^I;h[I;WI;�QI;KI;6DI;=I;�5I;�.I;�'I;Z!I;I;5I;�I;�
I;`I;NI;��H;m�H;��H;�H;��H;$�H;z�H;!�H;��H;��H;8�H;��H;)�H;��H;��H;��H;��H;��H;*�H;��H;5�H;��H;��H;�H;y�H; �H;��H;�H;��H;n�H;��H;JI;\I;�
I;�I;4I;I;W!I;�'I;�.I;�5I;=I;7DI;$KI;�QI;WI;a[I;�^I;�`I;�aI;obI;      OI;�NI;�MI;qKI;�HI;�DI;�@I;�;I;�6I;�1I;,I;�&I; !I;�I;�I;�I;I;�I;�I;I;��H;��H;V�H;��H;��H;��H;k�H;(�H;�H;��H;#�H;|�H;��H;��H;F�H; �H;�H; �H;A�H;��H;��H;{�H;#�H;��H;��H;%�H;e�H;��H;��H;��H;X�H;��H;��H;I;�I;�I;I;�I;�I;�I; !I;�&I;,I;�1I;�6I;�;I;�@I;�DI;�HI;uKI;�MI;�NI;      :I;�9I;�8I;%7I;�4I; 2I;�.I;H+I;P'I;6#I;�I;�I;NI;.I;I;!
I;�I;�I;��H;��H;?�H;��H;��H;��H;��H;u�H;&�H;�H;��H;)�H;��H;��H;\�H;	�H;��H;��H;��H;��H;��H;�H;\�H;��H;��H;&�H;��H;�H;"�H;v�H;��H;��H;��H;��H;9�H;��H;��H;�I;�I;"
I;I;+I;OI;�I;�I;6#I;R'I;E+I;�.I;2I;�4I;%7I;�8I;�9I;      �)I;�)I;�(I;�'I;�%I;�#I;=!I;mI;jI;EI;�I;�I;+I;�
I;|I;FI;[I;��H;�H;��H;�H;j�H;��H;��H;��H;@�H;	�H;�H;:�H;}�H;��H;t�H;��H;��H;v�H;M�H;8�H;P�H;q�H;��H;��H;t�H;��H;|�H;5�H;	�H;�H;A�H;��H;��H;��H;l�H;x�H;��H;�H;��H;\I;II;|I;�
I;(I;�I;�I;EI;gI;iI;D!I;�#I;�%I;�'I;�(I;�)I;      $I;�I;LI;?I;�I;9I;;I;I;�I;�I;\I;�
I;�I;'I;�I;��H;��H;K�H;#�H;�H;@�H;{�H;��H;��H;I�H;9�H;6�H;i�H;��H;��H;V�H;��H;��H;T�H;�H;�H;�H;�H;�H;W�H;��H;��H;V�H;��H;��H;g�H;4�H;7�H;L�H;��H;��H;{�H;9�H;�H;#�H;L�H;��H; I;�I;&I;�I;�
I;_I;�I;�I;	I;=I;4I;�I;:I;UI;�I;      vI;\I;�I;I;I;�I;I;<I;<I;	
I;�I;�I;UI;#I;��H;��H;��H;��H;��H;5�H;��H;�H;��H;��H;r�H;q�H;��H;��H;,�H;��H;�H;��H;W�H;�H;��H;��H;��H;��H;��H;�H;W�H;��H;�H;��H;&�H;��H;��H;s�H;w�H;��H;��H;�H;��H;-�H;��H;��H;��H;��H;��H;!I;RI;�I;�I;
I;>I;7I;
I;�I;I;I;�I;eI;      �I;�I;@I;�I;�I;WI;I;�	I;�I;I;?I;YI;[ I;w�H;��H;��H;��H;�H;��H;��H;��H;B�H;��H;��H;��H;��H;.�H;r�H;��H;D�H;��H;s�H;�H;��H;��H;��H;��H;��H;��H;��H;�H;w�H;��H;?�H;��H;o�H;0�H;��H;��H;��H;��H;@�H;��H;��H;�H;�H;��H;��H;��H;w�H;[ I;VI;?I;I;�I;�	I;I;WI;�I;�I;@I;�I;      ~I;dI;I;nI;�
I;�	I;TI;�I;mI;�I;$I;g I;��H;��H;�H;X�H;��H;�H;��H;4�H;��H;��H;��H;u�H;��H;��H;��H;>�H;��H;"�H;��H;M�H;�H;��H;��H;}�H;|�H;��H;��H;��H;�H;P�H;��H;�H;��H;;�H;��H;��H;��H;x�H;��H;��H;��H;2�H;��H;�H;��H;\�H;�H;��H;��H;d I;%I;�I;oI;�I;[I;�	I;�
I;oI; I;rI;      �I;WI;I;r
I;�	I;�I;�I;3I;�I;!I;oI;��H;�H;C�H;��H;��H;k�H;��H;A�H;��H;��H;g�H;]�H;[�H;a�H;r�H;��H;7�H;��H; �H;��H;8�H;�H;��H;��H;w�H;��H;z�H;��H;��H;�H;;�H;��H;�H;��H;3�H;��H;v�H;e�H;\�H;c�H;g�H;��H;��H;?�H;��H;j�H;��H;��H;E�H;��H;��H;oI;!I;�I;3I;�I;�I;�	I;w
I;I;dI;      ~I;eI; I;nI;�
I;�	I;SI;�I;mI;�I;"I;h I;��H;��H;�H;X�H;��H;�H;��H;4�H;��H;��H;��H;u�H;��H;��H;��H;>�H;��H;!�H;��H;M�H;�H;��H;��H;}�H;|�H;��H;��H;��H;�H;P�H;��H;�H;��H;:�H;��H;��H;��H;w�H;��H;��H;��H;2�H;��H;�H;��H;\�H;�H;��H;��H;d I;$I;�I;oI;�I;ZI;�	I;�
I;uI;I;lI;      �I;�I;;I;�I;�I;TI;I;�	I;�I;I;AI;YI;[ I;w�H;��H;��H;��H;�H;��H;��H;��H;C�H;��H;��H;��H;��H;.�H;r�H;��H;C�H;��H;s�H;�H;��H;��H;��H;��H;��H;��H;��H;�H;v�H;��H;=�H;��H;n�H;0�H;�H;��H;��H;��H;B�H;��H;��H;�H;�H;��H;��H;��H;u�H;[ I;XI;?I;I;�I;�	I;I;SI;�I;�I;AI;�I;      vI;[I;�I;I;I;�I;I;?I;?I;	
I;�I;�I;SI;#I;��H;��H;��H;��H;��H;4�H;��H;�H;��H;��H;u�H;s�H;��H;��H;-�H;��H;�H;��H;W�H;�H;��H;��H;��H;��H;��H;�H;X�H;��H;�H;��H;&�H;��H;��H;v�H;u�H;��H;��H;�H;��H;.�H;��H;��H;��H;��H;��H;!I;RI;�I;�I;	
I;>I;<I;I;�I;	I;I;�I;\I;      !I;�I;NI;8I;�I;=I;;I;I;�I;�I;_I;�
I;�I;'I;�I;  I;��H;K�H;!�H;�H;?�H;|�H;��H;��H;L�H;5�H;4�H;i�H;��H;��H;U�H;��H;��H;T�H;�H;�H;�H;�H;�H;U�H;��H;��H;V�H;��H;��H;e�H;4�H;9�H;I�H;��H;��H;|�H;8�H;�H; �H;K�H;��H; I;�I;&I;�I;�
I;\I;�I;�I;I;AI;8I;�I;CI;WI;�I;      �)I;�)I;�(I;�'I;�%I;�#I;B!I;kI;hI;FI;�I;�I;)I;�
I;I;FI;[I;��H;
�H;��H;�H;l�H;��H;��H;��H;A�H;�H;�H;<�H;|�H;��H;q�H;��H;��H;v�H;I�H;8�H;M�H;q�H;��H;��H;t�H;��H;{�H;5�H;�H;�H;B�H;��H;��H;��H;l�H;y�H;��H;
�H;��H;\I;HI;{I;�
I;)I;�I;�I;FI;hI;kI;C!I;�#I;�%I;�'I;�(I;�)I;      :I;�9I;�8I;7I;�4I;!2I;�.I;G+I;R'I;4#I;�I;�I;OI;/I;I;!
I;�I;�I;��H;��H;@�H;��H;��H;��H;��H;s�H;#�H;�H;��H;'�H;��H;��H;[�H;�H;��H;��H;��H;��H;��H;�H;\�H;��H;��H;%�H;��H;��H;#�H;w�H;��H;��H;��H;��H;9�H;��H;��H;�I;�I;!
I;I;,I;NI;�I;�I;4#I;R'I;G+I;�.I;2I;�4I;)7I;�8I;�9I;      $OI;�NI;�MI;zKI;xHI;�DI;�@I;�;I;�6I;�1I;,I;�&I;� I;�I;�I;�I;I;�I;�I;I;��H;��H;V�H;��H;��H;��H;k�H;&�H;�H;��H;#�H;{�H;��H;��H;C�H;�H;�H; �H;A�H;��H;��H;|�H;#�H;��H;��H;%�H;h�H;��H;��H;��H;Z�H;��H;��H;I;�I;�I;I;�I;�I;�I;� I;�&I;,I;�1I;�6I;�;I;�@I;�DI;�HI;�KI;�MI;�NI;      �bI;obI;�aI;�`I;x^I;l[I;�VI;�QI;)KI;3DI;=I;�5I;�.I;�'I;^!I;I;4I;�I;�
I;]I;OI;��H;m�H;��H;�H;��H;$�H;z�H;!�H;��H;��H;7�H;��H;)�H;��H;��H;��H;��H;��H;)�H;��H;7�H;��H;��H;�H;w�H;!�H;��H;�H;��H;o�H;��H;KI;\I;�
I;�I;4I;I;Z!I;�'I;�.I;�5I;=I;3DI;#KI;�QI;WI;h[I;�^I;�`I;�aI;lbI;      �GI;II;MI;�RI;$YI;�^I;�aI;sbI;�_I;GZI;mRI;�II;]@I;v7I;/I;#'I;�I;�I;�I;�I;�I;dI;E�H;��H;��H;O�H;�H;�H;}�H;#�H;��H;	�H;b�H;��H;r�H;;�H;4�H;>�H;q�H;��H;e�H;�H;�H;%�H;w�H;�H;
�H;U�H;��H;��H;H�H;cI;�I;�I;�I;�I;�I;!'I;/I;r7I;]@I;�II;mRI;DZI;�_I;lbI;�aI;|^I;6YI;�RI;MI;II;      ��H;ėH;A�H;��H;��H;�I;�%I;�@I;HTI;$_I;�aI;^I;�UI;	KI;A@I;6I;�,I;�#I;�I;�I;�I;	I;)I;��H;.�H;�H;F�H;�H;.�H;k�H;&�H;�H;6�H;��H;5�H;��H;��H;��H;4�H;��H;6�H;�H;(�H;k�H;(�H;�H;D�H;�H;,�H;��H;-I;	I;�I;�I;�I;�#I;�,I;6I;>@I;KI;�UI;^I;�aI;#_I;ETI;�@I;�%I;�I;��H;��H;E�H;��H;      <VF;(hF;��F;��F;1MG;��G;D#H;��H;T�H;I;Y@I;�XI;RaI;�^I;�TI;�HI;�<I;�1I;�'I;�I;�I;I;�	I;�I; I;;�H;�H;\�H;��H;��H;w�H;G�H;<�H;z�H;�H;��H;~�H;��H;�H;x�H;=�H;G�H;z�H;��H;��H;X�H;�H;B�H; I;�I;�	I;I;�I;�I;�'I;�1I;�<I;�HI;�TI;�^I;PaI;�XI;Z@I;I;L�H;��H;H#H;��G;@MG;��F;��F;hF;      a�@;:�@;�`A;Q&B;C;4D;�ME;�VF;�?G;#�G;ڐH;��H;�6I;�WI;.aI;+\I;�OI;EBI;�5I;�*I;� I;4I;�I;b
I;�I; I;-�H;��H;"�H;��H;��H;��H;H�H;z�H;��H;��H;e�H;��H;��H;{�H;I�H;��H;�H;��H;�H;��H;-�H; I;�I;`
I;�I;5I;� I;�*I;�5I;ABI;�OI;*\I;-aI;�WI;�6I;��H;֐H;%�G;�?G;�VF;�ME;�3D; C;X&B;�`A;8�@;      2Y4;.�4;��5;�7;��9;�<;��>;�A;!@C;9E;��F;.�G;b}H;c�H;�?I;�\I;`I;�UI;�FI;�8I;�,I;("I;�I;!I;\
I;�I;��H;��H;��H;��H;��H;��H;��H;��H;��H;��H;g�H;��H;��H;��H;��H;��H;��H;��H;��H;��H;��H;�I;X
I;#I;�I;+"I;�,I; 9I;�FI;�UI;`I;�\I;�?I;a�H;`}H;+�G;��F;9E;@C;�A;��>;�<;ɫ9;%�7;��5;�4;      �;۔;h�;�/";��&;��+;��0;��5;��:;B�>;q B;��D;��F;��G;��H;�I;SI;�`I;qYI; JI;;I;�-I;�"I;�I;�I;�	I;'I;K�H;q�H;T�H;��H;��H;��H;��H;��H;��H;d�H;��H;��H;��H;��H;��H;��H;X�H;k�H;H�H;)I;�	I;�I;�I;�"I;�-I;;I;!JI;qYI;�`I;SI;�I;��H;��G;��F;��D;q B;A�>;��:;��5;��0;��+;��&;�/";f�;;      ���:d��:��:��:��;IN;\L;�, ;�f);��1;�w8;��=;]&B;�E;&G;KH;x�H;SGI;/`I;�[I;�KI;�;I;�-I;."I;3I;
I;	I;dI;��H;��H;��H;j�H;y�H;�H;B�H;��H;g�H;��H;B�H;�H;y�H;i�H;��H;��H;��H;aI;	I;I;-I;2"I;�-I;�;I;�KI;�[I;/`I;RGI;v�H;KH;"G;�E;]&B;��=;�w8;��1;�f);�, ;WL;4N;��;��:��:P��:      ���9`�:X�":�Q:��:r��:|?�:R��:�M
;��;%�&;'1;c`9;�m?;T�C;>VF;&�G;��H;�=I;N_I;\I;�KI;;I;�,I;� I;�I;�I;�I;HI;��H;6�H;x�H;5�H;��H;��H;��H;��H;��H;��H;��H;5�H;u�H;7�H;��H;FI;�I;�I;�I;� I;�,I;;I;�KI;\I;O_I;�=I;��H;%�G;<VF;R�C;�m?;``9;'1;%�&;��;�M
;Z��:�?�:j��:��:�Q:t�":$�:      ��Ѻ �Ⱥj������p��`(��9��Z:���:���:"0;S;3f);�4;��<;�KB;��E;$�G;v�H;]:I;U_I;�[I;!JI;9I;�*I;�I;�I;�I;]I;I;��H;��H;�H;2�H;��H;3�H;��H;6�H;��H;-�H;�H;��H;��H;I;[I;�I;�I;�I;�*I;9I; JI;[I;Q_I;\:I;u�H; �G;��E;�KB;��<;�4;0f);S;"0;���:���:��Z:ؓ�9�(�`�����n����Ⱥ      �5���R��f ��'6��W�X�E�$�<ۺ�H[� 
Q��c,:��:�:�>;D1";��0;��:;DaA;�cE;��G;v�H;�=I;.`I;qYI;�FI;�5I;�'I;�I;�I;�
I;�I;��H;�H;�H;��H;�H;��H;>�H;��H;{�H;��H;�H;�H;��H;�I;�
I;�I;�I;�'I;�5I;�FI;nYI;+`I;�=I;u�H;��G;�cE;BaA;��:;��0;A1";�>;�:��:�c,:�
Q��H[�>ۺI�$�X�X�&6��i ���R��      H",���(�>H�FG��.���jλ*R���^e�\��(�� TX���Z:B��:2�;o�;��-;ƫ9;tA;�cE;"�G;��H;RGI;�`I;�UI;?BI;�1I;�#I;�I;�I;�I;�I;��H;H�H;��H;
�H;�H;��H;�H;�H;��H;H�H;�H;�I;�I;�I;�I;�#I;�1I;7BI;�UI;�`I;QGI;��H; �G;�cE;sA;ë9;��-;l�;.�;<��:��Z: TX�0��_���^e�,R���jλ�.��GG�@H���(�      �d��B��������)���zl�RH��k"�{.���W��g�k��� ������9���:g��:�;�-;ɫ9;BaA;��E;,�G;x�H;�RI;`I;�OI;�<I;�,I;�I;4I;I;~I;UI;��H;��H;��H;��H;c�H;��H;��H;��H;��H;QI;~I;I;/I;�I;�,I;�<I;�OI;`I;SI;u�H;"�G;��E;AaA;ȫ9;�-;�;c��:���:��9����� �j�k��W��|.���k"�RH��zl��)������B���      ���i9�[5��:��Ub̼|֮�u��� d�",�����Q��JG5��#��p�f9|��:��:�;��-;��:;�KB;@VF;KH;�I;�\I;#\I;�HI;6I;'I;I;�I;
I;CI;��H;��H;��H;X�H;��H;X�H;��H;��H;��H;?I;
I;�I;I;'I;6I;�HI;\I;�\I;�I;KH;4VF;�KB;��:;��-;�;��:t��:`�f9�#��QG5��Q�����",�� d�v��}֮�Vb̼;��\5��i9�      �]��IY��ZN��`=���'�m����᷾������W��$�h��u�X�����`9|��:]��:l�;��0;��<;W�C;#G; �H;�?I;*aI;�TI;<@I;/I;\!I;�I;I;yI;�I;��H;}�H;�H;��H;�H;z�H;��H;�I;uI;I;�I;[!I;/I;;@I;�TI;%aI;�?I;��H;"G;K�C;��<;��0;f�;]��:n��:�9����y�X�j���$��W�����ⷾ����m���'��`=��ZN��IY�      �A��!��c���*��潅�>�d��`=����]��d֮�N�y�|�(��һ�]e�ꄮ���f9���:2�;D1";�4;�m?;�E;��G;j�H;�WI;�^I;
KI;t7I;�'I;�I;)I;�
I;!I;I;m�H;��H;;�H;��H;j�H;I;!I;�
I;%I;�I;�'I;r7I;	KI;|^I;�WI;g�H;��G;�E;�m?;�4;@1";0�;���:`�f9�����]e��һ~�(�N�y�d֮�^�꼘���`=�>�d�罅��*��c��!��      ���GE	��������Wн�A�����h���3���� ¼�)��1x/��һr�X�t#����9F��:�>;2f);j`9;_&B;��F;j}H;�6I;PaI;�UI;a@I;�.I;� I;JI;(I;�I;PI;Q I;��H;��H;��H;P I;NI;�I;%I;HI; !I;�.I;`@I;�UI;LaI;�6I;d}H;��F;]&B;_`9;3f);�>;<��:��9|#��u�X��һ2x/��)��!¼�����3��h��󑽡A���Wн��콺��GE	�      ~^Z�`
V��I��6�������ܽ!��ڽ���aG�Z�
�ȼ�)��}�(�h��KG5������Z:�:S;'1;��=;��D;2�G;��H;�XI;^I;~II;�5I;�&I;�I;�I;�
I;�I;MI;` I;��H;a I;KI;�I;�
I;�I;�I;�&I;�5I;~II;^I;�XI;��H;.�G;��D;��=;'1;S;�:��Z:���QG5�i��~�(��)���ȼ[��aG�ڽ��!���ܽ������6��I�`
V�      � ���e�����ە����q��I���"���������k���ZN�[�!¼P�y��$��Q���� � pX���:0;,�&;�w8;r B;��F;ؐH;Y@I;�aI;oRI;=I;,I;�I;�I;\I;�I;4I;I;eI;I;4I;�I;\I;�I;�I;,I;=I;oRI;�aI;T@I;ҐH;��F;s B;�w8;�&;0;��: tX��� ��Q���$�P�y�!¼[��ZN�k������������"��I���q�ە������e��      d5�������W�Ҿ�a��z����l�	�6�DE	���Ƚk���aG����d֮��W����l�k�6���c,:���:��;��1;A�>;AE;&�G;I;&_I;CZI;9DI;�1I;3#I;EI; I;
I;	I;�I;I;�I;	I;
I;�I;BI;2#I;�1I;:DI;EZI;#_I;I; �G;>E;E�>;��1;�;���:�c,:8��m�k�����W�d֮�����aG�k����ȽDE	�	�6��l�z����a��W�Ҿ������      {A��q<�ea/����:�{]׾� ��w��>�DE	�����ڽ����3�^�꼙���",��W��f���Q�~��:�M
;�f);��:;%@C;�?G;P�H;HTI;�_I;*KI;�6I;R'I;gI;�I;>I;�I;oI;�I;mI;�I;<I;�I;gI;O'I;�6I;*KI;�_I;GTI;R�H;�?G;'@C;��:;�f);�M
;���:�Q�f���W��",�����^�꼘�3�ڽ������DE	�>�w��� ��{]׾�:���ea/��q<�      u�������a�{�l$_��q<�������}��w��	�6�����!���h����㷾�� d��.���^e�I[���Z:b��:�, ;��5;�A;�VF;��H;�@I;pbI;�QI;�;I;>+I;kI;I;9I;~	I;�I;.I;�I;~	I;6I;I;jI;>+I;�;I;�QI;rbI;�@I;��H;�VF;�A;��5;�, ;R��:��Z:I[��^e��.��� d�㷾�����h�!������	�6�w���}��������q<�l$_�a�{�����      <��������欿��� ����O��x����� ���l���"��ܽ���`=����v���k"�0R��Fۺ���9�?�:[L;�0;��>;�ME;J#H;�%I;�aI;�VI;�@I;�.I;<!I;@I;I;
I;MI;�I;JI;
I;I;>I;<!I;�.I;�@I; WI;�aI;�%I;P#H;�ME;��>;��0;ZL;z?�:Г�9Jۺ0R���k"�v������`=����ܽ��"��l�� ����뾁x���O� ������欿����      �������L��jȿk���������O���{]׾z����I�����A��>�d�n�~֮�RH��jλQ�$��(�r��:BN;��+;�<;�3D;��G;�I;�^I;k[I;�DI;%2I;�#I;BI;�I;^I;�	I;�I;�	I;]I;�I;BI;�#I; 2I;�DI;l[I;�^I;�I;��G;�3D;�<;��+;CN;f��:�(�T�$��jλRH�~֮�n�>�d��A������I�z���{]׾����O�����k���jȿL�Ῡ��      @�1i�������I�ѿk��� ���q<��:��a����q����Wн罅���'�Ub̼�zl��.��P�X�\����:��;Ύ&;ū9;$C;7MG;��H;6YI;�^I;�HI;�4I;�%I;�I;
I;�I;�
I;�	I;�
I;�I;I;�I;�%I;�4I;�HI;�^I;9YI;��H;@MG;!C;ƫ9;ώ&;��;��:T��Q�X��.���zl�Ub̼��'�罅��Wн����q��a���:��q<� ��k���I�ѿ������1i�      F:�.5�.�'��������jȿ���l$_���W�Ҿܕ���6�����*���`=�=�漮)��JG�(6�����,�Q:��:�/";�7;^&B;��F;��H;�RI;�`I;sKI;7I;�'I;;I;I;�I;nI;p
I;kI;�I;I;<I;�'I;7I;zKI;�`I;�RI;��H;��F;[&B;	�7;�/";��:�Q:���)6��IG��)��<���`=��*������6�ܕ��W�Ҿ��l$_����jȿ�������.�'�.5�      ��U�Z�O�H-?�.�'���M�ῴ欿a�{�ea/���뾝���I����d���ZN�\5������>H�f ��n�����":��:x�;��5;�`A;��F;H�H;MI;�aI;�MI;�8I;�(I;@I;�I;6I;I;I; I;7I;�I;BI;�(I;�8I;�MI;�aI;MI;N�H;��F;�`A;��5;w�;��:t�":d���g ��=H�����\5���ZN�d������I�������ea/�a�{��欿M����.�'�H-?�Z�O�      ��i���b�Z�O�.5�1i�������������q<�����e��`
V�GE	�!���IY�j9�D�����(��R���ȺX�:N��:�;?�4;>�@;hF;��H;II;ubI;�NI;�9I;�)I;�I;ZI;�I;ZI;ZI;XI;�I;[I;�I;�)I;�9I;�NI;zbI;II;��H;*hF;;�@;?�4;ޔ;J��:L�:��Ⱥ�R����(�D���j9��IY�!��GE	�`
V��e������q<������������1i�.5�Z�O���b�      ඕ�S���Ѭ��.�_���7�{�}߿����,b��V�-l¾Hx�c.���Ž��t�*��f����?�N��(��`�x9���:P�;��2;5@@;_fF;6�H;}�I;O�I;|I;�[I;�CI;2I;�%I;ZI;�I;/I;�I;XI;�%I;2I;�CI;�[I;!|I;Q�I;��I;=�H;nfF;2@@;��2;L�;���:@�x9%��N����?�f��*����t���Žc.�Hx�-l¾�V��,b����}߿{���7�.�_�Ѭ��S���      S���D���#}��+Y��3�����$ڿ%��Ľ\����(���s��3�5����p�c�T���<<�<������`��9I��:ϻ;O%3;Gp@;�yF;��H;��I;��I;�{I;H[I;KCI;�1I;N%I;I;TI; I;PI;I;N%I;�1I;NCI;G[I;�{I;�I;��I;��H;�yF;Gp@;O%3;̻;C��:P��9����<���<<�T��c��p�5����3��s�(�����Ľ\�%���$ڿ����3��+Y�#}�D���      Ѭ��#}�>tf��lG�ע%��p�.�ʿZ����>M����T�����d�Ȥ�̷�.�d��
��I���1�h���d�ຘ��9���:;�U4;��@;ұF;1�H;َI;��I;�yI;�YI;5BI;�0I;�$I;�I;�I;~I;�I;�I;�$I;�0I;7BI;�YI;�yI;��I;ݎI;5�H;�F;��@;�U4;;���:���9Z��i����1��I���
�.�d�̷�Ȥ���d�T�������>M�Z���.�ʿ�p�ע%��lG�>tf�#}�      .�_��+Y��lG�f.�{���꿲���M䂿��5���󾍰��N�N�V��R��!�Q����}���i!��g��p�d	:W
�:��;Z16;��A;9G;�I;5�I;u�I;jvI;HWI;g@I;j/I;�#I;�I;	I;�I;I;�I;�#I;k/I;k@I;GWI;nvI;x�I;6�I;I;CG;��A;Z16;��;Q
�:\	:h񳺊g��i!�}������!�Q�R��V��N�N���������5�M䂿�������{�f.��lG��+Y�      ��7��3�ע%�{��<����ſ	���½\�<����Ͼ����`�3��轻z��}�9�^�Ἓ���z��7}��dt��^:Y+�:��#;��8;��B;sG;n%I;��I;�I;rI;TI;�=I;o-I;"I;GI;�I;yI;�I;JI;"I;p-I;�=I;TI;
rI;�I;��I;r%I;sG;��B;��8;��#;]+�:�^:�dt��7}��z����^��}�9��z����`�3�������Ͼ<��½\�	�����ſ�<��{�ע%��3�      {�����p������ſ$���Ps���1�1r���d���d�}I�ΈŽ��}�`*�KC���^��B黀�D�G๊ �:��;l);7;;'D;1�G;SHI;��I;��I;�lI;�OI;�:I;+I; I;�I;wI;*I;uI;�I; I;+I;�:I;�OI;�lI;��I;��I;THI;:�G;)D;7;;l);��;� �:�F�~�D��B��^�KC��_*���}�ΈŽ|I��d��d��1r����1��Ps�$����ſ��꿃p����      }߿�$ڿ.�ʿ����	����Ps�QX:����%l¾�ǆ���7����85���Q�����t���75�n����� �8�ɼ:��;��.;��=;�EE;�YH;�hI;!�I;��I;$fI;KI;"7I;C(I;�I;�I;�I;wI;�I;�I;�I;E(I;#7I;KI;)fI;��I;$�I;�hI;�YH;�EE;��=;��.;��;�ɼ:��8���n���75��t������Q�85�������7��ǆ�%l¾���QX:��Ps�	�������.�ʿ�$ڿ      ���$��Z���M䂿½\���1�����J˾青�D�N�x��H������V�'�d�Ҽ��|��z��n��Tx����&:�P�:��;�W4;͠@;!gF;^�H;�I;�I;.�I;_I;�EI;3I;%I;AI;�I;�I;�I;�I;�I;BI;!%I;3I;�EI;_I;2�I;"�I;�I;c�H;&gF;ˠ@;�W4;��;�P�:��&:Px���n���z���|�d�ҼV�'����H���x��D�N�青��J˾�����1�½\�M䂿Z���$��      �,b�ý\��>M���5�<��1r��%l¾青�"&W��3�8Sؽ�z��ZG����}I����?���̻��-��
����:��;��&;|9;�C;�dG;HI;=�I;N�I;LvI;yWI;'@I;�.I;�!I;~I;UI;�I;�I;�I;VI;�I;�!I;�.I;,@I;WI;RvI;T�I;@�I;MI;�dG;�C;|9;��&;��;��:�
����-���̻��?�|I�����ZG��z��8Sؽ�3�"&W�青�%l¾1r��<����5��>M�ý\�      �V������������Ͼ�d���ǆ�D�N��3��c�[����\�3��*C���o���	�숻b�h��9��:�h;K�/;2�=;EE;�2H;�WI;��I;�I;�kI;�OI;!:I;�)I;"I;�I;�I;�I;xI;�I;�I;�I;"I;�)I;$:I;�OI;�kI;��I;��I;�WI;�2H;EE;7�=;R�/;�h;��:���9\��눻��	��o�)C��3����\�[���cཱ3�D�N��ǆ��d����Ͼ���������      ,l¾(��T������������d���7�x��8Sؽ[���d�D*�dkּ-\����'�/���R��~��h�:�Z;̣#;5=7;&�A;�F;S�H;n�I;�I;��I;�`I;�GI;�3I;&%I;rI;�I;SI;K
I;J	I;M
I;TI;�I;rI;&%I;�3I;�GI;�`I;��I;�I;l�I;Z�H;�F;(�A;:=7;У#;�Z;r�:`~���R�,����'�,\��dkּC*��d�[��8Sؽx����7��d���������T���(��      Hx��s���d�N�N�`�3�|I����H����z����\�C*��ݼJ���1<<��ڻ�V�`dt��&:z��:6C;�</;ID=;ЈD;��G;�8I;ŘI;��I;tI;$VI;Z?I;�-I;d I;�I;ZI;�
I;�I;I;�I;�
I;]I;�I;b I;�-I;`?I;.VI;tI;��I;ŘI;�8I;��G;׈D;PD=;�</;DC;���:�&:<dt��V�
�ڻ/<<�I����ݼC*���\��z��H������|I�`�3�N�N���d��s�      c.��3�Ȥ�V����ΈŽ85�����ZG�3��dkּI���yC��>�p6}����p�x9\��:	;'�&;�;8;��A;��F;��H;/yI;��I;�I;0fI;�KI;K7I;|'I;�I;�I;XI;I;�I;�I;�I;I;XI;�I;�I;�'I;R7I;�KI;4fI;��I;��I;6yI;��H;��F;��A;�;8;5�&;	;^��:��x9���j6}��>�yC�H���ckּ3��ZG����85��ΈŽ��V��Ȥ��3�      ��Ž5���̷�Q���z����}��Q�U�'����)C��-\��0<<��>n��R��@�"��:&��:
�;�'3;��>;�E;bH;]<I;ȗI;��I;�vI;�XI;�AI;u/I;�!I;�I;�I;S	I;cI;%I;tI;#I;bI;T	I;�I;�I;�!I;}/I;�AI;�XI;�vI;��I;їI;^<I;gH;�E;��>;�'3;�;*��:6��:��D�ຆn���>�/<<�,\��)C�����U�'��Q���}��z��R��̷�4���      ��t��p�.�d� �Q�}�9�_*����c�Ҽ|I���o���'��ڻp6}�R���9���:Jm�:��;��.;<;�oC;67G;��H;сI;ќI;хI;fI;<LI;�7I;�'I;�I;uI;NI;HI;�I;� I;Q I;� I;�I;JI;OI;tI;�I;�'I;�7I;ELI;fI;΅I;֜I;ҁI;��H;?7G;�oC;<;��.;��;Zm�:��:�9�F��l6}�	�ڻ��'��o�|I��c�Ҽ���^*�}�9�!�Q�.�d��p�      (��c��
����^��KC���t����|���?���	�.���V�&���@���:��:�h;�+;��9;��A;ufF;Q�H;q_I;��I;��I;sI;�VI;r@I;�.I;� I;TI;I;�I;jI;O I;�H;�H;~�H;L I;jI;�I;I;[I;� I;�.I;w@I;�VI;�rI;��I;��I;r_I;X�H;{fF;��A;��9;�+;�h;��:��:�� ����V�+����	���?���|��t��JC��_������
�b�      c��R���I��}�������^��75��z���̻�눻�R�Pdt���x90��:Tm�:�h;W�*;ٍ8;��@;ڼE;3(H;b8I;��I;�I;G~I;�`I;�HI;�5I;Y&I;tI;2I;�	I;�I;� I;��H;W�H;��H;T�H;��H;� I;�I;�	I;8I;wI;_&I;�5I;�HI;�`I;N~I;�I;��I;g8I;9(H;�E;��@;Ս8;\�*;�h;Zm�:4��:��x9Ddt��R��눻��̻�z��75��^����~����I��Q��      ��?��<<��1��h!��z��B�i���n����-�V�`~���&:P��:"��:��;�+;э8;;�@;�]E;a�G;BI;�I;N�I;3�I;hiI;8PI;<I;�+I;�I;lI;PI;+I;sI;��H;��H;R�H;��H;Q�H;��H;��H;qI;+I;VI;sI;�I;�+I;<I;3PI;oiI;3�I;J�I;�I;FI;j�G;�]E;:�@;Ս8;�+;��;"��:R��:�&:0~��T𳺋�-��n��k���B黶z��h!��1��<<�      N��B��h����g���7}�r�D����Dx���
�����9|�:���:	;�;��.;��9;��@;�]E;g�G;8I;�I; �I;J�I;�pI;VI;�AI;z0I;�"I;�I;�I;�I;�I;��H;^�H;w�H;a�H;��H;`�H;v�H;]�H;��H;�I;�I;�I;�I;�"I;y0I;�AI;�VI;�pI;F�I;�I;�I;?I;j�G;�]E;��@;��9;��.;�;	;���:��:���9�
��Dx�����y�D��7}��g��h���B��      *������X��T񳺴dt�G� �8��&:��:��:�Z;=C;,�&;�'3;<;��A;߼E;j�G;<I;U|I;��I;��I;}uI;n[I;FI;�4I;(&I;�I;GI;�	I;�I;9�H;��H;6�H;u�H;�H;�H;{�H;r�H;6�H;��H;9�H;�I;�	I;GI;�I;'&I;�4I;	FI;o[I;yuI;��I;ŜI;X|I;?I;g�G;�E;��A;<;�'3;,�&;AC;�Z;��:��:��&:��8�F๜dt�n�n��Ԏ��      ��x9Ж�9ȫ�9H	:��^:� �:�ɼ:�P�:��;�h;̣#;�</;�;8;��>;�oC;{fF;6(H;II;�I;��I;��I;�wI;m^I;6II;�7I;)I;I;�I;�I;GI;L I;I�H;S�H;:�H;��H;��H;��H;��H;��H;:�H;S�H;E�H;P I;JI;�I;�I;I;)I;�7I;5II;i^I;�wI;��I;��I;�I;EI;7(H;zfF;�oC;��>;�;8;�</;ѣ#;�h;��;�P�:�ɼ:z �:��^:<	:��9Ж�9      z��:]��:���:q
�:I+�:��;��;��;��&;P�/;<=7;MD=;��A;�E;=7G;X�H;h8I;�I;�I;��I;�wI;�_I;�JI;�9I;�*I;�I;4I;9I;~I;9I;��H;��H;�H;=�H;��H;�H;��H;�H;��H;=�H;�H;��H;�H;9I;~I;<I;/I;�I;�*I;�9I;�JI;�_I;�wI;��I;�I;�I;h8I;W�H;=7G;�E;��A;OD=;==7;L�/;��&;��;��;��;y+�:[
�:���:A��:      b�;˻;;��;��#;r);��.;�W4;!|9;9�=;-�A;ڈD;��F;mH;��H;w_I;��I;R�I;J�I;{uI;k^I;�JI;%:I;,I;4 I;~I;MI;�I;!I;��H;��H;4�H;�H;k�H;d�H;��H;T�H;��H;`�H;m�H;�H;2�H;�H;��H;I;�I;KI;�I;; I;,I;:I;�JI;n^I;{uI;K�I;N�I;��I;u_I;��H;iH;��F;ڈD;1�A;5�=;!|9;�W4;��.;l);��#;��;
;��;      ��2;V%3;�U4;S16;��8;7;;��=;Ƞ@;�C;CE;�F;��G;��H;^<I;ρI;��I;�I;6�I;�pI;k[I;5II;�9I;,I;� I;I;I;QI;�I;H�H;c�H;\�H;*�H;;�H;��H;��H;`�H; �H;[�H;��H;��H;9�H;(�H;^�H;b�H;F�H;�I;MI;I;I;� I;,I;�9I;5II;j[I;�pI;2�I;�I;��I;ρI;Z<I;��H;��G;�F;BE;�C;͠@;��=;7;;��8;O16;�U4;L%3;      P@@;Ap@;��@;��A;��B;1D;�EE;!gF;�dG;�2H;X�H;�8I;0yI;ԗI;ٜI;��I;R~I;siI;�VI;FI;�7I;�*I;< I;!I;\I;�I;=I;��H;��H;��H;�H;"�H;��H;o�H;��H;%�H;��H;�H;��H;p�H;��H;�H;�H;��H;��H;��H;7I;�I;^I;I;8 I;�*I;�7I;FI;�VI;qiI;S~I;��I;؜I;їI;2yI;�8I;[�H;�2H;�dG;gF;�EE;&D;��B;��A;��@;Cp@;      ]fF;�yF;ϱF;9G;�rG;;�G;�YH;l�H;MI;�WI;q�I;˘I;��I;��I;҅I;sI;�`I;8PI;�AI;�4I;)I;�I;~I;I;�I;RI;��H;��H;��H;T�H;-�H;c�H;�H;,�H;t�H;�H;�H;�H;p�H;,�H;�H;b�H;/�H;S�H;��H; �H;��H;VI;�I;I;|I;�I;)I;�4I;�AI;4PI;�`I;sI;ЅI;��I;��I;ʘI;u�I;�WI;MI;j�H;�YH;/�G;sG;BG;αF;�yF;      I�H;��H;(�H;I;c%I;QHI;�hI;�I;@�I;��I;�I;��I;��I;�vI;fI;�VI;�HI;<I;�0I;,&I;I;1I;OI;TI;:I;��H;�H;��H;i�H;2�H;l�H;��H;��H;�H;j�H;�H;�H;�H;h�H;	�H;��H;��H;m�H;0�H;c�H;��H;��H;��H;>I;SI;OI;5I;I;(&I;}0I; <I;�HI;�VI;fI;�vI;�I;��I;�I;��I;=�I;�I;�hI;MHI;y%I;�I;'�H;��H;      {�I;��I;ՎI;<�I;��I;��I;+�I;�I;P�I;��I;��I;tI;.fI;�XI;<LI;v@I;�5I;�+I;�"I;�I;�I;8I;�I;�I;��H;��H;��H;^�H;G�H;\�H;��H;��H;��H;��H;��H;A�H;&�H;>�H;��H;��H;��H;��H;��H;[�H;D�H;^�H;��H;��H;��H;�I;�I;9I;�I;�I;�"I;�+I;�5I;w@I;;LI;�XI;-fI;tI;��I;��I;N�I;�I;(�I;��I;��I;<�I;ՎI;�I;      N�I;ٛI;��I;��I;ٔI;��I;��I;4�I;HvI;�kI;�`I;,VI;�KI;�AI;�7I;�.I;b&I;�I;�I;LI;�I;{I; I;G�H;��H;��H;b�H;E�H;a�H;��H;��H;��H;��H;%�H;��H;��H;P�H;�H;��H;'�H;��H;��H;��H;��H;\�H;G�H;^�H;��H;��H;C�H; I;{I;�I;GI;�I;�I;b&I;�.I;�7I;�AI;�KI;)VI;�`I;�kI;KvI;2�I;��I;��I;�I;��I;��I;כI;      |I;�{I;�yI;evI;rI;�lI;'fI;!_I;{WI;�OI;�GI;d?I;O7I;/I;�'I;� I;{I;lI;�I;�	I;NI;6I;��H;b�H;��H;L�H;/�H;_�H;��H;��H;��H;��H;��H;��H;�H;��H;��H;��H;
�H;��H;��H;��H;��H;��H;��H;^�H;*�H;P�H;��H;_�H;��H;8I;II;�	I;�I;kI;zI;� I;�'I;{/I;N7I;`?I;�GI;�OI;{WI;_I;+fI;�lI;rI;lvI;�yI;{I;      �[I;c[I;�YI;RWI;TI;�OI;KI;�EI;.@I;(:I;�3I;�-I;�'I;�!I;�I;[I;<I;VI;�I;�I;V I;�H;�H;]�H;�H;*�H;l�H;��H;��H;��H;~�H;��H;V�H;��H;x�H;[�H;T�H;Y�H;t�H;��H;W�H;��H;~�H;��H;��H;��H;i�H;-�H; �H;\�H;�H; �H;P I;�I;�I;TI;<I;\I;�I;�!I;�'I;�-I;�3I;(:I;-@I;�EI;#KI;�OI;TI;RWI;�YI;`[I;      �CI;VCI;5BI;a@I;�=I;�:I;%7I;3I;�.I;�)I;(%I;i I;�I;�I;wI;I;
I;.I;�I;>�H;P�H;��H;3�H;'�H;�H;\�H;��H;��H;��H;��H;��H;A�H;��H;N�H;�H;��H;��H;��H;�H;Q�H;��H;@�H;��H;��H;��H;��H;��H;_�H;#�H;!�H;7�H;��H;J�H;:�H;�I;/I;
I;I;wI;�I;�I;e I;(%I;�)I;�.I;3I;)7I;�:I;�=I;g@I;<BI;WCI;      	2I;�1I;�0I;m/I;q-I;+I;A(I; %I;�!I; I;uI;�I;�I;�I;RI;�I;�I;vI;��H;��H;^�H;�H;�H;4�H;��H;�H;��H;��H;��H; �H;S�H;��H;3�H;��H;��H;�H;o�H;�H;��H;��H;2�H;��H;R�H;��H;��H;��H;��H;�H;��H;7�H;�H;�H;W�H;��H;��H;vI;�I;�I;RI;�I;�I;�I;wI; I;�!I;%I;B(I;+I;v-I;h/I;�0I;�1I;      �%I;Q%I;�$I;�#I;"I; I;�I;II;�I;�I;�I;dI;aI;[	I;OI;oI;� I;��H;a�H;;�H;A�H;=�H;h�H;��H;h�H;#�H;�H; �H;'�H;��H;��H;N�H;��H;��H;\�H;9�H;&�H;9�H;\�H;��H;��H;O�H;��H;}�H;"�H;��H;�H;#�H;n�H;��H;n�H;<�H;;�H;5�H;`�H;��H;� I;qI;NI;[	I;]I;`I;�I;�I;�I;EI;�I; I;"I;�#I;�$I;[%I;      NI;4I;�I;�I;UI;�I;�I;�I;\I;�I;_I;�
I;I;lI;�I;S I;��H;��H;x�H;v�H;��H;��H;_�H;��H;��H;f�H;a�H;��H;��H;�H;n�H;�H;��H;[�H;�H;�H;�H;�H;�H;^�H;��H;�H;n�H;�H;��H;��H;a�H;g�H;��H;��H;c�H;��H;��H;r�H;w�H;��H;��H;W I;�I;mI;I;�
I;aI;�I;]I;�I;�I;�I;QI;�I;�I;5I;      �I;^I;�I;I;�I;uI;�I;�I;�I;�I;T
I;I;�I;)I;� I;~�H;X�H;N�H;b�H;|�H;��H;�H;��H;M�H;�H;�H;�H;?�H;��H;��H;V�H;��H;��H;8�H;	�H;��H;��H;��H;�H;=�H;��H;��H;V�H;��H;��H;>�H;�H;�H;�H;Q�H;��H;�H;��H;x�H;a�H;T�H;[�H;��H;� I;)I;�I;�I;T
I;�I;�I;�I;�I;sI;�I;	I;�I;kI;      7I;�I;�I;�I;uI;&I;{I;�I;�I;yI;W	I;I;�I;~I;Z I;�H;��H;��H;��H; �H;��H;��H;S�H;��H;��H;�H;	�H;*�H;V�H;��H;M�H;��H;q�H;!�H;�H;��H;��H;��H;�H;#�H;s�H;��H;N�H;��H;P�H;&�H;�H;�H;��H;��H;W�H;��H;��H;�H;��H;��H;��H;�H;X I;~I;�I;I;W	I;yI;�I;�I;�I;%I;sI;�I;�I;I;      �I;`I;�I;I;�I;wI;�I;�I;�I;�I;R
I;I;�I;*I;� I;~�H;X�H;N�H;b�H;|�H;��H;�H;��H;M�H;�H;�H;�H;?�H;��H;��H;V�H;��H;��H;9�H;	�H;��H;��H;��H;�H;<�H;��H;��H;V�H;��H;��H;<�H;�H;�H;�H;P�H;��H;�H;��H;x�H;a�H;T�H;Z�H;��H;� I;(I;�I;�I;T
I;�I;�I;�I;�I;vI;�I;I;�I;eI;      DI;4I;�I;�I;UI;�I;�I;�I;\I;�I;aI;�
I;I;mI;�I;S I;��H;��H;x�H;v�H;��H;��H;_�H;��H;��H;d�H;a�H;��H;��H;�H;m�H;�H;��H;[�H;�H;�H;�H;�H;�H;^�H;��H;�H;n�H;�H;��H;��H;a�H;j�H;��H;��H;c�H;��H;��H;r�H;x�H;��H;��H;V I;�I;lI;I;�
I;_I;�I;]I;�I;�I;�I;UI;�I;�I;;I;      �%I;P%I;�$I;�#I;"I; I;�I;LI;�I;�I;�I;cI;^I;[	I;QI;oI;� I;��H;a�H;9�H;A�H;?�H;j�H;��H;l�H;%�H;�H; �H;)�H;��H;��H;N�H;��H;��H;^�H;8�H;'�H;;�H;[�H;��H;��H;Q�H;��H;}�H;"�H;��H;�H;(�H;o�H;��H;n�H;=�H;;�H;6�H;c�H;��H;� I;qI;OI;Z	I;]I;`I;�I;�I;�I;HI;�I; I;"I;�#I;�$I;S%I;      2I;�1I;�0I;e/I;o-I;+I;A(I;$%I;�!I; I;uI;�I;�I;�I;UI;�I;�I;vI;��H;��H;\�H;�H;�H;7�H;��H;�H;��H;��H;��H;��H;R�H;��H;2�H;��H;��H;�H;o�H;�H;��H;��H;0�H;��H;R�H;��H;��H;��H;��H;�H;��H;4�H;�H;�H;U�H;��H;��H;vI;�I;�I;PI;�I;�I;�I;tI;I;�!I; %I;F(I;
+I;t-I;r/I;�0I;�1I;      �CI;WCI;)BI;`@I;�=I;�:I;)7I;3I;�.I;�)I;-%I;i I;�I;�I;zI;I;
I;/I;�I;=�H;Q�H;��H;4�H;&�H;#�H;^�H;��H;��H;��H;��H;��H;>�H;��H;M�H;�H;��H;��H;��H;�H;N�H;��H;@�H;��H;��H;��H;��H;��H;a�H;!�H;�H;9�H;��H;I�H;:�H;�I;/I;
I;I;uI;�I;�I;h I;(%I;�)I;�.I;3I;(7I;�:I;�=I;h@I;.BI;UCI;      �[I;d[I;�YI;KWI;TI;�OI;KI;�EI;.@I;(:I;�3I;�-I;�'I;�!I;�I;\I;=I;TI;�I;�I;W I;�H;�H;]�H; �H;)�H;j�H;��H;��H;��H;|�H;��H;V�H;��H;x�H;Y�H;R�H;[�H;t�H;��H;W�H;��H;}�H;��H;��H;��H;h�H;/�H;�H;Y�H;�H;�H;P I;�I;�I;TI;?I;]I;�I;�!I;�'I;�-I;�3I;':I;.@I;�EI;"KI;�OI;TI;WWI;�YI;c[I;      (|I;�{I;�yI;ovI;�qI;�lI;'fI;#_I;}WI;�OI;�GI;e?I;P7I;}/I;�'I;� I;{I;nI;�I;�	I;PI;9I;��H;`�H;��H;L�H;/�H;a�H;��H;��H;��H;��H;��H;�H;�H;��H;��H;��H;
�H;��H;��H;��H;��H;��H;��H;\�H;-�H;Q�H;��H;\�H;��H;9I;JI;�	I;�I;lI;zI;� I;�'I;|/I;N7I;`?I;�GI;�OI;yWI;!_I;(fI;�lI;rI;xvI;�yI;�{I;      V�I;ۛI;��I;��I;ɔI;��I;��I;2�I;RvI;�kI;�`I;.VI;�KI;�AI;�7I;�.I;b&I;�I;�I;II;�I;|I;I;H�H;��H;��H;a�H;H�H;a�H;��H;��H;��H;��H;%�H;��H;��H;O�H;��H;��H;%�H;��H;��H;��H;��H;[�H;A�H;^�H;��H;��H;@�H;!I;|I;�I;II;�I;�I;`&I;�.I;�7I;�AI;�KI;(VI;�`I;�kI;LvI;4�I;��I;��I;ܔI;��I;��I;՛I;      ��I;�I;ɎI;9�I;��I;��I;+�I;#�I;Q�I;��I;��I;tI;-fI;�XI;?LI;w@I;�5I;�+I;�"I;�I;�I;;I;�I;�I;��H;��H;��H;_�H;I�H;Z�H;��H;��H;��H;��H;��H;>�H;'�H;?�H;��H;��H;��H;��H;��H;[�H;B�H;Z�H;��H;��H;��H;�I;�I;9I;�I;�I;�"I;�+I;�5I;w@I;<LI;�XI;-fI;tI;��I;��I;P�I;�I;+�I;��I;��I;<�I;׎I;�I;      8�H;��H;'�H;I;q%I;WHI;�hI;�I;@�I;��I;�I;��I;�I;�vI; fI;�VI;�HI;<I;~0I;)&I;I;5I;MI;XI;=I;��H;�H;��H;i�H;/�H;j�H;��H;��H;�H;i�H;�H;�H;�H;f�H;�H;��H;��H;l�H;/�H;e�H;��H;��H;��H;:I;QI;QI;5I;I;+&I;~0I;<I;�HI;�VI;fI;�vI;�I;��I;�I;��I;=�I;�I;�hI;SHI;v%I;
I;*�H;��H;      UfF;�yF;ڱF;1G;sG;A�G;�YH;l�H;QI;�WI;r�I;ΘI;��I;��I;ՅI;sI;�`I;:PI;�AI;�4I;)I;�I;|I;I;�I;OI;��H;�H;��H;Q�H;-�H;c�H;�H;,�H;r�H;�H;�H;�H;p�H;*�H;�H;c�H;0�H;Q�H;��H;��H;��H;VI;�I;I;~I;�I;)I;�4I;�AI;5PI;�`I;sI;ԅI;��I;��I;ȘI;t�I;�WI;GI;e�H;�YH;1�G;sG;6G;ñF;�yF;      M@@;Ap@;��@;��A;��B;3D;�EE;!gF;�dG;�2H;[�H;�8I;0yI;җI;ܜI;��I;S~I;uiI;�VI;FI;�7I;�*I;: I;"I;^I;�I;:I;��H;��H;��H;�H;!�H;��H;o�H;��H;!�H;��H;!�H;��H;p�H;��H;!�H;�H;��H;��H;��H;:I;�I;ZI;I;; I;�*I;�7I;FI;�VI;qiI;S~I;��I;ۜI;їI;2yI;�8I;V�H;�2H;�dG;"gF;�EE;'D;��B;��A;��@;@p@;      }�2;A%3;�U4;Y16;��8;#7;;��=;ɠ@;�C;BE;�F;��G;��H;[<I;ҁI;��I;�I;8�I;�pI;k[I;8II;�9I;,I;� I;I;I;PI;�I;H�H;`�H;]�H;*�H;:�H;��H;��H;]�H;�H;^�H;��H;��H;=�H;*�H;`�H;b�H;F�H;�I;PI;I;I;� I;,I;�9I;6II;k[I;�pI;3�I;�I;��I;ρI;X<I;��H;��G;�F;AE;�C;Ġ@;��=;7;;��8;u16;�U4;+%3;      T�;̻;;��;��#;p);��.;�W4;$|9;9�=;(�A;ڈD;��F;kH;��H;y_I;I;S�I;K�I;}uI;n^I;�JI;":I; ,I;: I;xI;MI;�I;$I;��H;�H;6�H;�H;k�H;c�H;��H;U�H;��H;`�H;j�H;�H;4�H;�H;��H;I;�I;NI;I;5 I;,I;!:I;�JI;n^I;}uI;M�I;L�I;��I;x_I;��H;gH;��F;׈D;*�A;9�=;"|9;�W4;��.;p);��#;�;;��;      z��:Y��:���:Q
�:G+�:��;��;��;��&;M�/;<=7;QD=;��A;�E;A7G;[�H;h8I;�I;�I;��I;�wI;�_I;�JI;�9I;�*I;�I;2I;<I;I;9I; �H;��H;�H;=�H;��H;�H;��H;�H;��H;;�H;�H;��H;�H;<I;|I;9I;4I;�I;�*I;�9I;�JI;�_I;�wI;��I;�I;�I;g8I;X�H;<7G;�E;��A;MD=;==7;M�/;��&;��;��;x�;y+�:C
�:���:I��:      ��x9x��9P��9H	:��^:� �:�ɼ:�P�:��;~h;У#;�</;�;8;��>;�oC;|fF;7(H;II;�I;��I;��I;�wI;k^I;8II;�7I;)I;I;�I;�I;GI;M I;I�H;S�H;>�H;��H;��H;��H;��H;��H;9�H;S�H;F�H;O I;JI;�I;�I;I;)I;�7I;8II;j^I;�wI;��I;��I;�I;FI;6(H;zfF;�oC;��>;�;8;�</;ѣ#;h;��;�P�:�ɼ:� �:�^:T	:���9���9      ������Z��T񳺴dt��F���8��&:��:��:�Z;AC;/�&;�'3;<;��A;�E;j�G;=I;X|I;ŜI;��I;}uI;o[I;	FI;~4I;%&I;�I;LI;�	I;�I;:�H;��H;8�H;u�H;{�H;�H;{�H;q�H;2�H;��H;7�H;�I;�	I;II;�I;(&I;�4I;FI;r[I;}uI;��I;ÜI;W|I;=I;f�G;߼E;��A;<;�'3;,�&;=C;�Z;	��:��:��&:��8(G๨dt�h�`�ຬ���      N��B��f����g���7}�r�D����Dx���
�����9~�:���:	;�;��.;��9;��@;�]E;j�G;=I;�I;�I;K�I;�pI;�VI;�AI;y0I;�"I;�I;�I;�I;�I;��H;^�H;x�H;a�H;��H;a�H;t�H;\�H;��H;�I;�I;�I;�I;�"I;z0I;�AI;VI;�pI;J�I;�I;�I;=I;g�G;�]E;��@;��9;��.;�;	;���:|�:���9�
��Dx�����s�D��7}��g��j���>��      ��?��<<��1��h!��z��B�h���n����-�R�8~���&:R��:&��:��;�+;Ս8;;�@;�]E;h�G;FI;�I;R�I;6�I;qiI;5PI;<I;�+I;�I;nI;TI;,I;sI;��H;��H;Q�H;��H;R�H;��H;��H;sI;(I;TI;nI;�I;�+I;<I;4PI;hiI;5�I;O�I;�I;BI;h�G;�]E;:�@;ҍ8;�+;��; ��:P��:�&:0~��V𳺍�-��n��j���B黷z��h!��1��<<�      c��R���I��|�������^��75��z���̻�눻�R�8dt���x94��:^m�:�h;\�*;؍8;��@;�E;:(H;g8I;��I;�I;Q~I;�`I;�HI;�5I;b&I;tI;6I;�	I;�I;� I;��H;W�H;��H;W�H;��H;� I;�I;�	I;6I;tI;]&I;�5I;�HI;�`I;H~I;�I;��I;e8I;3(H;߼E;��@;ԍ8;Y�*;�h;Xm�:0��:��x9Hdt��R��눻��̻�z��75��^����}����I��Q��      (��c��
����^��JC���t����|���?���	�+���V��������:��:�h;�+;��9;��A;~fF;Z�H;y_I;��I;��I;sI;�VI;u@I;�.I;� I;YI;I;�I;nI;S I;�H;�H;~�H;L I;hI;�I;	I;VI;� I;�.I;u@I;�VI;�rI;��I;��I;w_I;W�H;tfF;��A;��9;�+;�h;��:��:@�"����V�-����	���?���|��t��JC��_������
�b�      ��t��p�/�d� �Q�}�9�_*����c�Ҽ|I���o���'�
�ڻl6}�F�ຐ9���:Zm�:��;��.;<;�oC;?7G;��H;ՁI;ٜI;ԅI;fI;ALI;�7I;�'I;�I;uI;OI;MI;�I;� I;P I;� I;�I;JI;NI;qI;�I;�'I;�7I;>LI;fI;ЅI;ќI;ՁI;��H;=7G;�oC;<;��.;��;Xm�:��:�9�L��o6}��ڻ��'��o�|I��c�Ҽ���_*�~�9�!�Q�/�d��p�      ��Ž4���̷�Q���z����}��Q�U�'����)C��,\��/<<��>n��@�຀�.��:(��:�;�'3;��>;�E;iH;b<I;ԗI;��I;�vI;�XI;�AI;y/I;�!I;�I;�I;T	I;cI;"I;tI;%I;aI;T	I;�I;�I;�!I;y/I;�AI;�XI;�vI;��I;ʗI;a<I;kH;�E;��>;�'3;
�;&��:.��:@�L�ຆn���>�0<<�,\��)C�����U�'��Q���}��z��Q��̷�4���      c.��3�Ȥ�V����ΈŽ85�����ZG�3��ckּI��� yC��>�h6}������x9^��:		;/�&;�;8;��A;��F;��H;6yI;��I;�I;1fI;�KI;O7I;�'I;�I;�I;[I;I;�I;�I;�I;I;XI;�I;�I;}'I;N7I;�KI;0fI;�I;��I;/yI;��H;��F;��A;�;8;/�&;	;V��:��x9���l6}��>�yC�I���ckּ3��ZG����85��ΈŽ��V��Ȥ��3�      Hx��s���d�N�N�`�3�|I����H����z����\�C*��ݼI���0<<�	�ڻ�V�Hdt��&:���:>C;�</;PD=;وD;��G;�8I;ȘI;��I;tI;+VI;\?I;�-I;d I;�I;]I;�
I;�I;I;�I;�
I;\I;�I;a I;�-I;\?I;+VI;tI;��I;ØI;�8I;��G;ڈD;MD=;�</;>C;z��:�&:Pdt��V�
�ڻ0<<�J����ݼC*���\��z��H������|I�`�3�N�N���d��s�      ,l¾(��T������������d���7�x��8Sؽ[���d�D*�ckּ-\����'�-���R�h~��p�:�Z;գ#;<=7;-�A;�F;X�H;q�I;�I;��I;�`I;�GI;�3I;'%I;rI;�I;TI;M
I;L	I;M
I;TI;�I;rI;$%I;�3I;�GI;�`I;��I;�I;l�I;T�H;�F;-�A;8=7;ǣ#;�Z;h�:p~���R�.����'�-\��dkּD*��d�[��8Sؽx����7��d���������T���(��      �V������������Ͼ�d���ǆ�D�N��3��c�[����\�3��)C���o���	��눻`𳺈��9��:�h;P�/;9�=;JE;�2H;�WI;��I;��I;�kI;�OI;%:I;�)I;$I;�I;�I;�I;xI;�I;�I;�I;"I;�)I;":I;�OI;�kI;��I;��I;�WI;�2H;HE;:�=;M�/;zh;��:h��9b��눻��	��o�)C��3����\�[���cཱ3�D�N��ǆ��d����Ͼ���������      �,b�ý\��>M���5�<��1r��%l¾青�"&W��3�8Sؽ�z��ZG����|I����?���̻��-��
����:��;��&;|9;�C;�dG;MI;?�I;Q�I;SvI;}WI;-@I;�.I;�!I;�I;UI;�I;�I;�I;VI;�I;�!I;�.I;)@I;yWI;RvI;Q�I;?�I;KI;�dG;�C;|9;��&;��;��:�
����-���̻��?�}I�����ZG��z��8Sؽ�3�"&W�青�%l¾1r��<����5��>M�ý\�      ���$��Z���M䂿½\���1�����J˾青�D�N�x��H������V�'�d�Ҽ��|��z��n��Lx����&:�P�:��;�W4;Р@;&gF;a�H;�I;�I;2�I;_I;�EI;3I;!%I;DI;�I;�I;�I;�I;�I;DI; %I;3I;�EI;_I;1�I;�I;�I;a�H;"gF;͠@;�W4;��;�P�:��&:Rx���n���z���|�d�ҼV�'����H���x��D�N�青��J˾�����1�½\�M䂿Z���$��      }߿�$ڿ.�ʿ����	����Ps�QX:����%l¾�ǆ���7����85���Q�����t���75�n�������8�ɼ:��;��.;��=;�EE;�YH;�hI;!�I;��I;(fI;KI;#7I;E(I;�I;�I;�I;wI;�I;�I;�I;E(I;%7I;KI;(fI;��I;$�I;�hI;�YH;�EE;��=;��.;��;�ɼ:��8���n���75��t������Q�85�������7��ǆ�%l¾���QX:��Ps�	�������.�ʿ�$ڿ      {�����p������ſ$���Ps���1�1r���d���d�|I�ΈŽ��}�_*�KC���^��B�}�D��F๐ �:��;n);7;;)D;1�G;SHI;��I;��I;�lI;�OI;�:I;+I; I;�I;yI;-I;yI;�I; I;+I;�:I;�OI;�lI;��I;��I;UHI;:�G;'D;7;;p);��;� �:�Fแ�D��B��^�JC��`*���}�ΈŽ|I��d��d��1r����1��Ps�$����ſ��꿃p����      ��7��3�ע%�{��<����ſ	���½\�<����Ͼ����`�3��轻z��}�9�^�Ἓ���z��7}��dt��^:]+�:��#;��8;��B;	sG;n%I;��I;�I;rI;TI;�=I;p-I;"I;GI;�I;yI;�I;HI;"I;p-I;�=I;TI;	rI;�I;��I;t%I;sG;��B;��8;��#;]+�:��^:�dt��7}��z����^��}�9��z����`�3�������Ͼ<��½\�	�����ſ�<��{�ע%��3�      .�_��+Y��lG�f.�{���꿲���M䂿��5���󾍰��N�N�V��R��!�Q����}���i!��g��h�p	:U
�:��;Y16;��A;8G;�I;5�I;w�I;jvI;KWI;i@I;j/I;�#I;�I;	I;�I;I;�I;�#I;m/I;k@I;IWI;ovI;x�I;8�I;I;CG;��A;\16;��;Q
�:T	:h񳺌g��i!�}������!�Q�R��V��N�N���������5�M䂿�������{�f.��lG��+Y�      Ѭ��#}�>tf��lG�ע%��p�.�ʿZ����>M����T�����d�Ȥ�̷�.�d��
��I���1�h���`�ະ��9���:;�U4;��@;ұF;1�H;ڎI;��I;�yI;�YI;6BI;�0I;�$I;�I;�I;I;�I;�I;�$I;�0I;7BI;�YI;�yI;��I;ގI;6�H;�F;��@;�U4;;���:���9X��h����1��I���
�.�d�̷�ɤ���d�U�������>M�Z���.�ʿ�p�ע%��lG�>tf�#}�      S���D���#}��+Y��3�����$ڿ%��Ľ\����(���s��3�5����p�c�T���<<�<������h��9I��:ϻ;N%3;Gp@;�yF;��H;��I;��I;�{I;I[I;LCI;�1I;P%I;I;SI;I;PI;I;P%I;�1I;OCI;G[I;�{I;�I;��I;��H;�yF;Ep@;O%3;̻;C��:@��9����=���<<�T��c��p�5����3��s�(�����Ľ\�%���$ڿ����3��+Y�#}�D���      ����,������T���J�Q�ř$�4�����<�}�H(�@�׾�T���L+���սk����L���iO���ͻ���� m8jo�:[�;U�1;��?;�uF;g I;f�I;��I;��I;VvI;�WI;�AI;�1I;�'I;�!I;�I;�!I;�'I;�1I;�AI;�WI;VvI;��I;��I;k�I;j I;�uF;��?;S�1;Z�;do�:�m8�����ͻ�iO�L����k����ս�L+��T��@�׾H(�<�}���4���ƙ$�J�Q�T��������,��      �,��a��#P���{���K��x �����p�����w��$���Ҿf���  (���ѽҷ��'�����K�Fɻ,��`��8x��:z�;��1;�@;k�F;I;ݿI;�I;��I;�uI;#WI;fAI;�1I;�'I;�!I;�I;�!I;�'I;�1I;hAI;%WI;�uI;��I;�I;�I;"I;y�F;�@;��1;z�;v��:���8)��Fɻ�K����'�ҷ����ѽ  (�f�����Ҿ�$���w�p��������x ���K��{�#P��a��      ����#P�������d���;�#���㿲���#f�d��ž��z���<�ƽ%0v�T5�2����o@�����i��`u9AK�:];�73;"�@;��F;FI;��I;M�I;S�I;�sI;�UI;A@I;�0I;�&I;!I;0I;!I;�&I;�0I;A@I;�UI;�sI;Y�I;O�I;��I;JI;��F;"�@;�73;];=K�:�`u9zi������o@�2���T5�%0v�<�ƽ����z�žd��#f�������#����;���d����#P��      T����{���d��F�ř$�:����ɿ.蒿��K�P���j���Yb�F�1���s�a����@�����.��d��r�غ���9�Y�:.X;�25;#�A;Y!G;I7I;s�I;B�I;R�I;�pI;�SI;>I;y/I;�%I;" I;/I; I;�%I;v/I;>I;�SI;�pI;T�I;C�I;t�I;J7I;d!G;!�A;�25;.X;�Y�:���9j�غ�d����.�@������s�a�1���F��Yb��j��P����K�.蒿��ɿ:��ř$��F���d��{�      J�Q���K���;�ř$��;
��޿�����w�r,���澝���'�D������I��$�G�����N��������X�����9:Z��:�n!;��7;��B;J�G;�YI;*�I;W�I;��I;�lI;sPI;<I;�-I;$I;�I;�I;�I;$I;�-I;<I;uPI;�lI;��I;Z�I;/�I;�YI;T�G;��B;��7;�n!;\��:��9:P����������N�����$�G��I������'�D��������r,���w�����޿�;
�ř$���;���K�      ř$��x �#��:���޿o���ʅ���F�}�
��~����z��$���ս���A2+���ϼPp�����P�]� �*���:�;�8';��:;��C;�H;�}I;�I;o�I;׋I;kgI;�LI;9I;7+I;!"I;�I;)I;�I; "I;4+I;9I;�LI;jgI;ۋI;s�I;"�I;�}I;H;��C;��:;�8';�;��:�*�N�]�����Pp���ϼA2+������ս�$���z��~��}�
��F�ʅ��o����޿:��"���x �      4��������㿊�ɿ���ʅ����P�d��;�׾�`��S�H����@��R�a���͡���D��ɻ� ��ح��W�:�;`I-;7|=;CE;��H;�I;��I;s�I;��I;haI;"HI;�5I;p(I;�I;�I;QI;�I;�I;p(I;�5I;#HI;haI;��I;v�I;��I;�I;��H;#CE;8|=;bI-;�;�W�:�׭�� ��ɻ�D�͡����R�a��@����S�H��`��;�׾d����P�ʅ�������ɿ�㿳���      ��p�������.蒿��w��F�d��ʰ� ����Yb�)����ѽ�%��D4�ٟ�X�����H���潺���9Br�:��;�93;%Q@;zvF;�H;�I;��I;��I;�zI;�ZI;CI;�1I;b%I;?I;�I;"I;�I;BI;c%I;�1I;CI;�ZI;�zI;��I;��I;	�I;�H;�vF;$Q@;�93;��;@r�:���9�潺H�����X��؟�D4��%����ѽ)���Yb� ���ʰ�d���F���w�.蒿����p���      <�}���w�#f���K�r,�}�
�;�׾ �����k���'�ez꽝I���;V�=M�
����iO�mG�soE�̱�2��:B� ;��$;��8;[�B;��G;,KI;�I;�I;@�I;qI;�SI;�=I;�-I;"I;jI;I;�I;I;mI;"I;�-I;�=I;�SI;qI;D�I;�I;�I;.KI;��G;\�B;��8;��$;A� ;D��:���poE�jG໫iO�	���<M��;V��I��ez���'���k� ���;�׾}�
�r,���K�#f���w�      H(��$�d��P������~���`���Yb���'��U�G$��D�m�&����ϼ�/��>��������غ08�94��:�F;�G.;|=;GE;�\H;�I;s�I;y�I;��I;gI; LI;�7I;)I;pI;rI;rI;'I;qI;rI;pI;)I;�7I;LI;	gI;��I;�I;s�I;�I;�\H;IE;|=;�G.;�F;H��:P8�9��غ����>���/����ϼ&��D�m�G$���U���'��Yb��`���~�����P��d���$�      ?�׾��Ҿž�j��������z�S�H�)��ez�G$���/v�2+�ߐ�����5��ɻ<4�P(��~��:T��:5o!;P6;lA;��F;p�H;��I;��I;ߦI;F}I;�\I;[DI;	2I;r$I;�I;HI;�I;�I;�I;II;�I;s$I;2I;`DI;�\I;M}I;�I;��I;��I;x�H;��F;
lA;P6;8o!;n��:���:8(��34��ɻ��5���ސ�2+��/v�G$��ez�)��S�H���z������j��ž��Ҿ      �T��f�����z��Yb�&�D��$�����ѽ�I��D�m�2+�������L�K�ﻛ�p�P������9!T�:�/;o�-;d�<;BzD;ZH;�mI;��I;|�I;��I;�oI;�RI;�<I;,I;�I;I;/I;�I;�I;�I;.I;I;�I;,I;�<I;�RI;�oI;��I;}�I;��I;�mI;]H;IzD;m�<;r�-;�/;-T�:���9>�����p��K�K�������2+�D�m��I����ѽ���$�'�D��Yb���z�f���      �L+�  (���F�������ս�@���%���;V�%��ސ������MS�N��(��~D� �n8q�:�;a�$;�^7;(�A;d�F;��H;_�I;b�I;��I;��I;QbI;�HI;5I;(&I;/I;>I;�I;�
I;
I;�
I;�I;>I;/I;'&I;5I;�HI;YbI;�I;��I;`�I;f�I;��H;h�F;1�A;_7;n�$;�; q�:��n8tD�&��L���MS�����ސ�%���;V��%���@����ս����F���  (�      ��ս��ѽ;�ƽ1����I�����R�a�D4�<M���ϼ��L�K�O��OG��df���o���:�B�:�Y;��1;Ol>;�E;�/H;qI;��I;��I;ژI;�rI;�UI;�>I;�-I;b I;�I;�I;�
I;I;0I;I;�
I;�I;�I;a I;�-I;�>I;�UI;sI;ژI;��I;�I; qI;�/H;�E;Rl>;��1;�Y;�B�:��:��o�^f�LG��N��K�K�����ϼ<M�D4�Q�a�����I��1���;�ƽ��ѽ      j��ҷ��%0v�r�a�$�G�@2+���ן�	����/����5��(��bf��ج���g:3�:�;I-;g;;�NC;SG;�I;ɶI;�I;��I;	�I;
cI;~II;�5I;n&I;�I;7I;�I;�I;PI;XI;NI;�I;�I;9I;�I;u&I;�5I;�II;cI;	�I;��I;�I;ʶI;�I;SG;OC;g;;I-;�;A�:�g:�ج�]f�&�����5��/�����؟���@2+�%�G�r�a�%0v�ҷ��      
��'�T5���������ϼ̡��X���iO�>���ɻ��p��D���o���g:�_�:@G;n*;o9;��A;�uF;�H;��I;��I;��I;H�I;�pI;3TI;M>I;-I;�I;}I;�I;VI;�I;�I;�I;�I;�I;VI;�I;{I;�I; -I;T>I;:TI;�pI;B�I;��I;��I;ÔI;!�H;�uF;��A;s9;l*;EG;�_�:�g:��o��D⺙�p��ɻ>���iO�X��͡����ϼ������T5�&�      L�����2���@����N��Pp��D����hG�����64�D��� �n8��:9�:GG;�(;��7;Y�@;��E;KQH;mI;��I;��I;��I;#}I;�^I;�FI;�3I;�$I;\I;�I;�	I;I;�I;��H;P�H;��H;�I;I;�	I;�I;bI;�$I;�3I;�FI;�^I; }I;��I;��I;��I;mI;QQH;��E;]�@;��7;�(;HG;E�:��:��n8B���04�����hG໇���D�Pp��N��@���4������      �iO��K��o@���.���������ɻH��ooE���غ8(�����9�p�:�B�:�;j*;��7;�P@;�\E;�H;�II;~�I;h�I;�I;V�I;<hI;�NI;b:I;9*I;xI;�I;�I;I;I;2�H;b�H;��H;^�H;/�H;I;I;�I;�I;}I;:*I;f:I;�NI;:hI;_�I;�I;d�I;��I;�II;�H;�\E;�P@;��7;l*;�;�B�:�p�:���9 (����غioE� H���ɻ���������.��o@��K�      ��ͻMɻ�����d�����B�]�� ��潺���X8�9���:)T�:�;�Y;I-;s9;Z�@;�\E;��G;/5I;��I;C�I;ڵI;R�I;bpI;�UI;T@I;3/I;{!I;�I;@I;�I;�I;"�H;��H;�H;��H;�H;��H;!�H;�I;�I;DI;�I;}!I;9/I;Q@I;�UI;kpI;V�I;յI;G�I;��I;55I;��G;�\E;_�@;r9;I-;�Y;�;-T�:���:h8�9����潺� �I�]�����d������Mɻ      ���.��xi�\�غh����*�`׭����9<��:B��:f��:�/;g�$;��1;g;;��A;��E;�H;25I;9�I;��I;L�I;��I;�vI;L[I;^EI;�3I;5%I;�I;�I;P	I;�I;}�H;a�H;'�H;��H;n�H;��H;"�H;a�H;�H;�I;S	I;�I;�I;9%I;�3I;\EI;U[I;�vI;��I;M�I;��I;;�I;65I;�H;��E;��A;g;;��1;e�$;�/;n��:B��:@��:���9�׭� �*�X���t�غ�i�<��      @)m8���8_u9x��9P�9:��:�W�:Dr�:=� ;�F;4o!;q�-;�^7;Pl>;�NC;�uF;PQH;�II;��I;��I;��I;��I;|zI;_I;<II;K7I;a(I;`I;�I;I;�I;, I;u�H;��H;�H;��H;w�H;��H;�H;��H;r�H;' I;�I;I;�I;dI;`(I;I7I;CII;_I;xzI;��I;��I;��I;��I;�II;QQH;�uF;�NC;Kl>;�^7;o�-;;o!;�F;;� ;<r�:�W�:��:x�9:h��9�_u9���8      Vo�:���:QK�:�Y�:@��:�;�;��;��$;�G.;P6;i�<;*�A;�E;SG;!�H;mI;��I;H�I;P�I;��I;�{I;vaI;�KI;�9I;�*I;�I;�I;�I;%I;� I;��H;��H;k�H;��H;�H;��H;�H;��H;k�H;��H;��H;� I;(I;�I;�I;�I;�*I;�9I;�KI;paI;�{I;��I;O�I;J�I;��I;mI; �H;SG;�E;+�A;j�<;P6;�G.;��$;��;�;�;r��:�Y�:=K�:p��:      n�;x�;];:X;�n!;�8';jI-;�93;��8;|=;lA;MzD;f�F;�/H;�I;ȔI;��I;k�I;ڵI;��I;|zI;saI;vLI;;I;^,I;0 I;I;�I;;I;�I;v�H;��H;g�H;o�H;
�H;V�H;#�H;P�H;�H;q�H;g�H;��H;z�H;�I;9I;�I;I;1 I;e,I;;I;pLI;vaI;zI;��I;ܵI;g�I;��I;ǔI;�I;�/H;f�F;MzD;lA;|=;��8;�93;hI-;�8';�n!;8X;];X�;      O�1;��1;�73;�25;}�7;��:;1|=;!Q@;R�B;HE;��F;ZH;��H; qI;ȶI;��I;��I;�I;R�I;�vI;|_I;�KI;;I;�,I;� I;I;�I;I;tI;��H;q�H;m�H;#�H;��H;r�H;��H;��H;��H;p�H;��H;#�H;m�H;w�H;��H;qI;I;�I;I;� I;�,I;;I;�KI;}_I;�vI;Q�I;�I;��I;��I;ɶI;qI;��H;ZH;��F;EE;V�B;(Q@;.|=;��:;��7;�25;�73;��1;      ��?;�@;�@;�A;��B;��C;#CE;zvF;��G;�\H;x�H;�mI;b�I;�I;�I;��I;��I;a�I;opI;W[I;GII;�9I;e,I;� I;oI;^I;�I;�I;g�H;��H;��H;-�H;V�H;��H;��H;`�H;4�H;Z�H;��H;��H;U�H;(�H;��H;��H;d�H;�I;�I;^I;rI;� I;a,I;�9I;III;U[I;opI;_�I;��I;��I; �I;�I;b�I;�mI;x�H;�\H;��G;zvF;$CE;��C;��B;�A;�@;�@;      �uF;w�F;��F;Y!G;=�G;H;��H;�H;0KI;'�I;��I;��I;b�I;��I;��I;I�I;'}I;<hI;�UI;[EI;L7I;�*I;- I;I;\I;�I;GI;��H;��H;��H;&�H;>�H;��H;]�H;��H;�H;��H;�H;��H;`�H;��H;:�H;&�H;��H;��H;��H;@I;�I;^I;I;, I;�*I;L7I;ZEI;�UI;;hI;'}I;L�I;��I;��I;b�I;��I;��I;$�I;0KI;�H;��H;�H;T�G;d!G;��F;u�F;      t I;(I;>I;J7I;�YI;�}I;�I;�I;�I;v�I;��I;}�I;��I;ܘI;�I;�pI;�^I;�NI;W@I;�3I;i(I;�I;"I;�I;�I;EI;��H;#�H;��H;1�H;"�H;i�H;�H;�H;��H;�H;��H;�H;�H;�H;�H;e�H;"�H;/�H;��H;"�H;��H;GI;�I;�I; I;�I;g(I;�3I;V@I;�NI;�^I;�pI;�I;טI;��I;|�I;��I;r�I;�I;	�I;�I;�}I;�YI;?7I;<I;I;      a�I;�I;��I;w�I;�I;�I;��I;��I;�I;}�I;�I;��I;݃I;sI;	cI;5TI;�FI;_:I;4/I;4%I;dI;�I;�I;I;�I;��H;#�H;��H;D�H;!�H;W�H;��H;��H;�H;Z�H;�H;��H;��H;X�H;�H;��H;��H;W�H;�H;?�H;��H;�H;��H;�I;I;�I;�I;dI;2%I;3/I;\:I;�FI;7TI;	cI; sI;݃I;��I;�I;}�I;�I;��I;��I;�I;$�I;y�I;��I;׿I;      ��I;��I;D�I;P�I;L�I;p�I;v�I;��I;:�I;��I;L}I;�oI;TbI;�UI;�II;Q>I;�3I;=*I;�!I;�I;�I;�I;7I;pI;c�H;��H;��H;C�H;2�H;U�H;��H;��H;��H;��H;z�H;4�H;-�H;0�H;y�H;��H;��H;��H;��H;S�H;,�H;B�H;��H;��H;f�H;mI;9I;�I;�I;�I;�!I;:*I;�3I;T>I;�II;�UI;QbI;�oI;N}I;��I;=�I;��I;w�I;h�I;V�I;S�I;H�I;��I;      ��I;��I;_�I;O�I;��I;׋I;��I;�zI;	qI;
gI;�\I;�RI;�HI;�>I;�5I;-I;�$I;vI;�I;�I;#I;"I;�I;��H;��H;��H;1�H;#�H;[�H;��H;��H;��H;��H;�H;��H;{�H;\�H;y�H;��H;�H;��H;��H;��H;��H;W�H;#�H;+�H;��H;��H;��H;�I;$I;I;�I;�I;tI;�$I;-I;�5I;�>I;�HI;�RI;�\I;
gI;qI;�zI;��I;׋I;��I;T�I;\�I;��I;      UvI;�uI;�sI;�pI;�lI;kgI;haI;�ZI;�SI;LI;aDI;�<I;5I;�-I;w&I;�I;eI;�I;FI;W	I;�I;� I;v�H;r�H;��H;!�H;!�H;[�H;��H;��H;��H;��H;��H;Z�H;�H;��H;��H;��H;	�H;]�H;��H;��H;��H;��H;��H;Z�H;�H;$�H;��H;q�H;z�H;� I;�I;S	I;FI;�I;eI;�I;u&I;�-I;5I;�<I;^DI;LI;�SI;�ZI;oaI;cgI;�lI;�pI;�sI;�uI;      �WI;-WI;�UI;�SI;ePI;�LI;"HI;CI;�=I;�7I;	2I;,I;(&I;h I;�I;}I;�I;�I;�I;�I;3 I;��H;��H;j�H;*�H;4�H;c�H;��H;��H;��H;��H;��H;D�H;��H;{�H;@�H;K�H;A�H;x�H;��H;G�H;��H;��H;��H;��H;��H;b�H;6�H;.�H;d�H;�H;��H;, I;�I;�I;�I;�I;~I;�I;e I;'&I;,I;2I;�7I;�=I;CI;&HI;�LI;oPI;�SI;�UI;-WI;      �AI;tAI;C@I;�>I;<I;9I;�5I;�1I;�-I;)I;s$I;�I;0I;�I;:I;�I;�	I;I;�I;��H;}�H;��H;d�H;�H;S�H;��H;�H;��H;��H;��H;��H;B�H;��H;\�H;�H;��H;��H;��H;�H;_�H;��H;E�H;��H;��H;��H;��H;�H;��H;Y�H;�H;h�H;��H;w�H;�H;�I;I;�	I;�I;:I;�I;/I;�I;u$I;)I;�-I;�1I;�5I;9I;<I;~>I;P@I;tAI;      �1I;�1I;�0I;q/I;�-I;*+I;r(I;i%I;	"I;zI;�I;I;DI;�I;�I;[I;I;I;%�H;e�H;��H;j�H;l�H;��H;��H;T�H;�H;�H;��H;�H;W�H;��H;]�H;��H;��H;��H;~�H;��H;��H;��H;_�H;��H;V�H;�H;��H;�H;�H;V�H;��H;��H;q�H;h�H;��H;^�H;#�H;I;I;ZI;�I;�I;BI;I;�I;xI;	"I;e%I;v(I;*+I;�-I;t/I;�0I;�1I;      �'I;�'I;�&I;�%I;$I;"I;�I;MI;rI;�I;TI;?I;�I;�
I;�I;�I;�I;0�H;��H;(�H;�H;��H;�H;b�H;��H;��H;w�H;[�H;~�H;��H;�H;{�H;�H;��H;��H;\�H;X�H;a�H;~�H;��H;�H;|�H;�H;��H;w�H;X�H;x�H;��H;��H;c�H;
�H;��H;�H;"�H;��H;3�H;�I;�I;�I;�
I;�I;<I;TI;�I;qI;JI;�I;"I;$I;�%I;�&I;�'I;      �!I;�!I;	!I; I;�I;�I;�I;�I;I;|I;�I;�I;�
I;I;TI;�I;��H;\�H;�H;��H;��H;�H;N�H;��H;T�H;�H;�H; �H;;�H;�H;��H;C�H;��H;��H;a�H;+�H;.�H;/�H;_�H;��H;��H;D�H;��H;x�H;5�H; �H;�H;�H;W�H;��H;R�H;�H;��H;��H;�H;b�H;��H;�I;TI;I;�
I;�I;�I;yI;I;�I;�I;�I;�I;" I;!I;�!I;      �I;�I;@I;+I;�I;#I;WI;*I;�I;+I;�I;�I;
I;;I;bI;�I;Y�H;��H;��H;s�H;��H;��H;�H;��H;-�H;��H;��H;��H;1�H;`�H;��H;J�H;��H;{�H;W�H;(�H;�H;-�H;T�H;~�H;��H;K�H;��H;Y�H;,�H;��H;��H;��H;.�H;��H;"�H;��H;x�H;o�H;��H;��H;W�H;�I;aI;;I;	
I;�I;�I;)I;�I;(I;ZI;"I;�I;0I;=I;�I;      �!I;�!I;!I; I;�I;�I;�I;�I;I;{I;�I;�I;�
I;I;TI;�I;��H;\�H;�H;��H;��H;�H;N�H;��H;T�H;�H;�H;�H;<�H;}�H;��H;D�H;��H;��H;b�H;+�H;.�H;.�H;_�H;��H;��H;D�H;��H;v�H;5�H;��H;�H;�H;W�H;��H;R�H;�H;��H;��H;�H;b�H;��H;�I;SI;I;�
I;�I;�I;vI;I;�I;�I;�I;�I;& I;	!I;�!I;      �'I;�'I;�&I;�%I;$I;"I;�I;PI;rI;�I;VI;?I;�I;�
I;�I;�I;�I;2�H;��H;(�H;�H;��H;�H;`�H;��H;��H;x�H;\�H;~�H;��H;�H;z�H;�H;��H;��H;^�H;X�H;a�H;�H;��H;�H;{�H;�H;��H;w�H;W�H;x�H;��H;��H;b�H;
�H;��H;�H;"�H;��H;3�H;�I;�I;�I;�
I;�I;=I;TI;I;qI;NI;�I;"I;$I;�%I;�&I;�'I;      �1I;�1I;�0I;r/I;�-I;0+I;p(I;l%I;"I;xI;�I;I;DI;�I;�I;ZI;I;I;%�H;d�H;��H;k�H;l�H;��H;��H;V�H;�H;�H; �H;�H;U�H;��H;]�H;��H;��H;��H;~�H;��H;��H;��H;]�H;��H;U�H;�H;��H;��H;�H;W�H;��H;��H;q�H;k�H;��H;`�H;&�H;I;I;[I;�I;�I;BI;I;�I;wI;	"I;f%I;y(I;-+I;�-I;v/I;�0I;�1I;      �AI;zAI;H@I;{>I;<I;9I;�5I;�1I;�-I;)I;u$I;�I;0I;�I;=I;�I;�	I;I;�I;��H;}�H;��H;c�H;�H;V�H;��H;�H;��H;��H;��H;��H;A�H;��H;[�H;�H;��H;��H;��H;�H;\�H;��H;D�H;��H;��H;��H;��H;�H;��H;V�H;�H;j�H;��H;v�H;��H;�I;I;�	I;�I;:I;�I;0I;�I;s$I;)I;�-I;�1I;�5I;9I;<I;�>I;T@I;vAI;      �WI;/WI;�UI;�SI;ePI;�LI;%HI;CI;�=I;�7I;2I;
,I;)&I;g I;�I;I;�I;�I;�I;�I;4 I;��H;��H;g�H;.�H;6�H;c�H;��H;��H;��H;��H;��H;B�H;��H;|�H;@�H;K�H;D�H;x�H;��H;D�H;��H;��H;��H;��H;��H;a�H;7�H;+�H;a�H;�H;��H;, I;�I;�I;�I;�I;I;�I;g I;)&I;,I;2I;�7I;�=I;CI;'HI;�LI;gPI;�SI;�UI;,WI;      MvI;�uI;�sI;�pI;�lI;jgI;iaI;�ZI;�SI;LI;bDI;�<I;5I;�-I;x&I;�I;hI;�I;GI;U	I;�I;� I;w�H;r�H;��H; �H;�H;\�H;��H;��H;��H;��H;��H;Y�H;�H;��H;��H;��H;	�H;\�H;��H;��H;��H;��H;��H;X�H;�H;&�H;��H;n�H;{�H;� I;�I;T	I;GI;�I;hI;�I;x&I;�-I;5I;�<I;aDI;LI;�SI;�ZI;oaI;ggI;�lI;�pI;�sI;�uI;      ��I;��I;Y�I;V�I;��I;�I;��I;�zI;qI;gI;�\I;�RI;�HI;�>I;�5I;-I;�$I;wI;�I;�I;%I;%I;�I;��H;��H;��H;/�H;%�H;[�H;��H;��H;��H;��H;�H;��H;y�H;\�H;{�H;��H;�H;��H;��H;��H;��H;U�H;�H;-�H;��H;��H;��H;�I;%I;I;�I;�I;vI;�$I;-I;�5I;�>I;�HI;�RI;�\I;gI;qI;�zI;��I;ԋI;��I;`�I;c�I;��I;      ��I;��I;T�I;K�I;=�I;v�I;s�I;��I;B�I;��I;M}I;�oI;TbI;�UI;�II;T>I;�3I;?*I;~!I;�I;�I;�I;9I;qI;f�H;��H;��H;C�H;0�H;Q�H;��H;��H;��H;��H;y�H;3�H;,�H;3�H;y�H;��H;��H;��H;��H;S�H;)�H;=�H;��H;��H;c�H;iI;:I;�I;�I;�I;�!I;9*I;�3I;V>I;�II;�UI;TbI;�oI;L}I;��I;>�I;��I;y�I;p�I;N�I;N�I;V�I;��I;      m�I;׿I;��I;v�I;�I;)�I;��I;��I;�I;}�I;�I;��I;߃I;sI;cI;7TI;�FI;`:I;4/I;4%I;eI;�I;�I;I;�I;��H;�H;��H;D�H;�H;U�H;��H;��H;��H;[�H;��H;��H;��H;X�H;�H;��H;��H;W�H;�H;?�H;��H;�H;��H;�I;I;�I;�I;aI;2%I;4/I;\:I;�FI;8TI;cI;sI;݃I;��I;�I;�I;�I;��I;��I;�I;$�I;y�I;��I;׿I;      a I;0I;<I;Q7I;�YI;�}I;�I;�I;�I;u�I;��I;��I;��I;ܘI;	�I;�pI;�^I;�NI;V@I;�3I;k(I;�I; I;�I;�I;@I;��H;#�H;��H;.�H;!�H;h�H;�H;�H;�H;�H;��H;�H;|�H;�H;�H;f�H;"�H;.�H;��H;�H;��H;II;�I;�I;"I;�I;g(I;�3I;V@I;�NI;�^I;�pI;�I;טI;��I;y�I;��I;r�I;�I;�I;�I;�}I;�YI;T7I;>I;I;      �uF;w�F;��F;R!G;C�G;H;��H; �H;5KI;"�I;��I;��I;c�I;��I;�I;M�I;'}I;AhI;�UI;[EI;P7I;�*I;- I;I;^I;�I;DI;��H;��H;��H;$�H;=�H;��H;[�H;��H;�H;��H;�H;��H;[�H;��H;;�H;&�H;��H;��H;��H;DI;�I;\I;I;- I;�*I;L7I;[EI;�UI;:hI;(}I;M�I;��I;��I;`�I;��I;��I;%�I;+KI;�H;��H;�H;N�G;X!G;��F;i�F;      ��?;�@;�@;�A;��B;�C;$CE;|vF;��G;�\H;x�H;�mI;b�I;�I;#�I;��I;��I;c�I;ppI;V[I;III;�9I;d,I;� I;tI;YI;�I;�I;j�H;��H;��H;-�H;S�H;��H;��H;Z�H;1�H;Z�H;��H;��H;V�H;+�H;��H;��H;c�H;�I;�I;`I;oI;� I;e,I;�9I;GII;V[I;rpI;_�I;��I;��I; �I;�I;b�I;�mI;t�H;�\H;��G;zvF;&CE;��C;��B;�A;�@;�@;      0�1;��1;�73;�25;z�7;��:;.|=;!Q@;Y�B;BE;��F;]H;��H;qI;̶I;��I;��I;�I;R�I;�vI;�_I;�KI;;I;�,I;� I;I;�I;I;uI;��H;t�H;o�H;#�H;��H;n�H;��H;��H;��H;m�H;��H;$�H;n�H;u�H;��H;qI;I;�I;I;� I;�,I;;I;�KI;_I;�vI;S�I;�I;��I;��I;ƶI;qI;��H;YH;��F;DE;U�B;Q@;1|=;��:;��7;�25;�73;��1;      d�;x�; ];@X;�n!;�8';dI-;�93;��8;|=;
lA;LzD;f�F;�/H;�I;ʔI;��I;n�I;ܵI;��I;zI;vaI;sLI;;I;d,I;) I;I;�I;>I;�I;x�H;��H;g�H;o�H;�H;V�H;&�H;S�H;�H;l�H;e�H;��H;{�H;�I;7I;�I; I;. I;`,I;;I;sLI;taI;zI;��I;ݵI;g�I;��I;ǔI;�I;�/H;f�F;IzD;lA;|=;��8;�93;dI-;�8';�n!;BX;�\;b�;      Zo�:���:CK�:�Y�:F��:�;�;��;��$;�G.;P6;m�<;+�A;�E;SG;"�H;mI;��I;H�I;Q�I;��I;�{I;saI;�KI;�9I;�*I;�I;�I;�I;%I;� I;��H;��H;m�H;��H;�H;��H;�H;��H;h�H;��H;��H;� I;(I;�I;�I;�I;�*I;�9I;�KI;saI;�{I;��I;P�I;H�I;�I;mI; �H;
SG;�E;*�A;i�<;P6;�G.;��$;��;�;�;p��:�Y�:=K�:x��:       &m8���80`u9���9H�9:��:�W�:@r�:A� ;�F;9o!;q�-;�^7;Ol>;OC;�uF;PQH;�II;��I;��I;��I;��I;{zI;�_I;BII;G7I;`(I;bI;�I;I;�I;, I;u�H;��H;�H;��H;w�H;��H; �H;��H;s�H;) I;�I;I;�I;`I;`(I;I7I;=II;�_I;zzI;��I;��I;��I;��I;�II;NQH;�uF;�NC;Ol>;�^7;n�-;;o!;�F;=� ;Dr�:�W�:��:��9:���9�`u9���8      {��%��yi�V�غh����*��׭���9J��:>��:n��:�/;h�$;��1;g;;��A;��E;�H;35I;;�I;��I;P�I;��I;�vI;S[I;ZEI;�3I;5%I;�I;�I;S	I;�I;�H;d�H;(�H;��H;o�H;��H;"�H;]�H;|�H;�I;T	I;�I;�I;4%I;�3I;[EI;N[I;�vI;��I;M�I;��I;9�I;35I;�H;��E;��A;g;;��1;g�$;�/;n��:<��:F��:���9�׭� �*�\���l�غzi�)��      ��ͻLɻ�����d�����B�]�� ��潺���h8�9���:-T�:�;�Y;I-;v9;\�@;�\E;��G;35I;��I;G�I;ܵI;S�I;kpI;�UI;Q@I;6/I;!I;�I;CI;�I;�I;"�H;��H;�H;��H;�H;��H;�H;�I;�I;DI;�I;{!I;3/I;Q@I;�UI;dpI;V�I;ٵI;G�I;��I;25I;��G;�\E;Z�@;p9;I-;�Y;�;-T�:���:X8�9����潺� �C�]�����d������Hɻ      �iO�ߔK��o@���.���������ɻ�G��joE���غ(�����9�p�:�B�:�;n*;��7;�P@;�\E;�H;�II;��I;n�I;�I;`�I;;hI;�NI;d:I;?*I;xI;�I;�I;I;I;2�H;a�H;��H;b�H;-�H;I;I;�I;�I;xI;:*I;b:I;�NI;:hI;V�I;�I;g�I;��I;�II;�H;�\E;�P@;��7;l*;�;�B�:�p�:���9(����غjoE��G���ɻ���������.��o@�ߔK�      L�����2���?����N��Pp��D����hG�����34�>��� �n8��:G�:JG;�(;��7;Z�@;��E;TQH;mI;��I;��I;��I;#}I;�^I;�FI;�3I;�$I;aI;�I;�	I;I;�I;��H;P�H;��H;�I;I;�	I;�I;aI;�$I;�3I;�FI;�^I; }I;��I;��I;��I;mI;JQH;��E;Y�@;��7;�(;GG;A�:��: �n8D���24�����hG໇���D�Pp��N��@���3������      
��'�T5���������ϼ̡��X���iO�>���ɻ��p��D���o���g:�_�:CG;n*;r9;��A;�uF;$�H;ʔI;��I;��I;I�I;�pI;5TI;U>I;-I;�I;~I;�I;]I;�I;�I;�I;�I;�I;TI;�I;xI;�I;-I;Q>I;4TI;�pI;B�I;��I;��I;ǔI; �H;�uF;��A;o9;j*;CG;�_�:�g:��o��D⺙�p��ɻ>���iO�X��͡����ϼ������T5�&�      j��ѷ��%0v�r�a�$�G�@2+���ן�	����/����5��&��^f��ج���g:?�:
�;I-;g;;OC;SG;�I;ͶI; �I; �I;�I;cI;�II;�5I;t&I;�I;9I;�I;�I;MI;XI;NI;�I;�I;6I;�I;q&I;�5I;�II;
cI;�I;��I;�I;̶I;�I;SG;�NC;g;;I-;�;;�:��g:�ج�_f�(�����5��/��	���؟���@2+�%�G�s�a�%0v�ѷ��      ��ս��ѽ;�ƽ1����I�����Q�a�D4�<M���ϼ��K�K�N��LG��Zf���o���:�B�:�Y;��1;Wl>;�E;�/H;$qI;�I;��I;ܘI;sI;�UI;�>I;�-I;d I;�I;�I;�
I;I;/I;I;�
I;�I;�I;^ I;�-I;�>I;�UI; sI;טI;��I;��I;"qI;�/H;�E;Il>;��1;�Y;�B�:��:��o�bf�LG��N��K�K�����ϼ<M�D4�R�a�����I��1���;�ƽ��ѽ      �L+�  (���F�������ս�@���%���;V�%��ސ������MS�M��$��tD⺀�n8 q�:�;i�$;_7;/�A;n�F; �H;h�I;d�I;��I;�I;[bI;�HI;5I;(&I;0I;AI;�I;�
I;
I;�
I;�I;>I;/I;"&I;5I;�HI;YbI;��I;��I;_�I;a�I;��H;k�F;-�A;�^7;i�$;�;�p�: �n8|D�&��M���MS�����ސ�&���;V��%���@����ս����F���  (�      �T��f�����z��Yb�&�D��$�����ѽ�I��D�m�2+�������K�K�ﻕ�p�H������9-T�:�/;x�-;j�<;LzD;`H;�mI;��I;|�I;��I;�oI;�RI;�<I;,I;�I;I;/I;�I;�I;�I;/I;I;�I; ,I;�<I;�RI;�oI;��I;z�I;��I;�mI;]H;MzD;i�<;k�-;�/;#T�:���9H�����p��L�K�������2+�D�m��I����ѽ���$�'�D��Yb���z�f���      ?�׾��Ҿž�j��������z�S�H�)��ez�G$���/v�2+�ސ�����5��ɻ74�H(�����:b��:?o!;P6;lA;��F;w�H;��I;��I;�I;M}I;�\I;aDI;2I;s$I;�I;HI;�I;�I;�I;HI;�I;r$I;2I;]DI;�\I;M}I;�I;��I;��I;s�H;��F;lA;P6;1o!;`��:~��:P(��94��ɻ��5���ސ�2+��/v�G$��ez�)��S�H���z������j��ž��Ҿ      H(��$�d��P������~���`���Yb���'��U�G$��D�m�&����ϼ�/��=��������غP8�9B��:�F;�G.;|=;LE;�\H;!�I;v�I;|�I;��I;gI;LI;�7I;)I;rI;rI;rI;'I;qI;rI;pI;)I;�7I;LI;gI;��I;z�I;s�I;�I;�\H;KE;|=;�G.;�F;>��:88�9��غ����>���/����ϼ&��D�m�G$���U���'��Yb��`���~�����P��d���$�      <�}���w�#f���K�r,�}�
�;�׾ �����k���'�ez꽝I���;V�<M�	����iO�lG�qoE����@��:G� ;��$;��8;]�B; �G;0KI;�I;�I;E�I;qI;�SI;�=I;�-I;	"I;kI;I;�I;I;kI;"I;�-I;�=I;�SI;qI;B�I;�I;�I;/KI;��G;b�B;��8;��$;;� ;@��:ȱ�soE�lG໫iO�	���<M��;V��I��ez���'���k� ���;�׾}�
�r,���K�#f���w�      ��p�������.蒿��w��F�d��ʰ� ����Yb�)����ѽ�%��D4�؟�X�����H���潺В�9Nr�:��;�93;+Q@;~vF;�H;	�I;��I;��I;�zI;�ZI;CI;�1I;c%I;?I;�I;"I;�I;BI;b%I;�1I;CI;�ZI;�zI;��I;��I;�I;�H;|vF;*Q@;�93;��;6r�:В�9�潺H�����X��ٟ�D4��%����ѽ)���Yb� ���ʰ�d���F���w�.蒿����p���      4��������㿊�ɿ���ʅ����P�d��;�׾�`��S�H����@��R�a���͡���D��ɻ� ��׭��W�:�;bI-;8|=;!CE;��H;�I;��I;w�I;��I;jaI;#HI;�5I;r(I;�I;�I;SI;�I;�I;p(I;�5I;"HI;haI;��I;v�I;��I;�I;��H; CE;;|=;fI-;�;�W�:�׭�� ��ɻ�D�͡����R�a��@����S�H��`��;�׾d����P�ʅ�������ɿ�㿳���      ř$��x �"��:���޿o���ʅ���F�}�
��~����z��$���ս���A2+���ϼPp�����M�]��*���:�;�8';��:;��C;�H;�}I;�I;t�I;ۋI;ogI;�LI;9I;9+I;!"I;�I;*I;�I;""I;7+I;9I;�LI;jgI;ًI;s�I;"�I;�}I;H;��C;��:;�8';�;��:�*�Q�]�����Pp���ϼA2+������ս�$���z��~��}�
��F�ʅ��o����޿:��"���x �      J�Q���K���;�ř$��;
��޿�����w�r,���澝���'�D������I��$�G�����N��������P�����9:\��:�n!;��7;��B;I�G;�YI;+�I;Z�I;��I;�lI;sPI;<I;�-I;
$I;�I;�I;�I;$I;�-I;<I;sPI;�lI;��I;Z�I;.�I;�YI;Q�G;��B;��7;�n!;V��:x�9:T����������N�����$�G��I������'�D��������r,���w�����޿�;
�ř$���;���K�      T����{���d��F�ř$�:����ɿ.蒿��K�P���j���Yb�F�1���s�a����?�����.��d��j�غ��9�Y�:.X;�25;#�A;X!G;H7I;s�I;C�I;R�I;�pI;�SI;~>I;y/I;�%I;" I;0I; I;�%I;v/I;�>I;�SI;�pI;T�I;B�I;v�I;L7I;c!G;!�A;�25;.X;�Y�:���9f�غ�d����.�?������s�a�1���F��Yb��j��P����K�.蒿��ɿ:��ř$��F���d��{�      ����#P�������d���;�#���㿲���#f�d��ž��z���<�ƽ%0v�T5�2����o@�����|i��`u9AK�:];�73;%�@;��F;FI;��I;P�I;S�I;�sI;�UI;?@I;�0I;�&I;!I;0I;!I;�&I;�0I;A@I;�UI;�sI;X�I;M�I;��I;LI;��F;"�@;�73;];;K�:p`u9yi������o@�2���T5�%0v�<�ƽ����z�žd��#f�������#����;���d����#P��      �,��a��#P���{���K��x �����p�����w��$���Ҿf���  (���ѽҷ��'�����K�Fɻ)�����8x��:z�;��1;�@;k�F;I;޿I;�I;��I;�uI;%WI;fAI;�1I;�'I;�!I;�I;�!I;�'I;�1I;hAI;&WI;�uI;��I;�I;�I;#I;{�F;�@;��1;z�;r��:���8'��Hɻ�K����'�ҷ����ѽ  (�f�����Ҿ�$���w�p��������x ���K��{�#P��a��      D(��q'���o��N�d��X1�~x�	Ŀ����3�w���x����4�k��Y+���'���ü:yY��kٻp&���p�N��:;;��0;��?;��F;j I; �I;��I;,�I;g�I;LdI;�KI;�9I;m.I;�'I;�%I;�'I;k.I;�9I;�KI;MdI;g�I;0�I;��I;�I;j I;΀F;��?;��0;6;B��:��p�p&��kٻ:yY���ü�'�Y+��k�ཽ�4��x��w���3����	Ŀ~x��X1�d�N��o��q'��      q'���X��f^�������]]���,�P9�6g��T�����/����o��g1��hܽ���-$�_l���|U�f�Ի�!� �,�{�:�;�51;��?;7�F;A'I;b�I;�I;=�I;��I;�cI;>KI;x9I;.I;{'I;�%I;v'I; .I;w9I;@KI;�cI;��I;A�I;�I;d�I;A'I;B�F;��?;�51;�;s�: �,�~!�f�Ի�|U�_l���-$����hܽg1��o���ྚ�/�T���6g��P9���,��]]�����f^���X��      �o��f^���ē��4z�5K�h��R��&ﱿT�v��X#���Ѿń��&�p�нc̀�_��v���L�I��ǻ�4��"9��:6�; �2;��@;��F;�:I;��I;��I;��I;u�I;KbI;�II;�8I;Z-I;�&I;�$I;�&I;[-I;�8I;�II;KbI;r�I;��I;��I;��I;�:I;��F;��@;�2;6�;��:@"9�4��ǻM�I�v���_��c̀�p�н�&�ń���Ѿ�X#�T�v�&ﱿR��h��5K��4z��ē�f^��      N������4z���V��X1��<�tؿ����RZ��	�(���IUo����^y��.l�Y��R��B�7�������ų9��:��;X�4;jtA;_2G;�XI;��I;J�I;�I;�I;�_I;�GI;"7I;�+I;�%I;�#I;�%I;�+I;!7I;�GI;�_I;�I;�I;M�I;��I;�XI;i2G;jtA;Y�4;��;���:�ų9�����B�7��R��Y�.l�^y�����IUo�(����	��RZ����tؿ�<��X1���V��4z�����      d��]]�5K��X1�Zf��nQ��S���[58��A���נ���O���_什�Q����@ߓ��� ��V���氺��":Ը�: ;�07;�B;0�G;�{I;��I;��I;��I;:|I;7\I;LEI;5I;3*I;1$I;)"I;-$I;5*I;5I;MEI;8\I;7|I;��I;��I;��I;�{I;:�G;�B;�07; ;Ը�:�":�氺�V���� �@ߓ�����Q�_什����O��נ��A��[58�S���nQ���Zf��X1�5K��]]�      �X1���,�h���<��5g��e_���U�͂�֌Ⱦń�*�-�i��P ��&�2�?ټb�{�"��n�(�O���u:�P ;�&;+#:;=�C;�%H;�I;!�I;��I;�I;]vI;�WI;�AI;z2I;(I;D"I;^ I;@"I;(I;w2I;�AI;�WI;\vI;�I;��I;'�I;�I;�%H;@�C;)#:;�&;�P ;��u:�O��n�"�b�{�?ټ&�2�P ��i��*�-�ń�֌Ⱦ͂��U�e_��5g��<�h����,�      ~x�P9�R��sؿnQ��e_��6�_��X#�p���f��9�S�{�����l�B�	w�� �M���Ի��+�0=T���:�e;�\,;�/=;�BE;Q�H;z�I;��I;��I;��I;�oI;�RI;>I;]/I;}%I;�I;FI;�I;~%I;^/I;>I;�RI;�oI;��I;��I;��I;x�I;Z�H;�BE;�/=;�\,;�e;��:�<T���+���Ի�M�	w��B�l�����{�9�S��f��p���X#�6�_�e_��nQ��sؿR��P9�      	Ŀ6g��&ﱿ���S����U��X#�t��d���IUo��#��hܽ����n<����<����� ��᝻F�Ժxt�9`��:�V;̇2;� @;T�F;�I;��I;C�I;)�I;i�I; hI;MI;�9I;�+I;�"I;jI;�I;iI;�"I;�+I;�9I;MI;�gI;o�I;,�I;G�I;��I;�I;Y�F;� @;Ї2;�V;Z��:�t�9D�Ժ�᝻�� �;�������n<�����hܽ�#�IUo�d���t���X#��U�S������&ﱿ6g��      ���T���T�v��RZ�[58�͂�p��d���foy�]1�_O��\什�`�M�����pyY�$�컘�T��1�x�u:���:F#;98;	�B;f�G;�lI;�I;�I;-�I;v�I;�_I;GI;�4I;%(I;�I;�I;I;�I;�I;&(I;�4I;GI;�_I;z�I;/�I;�I;�I;�lI;p�G;�B;98;J#;���:��u:�1���T�"��pyY����M���`�[什_O��]1�foy�d���p��͂�[58��RZ�T�v�T���      �3���/��X#��	��A��֌Ⱦ�f��HUo�^1�˰��|n��Ҽx��'��>ټ�@���k�м��"����39�#�:.R;	e-;�/=;�	E;\xH;��I;�I;p�I;��I;vI;aWI;�@I;�/I;#$I;;I;�I;6I;�I;<I;%$I;�/I;�@I;eWI;vI;�I;v�I;�I;��I;dxH;�	E;�/=;e-;,R;�#�:��39��μ���k��@���>ټ�'�Ѽx�|n��˰��]1�HUo��f��֌Ⱦ�A���	��X#���/�      v���ྃ�Ѿ(����נ�ń�9�S��#�_O��|n��J̀���2���𛼃�>� �Ի��B��#�4m:�G�:^ ;��5;�FA;��F;�I;N�I;Q�I;��I;j�I;njI;�NI;:I;�*I;�I;�I;�I;KI;�I;�I;�I;�*I;:I;�NI;rjI;o�I;��I;U�I;N�I;�I;��F;�FA;��5;^ ;�G�:Dm:�#���B���Ի��>�������2�J̀�|n��_O���#�9�S�ń��נ�(�����Ѿ��      �x���o��ń�IUo���O�*�-�{��hܽ\什Ҽx���2�tb��VR��X|U�Z2��:��$갺�u�9��:D;��,;�h<;crD;N%H;��I;g�I;��I;�I;�I;�^I;FI;V3I;�%I;�I;^I;hI;4I;hI;^I;�I;�%I;U3I;FI;�^I;�I;�I;��I;g�I;ʏI;S%H;jrD;�h<;��,;D;��:�u�9갺8��Y2��V|U�UR��tb����2�Ҽx�[什�hܽ{�*�-���O�IUo�ń��o��      ��4�f1��&������i�ཅ�������`��'���UR��F�]����#V���X�� Io����:h�;$#;�6;QtA;R�F;�	I;r�I;��I;p�I;�I;�pI;�SI;�=I;�,I;w I;�I;�I;GI;9I;FI;�I;�I;y I;�,I;�=I;�SI;�pI;�I;p�I;��I;|�I;�	I;W�F;VtA;�6;1#;n�;���: Go��X��!V��~��D�]�TR����'��`��������h��������&�f1�      j�ྲྀhܽo�н^y��_什P ��l��n<�M���>ټ��W|U���������1�������u:Wl�:�;b71;S)>;S	E;
JH;T�I;��I;��I;�I;׃I;YbI;�HI;&5I;c&I;gI;qI;<I;%I;
I;%I;:I;rI;hI;`&I;-5I;�HI;bbI;��I;�I;��I;��I;W�I;JH;Z	E;S)>;n71;
�;Sl�:��u:�����1��������V|U����>ټM���n<�l�P ��_什^y��o�н�hܽ      Y+����c̀�-l��Q�&�2�B��������@����>�Z2��$V���1�����#R:���:�;t\,;1;;�;C;�eG;U9I;��I;/�I;��I;C�I;�qI;�TI;b>I;8-I;3 I;zI;rI;�
I;I;I;I;�
I;tI;~I;0 I;<-I;f>I;�TI;�qI;C�I;��I;7�I;��I;W9I;�eG;�;C;=;;z\,;�;���: $R:���1�"V��X2����>��@��������B�%�2��Q�-l�c̀���      �'��-$�_��Y����?ټw��;���pyY��k� �Ի:��
Y�������#R:���:�R;�);܍8;��A;��F;3�H;)�I;��I;��I;��I;�I;�`I;�GI;�4I;�%I;JI;�I;�I;qI;I;FI;I;mI;�I;�I;HI;�%I;�4I;�GI;�`I;�I;��I;��I;��I;*�I;;�H;��F;��A;��8;�);�R;���:$R:����Y��:����Ի�k�oyY�;���	w��	?ټ���Y�^���-$�      ��ü^l��w����R��?ߓ�b�{��M��� �"��˼����B�갺@Ho���u:���:�R;/�';17;��@;��E;�lH;.�I;h�I;��I;�I;x�I;�lI;�QI;&<I;�+I;�I;�I;eI;�I;CI;0I;�I;,I;AI;�I;eI;�I;�I;�+I;*<I;�QI;�lI;s�I;�I;��I;h�I;2�I;�lH;��E;��@;17;3�';�R;���:��u: Ho�갺��B�˼�� �컌� ��M�a�{�@ߓ��R��x���\l��      4yY��|U�M�I�@�7��� �"���Ի�᝻��T���#��u�9���:Ql�:�;�);17;/ @;:]E;�$H;dkI;
�I;U�I;��I;'�I;�wI;�ZI;�CI;w1I;N#I;%I;�I;-	I;rI;9I;m�H;��H;j�H;6I;rI;.	I;�I;,I;S#I;z1I;�CI;�ZI;�wI;.�I;��I;R�I;�I;hkI;�$H;>]E;. @;17;�);�;Sl�:���:�u�9�#����T��᝻��Ի"��� �A�7�K�I��|U�      �kٻn�Ի�ǻ����V���n���+�6�Ժ��1�0�39Tm:��:l�;�;z\,;��8;��@;A]E;�
H;LVI;q�I;��I;��I;c�I;��I;�bI;bJI;%7I;�'I;�I;.I;�
I;8I;;I;i�H;��H;y�H;��H;f�H;;I;9I;�
I;3I;�I;�'I;*7I;`JI;�bI;�I;g�I;��I;��I;v�I;PVI;�
H;<]E;��@;ݍ8;{\,;�;l�;��:`m: �39�1�8�Ժ��+��n��V������ǻl�Ի      p&��!��4���氺�O��<T�ht�9��u:�#�:�G�:D;*#;i71;;;;��A;��E;�$H;MVI;�I;��I;�I;��I;��I;iI;'PI;<I;�+I;I;�I;�I;�I;�I;5�H;��H;��H;�H;��H;��H;3�H;�I;�I;�I;�I;I;�+I;<I;&PI;iI;��I;��I;�I;��I;�I;PVI;�$H;��E;��A;=;;g71;)#;D;�G�:�#�:��u:�t�9�<T��O��氺���4��!�       �p� �,�� 9�ų9Č":��u:��:`��:���:.R;\ ;��,;�6;S)>;�;C;��F;�lH;lkI;t�I;��I;��I;�I;r�I;�mI;wTI;%@I;�/I;""I;WI;�I;�I;�I;u�H;u�H;��H;X�H;��H;Q�H;��H;u�H;u�H;�I;�I;�I;WI;'"I;�/I;%@I;~TI;�mI;n�I;�I;��I;��I;v�I;ikI;�lH;��F;�;C;P)>;�6;��,;` ;.R;���:Z��:��:|�u:�":�ų9p!9 �,�      4��:��:��:��:���:�P ;�e;�V;J#;e-;��5;�h<;RtA;X	E;�eG;8�H;2�I;�I;��I;�I;�I;�I;pI;LWI;�BI;@2I;�$I;sI;oI;B	I;tI;��H;��H;�H;\�H;6�H;��H;0�H;Y�H;�H;��H;��H;yI;D	I;oI;wI;�$I;A2I;�BI;KWI;pI;��I;�I;�I;��I;�I;3�I;8�H;�eG;V	E;StA;�h<;��5;e-;L#;�V;�e;�P ;��:���:��:s�:      G;�;,�;��;� ;�&;�\,;ۇ2;98;�/=;�FA;orD;U�F;JH;[9I;.�I;n�I;Z�I;��I;��I;p�I;pI;IXI;�DI;�3I;]&I;I;�I;�
I;oI;��H;��H;��H;��H;<�H;J�H;�H;E�H;9�H;��H;��H;��H;��H;oI;~
I;�I;I;_&I;�3I;�DI;EXI;pI;s�I;��I;��I;U�I;n�I;.�I;[9I;JH;U�F;orD;�FA;�/=;98;ׇ2;�\,;�&; ;��;(�;�;      ��0;�51;
�2;Q�4;�07;-#:;�/=;� @;�B;�	E;��F;P%H;�	I;U�I;��I;��I;��I;��I;c�I;��I;�mI;DWI;�DI;�4I;='I;-I;�I;{I;;I;. I;,�H;��H;|�H;��H;e�H;��H;k�H;��H;c�H;��H;|�H;��H;1�H;. I;8I;I;�I;1I;B'I;�4I;�DI;HWI;�mI;��I;c�I;��I;��I;��I;��I;R�I;�	I;Q%H;��F;�	E;�B;� @;�/=;#:;�07;M�4;	�2;�51;      ��?;��?;��@;_tA;�B;F�C;�BE;W�F;j�G;`xH;�I;ˏI;u�I;��I;7�I;��I;�I;1�I;�I;iI;�TI;�BI;�3I;G'I;�I;|I;I;�I;� I;~�H;�H;k�H;a�H;��H;��H;/�H;��H;*�H;��H;��H;a�H;i�H;�H;��H;� I;�I;I;�I;�I;D'I;�3I;�BI;�TI;iI;�I;.�I;�I;��I;6�I;��I;x�I;͏I;�I;`xH;h�G;T�F;�BE;:�C;�B;]tA;�@;��?;      ��F;@�F;��F;\2G;%�G;�%H;Y�H;�I;�lI;��I;T�I;p�I;��I;��I;��I;��I;x�I;�wI;�bI;&PI;'@I;:2I;\&I;0I;yI;:I;I; I;��H;F�H;x�H;V�H;|�H;'�H;^�H;��H;��H;��H;[�H;(�H;~�H;S�H;z�H;F�H;��H; I;I;<I;�I;0I;[&I;@2I;'@I;%PI;�bI;�wI;{�I;��I;��I;��I;��I;p�I;X�I;��I;�lI;�I;Z�H;�%H;:�G;j2G;��F;@�F;      t I;H'I;�:I;�XI;�{I;�I;}�I;�I;�I;�I;U�I;��I;m�I;�I;C�I;�I;�lI;�ZI;cJI; <I;�/I;�$I;"I;I;I;I;I;��H;v�H;��H;L�H;T�H;��H;��H;�H;��H;q�H;��H;�H;��H;��H;R�H;P�H;��H;p�H;��H;I;I;I;�I;"I;�$I;�/I;<I;cJI;�ZI;�lI;�I;@�I;�I;m�I;��I;U�I;�I;�I;��I;v�I;�I;�{I;�XI;�:I;2'I;      ��I;d�I;��I;��I;��I;"�I;��I;C�I;�I;v�I;��I;�I;�I;ރI;�qI;�`I;�QI;�CI;%7I;�+I;'"I;oI;�I;}I;�I;� I;��H;l�H;��H;V�H;T�H;��H;��H;��H;��H;��H;q�H;��H;��H;��H;��H;��H;T�H;T�H;��H;j�H;��H;� I;�I;|I;�I;qI;%"I;�+I;#7I;�CI;�QI;�`I;�qI;݃I;�I;�I;��I;t�I;��I;@�I;��I;�I;��I;��I;��I;[�I;      ��I;��I;��I;[�I;��I;��I;��I;-�I;'�I;�I;n�I;�I;�pI;bbI;�TI;�GI;-<I;{1I;�'I;I;^I;iI;~
I;6I;� I;��H;m�H;��H;P�H;O�H;��H;P�H;@�H;��H;��H;��H;��H;��H;��H;��H;A�H;L�H;��H;M�H;L�H;��H;i�H;��H;� I;1I;{
I;iI;ZI;I;�'I;x1I;*<I;�GI;�TI;_bI;�pI;
�I;q�I;�I;(�I;,�I;��I;��I;��I;\�I;��I;��I;      ,�I;9�I;��I;
�I;��I;�I;��I;r�I;w�I;vI;ujI;�^I;�SI;�HI;d>I;�4I;�+I;N#I;�I;�I;�I;?	I;lI;, I;��H;?�H;��H;X�H;U�H;��H;*�H;�H;8�H;��H;�H;��H;��H;��H;�H;��H;6�H;�H;*�H;��H;O�H;X�H;��H;@�H;��H;) I;oI;@	I;�I;�I;�I;L#I;�+I;�4I;c>I;�HI;�SI;�^I;rjI;vI;v�I;k�I;��I;�I;��I;�I;��I;6�I;      d�I;��I;w�I;��I;4|I;]vI;�oI;hI;�_I;jWI;�NI;FI;�=I;.5I;@-I;�%I;�I;,I;2I;�I;�I;vI;��H;-�H;�H;w�H;M�H;Y�H;��H;-�H;	�H;�H;T�H;��H;u�H;-�H;��H;,�H;t�H;��H;W�H;�H;�H;*�H;��H;V�H;J�H;w�H;�H;,�H;��H;vI;�I;�I;5I;)I;�I;�%I;?-I;-5I;�=I;FI;�NI;jWI;�_I;hI;�oI;VvI;<|I;��I;v�I;��I;      JdI;�cI;DbI;�_I;)\I;�WI;�RI;MI;	GI;�@I;:I;]3I;�,I;i&I;5 I;MI;�I;�I;�
I;�I;�I;��H;��H;��H;k�H;O�H;Q�H;��H;U�H;�H;�H;M�H;��H;%�H;��H;��H;��H;��H;��H;&�H;��H;M�H;�H;�H;O�H;��H;O�H;O�H;n�H;��H;��H;��H;�I;�I;�
I;�I;�I;OI;3 I;g&I;�,I;Y3I;:I;�@I;GI;MI;�RI;�WI;1\I;�_I;NbI;�cI;      �KI;LKI;�II;�GI;IEI;�AI;>I;�9I;�4I;�/I;�*I;�%I;z I;mI;~I;�I;iI;.	I;=I;�I;~�H;��H;��H;u�H;a�H;t�H;��H;��H;H�H;;�H;Q�H;��H;�H;��H;J�H;�H;.�H;�H;H�H;��H;�H;��H;P�H;4�H;C�H;��H;��H;u�H;d�H;u�H;��H;��H;x�H;�I;?I;-	I;iI;�I;I;kI;y I;�%I;�*I;�/I;�4I;�9I;>I;�AI;LEI;�GI;JI;LKI;      �9I;x9I;�8I;7I;5I;k2I;]/I;�+I;'(I;-$I; I;�I;�I;xI;{I;�I;�I;sI;?I;7�H;|�H;�H;��H;��H;��H;�H;��H;��H;��H;��H;��H;%�H;��H;5�H;��H;��H;��H;��H;��H;9�H;��H;%�H;��H;��H;�H;��H;��H;�H;��H;��H;��H;�H;u�H;/�H;=I;vI;�I;�I;yI;xI;�I;�I; I;-$I;'(I;�+I;c/I;k2I;5I;7I;�8I;�9I;      ].I;9.I;_-I;�+I;?*I;
(I;�%I;�"I;�I;JI;�I;oI;�I;FI;�
I;uI;LI;8I;k�H;��H;��H;U�H;5�H;U�H;��H;P�H;�H;��H;��H;�H;o�H;��H;J�H;��H;��H;��H;}�H;��H;��H;��H;J�H;��H;m�H;�H;��H;��H;�H;P�H;��H;V�H;8�H;U�H;��H;��H;j�H;9I;LI;vI;�
I;FI;�I;jI;�I;JI;�I;�"I;�%I;(I;9*I;,I;\-I;:.I;      �'I;�'I;�&I;�%I;#$I;@"I;�I;sI;�I;�I;�I;sI;KI;)I;I;I;3I;h�H;��H;��H;^�H;.�H;B�H;��H;&�H;��H;��H;��H;��H;��H;,�H;��H;�H;��H;��H;c�H;q�H;f�H;��H;��H;�H;��H;)�H;��H;��H;��H;��H;��H;'�H;��H;F�H;/�H;W�H;��H;��H;m�H;3I;I;I;*I;HI;mI;�I;�I;�I;mI;  I;="I;&$I;�%I;�&I;�'I;      �%I;�%I;�$I;�#I;!"I;W I;JI;�I;I;:I;VI;?I;BI;'
I;I;JI;�I; �H;}�H;	�H;��H;��H;�H;[�H;��H;��H;i�H;s�H;��H;��H;��H;��H;/�H;��H;}�H;m�H;v�H;o�H;z�H;��H;0�H;��H;��H;��H;~�H;p�H;j�H;��H;��H;\�H;�H;��H;��H;�H;}�H; �H;�I;LI;I;'
I;@I;<I;YI;:I;I;�I;NI;W I;"I;�#I;�$I;�%I;      �'I;�'I;�&I;�%I;%$I;A"I;�I;pI;�I;�I;�I;sI;KI;,I;I;I;3I;g�H;��H;��H;`�H;/�H;B�H;��H;&�H;��H;��H;��H;��H;��H;,�H;��H; �H;��H;��H;c�H;q�H;f�H;��H;��H;�H;��H;)�H;��H;��H;��H;��H;��H;'�H;��H;F�H;.�H;W�H;��H;��H;m�H;2I;I;I;(I;HI;mI;�I;�I;�I;oI;�I;@"I;&$I;�%I;�&I;�'I;      T.I;:.I;Z-I;�+I;=*I;(I;�%I;�"I;�I;JI;�I;oI;�I;FI;�
I;tI;JI;;I;k�H;��H;��H;W�H;5�H;S�H;��H;O�H;�H;��H;��H;�H;n�H;��H;H�H;��H;��H;��H;}�H;��H;��H;��H;K�H;��H;m�H;�H;��H;��H;�H;Q�H;��H;S�H;9�H;V�H;��H;��H;j�H;9I;LI;uI;�
I;FI;�I;lI;�I;II;�I;�"I;�%I;
(I;<*I;,I;\-I;?.I;      �9I;x9I;�8I;7I;5I;r2I;]/I;�+I;)(I;-$I; I;�I;�I;xI;|I;�I;�I;uI;?I;5�H;|�H;�H;��H;��H;��H;�H;��H;��H;��H;��H;��H;#�H;��H;5�H;��H;��H;��H;��H;��H;6�H;��H;#�H;��H;��H;~�H;��H;��H;!�H;��H;��H;��H;�H;q�H;3�H;?I;uI;�I;�I;yI;xI;�I;�I; I;-$I;)(I;�+I;e/I;n2I;5I;7I;�8I;}9I;      �KI;RKI;�II;�GI;FEI;�AI;>I;�9I;�4I;�/I;�*I;�%I;z I;jI;I;�I;iI;/	I;?I;�I;~�H;��H;��H;u�H;d�H;r�H;��H;��H;H�H;9�H;O�H;��H;�H;��H;J�H;�H;.�H;�H;J�H;��H;�H;��H;O�H;2�H;A�H;��H;��H;u�H;a�H;r�H;��H;��H;w�H;�I;=I;-	I;hI;�I;I;kI;z I;�%I;�*I;�/I;�4I;�9I;>I;�AI;JEI;HI;JI;OKI;      CdI;�cI;9bI;�_I;)\I;�WI;�RI;MI;GI;�@I;:I;]3I;�,I;i&I;7 I;MI;�I;�I;�
I;�I;�I;��H;��H;��H;n�H;O�H;Q�H;��H;V�H;�H;�H;L�H;��H;"�H;��H;��H;��H;��H;��H;%�H;��H;L�H;�H;�H;N�H;��H;N�H;P�H;k�H;��H;��H;��H;�I;�I;�
I;�I;�I;OI;5 I;g&I;�,I;\3I;:I;�@I;GI;MI;�RI;�WI;)\I;�_I;?bI;�cI;      Z�I;��I;y�I;��I;8|I;]vI;�oI;hI;�_I;jWI;�NI;FI;�=I;/5I;@-I;�%I;�I;)I;3I;�I;�I;yI;��H;,�H;�H;r�H;J�H;X�H;��H;,�H;�H;�H;T�H;��H;v�H;,�H;��H;-�H;r�H;��H;T�H;�H;�H;)�H;��H;R�H;I�H;x�H;�H;)�H;��H;xI;�I;�I;6I;)I;�I;�%I;?-I;/5I;�=I;FI;�NI;hWI;�_I;hI;�oI;[vI;B|I;�I;}�I;��I;      5�I;@�I;��I;�I;��I;�I;��I;s�I;z�I;vI;pjI;�^I;�SI;�HI;g>I;�4I;�+I;O#I;�I;�I;�I;B	I;lI;* I;��H;;�H;��H;Z�H;U�H;��H;)�H;�H;4�H;��H;�H;��H;��H;��H;�H;��H;6�H;�H;)�H;��H;N�H;V�H;��H;@�H;��H;& I;pI;@	I;�I;�I;�I;L#I;�+I;�4I;d>I;�HI;�SI;�^I;pjI;vI;t�I;o�I;��I;ޟI;��I;�I;��I;9�I;      ��I;�I;��I;R�I;��I;��I;��I;,�I;/�I; �I;n�I;�I;�pI;`bI;�TI;�GI;*<I;}1I;�'I;I;`I;kI;|
I;5I;� I;��H;j�H;��H;P�H;J�H;��H;P�H;?�H;��H;��H;��H;��H;��H;��H;�H;@�H;N�H;��H;K�H;J�H;��H;i�H;��H;� I;/I;
I;kI;ZI;I;�'I;x1I;*<I;�GI;�TI;`bI;�pI;
�I;n�I;��I;*�I;-�I;��I;��I;��I;V�I;��I;��I;      �I;\�I;��I;��I;��I;.�I;��I;G�I;�I;v�I;��I;�I;�I;ރI;�qI;�`I;�QI;�CI;#7I;�+I;("I;qI;�I;I;�I;� I;��H;j�H;��H;Q�H;U�H;��H;��H;��H;��H;��H;q�H;��H;��H;��H;��H;��H;T�H;Q�H;��H;f�H;��H;� I;�I;xI;�I;oI;""I;�+I;&7I;�CI;�QI;�`I;�qI;݃I;�I;	�I;��I;v�I; �I;@�I;��I;�I;��I;��I;��I;\�I;      a I;O'I;�:I;�XI;�{I;�I;z�I;�I;�I;�I;U�I;��I;j�I;�I;C�I;�I;�lI;�ZI;cJI;<I;�/I;�$I;I;I;I;I;I;��H;w�H;��H;L�H;T�H;��H;��H;�H;��H;q�H;��H;�H;��H;��H;T�H;L�H;��H;p�H;��H;I;I;I;�I;"I;�$I;�/I;<I;fJI;�ZI;�lI;	�I;C�I;�I;k�I;��I;U�I;�I;�I;��I;~�I;�I;�{I;�XI;�:I;:'I;      ��F;?�F;��F;Y2G;*�G;&H;T�H;�I;�lI;��I;U�I;s�I;��I;��I;��I;��I;x�I;�wI;�bI;&PI;,@I;=2I;[&I;3I;I;7I;I;I;��H;C�H;z�H;W�H;{�H;'�H;]�H;��H;��H;��H;Z�H;'�H;|�H;V�H;{�H;B�H;��H;� I;I;;I;{I;.I;[&I;=2I;'@I;&PI;�bI;�wI;{�I;��I;��I;��I;��I;m�I;X�I;��I;�lI;�I;Y�H;�%H;4�G;^2G;��F;2�F;      ��?;��?;��@;]tA;��B;I�C;�BE;U�F;l�G;axH;�I;ϏI;v�I;��I;:�I;��I;�I;2�I;�I;iI;�TI;�BI;�3I;H'I;�I;yI;I;�I;� I;}�H;�H;n�H;`�H;��H;��H;*�H;��H;+�H;��H;��H;a�H;k�H;�H;~�H;� I;�I;I;I;�I;D'I;�3I;�BI;�TI;iI;�I;.�I;�I;��I;:�I;��I;v�I;ʏI;�I;axH;h�G;R�F;�BE;<�C;�B;_tA;�@;��?;      ��0;w51;�2;W�4;�07;3#:;�/=;� @;�B;�	E;��F;Q%H;�	I;T�I;��I;��I;��I;��I;c�I;��I;�mI;GWI;�DI;�4I;B'I;*I;�I;I;;I;- I;.�H;��H;|�H;��H;d�H;��H;m�H;��H;`�H;��H;~�H;��H;1�H;0 I;6I;{I;�I;.I;>'I;�4I;�DI;EWI;�mI;��I;g�I;��I;��I;��I;��I;Q�I;�	I;M%H;��F;�	E;�B;� @;�/=;*#:;�07;p�4;�2;`51;      C;�;"�;��;� ;�&;�\,;և2;98;�/=;�FA;orD;R�F;JH;^9I;0�I;l�I;Z�I;��I;��I;s�I;pI;FXI;�DI;�3I;X&I;I;�I;�
I;lI;��H;��H;��H;��H;<�H;J�H;�H;H�H;8�H;��H;��H;��H;��H;oI;|
I;�I;I;\&I;�3I;�DI;EXI;pI;s�I;��I;��I;S�I;o�I;.�I;^9I;JH;T�F;krD;�FA;�/=;98;Ӈ2;�\,;�&;� ;��; �;�;      <��:��:��:���:���:�P ;�e;�V;L#;e-;��5;�h<;RtA;W	E;�eG;:�H;1�I;�I;��I;�I;�I;��I;pI;KWI;�BI;=2I;�$I;vI;pI;B	I;xI;��H;��H;�H;Y�H;2�H;��H;3�H;W�H;�H;��H;��H;{I;D	I;lI;qI;�$I;A2I;�BI;NWI;pI;��I;�I;�I;��I;�I;/�I;8�H;�eG;V	E;RtA;�h<;��5;e-;L#;�V;�e;�P ;��:��:��:y�:      ��p� �,��!9�ų9��":��u:��:Z��:���:*R;_ ;��,;�6;S)>;�;C;��F;�lH;kkI;t�I;��I;��I;�I;r�I;�mI;~TI;"@I;�/I;%"I;YI;�I;�I;�I;u�H;u�H;��H;T�H;��H;V�H;��H;o�H;u�H;�I;�I;�I;VI;""I;�/I;#@I;yTI;�mI;n�I;�I;��I;��I;t�I;fkI;�lH;��F;�;C;R)>;�6;��,;` ;.R;���:`��:��:��u:�":�ų9�"9 �,�      p&�~!��4����氺�O��<T��t�9��u:�#�:�G�:D;,#;i71;?;;��A;��E;�$H;MVI;�I;��I;�I;��I;��I;iI;'PI;<I;�+I;I;�I;�I;�I;�I;6�H;��H;��H;�H;��H;��H;0�H;�I;�I;�I;�I;I;�+I;<I;&PI;	iI; �I;��I;�I;��I;�I;MVI;�$H;��E;��A;;;;g71;)#;D;�G�:�#�:��u:�t�9�<T�(�O��氺���4��!�      �kٻl�Ի�ǻ����V���n���+�8�Ժ�1�0�39\m:��:n�;
�;~\,;�8;��@;?]E;�
H;OVI;x�I;��I;��I;f�I;�I;�bI;`JI;)7I;�'I;�I;0I;�
I;9I;<I;k�H;��H;z�H;��H;d�H;8I;8I;�
I;2I;�I;�'I;%7I;`JI;�bI;��I;i�I;��I;��I;t�I;OVI;�
H;;]E;��@;ߍ8;{\,;
�;l�;��:Tm:�39 �1�8�Ժ��+��n��V������ǻh�Ի      6yY��|U�N�I�@�7��� ��!���Ի�᝻��T���#��u�9���:Sl�:�;�);17;/ @;<]E;�$H;ikI;�I;Z�I;��I;1�I;�wI;�ZI;�CI;}1I;N#I;)I;�I;.	I;uI;9I;k�H;��H;m�H;5I;pI;-	I;�I;)I;P#I;x1I;�CI;�ZI;�wI;&�I;��I;U�I;�I;dkI;�$H;:]E;, @;17;�);�;Ql�:���:�u�9�#����T��᝻��Ի "��� �@�7�P�I��|U�      ��ü^l��w����R��?ߓ�a�{��M��� �!��˼����B�갺 Ho���u:���:�R;3�';17;��@;��E;�lH;5�I;n�I;��I;�I;x�I;�lI;�QI;-<I;�+I;�I;�I;fI;�I;FI;/I;�I;/I;AI;�I;bI;�I;�I;�+I;)<I;QI;�lI;s�I;�I;��I;k�I;1�I;�lH;��E;��@;17;0�';�R;���:��u:@Ho�갺��B�̼�� �컋� ��M�`�{�@ߓ��R��x���]l��      �'��-$�_��X����
?ټw��:���pyY��k���Ի8��Y������$R:���:�R;�);ߍ8;��A;��F;;�H;0�I;��I;��I;��I;�I;�`I;�GI;�4I;�%I;KI;�I;�I;tI;I;EI;I;nI;�I;�I;FI;�%I;�4I;�GI;�`I;�I;��I;��I;��I;-�I;7�H;��F;��A;ݍ8;�);�R;���:�#R:����Y��:����Ի�k�pyY�;���	w��
?ټ���Y�_���-$�      Y+����c̀�-l��Q�%�2�B��������@����>�Y2��"V���1�x��$R:���:�;z\,;:;;�;C;�eG;`9I;��I;7�I;��I;C�I;�qI;�TI;c>I;<-I;3 I;{I;vI;�
I;I;I;I;�
I;rI;zI;- I;9-I;`>I;�TI;�qI;@�I;��I;0�I;��I;[9I;�eG;�;C;:;;v\,;�;���:�#R:���1�$V��Z2����>��@��������B�%�2��Q�.l�c̀���      j�ྲྀhܽp�н]y��^什P ��l��n<�M���>ټ��V|U��������1�p�����u:Sl�:	�;i71;Z)>;Z	E;JH;X�I;��I;��I;�I;ۃI;`bI;�HI;-5I;d&I;gI;tI;<I;"I;
I;&I;9I;qI;gI;_&I;(5I;�HI;]bI;ڃI;�I;��I;��I;X�I;JH;X	E;L)>;k71;�;Ol�:��u:�����1��������W|U����>ټM���n<�l�P ��_什^y��o�н�hܽ      ��4�f1��&������i�ང�������`��'���UR��D�]�~�� V���X�� Ho����:l�;-#; �6;XtA;Y�F;�	I;|�I;��I;p�I;�I;�pI;�SI;�=I;�,I;y I;�I;�I;FI;9I;FI;�I;�I;y I;�,I;�=I;�SI;�pI;�I;n�I;��I;t�I;�	I;X�F;StA;�6;.#;h�;���: Ho��X��"V��~��F�]�UR����'��`��������h��������&�f1�      �x���o��ń�IUo���O�*�-�{��hܽ[什Ҽx���2�tb��UR��V|U�X2��8��갺�u�9��:D;��,;�h<;lrD;U%H;ˏI;j�I;��I;�I;
�I;�^I;FI;V3I;�%I;�I;^I;hI;5I;iI;\I;�I;�%I;R3I;FI;�^I;�I;�I;��I;f�I;ÏI;S%H;lrD;�h<;��,;D;��:xu�9"갺:��Z2��W|U�UR��tb����2�Ҽx�[什�hܽ{�*�-���O�IUo�ń��o��      v���ྃ�Ѿ(����נ�ń�9�S��#�_O��|n��J̀���2���𛼂�>���Ի��B��#�@m:�G�:f ;��5;�FA;��F;�I;R�I;S�I;��I;q�I;pjI;�NI;:I;�*I;  I;�I;�I;LI;�I;�I;�I;�*I;:I;�NI;pjI;o�I;��I;Q�I;M�I;�I;��F;�FA;��5;X ;�G�:,m:�#���B� �Ի��>�������2�J̀�|n��_O���#�9�S�ń��נ�(�����Ѿ��      �3���/��X#��	��A��֌Ⱦ�f��HUo�]1�˰��|n��Ѽx��'��>ټ�@���k�̼�� ����39�#�:4R;e-;�/=;�	E;cxH;��I;�I;s�I;�I;vI;gWI;�@I;�/I;'$I;<I;�I;6I;�I;<I;#$I;�/I;�@I;dWI;vI;�I;s�I;�I;��I;_xH;�	E;�/=;e-;&R;�#�:��39"��μ���k��@���>ټ�'�Ҽx�|n��˰��^1�HUo��f��֌Ⱦ�A���	��X#���/�      ���T���T�v��RZ�[58�͂�p��d���foy�]1�_O��[什�`�M�����oyY�#�컗�T��1���u:��:M#;98;�B;p�G;�lI;�I;�I;2�I;x�I;�_I;GI;�4I;'(I;�I;�I;I;�I;�I;%(I;�4I;GI;�_I;t�I;/�I;�I;�I;�lI;j�G;�B;98;F#;���:��u:$�1���T�$��pyY����M���`�\什_O��]1�foy�d���p��͂�[58��RZ�T�v�T���      	Ŀ6g��&ﱿ���S����U��X#�t��d���IUo��#��hܽ����n<����;����� ��᝻@�Ժ�t�9n��:�V;҇2;� @;[�F;�I;��I;D�I;,�I;k�I;hI;MI;�9I;�+I;�"I;jI;�I;iI;�"I;�+I;�9I;MI;hI;l�I;+�I;E�I;��I;�I;W�F;� @;Ӈ2;�V;X��:�t�9F�Ժ�᝻�� �<�������n<�����hܽ�#�IUo�d���t���X#��U�S������&ﱿ6g��      ~x�P9�R��sؿnQ��e_��6�_��X#�p���f��9�S�{�����l�B�w���M���Ի��+��<T���:�e;�\,;�/=;�BE;T�H;x�I;��I;��I;��I;�oI;�RI;>I;^/I;~%I;�I;FI;�I;%I;]/I;>I;�RI;�oI;��I;��I;��I;{�I;Y�H;�BE;�/=;�\,;�e;��:�<T���+���Ի�M�	w��B�l�����{�9�S��f��p���X#�6�_�e_��nQ��sؿR��P9�      �X1���,�h���<��5g��e_���U�͂�֌Ⱦń�*�-�i��P ��&�2�
?ټa�{�"��n��O���u:�P ;�&;-#:;?�C;�%H;�I;$�I;��I;�I;bvI;�WI;�AI;{2I;(I;C"I;` I;C"I;(I;x2I;�AI;�WI;]vI;�I;��I;)�I;�I;�%H;?�C;0#:;�&;�P ;��u:�O��n�"�b�{�?ټ&�2�P ��i��*�-�ń�֌Ⱦ͂��U�e_��5g��<�h����,�      d��]]�5K��X1�Zf��nQ��S���[58��A���נ���O���_什�Q����@ߓ��� ��V��|氺�":ظ�: ;�07;�B;.�G;�{I;��I;��I;��I;;|I;7\I;LEI;5I;0*I;1$I;+"I;-$I;5*I;5I;LEI;5\I;8|I;��I;��I;��I;�{I;8�G;�B;�07; ;Ը�:�":�氺�V���� �@ߓ�����Q�_什����O��נ��A��[58�S���nQ���Zf��X1�5K��]]�      N������4z���V��X1��<�sؿ����RZ��	�(���IUo����^y��.l�Y��R��B�7�������ų9��:��;Y�4;ktA;\2G;�XI;��I;N�I;�I;��I;�_I;�GI;"7I;�+I;�%I;�#I;�%I;�+I;7I;�GI;�_I;�I;�I;M�I;��I;�XI;h2G;jtA;[�4;��;���:�ų9
�����B�7��R��Y�.l�^y�����IUo�(����	��RZ����tؿ�<��X1���V��4z�����      �o��f^���ē��4z�5K�h��R��&ﱿT�v��X#���Ѿń��&�p�нc̀�_��v���M�I��ǻ�4��"9��:6�;!�2;��@;��F;�:I;��I;��I;��I;y�I;KbI;�II;�8I;X-I;�&I;�$I;�&I;[-I;�8I;�II;KbI;u�I;��I;��I;��I;�:I;��F;��@;!�2;6�;��: "9�4��ǻL�I�v���_��c̀�p�н�&�ń���Ѿ�X#�T�v�&ﱿR��h��5K��4z��ē�f^��      q'���X��f^�������]]���,�P9�6g��T�����/����o��g1��hܽ���-$�_l���|U�f�Ի~!� �,�{�:�;�51;��?;5�F;A'I;b�I;�I;?�I;��I;�cI;>KI;x9I; .I;y'I;�%I;v'I; .I;x9I;@KI;�cI;��I;A�I;�I;d�I;C'I;C�F;��?;�51;�;u�: �,�~!�g�Ի�|U�_l���-$����hܽg1��o���ྚ�/�T���6g��P9���,��]]�����f^���X��      l����������Т��/�j��5���	� �ȿ&8����7�D�꾂S���7�
3�~L���)���Ƽ��\� �ݻ�+�`Uɸ��:x;��0;��?;I�F;�+I;��I;��I;ԽI;!�I;�hI;�NI;�<I;�0I;�)I;�'I;�)I;�0I;�<I;�NI;�hI;�I;ؽI;��I;��I;�+I;W�F;��?;��0;x;��:@Vɸ�+� �ݻ��\���Ƽ�)�~L��
3��7��S��D�꾨�7�&8�� �ȿ��	��5�/�j�Т����������      ��������B��^�����c�621�%X��ÿiڇ�r�3��s��7��|74�a�>ى���&�Nü'�X���ػ��%�@�J�ʃ�:�b;|�0;u�?;�F;�2I;��I;9�I;�I;H�I;PhI;�NI;0<I;w0I;a)I;�'I;\)I;z0I;.<I;�NI;ShI;C�I;�I;9�I;��I;�2I;�F;u�?;y�0;�b;���: �J���%���ػ'�X�Nü��&�>ى�a�|74��7���s�r�3�iڇ��ÿ%X�621���c�^����B�����      �����B����F��x�P���#�M�������x|��'�YD־�X��o�)�Խ�Ă�J<�9_��}-M���ʻ[��`&�8ȓ�:�;K2;v@;O�F;�FI;j�I;�I;*�I;��I;�fI;=MI;B;I;�/I;�(I;�&I;�(I;�/I;A;I;?MI;�fI;��I;-�I;�I;m�I;�FI;[�F;v@;K2;�;���: &�8X����ʻ}-M�8_��J<��Ă�Խo�)��X��YD־�'��x|����M�����#�x�P�F�����B��      Т��^���F���/]��5�N���,ݿ+8��qm_��K��t��W�s�#>����9�o��3��۩���:�nT�����(�9�f�:�<;�_4;hA;8G;{dI;�I;*�I;]�I;_�I;&dI;KI;�9I;H.I;�'I;�%I;�'I;K.I;�9I;KI;)dI;[�I;^�I;+�I;�I;ydI;8G;hA;�_4;�<;�f�:�'�9���pT����:��۩��3�9�o����#>�W�s��t���K�qm_�+8���,ݿN���5��/]�F��^���      /�j���c�x�P��5���s��I���hڇ�Fv<�(���p���_S��������
+T��� �+$���G#�ђ��p1���:���:6�;17;q�B;|�G;ćI;�I;e�I;ʮI;��I;�`I;IHI;�7I;a,I;&I; $I;&I;e,I;�7I;LHI;�`I;��I;ϮI;d�I;�I;ćI;��G;r�B;/7;3�;���:��:h1��ђ���G#�+$���� �
+T���������_S�p��(���Fv<�hڇ�I���s�����5�x�P���c�      �5�621���#�N��r���ÿ�ҕ�Z������̾�X���0�3�.W����5��zܼA��Z��c�s��U\�h�n:���:ج%;��9;��C;�.H;�I;�I;�I;��I;x{I;\I;�DI;�4I;(*I;$I;"I;$I;+*I;�4I;�DI;\I;u{I;��I;�I;�I;�I;�.H;��C;��9;۬%;���:P�n:�U\�a�s�Y��@���zܼ��5�.W��3��0��X����̾���Z��ҕ��ÿs��N����#�621�      ��	�%X�M����,ݿI����ҕ��d��'�@��#���x�W����k���2�o��G��*���Q���ػ�0���~���:z�;0,;b=;7BE;��H;��I;��I;E�I;�I;btI;�VI;�@I;�1I;�'I;�!I;�I;�!I;�'I;�1I;�@I;�VI;`tI;�I;F�I;��I;�I;��H;;BE;c=;1,;{�;��:0�~��0���ػ�Q��*���G�2�o�k������x�W�#���@�꾌'��d��ҕ�I����,ݿM���%X�       �ȿ�ÿ���+8��hڇ�Z��'�����l8��W�s�,�&�X�/i??��V�琼WG#�c7��~Tܺh�9W�:��;L2;P@;�F;�I;��I;u�I;P�I;D�I;�lI;�PI;[<I;�-I;�$I;%I;GI;%I;�$I;�-I;]<I;�PI;�lI;H�I;R�I;w�I;��I;�I;�F;O@;L2;��;	W�:��9xTܺc7��VG#�琼�V�i??�/X�,�&�W�s�l8�������'�Z�hڇ�+8������ÿ      &8��iڇ��x|�qm_�Fv<����?��l8��$6~�o74��l��{���7nc�4���^����\��9�JZ���=���n:F��:�#;�8;��B;t�G;�xI;p�I;��I;��I;݆I;8dI;xJI;�7I;*I;5!I;PI;�I;OI;8!I;*I;�7I;zJI;8dI;��I;��I;��I;p�I;�xI;y�G;��B;�8;�#;B��:��n:��=�JZ��9���\��^��4��7nc�{����l��o74�$6~�l8��?�꾎��Fv<�qm_��x|�iڇ�      ��7�r�3��'��K�'�����̾#���W�s�o74����!N��·|���)�9zܼ�Y��@ ����D����S9Љ�:!�; -;=;�E;��H;J�I;1�I;��I;��I;{I;^[I;�CI;X2I;&I;�I;-I;�I;+I;�I;&I;Y2I;�CI;c[I;!{I;��I;��I;1�I;K�I;�H;�E;=;-; �;���:T9@������? ��Y��8zܼ��)�·|�!N�����o74�W�s�#�����̾'����K��'�r�3�      D���s�YD־�t��p���X��x�W�,�&��l��!N���Ă�j�5�����|Q����A�E�ػ��G�"/�f:�a�:��;`�5;�9A;E�F;�*I;��I;��I;
�I;Z�I;/oI;gRI;�<I;-I;�!I;AI;I;�I;I;CI;�!I;-I;�<I;kRI;4oI;a�I;�I;��I;��I;�*I;H�F;�9A;g�5;��;b�:,f:"/���G�D�ػ��A�|Q������i�5��Ă�!N���l��,�&�x�W��X��p���t��YD־�s�      �S���7���X��W�s��_S��0����W�{���·|�i�5�j���ک�5�X� c �z��3����9
��:�;��,;�L<;SoD;.H;I;��I;��I;S�I;N�I;7cI;[II;�5I;�'I;GI;�I;�I;�I;�I;�I;JI;�'I;�5I;_II;=cI;Z�I;Z�I;��I;��I;ɛI;.H;\oD;�L<;�,;�;��:��9�3��x� c �4�X��ک�i��i�5�·|�{���Wར��~�0��_S�W�s��X���7��      �7�|74�o�)�#>����3�k���/7nc���)������ک�va��Q�T���N���ȸ ��:��;�#;r�6;hA;��F;�I;4�I;]�I;�I;v�I;�uI;mWI;r@I;
/I;c"I;I;�I;gI;[I;gI;�I;I;f"I;	/I;y@I;tWI;�uI;}�I;�I;]�I;=�I;�I;��F;hA;t�6;�#;��;��:��ȸN�T����Q�va��ک�������)�7nc�/k���3����#>�o�)�|74�      	3�`�Խ�������/W��1�o�h??�4��8zܼ|Q��4�X��Q��6�������Ϲx�n:�m�:>;��0;�>;.E;MSH;J�I;��I;^�I;?�I;U�I;�fI;"LI;�7I;e(I;I;�I;^I;I;>I;I;]I;�I;I;b(I;�7I;*LI;�fI;\�I;@�I;]�I;��I;M�I;TSH;6E;�>;��0;>;�m�:��n:��Ϲ����6���Q�3�X�|Q��8zܼ4��h??�1�o�.W���������Խ`�      }L��>ى��Ă�8�o�
+T���5��G��V��^���Y����A� c �V���������4�J:Yl�:�e;,;��:;5C;lG;�DI; �I;��I;��I;��I;�vI;�XI;BAI;�/I;"I;�I;�I;�I;�I;HI;�I;�I;�I;�I;"I;�/I;IAI;�XI;�vI;��I;��I;��I;�I;�DI;lG;5C;��:;#,;�e;gl�:4�J:������T���c ���A��Y���^���V��G���5�+T�8�o��Ă�>ى�      �)���&�I<��3��� ��zܼ�*��琼��\�@ �E�ػ{�!N���Ϲ0�J:pj�:f�;t�(;�e8;��A;�F;��H;�I;j�I;��I;��I;]�I;\eI;�KI;7I;�'I;�I;I;�I;aI;�I;'I;�I;^I;�I;I;�I;�'I;7I;�KI;ceI;_�I;��I;�I;m�I;!�I;��H;�F;��A;�e8;q�(;l�;tj�:<�J:��Ϲ N�x�C�ػ? ���\�琼�*���zܼ�� ��3�I<���&�      ��ƼNü9_���۩�*$��A���Q�TG#��9�����G��3����ȸ��n:al�:m�;�';�7;qv@;�E;vH;�I;��I;��I;8�I;��I;�qI;qUI;*?I;�-I;y I;I;kI;�I;CI;�I;I;�I;@I;�I;mI;I;� I;�-I;/?I;wUI;�qI;��I;A�I;��I;��I;��I;vH;'�E;vv@;�7;�';n�;gl�:��n:@�ȸ�3����G�����9�TG#��Q�@��+$���۩�:_��Nü      ��\�%�X�~-M���:��G#�X����ػ`7��JZ�6���"/���9��:�m�:�e;q�(;7;�@;!]E;}-H;1wI;t�I;��I;��I;��I;�|I;�^I;�FI;�3I;J%I;�I;�I;D
I;?I;"I;- I;r�H;* I;!I;?I;F
I;�I;�I;P%I;�3I;�FI;�^I;�|I;��I;��I;��I;z�I;5wI;�-H;&]E;�@;�7;q�(;�e;�m�:��:��9�!/�6���BZ�`7����ػX���G#���:�|-M�%�X�      �ݻ��ػ��ʻnT��Ғ��S�s���0�jTܺ��=�@T9@f:��:��;>;",;�e8;qv@;(]E;/H;�aI;�I;��I;=�I;��I;Q�I;�fI;�MI;�9I;�)I;iI;mI;�I;2I;I;G�H;~�H;��H;}�H;E�H;I;3I;�I;rI;lI;�)I;�9I;�MI;�fI;[�I;��I;:�I;��I;�I;bI;1H;#]E;vv@;�e8;#,;>;��;��:Hf:0T9��=�jTܺ��0�Z�s�ђ��rT����ʻ��ػ      �+���%�T�� ����1���U\���~�P�9��n:ډ�:
b�:�;�#;��0;��:;��A;!�E;�-H; bI;��I;d�I;y�I;�I;��I;�mI;�SI;?I;2.I;� I;VI;�I;^I;uI;��H;r�H;�H;u�H;�H;o�H;��H;zI;]I;�I;VI;� I;9.I;?I;�SI;�mI;��I;�I;}�I;k�I;��I;bI;�-H;#�E;��A;��:;��0;�#;�;b�:މ�:��n:��9 �~��U\�t1�����b����%�      @Qɸ��J��#�8�'�9Ч:X�n:��:W�:@��: �;��;��,;p�6;�>;
5C;�F;vH;9wI;�I;d�I;3�I;��I;U�I;�rI;�XI;2CI;�1I;'$I;�I;�I;�I;EI;>�H;1�H;��H;��H;u�H;��H;��H;.�H;>�H;AI;�I;�I;�I;*$I;�1I;2CI;�XI;�rI;R�I;ŸI;:�I;e�I;�I;7wI;vH;�F;5C;�>;r�6;��,;��;!�;:��:	W�:��:H�n:��:�'�9�$�8 �J�      ��:؃�:ړ�:�f�:���:���:x�;��;�#;-;f�5;�L<;hA;3E;lG;��H;��I;w�I;��I;}�I;øI;�I;�tI;u[I;FFI;�4I;�&I;2I;�I;O
I;hI;��H;�H;v�H;��H;��H;g�H;��H;��H;v�H;�H;��H;nI;Q
I;�I;4I;�&I;�4I;KFI;u[I;�tI;�I;ƸI;}�I;��I;w�I;��I;��H;lG;0E;hA;�L<;i�5; -;�#;��;��;���:ͱ�:�f�:ȓ�:ă�:      *x;�b;�;�<;%�;�%;;,;+L2;�8;=;�9A;`oD;��F;\SH;�DI;$�I;��I;��I;=�I;�I;T�I;�tI;]\I;�GI;|6I;�(I;�I;=I;�I;MI;B I;r�H;M�H;�H;��H;��H;��H;��H;��H;�H;M�H;r�H;H I;MI;�I;BI;�I;�(I;�6I;�GI;X\I;�tI;V�I;�I;?�I;��I;��I;$�I;�DI;XSH;��F;_oD;�9A;=;�8;'L2;8,;۬%;6�;�<;�;�b;      ��0;��0;K2;�_4;"7;��9;[=;O@;��B;�E;A�F;.H;�I;K�I;��I;k�I;��I;��I;��I;��I;rI;m[I;�GI;7I;m)I;�I;PI;�I;0I;� I;��H;��H;��H;��H;��H;
�H;��H;�H;��H;��H;��H;��H;��H;� I;/I;�I;OI;�I;t)I;7I;�GI;q[I;�rI;��I;��I;��I;��I;j�I; �I;G�I;�I;.H;G�F;�E;��B;S@;Y=;��9;*7;�_4;K2;��0;      Ĥ?;q�?;v@;hA;`�B;��C;<BE;�F;u�G;�H;�*I;̛I;6�I;��I;��I;�I;B�I;��I;\�I;�mI;�XI;GFI;�6I;x)I;YI;�I;4I;�I;vI;2�H;��H;��H;��H;*�H;�H;o�H;2�H;i�H;�H;,�H;��H;��H;��H;5�H;qI;�I;1I;�I;]I;v)I;�6I;MFI;�XI;�mI;_�I;��I;E�I;�I;��I;��I;8�I;ΛI;�*I;�H;t�G;ބF;>BE;��C;n�B;hA;v@;q�?;      E�F;�F;E�F;8G;n�G;�.H;��H;I;�xI;S�I;��I;��I;b�I;h�I;��I;��I;��I;�|I;�fI;�SI;4CI;�4I;�(I;�I;�I;qI;-I;�I;o�H;��H;��H;��H;��H;��H;��H;��H;��H;��H;��H;��H;��H;��H;��H;��H;m�H;�I;*I;wI;�I;�I;�(I;�4I;4CI;�SI;�fI;�|I;��I;��I;��I;b�I;a�I;��I;��I;R�I;�xI; I;��H;�.H;��G;8G;G�F;�F;      �+I;�2I;�FI;ydI;��I;�I;��I;��I;p�I;1�I;��I;��I;�I;B�I;��I;_�I;�qI;�^I;�MI;?I;�1I;�&I;�I;TI;1I;,I;�I;��H;�H;��H;��H;��H;8�H;�H;,�H;��H;��H;��H;*�H;�H;9�H;��H;��H;��H;�H;��H;�I;0I;8I;QI;�I;�&I;�1I;?I;�MI;�^I;�qI;b�I;��I;=�I;�I;��I;��I;/�I;l�I;��I;~�I;�I;ʇI;pdI;�FI;�2I;      ��I;��I;d�I;�I;�I;�I;��I;u�I;��I;��I;�I;[�I;v�I;^�I;�vI;^eI;pUI;�FI;�9I;3.I;,$I;-I;=I;�I;�I;�I;��H;0�H;�H;��H;~�H;��H;��H;��H;"�H;��H;��H;��H;"�H;��H;��H;��H;��H;��H;�H;0�H;��H;�I;�I;�I;>I;/I;*$I;0.I;�9I;�FI;qUI;aeI;�vI;\�I;x�I;[�I;�I;��I;��I;p�I;��I;�I;�I;
�I;d�I;��I;      ��I;+�I;��I;8�I;W�I;�I;H�I;V�I;��I;��I;_�I;Z�I;�uI;�fI;�XI;�KI;2?I;�3I;�)I;� I;�I;�I;�I;.I;oI;h�H;�H;�H;��H;|�H;��H;��H;N�H;��H;;�H;��H;��H;��H;9�H;��H;Q�H;��H;��H;{�H;��H;�H;�H;f�H;qI;)I;�I;�I;�I;� I;�)I;�3I;0?I;�KI;�XI;�fI;�uI;X�I;c�I;��I;��I;U�I;I�I;��I;a�I;;�I;��I;'�I;      սI;�I;4�I;Y�I;ŮI;��I;�I;K�I;��I;"{I;7oI;GcI;tWI;-LI;IAI;7I;�-I;G%I;fI;VI;�I;K
I;JI;� I;5�H;��H;��H;��H;��H;��H;��H;F�H;\�H;��H;"�H;��H;��H;��H; �H;��H;\�H;F�H;��H;��H;|�H;��H;��H;��H;8�H;� I;LI;M
I;�I;TI;fI;F%I;�-I;7I;GAI;)LI;qWI;AcI;6oI;#{I;݆I;D�I;�I;��I;ŮI;a�I;2�I;�I;      �I;]�I;�I;f�I;��I;v{I;`tI;�lI;<dI;j[I;qRI;jII;|@I;�7I;�/I;�'I;� I;�I;tI;I;�I;iI;B I;��H;��H;��H;��H;��H;��H;��H;7�H;5�H;��H;��H;k�H;D�H;0�H;B�H;j�H;��H;��H;5�H;9�H;��H;��H;�H;��H;��H;��H;��H;F I;kI;�I;�I;rI;�I;� I;�'I;�/I;�7I;z@I;fII;nRI;h[I;:dI;�lI;htI;o{I;��I;g�I;��I;]�I;      �hI;ZhI;�fI;dI;|`I;�[I;�VI;�PI;JI;�CI;�<I;�5I;/I;l(I;"I;�I;I;�I;I;cI;NI;��H;p�H;��H;��H;��H;��H;�H;��H;H�H;2�H;��H;��H;0�H;��H;��H;��H;��H;��H;3�H;��H;~�H;1�H;D�H;��H;��H;��H;��H;��H;��H;s�H;��H;GI;^I; I;�I;I;�I;"I;i(I;/I;�5I;�<I;�CI;|JI;�PI;�VI; \I;�`I;%dI;�fI;[hI;      �NI;�NI;<MI;KI;FHI;�DI;�@I;Z<I;7I;U2I;-I;�'I;g"I;I;�I;I;rI;G
I;:I;{I;H�H;�H;I�H;��H;��H;��H;6�H;��H;V�H;_�H;��H;��H;�H;��H;w�H;3�H;.�H;3�H;u�H;��H;�H;��H;��H;W�H;Q�H;��H;5�H;��H;��H;��H;L�H;�H;B�H;wI;9I;F
I;tI;I;�I;I;d"I;�'I;!-I;V2I;�7I;T<I;�@I;�DI;IHI;KI;IMI;�NI;      �<I;.<I;;;I;�9I;�7I;�4I;�1I;.I;*I;&I;�!I;UI;I;�I;�I;�I;�I;?I;I; �H;7�H;t�H;��H;��H;%�H;��H;�H;��H;��H;��H;��H;2�H;��H;O�H;�H;��H;��H;��H;�H;O�H;��H;2�H;��H;��H;��H;��H;�H;��H;(�H;��H;�H;s�H;0�H;��H;I;@I;�I;�I;�I;�I;I;QI;�!I; &I;*I;�-I;�1I;�4I;�7I;�9I;E;I;;<I;      �0I;�0I;�/I;M.I;k,I;$*I;�'I;�$I;<!I;�I;NI;�I;	I;jI;�I;gI;JI;"I;K�H;s�H;��H;��H;��H;��H;�H;}�H;%�H;!�H;?�H;%�H;e�H;��H;w�H;�H;��H;��H;��H;��H;��H;�H;w�H;��H;c�H;�H;6�H;�H;%�H;|�H;�H;��H;��H;��H;��H;n�H;H�H;$I;JI;hI;�I;jI;	I;�I;QI;�I;<!I;�$I;�'I;%*I;e,I;U.I;�/I;�0I;      �)I;i)I;�(I;�'I;�%I;$I;�!I;,I;OI;6I;	I;�I;kI;%I;	I;�I;�I;* I;��H;�H;��H;��H;��H;��H;f�H;��H;��H;��H;��H;��H;B�H;��H;7�H;��H;��H;f�H;f�H;j�H;��H;��H;7�H;��H;@�H;��H;��H;��H;��H;��H;f�H;��H;��H;��H;��H;	�H;��H;- I;�I;�I;	I;'I;kI;�I;I;6I;PI;(I;�!I;$I;�%I;�'I;�(I;v)I;      �'I;�'I;�&I;�%I;�#I;"I;�I;NI;�I;�I;�I;�I;bI;II;TI;-I;(I;v�H;��H;{�H;~�H;g�H;��H;��H;.�H;��H;��H;��H;��H;��H;*�H;��H;.�H;��H;��H;c�H;I�H;e�H;��H;��H;/�H;��H;)�H;��H;��H;��H;��H;��H;.�H;��H;��H;f�H;v�H;w�H;��H;v�H;'I;/I;TI;KI;bI;�I;�I;�I;�I;MI;�I;"I;�#I;�%I;�&I;�'I;      �)I;j)I;�(I;�'I;�%I;$I;�!I;*I;OI;6I;	I;�I;mI;'I;	I;�I;�I;* I;��H;�H;��H;��H;��H;��H;f�H;��H;��H;��H;��H;��H;B�H;��H;9�H;��H;��H;f�H;f�H;j�H;��H;��H;7�H;��H;@�H;��H;��H;��H;��H;��H;f�H;��H;��H;��H;��H;
�H;��H;- I;�I;�I;	I;&I;kI;�I;I;4I;PI;*I;�!I;$I;�%I;�'I;�(I;q)I;      �0I;�0I;�/I;H.I;k,I;$*I;�'I;�$I;<!I;�I;NI;�I;	I;hI;�I;eI;II;$I;K�H;u�H;��H;��H;��H;��H;�H;|�H;%�H;!�H;=�H;"�H;d�H;��H;x�H;�H;��H;��H;��H;��H;��H;�H;w�H;��H;c�H;�H;8�H;�H;#�H;}�H;�H;��H;��H;��H;��H;n�H;H�H;$I;LI;hI;�I;jI;	I;�I;QI;�I;<!I;�$I;�'I;"*I;i,I;R.I;�/I;�0I;      �<I;0<I;:;I;�9I;�7I;�4I;�1I;.I;*I;&I;�!I;SI;I;�I;�I;�I;�I;BI;I; �H;7�H;t�H;��H;��H;(�H;��H;�H;��H;��H;��H;��H;0�H;��H;N�H;�H;��H;��H;��H;�H;N�H;��H;2�H;��H;��H;��H;��H;�H;��H;&�H;��H;�H;t�H;-�H;��H;I;@I;�I;�I;�I;�I;I;QI;�!I;&I;*I;.I;�1I;�4I;�7I;�9I;B;I;3<I;      �NI;�NI;?MI;KI;CHI;�DI;�@I;`<I;�7I;U2I;-I;�'I;d"I;I;�I;I;rI;F
I;7I;{I;I�H;�H;G�H;��H;��H;��H;4�H;��H;V�H;^�H;��H;��H;�H;��H;x�H;3�H;.�H;3�H;w�H;��H;�H;��H;��H;W�H;N�H;��H;4�H;��H;��H;��H;M�H;�H;>�H;xI;7I;D
I;qI;I;�I;I;g"I;�'I; -I;U2I;�7I;[<I;�@I;�DI;HHI;#KI;PMI;�NI;      �hI;]hI;�fI;dI;}`I;\I;�VI;�PI;|JI;�CI;�<I;�5I;/I;i(I;"I;�I;I;�I;�I;aI;OI;��H;o�H;��H;��H;��H;��H;�H;��H;F�H;/�H;}�H;��H;/�H;��H;��H;��H;��H;��H;0�H;��H;~�H;.�H;C�H;��H;��H;��H;��H;��H;��H;u�H;��H;DI;^I;�I;�I;I;�I;"I;k(I;/I;�5I;�<I;�CI;~JI;�PI;�VI;�[I;}`I;)dI;�fI;XhI;      �I;^�I;�I;_�I;��I;v{I;btI;�lI;;dI;g[I;mRI;iII;y@I;�7I;�/I;�'I;� I;�I;rI;�I;�I;kI;B I;��H;��H;��H;��H;��H;��H;��H;6�H;5�H;��H;��H;n�H;B�H;0�H;E�H;h�H;��H;��H;5�H;5�H;��H;��H;~�H;��H;��H;��H;��H;E I;iI;�I;�I;tI;�I;� I;�'I;�/I;�7I;z@I;fII;pRI;e[I;<dI;�lI;htI;t{I;��I;j�I;�I;`�I;      ۽I;�I;.�I;a�I;��I;��I;�I;N�I;��I;#{I;2oI;DcI;qWI;*LI;JAI;7I;�-I;I%I;fI;VI;�I;N
I;II;� I;8�H;��H;��H;��H;��H;��H;��H;F�H;X�H;��H; �H;��H;��H;��H;�H;��H;[�H;F�H;��H;��H;{�H;��H;��H;��H;4�H;� I;MI;K
I;�I;TI;iI;F%I;�-I;7I;JAI;*LI;qWI;AcI;3oI;%{I;܆I;J�I;�I;�I;îI;i�I;6�I;�I;      ��I;,�I;�I;.�I;H�I;�I;E�I;V�I;��I;��I;a�I;Z�I;�uI;�fI;�XI;�KI;0?I;�3I;�)I;� I;�I;�I;�I;.I;qI;c�H;�H;�H;��H;z�H;��H;��H;N�H;��H;9�H;��H;��H;��H;6�H;��H;N�H;��H;��H;x�H;��H;�H;�H;f�H;mI;%I;�I;�I;�I;� I;�)I;�3I;0?I;�KI;�XI;�fI;�uI;W�I;b�I;��I;��I;U�I;L�I;�I;W�I;1�I;�I;'�I;      ��I;��I;Y�I;�I;�I;�I;��I;w�I;��I;��I;�I;\�I;x�I;\�I;�vI;_eI;qUI;�FI;�9I;0.I;-$I;0I;=I;�I;�I;�I;��H;0�H;!�H;��H;�H;�H;��H;��H;"�H;��H;��H;��H;!�H;��H;��H;��H;~�H;��H;�H;,�H;��H;�I;�I;~I;@I;-I;'$I;0.I;�9I;�FI;tUI;aeI;�vI;[�I;x�I;Z�I;�I;��I;��I;p�I;��I;�I;�I;
�I;c�I;��I;      �+I;�2I;�FI;�dI;��I;�I;��I;��I;p�I;1�I;��I;��I;�I;@�I;��I;`�I;�qI;�^I;�MI;?I;�1I;�&I;�I;WI;6I;*I;�I;��H;�H;��H;��H;��H;6�H;�H;-�H;��H;��H;��H;*�H;�H;8�H;��H;��H;��H;�H;��H;�I;/I;2I;PI;�I;�&I;�1I;?I;NI;�^I;�qI;c�I;��I;@�I;�I;��I;��I;/�I;l�I;��I;��I;�I;ȇI;�dI;�FI;�2I;      ?�F;�F;S�F;8G;v�G;�.H;��H;I;�xI;R�I;��I;��I;b�I;e�I;��I;��I;��I;�|I;�fI;�SI;9CI;�4I;�(I;�I;�I;pI;-I;�I;s�H;��H;��H;��H;��H;��H;��H;��H;��H;��H;��H;��H;��H;��H;��H;��H;i�H;�I;,I;tI;�I;�I;�(I;�4I;3CI;�SI; gI;�|I;��I;��I;��I;d�I;a�I;��I;��I;R�I;�xI;�I;��H;�.H;~�G;8G;9�F;�F;      Ĥ?;q�?;	v@;hA;a�B;��C;<BE;߄F;x�G;�H;�*I;ϛI;6�I;��I;��I;�I;D�I;âI;_�I;�mI;�XI;KFI;�6I;z)I;]I;�I;2I;�I;wI;2�H;��H;��H;��H;*�H;�H;l�H;2�H;l�H;�H;)�H;��H;��H;��H;2�H;mI;�I;2I;�I;YI;t)I;�6I;JFI;�XI;�mI;b�I;��I;E�I;�I;��I;��I;8�I;˛I;�*I;�H;r�G;ބF;?BE;��C;l�B;hA;
v@;q�?;      f�0;o�0;K2;�_4;7;��9;X=;P@;��B;�E;D�F;.H;�I;H�I;�I;m�I;��I;��I;��I;��I;�rI;q[I;�GI;!7I;t)I;�I;PI;�I;2I;� I;��H;��H;��H;��H;��H;�H;��H;	�H;��H;��H;��H;��H;��H;� I;/I;�I;PI;�I;p)I;7I;�GI;n[I;�rI;��I;��I;��I;��I;m�I; �I;G�I;�I;.H;E�F;�E;��B;J@;\=;��9;/7;�_4;K2;Z�0;      &x;�b;~;�<;#�;ެ%;4,;'L2;�8;=;�9A;_oD;��F;ZSH;�DI;%�I;��I;��I;?�I;�I;X�I;�tI;[\I;�GI;�6I;�(I;�I;AI;�I;JI;E I;v�H;L�H;�H;��H;��H;��H;��H;��H;�H;L�H;s�H;H I;NI;�I;=I;�I;�(I;~6I;�GI;Z\I;�tI;U�I;�I;A�I;��I;��I;%�I;�DI;WSH;��F;]oD;�9A;=;�8;$L2;4,;߬%;"�;�<;};�b;      ��:؃�:̓�:�f�:���:���:��;��;�#; -;f�5;�L<;hA;0E;lG;��H;��I;x�I;��I;��I;ɸI;�I;�tI;v[I;NFI;�4I;�&I;3I;�I;O
I;kI;��H;�H;v�H;��H;��H;i�H;��H;��H;t�H;�H;��H;nI;Q
I;�I;2I;�&I;�4I;GFI;v[I;�tI;�I;øI;~�I;��I;u�I;��I;��H;lG;2E;hA;�L<;i�5; -;�#;��;z�;���:Ǳ�:�f�:Ɠ�:���:       Sɸ��J�`%�8�'�9̧:x�n:��:W�:F��:�;��; �,;r�6;�>;5C;�F;vH;8wI;�I;g�I;7�I;ŸI;U�I;�rI;�XI;0CI;�1I;*$I;�I;�I;�I;HI;>�H;3�H;��H;��H;v�H;��H;��H;-�H;@�H;EI;�I;�I;�I;'$I;�1I;0CI;�XI;�rI;Q�I;��I;6�I;h�I;�I;4wI;vH;�F;5C;�>;r�6;��,;��; �;:��:W�:��:\�n:�:�'�9�&�8��J�      {+���%�X�������1���U\� �~���9��n:މ�:b�:�;�#;��0;��:;��A;$�E;�-H;bI;��I;k�I;~�I;�I;��I;�mI;�SI;?I;5.I;� I;TI;�I;`I;zI;��H;s�H;�H;w�H;�H;o�H;��H;xI;]I;�I;TI;� I;2.I;?I;�SI;�mI;��I;�I;z�I;h�I;��I;bI;�-H;$�E;��A;��:;��0;�#;�;b�:؉�:��n:��9 �~��U\�v1�����[����%�      �ݻ��ػ��ʻlT��Ғ��R�s���0�jTܺ��=�0T9@f:��:��;>;',;�e8;sv@;(]E;0H;bI;�I;��I;?�I;��I;[�I;�fI;�MI;�9I;�)I;iI;oI;�I;3I;	I;I�H;~�H;��H;�H;G�H;I;5I;�I;qI;iI;�)I;�9I;�MI;�fI;R�I;��I;;�I;��I;�I;bI;/H;#]E;uv@;�e8;#,;>;��;��:@f:0T9��=�fTܺ��0�U�s�Ԓ��lT����ʻ��ػ      ��\�#�X�~-M���:��G#�U����ػ\7��CZ�6����!/���9��:�m�:�e;u�(;�7;�@;%]E;�-H;4wI;z�I;��I;��I;��I;�|I;�^I;�FI;�3I;J%I;�I;�I;F
I;BI;"I;- I;t�H;. I;I;?I;F
I;�I;�I;L%I;�3I;�FI;�^I;�|I;��I;��I;��I;u�I;1wI;�-H;#]E;�@;�7;q�(;�e;�m�:��:��9"/�:���FZ�^7����ػX���G#���:��-M�#�X�      ��ƼNü9_���۩�*$��@���Q�TG#��9�����G��3��`�ȸ��n:il�:q�;�';�7;sv@;$�E;vH;��I;��I;��I;B�I;��I;�qI;sUI;3?I;�-I;} I;I;nI;�I;DI;�I;!I;�I;?I;�I;jI;I;} I;�-I;-?I;pUI;�qI;�I;:�I;��I;��I;��I;vH;$�E;rv@;�7;�';m�;el�:��n:��ȸ�3����G�����9�TG#��Q�?��+$���۩�:_��Nü      �)���&�I<��3��� ��zܼ�*��琼��\�@ �C�ػx�N���Ϲ@�J:xj�:i�;u�(;�e8;��A;�F;��H;%�I;m�I;�I;��I;]�I;_eI;�KI;7I;�'I;�I;I;�I;dI;�I;'I;�I;^I;�I;I;�I;�'I;7I;�KI;\eI;[�I;��I;��I;k�I;"�I;��H;
�F;��A;�e8;q�(;j�;nj�:0�J:��Ϲ!N�{�E�ػ@ ���\�琼�*���zܼ�� ��3�J<���&�      }L��>ى��Ă�8�o�
+T���5��G��V��^���Y����A� c �T���������H�J:el�:�e;#,;��:;5C;lG;�DI;�I;��I;��I;��I;�vI;�XI;FAI;�/I;"I;�I;�I;�I;�I;HI;�I;�I;�I;�I;"I;�/I;BAI;�XI;�vI;��I;��I;��I;�I;�DI;lG;5C;��:;,;�e;el�:0�J:������V��� c ���A��Y���^���V��G���5�+T�9�o��Ă�>ى�      	3�`�Խ�������.W��1�o�h??�4��8zܼ|Q��3�X��Q��6�������Ϲ��n:�m�:>;��0;�>;5E;TSH;N�I;��I;b�I;@�I;Z�I;�fI;&LI;�7I;e(I;I;�I;`I;I;>I; I;\I;�I;I;a(I;�7I;%LI;�fI;X�I;=�I;]�I;��I;N�I;XSH;2E;�>;��0;>;�m�:��n:��Ϲ����6���Q�4�X�|Q��8zܼ4��h??�2�o�.W���������Խ`�      �7�|74�o�)�#>����3�k���/7nc���)������ک�va��Q�R���N�@�ȸ"��:��;�#;z�6;hA;��F;�I;=�I;`�I;�I;y�I;�uI;qWI;v@I;/I;d"I;I;�I;gI;[I;gI;�I;I;d"I;/I;s@I;nWI;�uI;x�I;�I;[�I;5�I;�I;��F;hA;l�6;�#;��;��:`�ȸN�T����Q�wa��ک�������)�7nc�/k���3����#>�o�)�|74�      �S���7���X��W�s��_S��0����W�{���·|�i�5�i���ک�4�X� c �x��3����9��:�;�,;�L<;\oD;.H;˛I;��I;��I;U�I;W�I;9cI;aII;�5I;�'I;MI;�I;�I;�I;�I;�I;II;�'I;�5I;^II;9cI;W�I;T�I;��I;��I;I;.H;]oD;�L<;��,;�;
��:��9�3��{� c �5�X��ک�i��i�5�·|�{���Wར��~�0��_S�W�s��X���7��      D���s�YD־�t��p���X��x�W�,�&��l��!N���Ă�i�5�����|Q����A�D�ػ��G�"/�,f:b�:��;g�5;�9A;J�F;�*I;��I;��I;�I;b�I;2oI;kRI;�<I;-I;�!I;CI;I;�I;I;CI;�!I;-I;�<I;iRI;0oI;a�I;�I;��I;��I;�*I;J�F;�9A;b�5;��;b�:f: "/���G�E�ػ��A�|Q������i�5��Ă�!N���l��,�&�y�W��X��p���t��YD־�s�      ��7�r�3��'��K�'�����̾#���W�s�o74����!N��·|���)�8zܼ�Y��> ����>���0T9���:(�;-;=;�E;�H;N�I;1�I;��I;��I;!{I;d[I;�CI;Y2I;&I;�I;-I;�I;-I;�I;&I;Y2I;�CI;c[I;{I;��I;��I;/�I;K�I;��H;�E;=;-;�;މ�:�S9F������@ ��Y��8zܼ��)�·|�!N�����o74�W�s�#�����̾'����K��'�r�3�      &8��iڇ��x|�qm_�Fv<����?��l8��$6~�o74��l��{���7nc�4���^����\��9�LZ���=���n:T��:�#;�8;��B;{�G;�xI;r�I;��I;��I;߆I;<dI;xJI;�7I;*I;5!I;PI;�I;OI;6!I;*I;�7I;xJI;7dI;܆I;��I;��I;o�I;�xI;w�G;��B;�8;�#;:��:��n:��=�MZ��9���\��^��4��7nc�{����l��o74�$6~�l8��?�꾎��Fv<�qm_��x|�iڇ�       �ȿ�ÿ���+8��hڇ�Z��'�����l8��W�s�,�&�X�/i??��V�琼VG#�d7��rTܺ��9W�:��;!L2;V@;�F;�I;��I;u�I;S�I;D�I;�lI;�PI;]<I;�-I;�$I;#I;GI;#I;�$I;�-I;]<I;�PI;�lI;F�I;S�I;u�I;��I;�I;�F;S@;!L2;��;W�:��9~Tܺd7��VG#�琼�V�i??�/X�,�&�W�s�l8�������'�Z�hڇ�+8������ÿ      ��	�%X�M����,ݿI����ҕ��d��'�@��#���x�W����k���2�o��G��*���Q���ػ �0� �~���:~�;3,;f=;<BE;��H;��I;��I;I�I;�I;dtI;�VI;�@I;�1I;�'I;�!I;�I;�!I;�'I;�1I;�@I;�VI;atI;�I;H�I;��I;��I;��H;9BE;f=;5,;z�;��: �~��0���ػ�Q��*���G�2�o�k������x�W�#���@�꾌'��d��ҕ�I����,ݿM���%X�      �5�621���#�N��r���ÿ�ҕ�Z������̾�X���0�3�.W����5��zܼ@��Z��_�s��U\�t�n:���:۬%;��9;��C;�.H;�I;�I;�I;��I;{{I;\I;�DI;�4I;)*I;$I;"I;$I;+*I;�4I;�DI;\I;v{I;��I;�I;�I;�I;�.H;��C;��9;ެ%;���:X�n:�U\�d�s�Z��A���zܼ��5�.W��3��0��X����̾���Z��ҕ��ÿr��N����#�621�      /�j���c�x�P��5���s��I���hڇ�Fv<�(���p���_S��������
+T��� �+$���G#�В��h1���:���:4�;07;s�B;z�G;I;�I;e�I;ʮI;��I;�`I;IHI;�7I;`,I;&I;$I;	&I;d,I;�7I;LHI;�`I;��I;ͮI;e�I;�I;ćI;��G;r�B;37;4�;���:�:l1��Ғ���G#�,$���� �+T���������_S�p��(���Fv<�hڇ�I���s�����5�x�P���c�      Т��^���F���/]��5�N���,ݿ+8��qm_��K��t��W�s�#>����9�o��3��۩���:�nT�����0(�9�f�:�<;�_4;hA;
8G;xdI;�I;+�I;Z�I;b�I;&dI;KI;�9I;J.I;�'I;�%I;�'I;K.I;�9I;KI;)dI;]�I;^�I;*�I;�I;ydI;8G;hA;�_4;�<;�f�:�'�9���pT����:��۩��3�9�o����#>�W�s��t���K�qm_�+8���,ݿN���5��/]�F��^���      �����B����F��x�P���#�M�������x|��'�YD־�X��o�)�Խ�Ă�J<�8_��}-M���ʻX���&�8ȓ�:�;K2;v@;N�F;�FI;j�I;�I;*�I;�I;�fI;=MI;B;I;�/I;�(I;�&I;�(I;�/I;B;I;?MI;�fI;��I;+�I;�I;n�I;�FI;[�F;v@;K2;�;���:�%�8X����ʻ~-M�8_��J<��Ă�Խo�)��X��YD־�'��x|����M�����#�x�P�F�����B��      ��������B��^�����c�621�%X��ÿiڇ�r�3��s��7��|74�a�>ى���&�Nü'�X���ػ��%���J�ʃ�:�b;|�0;u�?;�F;�2I;��I;9�I;�I;H�I;QhI;�NI;0<I;y0I;_)I;�'I;\)I;y0I;0<I;�NI;ThI;C�I;�I;9�I;��I;�2I;�F;s�?;z�0;�b;���: �J���%���ػ(�X�Nü��&�>ى�a�|74��7���s�r�3�iڇ��ÿ%X�621���c�^����B�����      D(��r'���o��N�d��X1�~x�	Ŀ����3�x���x����4�l��Z+���'���ü:yY��kٻp&� �p�J��:9;��0;��?;F;k I; �I;��I;/�I;k�I;OdI;�KI;�9I;n.I;�'I;�%I;�'I;n.I;�9I;�KI;PdI;g�I;0�I;��I;�I;h I;̀F;��?;��0;4;B��:��p�p&��kٻ;yY���ü�'�Z+��l�ཽ�4��x��x���3����	Ŀ~x��X1�d�N��o��r'��      q'���X��e^�������]]���,�P9�6g��U�����/����o��g1��hܽ���-$�_l���|U�g�Ի�!� �,�y�:�;�51;��?;7�F;A'I;d�I;�I;@�I;��I;�cI;AKI;{9I; .I;}'I;�%I;y'I;".I;z9I;BKI;�cI;��I;C�I;�I;d�I;@'I;B�F;��?;�51;�;o�: �,��!�h�Ի�|U�_l���-$����hܽg1��o���ྙ�/�U���6g��P9���,��]]�����e^���X��      �o��e^���ē��4z�5K�h��R��'ﱿU�v��X#���Ѿń��&�o�нc̀�_��v���J�I��ǻ�4�`"9��:6�;!�2;��@;��F;�:I;��I;��I;��I;w�I;NbI;�II;�8I;\-I;�&I;�$I;�&I;\-I;�8I;JI;NbI;r�I;��I;��I;��I;�:I;��F;��@;�2;2�;��:"9�4��ǻL�I�v���_��c̀�o�н�&�ń���Ѿ�X#�U�v�'ﱿR��h��5K��4z��ē�e^��      N������4z���V��X1��<�uؿ����RZ��	�(���HUo����^y��-l�Y��R��D�7�������ų9��:��;[�4;ktA;^2G;�XI;��I;M�I;�I;��I;�_I;�GI;%7I;�+I;�%I;�#I;�%I;�+I;"7I;�GI;�_I;�I;�I;M�I;��I;�XI;h2G;jtA;X�4;��;���:�ų9�����C�7��R��Y�-l�^y�����HUo�(����	��RZ����uؿ�<��X1���V��4z�����      d��]]�5K��X1�Zf��nQ��T���[58��A���נ���O���`什�Q����@ߓ��� ��V���氺��":Ը�: ;�07;�B;0�G;�{I;��I;��I;��I;:|I;:\I;MEI;5I;6*I;3$I;,"I;0$I;7*I;5I;NEI;8\I;7|I;��I;��I;��I;�{I;8�G;�B;�07; ;Ҹ�:�":�氺�V���� �@ߓ�����Q�`什����O��נ��A��[58�T���nQ���Zf��X1�5K��]]�      �X1���,�h���<��5g��e_���U�͂�֌Ⱦ	ń�*�-�j��P ��%�2�
?ټb�{�"��n�(�O���u:�P ;�&;+#:;?�C;�%H;�I;"�I;��I;�I;]vI;�WI;�AI;|2I;(I;F"I;a I;A"I;(I;x2I;�AI;�WI;]vI;�I;��I;(�I;�I;�%H;?�C;)#:;�&;�P ;��u:�O��n�"�b�{�?ټ%�2�P ��j��*�-�	ń�֌Ⱦ͂��U�e_��5g��<�h����,�      ~x�P9�R��uؿnQ��e_��6�_��X#�r���f��9�S�{�����l�B�	w�� �M���Ի��+�@=T���:�e;�\,;�/=;�BE;S�H;}�I;��I;��I;��I;�oI;�RI;>I;^/I;�%I;�I;GI;�I;�%I;^/I;>I;�RI;�oI;��I;��I;��I;x�I;Z�H;�BE;�/=;�\,;�e;��:�<T���+���Ի�M�	w��B�l�����{�9�S��f��r���X#�6�_�e_��nQ��uؿR��P9�      	Ŀ6g��'ﱿ���T����U��X#�t��d���HUo��#��hܽ����n<����=����� ��᝻F�Ժxt�9b��:�V;̇2;� @;U�F;�I;��I;C�I;+�I;l�I; hI;MI;�9I;�+I;�"I;lI;�I;iI;�"I;�+I;�9I;MI; hI;o�I;,�I;H�I;��I;�I;Y�F;� @;χ2;�V;Z��:�t�9D�Ժ�᝻�� �=�������n<�����hܽ�#�HUo�d���t���X#��U�T������'ﱿ6g��      ���U���U�v��RZ�[58�͂�q��d���foy�]1�_O��]什�`�M�����pyY�$�컗�T��1�t�u: ��:H#;98;�B;j�G;�lI;�I;�I;/�I;w�I;�_I;GI;�4I;%(I;�I;�I;I;�I;�I;&(I;�4I;GI;�_I;z�I;2�I;�I;�I;�lI;n�G;�B;98;I#;���:��u:�1���T�#��pyY����M���`�\什_O��]1�foy�d���q��͂�[58��RZ�U�v�U���      �3���/��X#��	��A��֌Ⱦ�f��GUo�^1�˰��|n��Լx��'��>ټ�@���k�м������39�#�:.R;e-;�/=;�	E;]xH;��I;�I;q�I;�I;vI;cWI;�@I;�/I;%$I;<I;�I;7I;�I;>I;%$I;�/I;�@I;eWI;vI;�I;v�I;�I;��I;axH;�	E;�/=;e-;.R;�#�:�39 ��μ���k��@���>ټ�'�Ӽx�|n��˰��]1�GUo��f��֌Ⱦ�A���	��X#���/�      w���ྃ�Ѿ(����נ�ń�9�S��#�`O��|n��J̀���2���𛼄�>� �Ի��B��#�4m:�G�:^ ;��5;�FA;��F;�I;R�I;U�I;��I;j�I;mjI;�NI;:I;�*I;�I;�I;�I;II;�I;�I;�I;�*I;:I;�NI;tjI;q�I;��I;W�I;P�I;�I;��F;�FA;��5;_ ;�G�:Dm:�#���B� �Ի��>�������2�J̀�|n��_O���#�9�S�ń��נ�(�����Ѿ��      �x���o��ń�HUo���O�*�-�{��hܽ]什Լx���2�tb��VR��X|U�^2��:��*갺�u�9��:
D;��,;�h<;crD;P%H;ÏI;j�I;��I;�I;�I;�^I;FI;W3I;�%I;�I;_I;iI;4I;hI;^I;�I;�%I;S3I;FI;�^I;�I;�I;��I;g�I;ʏI;Q%H;jrD;�h<;��,;D;��:�u�9갺:��\2��W|U�UR��tb����2�Լx�\什�hܽ{�*�-���O�HUo�ń��o��      ��4�g1��&������j�ཅ�������`��'���UR��F�]���!V���X���Io����:h�;&#;�6;RtA;Q�F;�	I;u�I;��I;q�I;�I;�pI;�SI;�=I;�,I;w I;�I;�I;GI;;I;GI;�I;�I;y I;�,I;�=I;�SI;�pI;�I;r�I;��I;}�I;�	I;U�F;ZtA;�6;3#;p�;���:@Go��X�� V��~��E�]�UR����'��`��������j��������&�f1�      k�ྲྀhܽn�н^y��`什P ��l��n<�M���>ټ��X|U���������1�������u:Sl�:�;b71;S)>;V	E;
JH;W�I;��I;��I;�I;׃I;YbI;�HI;$5I;c&I;gI;qI;<I;#I;
I;#I;:I;rI;gI;b&I;-5I;�HI;cbI;ރI;�I;��I;��I;W�I;JH;[	E;V)>;n71;�;Sl�:��u:�����1�������V|U����>ټM���n<�l�P ��`什^y��n�н�hܽ      Y+����c̀�,l��Q�%�2�B��������@����>�^2��"V���1�����#R:���:�;w\,;4;;�;C;�eG;X9I;��I;-�I;��I;D�I;�qI;�TI;`>I;5-I;1 I;zI;qI;�
I;I;I;I;�
I;rI;{I;1 I;<-I;g>I;�TI;�qI;F�I;��I;7�I;��I;Y9I;�eG;�;C;?;;}\,;�;���:�#R:���1� V��[2����>��@��������B�$�2��Q�-l�c̀���      �'��-$�_��Y����?ټw��<���pyY��k� �Ի<��Y�������#R:���:�R;�);ݍ8;��A;��F;4�H;)�I;��I;��I;��I;�I;�`I;�GI;�4I;�%I;JI;�I;�I;oI;I;FI;I;mI;�I;�I;HI;�%I;�4I;�GI;�`I;�I;��I;��I;��I;*�I;;�H;��F;��A;�8;�);�R;���: $R:����Y��8����Ի�k�oyY�<���	w��	?ټ���Y�_���-$�      ��ü^l��w����R��?ߓ�b�{��M��� � ��˼����B�"갺 Io���u:���:�R;/�';17;��@;��E;�lH;/�I;i�I;��I;�I;v�I;�lI;�QI;&<I;�+I;�I;�I;eI;�I;EI;0I;�I;,I;AI;�I;cI;�I;�I;�+I;)<I;�QI;�lI;t�I;�I;��I;h�I;5�I;�lH;�E;��@;17;3�';�R;���:��u:@Ho�갺��B�ʼ�� �컊� ��M�b�{�@ߓ��R��x���]l��      4yY��|U�K�I�@�7��� �"���Ի�᝻��T����#��u�9���:Ql�:�;�);17;0 @;;]E;�$H;ekI;
�I;V�I;��I;'�I;�wI;�ZI;�CI;w1I;N#I;%I;�I;-	I;rI;8I;m�H;��H;k�H;5I;rI;+	I;�I;,I;U#I;z1I;�CI;�ZI;�wI;0�I;��I;R�I;�I;kkI;�$H;?]E;/ @;17;�);�;Sl�:���:�u�9�#����T��᝻��Ի "��� �A�7�I�I��|U�      �kٻl�Ի�ǻ����V���n���+�8�Ժ��1��39Tm:��:j�;
�;z\,;�8;��@;A]E;�
H;LVI;q�I;��I;��I;c�I;��I;�bI;`JI;#7I;�'I;�I;,I;�
I;8I;;I;i�H;��H;z�H;��H;f�H;8I;8I;�
I;2I;�I;�'I;*7I;cJI;�bI;�I;i�I;��I;��I;x�I;QVI;�
H;<]E;Å@;�8;}\,;�;l�;��:dm:0�39��1�2�Ժ��+��n��V������ǻl�Ի      !p&��!��4���氺�O��<T�`t�9��u:�#�:�G�:D;)#;h71;;;;��A;��E;�$H;LVI;�I;��I;�I;��I;��I;iI;)PI;<I;�+I;I;�I;�I;�I;�I;3�H;��H;��H;�H;��H;��H;2�H;�I;�I;�I;�I;I;�+I;<I;)PI;iI;��I;��I;�I;��I;�I;SVI;�$H;��E;��A;>;;h71;*#;D;�G�:�#�:��u:�t�9�<T� �O��氺���4��!�      @�p� �,�� 9�ų9��":��u:��:b��:���:.R;\ ;��,;�6;U)>;�;C;��F;�lH;lkI;t�I;��I;��I;�I;r�I;�mI;wTI;&@I;�/I;!"I;VI;�I;�I;�I;t�H;t�H;��H;W�H;��H;P�H;��H;t�H;t�H;�I;�I;�I;WI;("I;�/I;%@I;~TI;�mI;n�I;�I;��I;��I;x�I;ikI;�lH;��F;�;C;R)>;�6;��,;` ;.R;���:X��:��:t�u:�":�ų9p!9 �,�      8��:��:�:��:���:�P ;�e;�V;L#;e-;��5;�h<;UtA;Z	E;�eG;8�H;2�I;�I;��I;�I;�I;�I;pI;LWI;�BI;@2I;�$I;qI;lI;B	I;tI;��H;��H;�H;Z�H;5�H;��H;/�H;W�H;�H;��H;��H;yI;D	I;oI;wI;�$I;D2I;�BI;LWI;pI;��I;�I;�I;��I;�I;3�I;7�H;�eG;V	E;StA;�h<;��5;e-;L#;�V;�e;�P ;��:���:��:{�:      I;�;.�;��;� ;�&;�\,;ڇ2;98;�/=;�FA;orD;U�F;JH;[9I;.�I;l�I;Y�I;��I;��I;r�I;pI;IXI;�DI;�3I;\&I;I;�I;
I;oI;��H;��H;��H;��H;;�H;J�H;�H;E�H;8�H;��H;��H;��H;��H;oI;~
I;�I;I;_&I;�3I;�DI;EXI;pI;u�I;��I;��I;U�I;o�I;.�I;[9I;JH;U�F;orD;�FA;�/=;98;ׇ2;�\,;�&; ;��;(�;�;      ��0;�51;�2;R�4;�07;-#:;�/=;� @;�B;�	E;��F;N%H;�	I;W�I;��I;��I;��I;��I;e�I;��I;�mI;DWI;�DI;�4I;;'I;-I;�I;|I;8I;. I;,�H;��H;{�H;��H;e�H;��H;j�H;��H;c�H;��H;|�H;��H;1�H;. I;8I;I;�I;1I;B'I;�4I;�DI;HWI;�mI;��I;c�I;��I;��I;��I;��I;R�I;�	I;Q%H;��F;�	E;�B;� @;�/=;#:;�07;P�4;�2;�51;      ��?;��?;��@;]tA;��B;F�C;�BE;X�F;l�G;axH;�I;ΏI;x�I;��I;7�I;��I;�I;2�I;�I;iI;�TI;�BI;�3I;G'I;�I;}I;I;�I;� I;}�H;�H;k�H;a�H;��H;��H;.�H;��H;(�H;��H;��H;a�H;g�H;�H;��H;� I;�I;I;�I;�I;D'I;�3I;�BI;�TI;iI;�I;.�I;�I;��I;6�I;��I;x�I;ϏI;�I;axH;j�G;U�F;�BE;<�C;�B;`tA;��@;��?;      ��F;?�F;��F;Y2G;%�G;�%H;Y�H;�I;�lI;��I;U�I;s�I;��I;��I;��I;��I;z�I;�wI;�bI;'PI;)@I;:2I;[&I;1I;{I;8I;I;� I;��H;C�H;x�H;V�H;|�H;(�H;]�H;��H;��H;��H;[�H;'�H;�H;S�H;z�H;F�H;��H;I;I;>I;�I;0I;[&I;@2I;)@I;&PI;�bI;�wI;}�I;��I;��I;��I;��I;p�I;[�I;��I;�lI;�I;[�H;�%H;:�G;l2G;��F;@�F;      r I;K'I;�:I;�XI;�{I;�I;~�I;�I;�I;�I;W�I;��I;m�I;�I;C�I;�I;�lI;�ZI;dJI;<I;�/I;�$I;!I;I;I;I;I;��H;s�H;��H;L�H;U�H;��H;��H;�H;��H;q�H;��H;�H;��H;��H;R�H;M�H;��H;q�H;��H;I;I;I;�I;"I;�$I;�/I;<I;cJI;�ZI;�lI;	�I;B�I;�I;m�I;��I;X�I;�I;�I;��I;x�I;�I;�{I;�XI;�:I;3'I;      ��I;f�I;��I;��I;��I;"�I;��I;C�I;�I;v�I;��I;�I;�I;ރI;�qI;�`I;�QI;�CI;#7I;�+I;'"I;mI;�I;|I;�I;� I;��H;j�H;��H;S�H;T�H;��H;��H;��H;��H;��H;p�H;��H;��H;��H;��H;��H;U�H;V�H;��H;l�H;��H;� I;�I;|I;�I;qI;'"I;�+I;%7I;�CI;�QI;�`I;�qI;݃I;�I;�I;��I;v�I;�I;C�I;��I;�I;��I;��I;��I;\�I;      ��I;��I;��I;[�I;��I;��I;��I;-�I;*�I;�I;q�I;�I;�pI;cbI;�TI;�GI;,<I;{1I;�'I;I;^I;gI;{
I;5I;� I;��H;l�H;��H;O�H;M�H;��H;P�H;?�H;��H;��H;��H;��H;��H;��H;��H;C�H;N�H;��H;N�H;O�H;��H;j�H;��H;� I;4I;|
I;iI;\I;I;�'I;x1I;,<I;�GI;�TI;bbI;�pI;�I;t�I;�I;+�I;-�I;��I;��I;��I;]�I;��I;��I;      .�I;<�I;��I;�I;��I;ߟI;��I;s�I;z�I;vI;ujI;�^I;�SI;�HI;d>I;�4I;�+I;N#I;�I;�I;�I;<	I;kI;* I;}�H;<�H;��H;V�H;R�H;��H;)�H;�H;8�H;��H;�H;��H;��H;��H;�H;��H;8�H;�H;,�H;��H;T�H;W�H;��H;@�H;��H;* I;nI;@	I;�I;�I;�I;K#I;�+I;�4I;d>I;�HI;�SI;�^I;ujI;vI;w�I;n�I;��I;�I;��I;�I;��I;<�I;      d�I;��I;w�I;��I;5|I;]vI;�oI;hI;�_I;mWI;�NI;FI;�=I;15I;?-I;�%I;�I;*I;2I;�I;�I;tI;��H;,�H;�H;t�H;L�H;X�H;��H;-�H;�H;�H;T�H;��H;v�H;/�H;��H;,�H;u�H;��H;W�H;�H;�H;,�H;��H;X�H;J�H;w�H;�H;,�H;��H;vI;�I;�I;2I;)I;�I;�%I;?-I;.5I;�=I;FI;�NI;mWI;�_I;hI;�oI;XvI;<|I;��I;v�I;��I;      MdI;�cI;CbI;�_I;)\I;�WI;�RI;MI;GI;�@I;:I;^3I;�,I;j&I;4 I;MI;�I;�I;�
I;�I;�I;��H;��H;��H;j�H;L�H;O�H;��H;R�H;�H;	�H;L�H;��H;#�H;��H;��H;��H;��H;��H;&�H;��H;O�H;	�H;�H;N�H;��H;O�H;M�H;m�H;��H;��H;��H;�I;�I;�
I;�I;�I;OI;7 I;j&I;�,I;\3I;:I;�@I;GI;MI;�RI;�WI;3\I;�_I;NbI;�cI;      �KI;NKI;�II;�GI;IEI;�AI;>I;�9I;�4I;�/I;�*I;�%I;| I;mI;I;�I;lI;.	I;=I;�I;��H;��H;��H;u�H;`�H;r�H;��H;��H;G�H;9�H;P�H;��H;�H;��H;G�H;�H;.�H;�H;F�H;��H;�H;��H;P�H;2�H;C�H;��H;��H;t�H;b�H;t�H;��H;��H;x�H;�I;?I;/	I;mI;�I;I;mI;z I;�%I;�*I;�/I;�4I;�9I;>I;�AI;MEI;�GI;JI;LKI;      �9I;w9I;�8I;7I;5I;m2I;]/I;�+I;)(I;0$I; I;�I;�I;{I;{I;�I;�I;sI;=I;7�H;}�H;�H;��H;��H;��H;�H;��H;��H;��H;��H;��H;%�H;��H;5�H;��H;��H;��H;��H;��H;6�H;��H;%�H;��H;��H;~�H;��H;��H;�H;��H;��H;��H; �H;u�H;2�H;=I;uI;�I;�I;{I;yI;�I;�I; I;.$I;)(I;�+I;e/I;k2I;5I;7I;�8I;�9I;      _.I;:.I;_-I;�+I;?*I;(I;�%I;�"I;�I;LI;�I;oI;�I;GI;�
I;vI;LI;9I;m�H;��H;��H;V�H;5�H;U�H;��H;O�H;�H;��H;��H;�H;n�H;��H;G�H;��H;��H;��H;z�H;��H;��H;��H;H�H;��H;m�H;�H;��H;��H;�H;P�H;��H;U�H;8�H;U�H;��H;��H;j�H;;I;MI;xI;�
I;FI;�I;lI;�I;LI;�I;�"I;�%I;(I;:*I;,I;^-I;<.I;      �'I;�'I;�&I;�%I;%$I;@"I;�I;sI;�I;�I;�I;sI;MI;*I;I;I;3I;j�H;��H;��H;^�H;/�H;B�H;��H;&�H;��H;��H;��H;��H;��H;*�H;��H;�H;��H;��H;a�H;p�H;c�H;��H;��H;�H;��H;)�H;��H;��H;��H;��H;��H;$�H;��H;F�H;/�H;W�H;��H;��H;m�H;5I;I;I;,I;MI;pI;�I;�I;�I;oI; I;@"I;&$I;�%I;�&I;�'I;      �%I;�%I;�$I;�#I;!"I;X I;JI;�I;I;:I;YI;BI;BI;'
I;I;JI;�I;��H;��H;�H;��H;��H;�H;\�H;��H;��H;i�H;q�H;��H;��H;��H;��H;.�H;��H;z�H;j�H;s�H;l�H;w�H;��H;0�H;��H;��H;��H;}�H;m�H;j�H;��H;��H;\�H;
�H;��H;��H;�H;��H; �H;�I;MI;I;)
I;@I;>I;ZI;:I;I;�I;OI;X I;"I;�#I;�$I;�%I;      �'I;�'I;�&I;�%I;&$I;C"I;�I;qI;�I;�I;�I;sI;NI;,I;I;I;3I;j�H;��H;��H;`�H;0�H;A�H;��H;&�H;��H;��H;��H;��H;��H;*�H;��H;�H;��H;��H;a�H;o�H;c�H;��H;��H;�H;��H;)�H;��H;��H;��H;��H;��H;$�H;��H;F�H;.�H;V�H;��H;��H;m�H;2I;I;I;*I;JI;pI;�I;�I;�I;pI;  I;A"I;&$I;�%I;�&I;�'I;      V.I;<.I;[-I;�+I;?*I;
(I;�%I;�"I;�I;JI;�I;mI;�I;FI;�
I;vI;JI;;I;m�H;��H;��H;V�H;4�H;S�H;��H;M�H;�H;��H;��H;�H;m�H;��H;G�H;��H;��H;��H;z�H;��H;��H;��H;J�H;��H;m�H;�H;��H;��H;�H;Q�H;��H;S�H;6�H;U�H;��H;��H;j�H;9I;LI;vI;�
I;FI;�I;oI;�I;JI;�I;�"I;�%I;(I;=*I;,I;_-I;=.I;      �9I;x9I;�8I;7I;5I;r2I;]/I;�+I;)(I;-$I; I;�I;�I;yI;{I;�I;�I;uI;?I;7�H;}�H;�H;��H;��H;��H;�H;��H;��H;��H;��H;��H;%�H;��H;5�H;��H;��H;��H;��H;��H;5�H;��H;%�H;��H;��H;~�H;��H;��H;�H;��H;��H;��H;�H;q�H;2�H;?I;sI;�I;�I;|I;{I;�I;�I; I;.$I;)(I;�+I;g/I;q2I;5I;7I;�8I;{9I;      �KI;SKI;JI;�GI;GEI;�AI;>I;�9I;�4I;�/I;�*I;�%I;y I;kI;�I;�I;jI;.	I;<I;�I;��H;��H;��H;t�H;b�H;q�H;��H;��H;J�H;9�H;O�H;��H;�H;��H;H�H;�H;,�H;�H;F�H;��H;�H;��H;O�H;4�H;@�H;��H;��H;t�H;`�H;q�H;��H;��H;t�H;�I;=I;-	I;jI;�I;I;kI;| I;�%I;�*I;�/I;�4I;�9I;>I;�AI;LEI;HI;JI;PKI;      BdI;�cI;9bI;�_I;*\I;�WI;�RI;MI;GI;�@I;:I;]3I;�,I;g&I;5 I;MI;�I;�I;�
I;�I;�I;��H;��H;��H;n�H;L�H;O�H;��H;U�H;�H;	�H;P�H;��H;"�H;��H;��H;��H;��H;��H;%�H;��H;L�H;�H;�H;O�H;��H;N�H;O�H;j�H;��H;��H;��H;�I;�I;�
I;�I;�I;OI;5 I;j&I;�,I;^3I;:I;�@I;GI;MI;�RI;�WI;*\I;�_I;?bI;�cI;      Z�I;��I;y�I;��I;:|I;]vI;�oI;hI;�_I;hWI;�NI;FI;�=I;.5I;=-I;�%I;�I;*I;2I;�I;�I;xI;��H;,�H;�H;r�H;L�H;X�H;��H;-�H;�H;�H;W�H;��H;x�H;,�H;��H;/�H;t�H;��H;T�H;�H;�H;)�H;��H;T�H;I�H;u�H;�H;'�H;��H;xI;�I;�I;3I;)I;�I;�%I;@-I;/5I;�=I;FI;�NI;hWI;�_I;hI;�oI;[vI;B|I;�I;|�I;��I;      3�I;A�I;��I;�I;��I;�I;��I;s�I;z�I;vI;njI;�^I;�SI;�HI;f>I;�4I;�+I;O#I;�I;�I;�I;@	I;kI;, I;��H;<�H;��H;X�H;U�H;��H;,�H;�H;8�H;��H;�H;��H;��H;��H;�H;��H;8�H;�H;)�H;��H;O�H;T�H;��H;?�H;}�H;& I;rI;?	I;�I;�I;�I;K#I;�+I;�4I;f>I;�HI;�SI;�^I;tjI;vI;w�I;r�I;��I;ޟI;��I;�I;��I;9�I;      ��I; �I;��I;R�I;��I;��I;��I;-�I;1�I; �I;m�I;�I;�pI;`bI;�TI;�GI;*<I;}1I;�'I;I;aI;iI;z
I;6I;� I;��H;l�H;��H;Q�H;N�H;��H;U�H;A�H;��H;��H;��H;��H;��H;��H;��H;C�H;P�H;��H;M�H;J�H;��H;i�H;��H;� I;/I;
I;iI;\I;I;�'I;x1I;*<I;�GI;�TI;_bI;�pI;�I;r�I; �I;+�I;0�I;��I;��I;��I;T�I;��I;��I;      �I;\�I;��I;��I;��I;.�I;��I;J�I;�I;v�I;��I;�I;�I;݃I;�qI;�`I;�QI;�CI;#7I;�+I;)"I;sI;�I;I;�I;� I;��H;l�H;��H;T�H;V�H;��H;��H;��H;��H;��H;q�H;��H;��H;��H;��H;��H;U�H;S�H;��H;f�H;��H;� I;�I;yI;�I;qI;$"I;�+I;&7I;�CI;�QI;�`I;�qI;݃I;�I;�I;��I;x�I;�I;C�I;��I;�I;��I;��I;��I;\�I;      a I;N'I;�:I;�XI;�{I;�I;{�I;�I;�I;�I;T�I;��I;j�I;�I;D�I;�I;�lI;�ZI;cJI;<I;�/I;�$I;I;I;I;I;I;��H;w�H;��H;L�H;X�H;��H;��H;�H;��H;p�H;��H;�H;��H;��H;U�H;M�H;��H;o�H;��H;I;I;I;�I;#I;�$I;�/I;<I;fJI;�ZI;�lI;	�I;D�I;�I;k�I;��I;W�I;�I;�I;�I;��I;�I;�{I;�XI;�:I;:'I;      ��F;>�F;��F;Y2G;*�G;&H;V�H;�I;�lI;��I;U�I;t�I;��I;��I;��I;��I;x�I;�wI;�bI;%PI;,@I;?2I;Y&I;3I;I;5I;I;I;��H;D�H;z�H;X�H;|�H;(�H;^�H;��H;��H;��H;Z�H;'�H;|�H;V�H;{�H;D�H;��H;� I;I;:I;}I;.I;\&I;?2I;)@I;'PI;�bI;�wI;}�I;��I;��I;��I;��I;n�I;Y�I;��I;�lI;�I;Y�H;�%H;4�G;\2G;��F;2�F;      ��?;��?;��@;atA;��B;K�C;�BE;U�F;j�G;`xH;�I;ΏI;v�I;��I;:�I;��I;�I;2�I;�I;iI;�TI;�BI;�3I;G'I;�I;yI;I;�I;� I;}�H;�H;n�H;`�H;��H;��H;+�H;��H;+�H;��H;��H;a�H;k�H;�H;}�H;� I;�I;I;}I;�I;E'I;�3I;�BI;�TI;iI;�I;-�I;�I;��I;8�I;��I;x�I;ˏI;�I;`xH;f�G;R�F;�BE;<�C; �B;`tA;��@;��?;      ��0;u51;�2;Y�4;�07;5#:;�/=;� @;	�B;�	E;��F;P%H;�	I;R�I;��I;��I;��I;��I;e�I;��I;�mI;HWI;�DI;�4I;B'I;*I;�I;I;<I;- I;0�H;��H;|�H;��H;d�H;��H;k�H;��H;a�H;��H;�H;��H;1�H;. I;8I;yI;�I;.I;>'I;�4I;�DI;GWI;�mI;��I;g�I;��I;��I;��I;��I;R�I;�	I;N%H;��F;�	E;�B;� @;�/=;*#:;�07;p�4;�2;`51;      D;�; �;��;� ;�&;�\,;ׇ2;98;�/=;�FA;orD;T�F;JH;_9I;1�I;n�I;Z�I;��I;��I;u�I;pI;FXI;�DI;�3I;X&I;I;�I;�
I;lI;��H;��H;��H;��H;;�H;I�H;�H;H�H;8�H;��H;��H;��H;��H;pI;~
I;�I;"I;\&I;�3I;�DI;FXI;pI;s�I;��I;��I;S�I;o�I;0�I;^9I;JH;U�F;lrD;�FA;�/=;98;և2;�\,;�&;� ;��;�;�;      <��:��:��:���:���:�P ;�e;�V;L#;e-;��5;�h<;UtA;X	E;�eG;;�H;3�I;�I;��I;�I;�I;��I;pI;LWI;�BI;?2I;�$I;wI;pI;B	I;xI;��H;��H;�H;W�H;0�H;��H;3�H;V�H;�H;��H;��H;{I;D	I;lI;sI;�$I;A2I;�BI;OWI;pI;��I;�I;�I;��I;�I;2�I;:�H;�eG;W	E;StA;�h<;��5;e-;O#;�V;�e;�P ;��:��:��:s�:      ��p� �,��!9�ų9Č":��u:��:`��:���:*R;_ ;��,;�6;S)>;�;C;��F;�lH;lkI;u�I;��I;��I;�I;r�I;�mI;~TI;"@I;�/I;%"I;ZI;�I;�I;�I;u�H;u�H;��H;T�H;��H;V�H;��H;o�H;u�H;�I;�I;�I;VI;""I;�/I;%@I;zTI;�mI;p�I;�I;��I;��I;v�I;hkI;�lH;��F;�;C;S)>;�6;��,;_ ;.R;���:`��:��:��u:�":�ų9�"9 �,�      	p&��!��4����氺�O��<T��t�9��u:�#�:�G�:D;*#;i71;?;;��A;��E;�$H;MVI;�I;��I;�I;��I;��I;iI;'PI;<I;�+I;I;�I;�I;�I;�I;7�H;��H;��H;�H;��H;��H;/�H;�I;�I;�I;�I;I;�+I;<I;'PI;	iI;�I;��I;�I;��I;�I;OVI;�$H;��E;��A;=;;g71;)#;D;�G�:�#�:��u:�t�9�<T� �O��氺���4��!�      �kٻl�Ի�ǻ����V���n���+�2�Ժ�1�0�39Tm:��:l�;
�;�\,;�8;��@;?]E;�
H;PVI;x�I;��I;��I;f�I;�I;�bI;`JI;&7I;�'I;�I;/I;�
I;9I;;I;j�H;��H;z�H;��H;f�H;8I;8I;�
I;0I;�I;�'I;"7I;cJI;�bI;��I;i�I;��I;��I;t�I;OVI;�
H;;]E;��@;��8;{\,;
�;l�;��:\m: �39��1�0�Ժ��+��n��V������ǻh�Ի      6yY��|U�L�I�@�7��� ��!���Ի�᝻��T���#��u�9���:Sl�:�;�);17;0 @;<]E;�$H;ikI;�I;Y�I;��I;2�I;�wI;�ZI;�CI;}1I;N#I;)I;�I;/	I;sI;9I;m�H;��H;n�H;4I;rI;-	I;�I;)I;P#I;x1I;�CI;�ZI;�wI;)�I;��I;V�I;�I;ekI;�$H;;]E;. @;17;�);�;Ql�:���:�u�9�#����T��᝻��Ի "��� �A�7�N�I��|U�      ��ü^l��w����R��?ߓ�b�{��M��� � ��ʼ����B�갺@Ho���u:���:�R;5�';17;��@;��E;�lH;5�I;l�I;��I;�I;x�I;�lI;�QI;,<I;�+I;�I;�I;hI;�I;EI;0I;�I;0I;?I;�I;cI;�I;�I;�+I;'<I;�QI;�lI;v�I;�I;��I;l�I;2�I;�lH;��E;��@;17;0�';�R;���:��u:@Ho�갺��B�˼���컊� ��M�a�{�@ߓ��R��x���]l��      �'��-$�_��X����
?ټw��<���oyY��k���Ի8��Y������$R:���:�R;�);ߍ8;��A;��F;;�H;0�I;��I;��I;��I;�I;�`I;�GI;�4I;�%I;KI;�I;�I;tI;I;FI;I;mI;�I;�I;GI;�%I;�4I;�GI;�`I;�I;��I;��I;��I;-�I;7�H;��F;��A;ݍ8;�);�R;���:�#R:����Y��:����Ի�k�pyY�<���	w��
?ټ���Y�`���-$�      Y+����c̀�,l��Q�$�2�B��������@����>�\2��!V���1����$R:���:�;z\,;:;;�;C;�eG;_9I;��I;7�I;��I;B�I;�qI;�TI;c>I;<-I;4 I;|I;xI;�
I;I;I;I;�
I;rI;zI;. I;8-I;`>I;�TI;�qI;C�I;��I;0�I;��I;[9I;�eG;�;C;;;;w\,;�;���:�#R:���1�!V��\2����>��@��������B�$�2��Q�-l�c̀���      k�ྲྀhܽo�н^y��`什P ��l��n<�M���>ټ��V|U��������1�x�����u:Wl�:
�;h71;Z)>;Z	E;JH;[�I;��I;��I;�I;ڃI;`bI;�HI;+5I;f&I;gI;tI;=I;#I;
I;%I;9I;qI;gI;_&I;&5I;�HI;]bI;ڃI;�I;��I;��I;X�I;JH;V	E;N)>;i71;�;Ql�:��u:�����1�������W|U����>ټM���n<�l�P ��`什^y��n�н�hܽ      ��4�f1��&������j�ཅ�������`��'���UR��E�]�~��V���X�� Ho����:l�;-#; �6;YtA;X�F;�	I;�I;��I;n�I;�I;�pI;�SI;�=I;�,I;y I;�I;�I;HI;<I;HI;�I;�I;y I;�,I;�=I;�SI;�pI;�I;n�I;��I;v�I;�	I;W�F;StA;�6;.#;h�;���:�Go��X�� V��~��F�]�UR����'��`��������j��������&�f1�      �x���o��ń�HUo���O�*�-�{��hܽ\什Լx���2�tb��UR��W|U�[2��8��갺�u�9��:D;��,;�h<;krD;U%H;ΏI;j�I;��I;�I;
�I;�^I;FI;W3I;�%I;�I;_I;hI;5I;iI;\I;�I;�%I;S3I;FI;�^I;�I;�I;��I;g�I;ÏI;Q%H;lrD;�h<;��,;D;��:�u�9갺:��\2��X|U�VR��tb����2�Լx�\什�hܽ{�*�-���O�HUo�ń��o��      w���ྃ�Ѿ(����נ�ń�9�S��#�_O��|n��J̀���2���𛼂�>� �Ի��B��#�Dm:�G�:e ;��5;�FA;��F;�I;R�I;S�I;��I;o�I;qjI;�NI;:I;�*I;�I;�I;�I;LI;�I;�I;�I;�*I;:I;�NI;pjI;o�I;��I;S�I;Q�I;�I;��F;�FA;��5;X ;�G�:4m:�#���B� �Ի��>�������2�J̀�|n��_O���#�9�S�ń��נ�(�����Ѿ��      �3���/��X#��	��A��֌Ⱦ�f��GUo�]1�˰��|n��Ӽx��'��>ټ�@���k�̼�� ���39�#�:4R;e-;�/=;�	E;fxH;��I;�I;q�I;�I;vI;hWI;�@I;�/I;'$I;>I;�I;7I;�I;>I;&$I;�/I;�@I;eWI;vI;�I;s�I;�I;��I;\xH;�	E;�/=;e-;&R;�#�:��39 ��̼���k��@���>ټ�'�Լx�|n��˰��^1�GUo��f��֌Ⱦ�A���	��X#���/�      ���U���U�v��RZ�[58�͂�q��d���foy�]1�_O��\什�`�M�����pyY�#�컘�T��1���u:��:L#;98;�B;p�G;�lI;�I;�I;2�I;x�I;�_I;GI;�4I;*(I;�I;�I;I;�I;�I;%(I;�4I;GI;�_I;v�I;1�I;�I;�I;�lI;j�G;�B;98;E#;���:��u:�1���T�#��pyY����M���`�]什_O��]1�foy�d���q��͂�[58��RZ�U�v�U���      	Ŀ6g��&ﱿ���T����U��X#�t��d���GUo��#��hܽ����n<����<����� ��᝻@�Ժ�t�9n��:�V;҇2;� @;[�F;�I;��I;C�I;+�I;k�I;hI;MI;�9I;�+I;�"I;lI;�I;iI;�"I;�+I;�9I;MI;hI;l�I;+�I;D�I;��I;�I;U�F;� @;Ї2;�V;R��:�t�9J�Ժ�᝻�� �=�������n<�����hܽ�#�HUo�d���t���X#��U�T������'ﱿ6g��      ~x�P9�R��uؿnQ��e_��6�_��X#�q���f��9�S�{�����l�B�	w���M���Ի��+��<T���:�e;�\,;�/=;�BE;T�H;z�I;��I;��I;��I;�oI;�RI;>I;^/I;~%I;�I;GI;�I;�%I;^/I;>I;�RI;�oI;��I;��I;��I;z�I;Z�H;�BE;�/=;�\,;�e;��:�<T���+���Ի�M�	w��B�l�����{�9�S��f��r���X#�6�_�e_��nQ��uؿR��P9�      �X1���,�h���<��5g��e_���U�͂�֌Ⱦ	ń�*�-�j��P ��%�2�
?ټa�{�"��n��O���u:�P ;�&;-#:;?�C;�%H;�I;$�I;��I;�I;bvI;�WI;�AI;{2I;(I;D"I;a I;D"I;(I;{2I;�AI;�WI;]vI;�I;��I;(�I;�I;�%H;?�C;.#:;�&;�P ;|�u:�O��n�"�b�{�?ټ&�2�P ��j��*�-�	ń�֌Ⱦ͂��U�e_��5g��<�h����,�      d��]]�5K��X1�Zf��nQ��T���[58��A���נ���O���`什�Q����@ߓ��� ��V���氺�":Ը�: ;�07;�B;0�G;�{I;��I;��I;��I;;|I;8\I;LEI;5I;3*I;4$I;,"I;0$I;6*I;5I;MEI;8\I;8|I;��I;��I;��I;�{I;8�G;�B;�07; ;Ը�:��":�氺�V���� �@ߓ�����Q�`什����O��נ��A��[58�T���nQ���Zf��X1�5K��]]�      N������4z���V��X1��<�uؿ����RZ��	�(���HUo����^y��-l�Y��R��C�7������ Ƴ9��:��;Y�4;ktA;\2G;�XI;��I;N�I;�I;��I;�_I;�GI;#7I;�+I;�%I;�#I;�%I;�+I;"7I;�GI;�_I;��I;�I;K�I;��I;�XI;f2G;jtA;[�4;��;���:�ų9�����D�7��R��Y�-l�^y�����HUo�(����	��RZ����uؿ�<��X1���V��4z�����      �o��e^���ē��4z�5K�h��R��'ﱿU�v��X#���Ѿń��&�o�нc̀�_��v���J�I��ǻ�4��"9��:4�;"�2;��@;��F;�:I;��I;��I;��I;z�I;NbI;�II;�8I;Z-I;�&I;�$I;�&I;\-I;�8I;JI;NbI;s�I;��I;��I;��I;�:I;��F;��@; �2;2�;��:�!9�4��ǻK�I�v���_��c̀�o�н�&�ń���Ѿ�X#�U�v�'ﱿR��h��5K��4z��ē�e^��      q'���X��e^�������]]���,�P9�6g��U�����/����o��g1��hܽ���-$�_l���|U�f�Ի!� �,�y�:�;�51;��?;5�F;A'I;c�I;�I;@�I;��I;�cI;AKI;{9I;!.I;|'I;�%I;y'I;".I;{9I;BKI;�cI;��I;C�I;�I;d�I;A'I;B�F;��?;�51;�;o�: �,�!�h�Ի�|U�_l���-$����hܽg1��o���ྙ�/�U���6g��P9���,��]]�����e^���X��      ����,������T���J�Q�Ǚ$�3�����;�}�H(�A�׾�T���L+���սk���� L���iO���ͻ���� m8do�:]�;U�1;��?;�uF;j I;i�I;��I;��I;YvI;�WI;�AI;�1I;�'I;�!I;�I;�!I;�'I;�1I;�AI;�WI;VvI;��I;��I;k�I;g I;�uF;��?;R�1;V�;`o�:�m8�����ͻ�iO� L����k����ս�L+��T��A�׾H(�;�}���3���Ǚ$�J�Q�T��������,��      �,��a��#P���{���K��x �����q�����w��$���Ҿg���  (���ѽҷ��(�����K�Fɻ,�����8v��:z�;��1;�@;m�F;!I;߿I;�I;��I;�uI;(WI;iAI;�1I;�'I;�!I;�I;�!I;�'I;�1I;jAI;)WI;�uI;��I;�I;�I;I;w�F;�@;��1;t�;l��:���8*��Fɻ�K����(�ҷ����ѽ  (�g�����Ҿ�$���w�q��������x ���K��{�#P��a��      ����#P�������d���;�#���㿳���#f�d��ž��z���=�ƽ%0v�T5�2����o@�����i��`u9AK�:];�73;�@;��F;JI;��I;R�I;V�I;�sI;�UI;E@I;�0I;�&I;!I;4I;!I;�&I;�0I;C@I;�UI;�sI;Z�I;P�I;��I;FI;��F;!�@;�73;];7K�:``u9zi������o@�2���T5�&0v�=�ƽ����z�žd��#f�������#����;���d����#P��      T����{���d��F�Ǚ$�:����ɿ.蒿��K�Q���j���Yb�E�1���s�a����?�����.��d��r�غذ�9�Y�:.X;�25;!�A;\!G;J7I;v�I;D�I;T�I;�pI;�SI;�>I;|/I;�%I;' I;2I;" I;�%I;{/I;�>I;�SI;�pI;V�I;D�I;v�I;I7I;b!G; �A;�25;(X;�Y�:���9p�غ�d����.�?������s�a�1���E��Yb��j��Q����K�.蒿��ɿ:��Ǚ$��F���d��{�      J�Q���K���;�Ǚ$��;
��޿�����w�q,���澝���'�D������I��#�G�����N��������X�����9:V��:�n!;��7;��B;M�G;�YI;,�I;Z�I;��I;�lI;wPI;<I;�-I;$I;�I;�I;�I;$I;�-I;<I;vPI;�lI;ÒI;Z�I;/�I;�YI;S�G;��B;��7;�n!;T��:��9:T����������N�����$�G��I������'�D��������q,���w�����޿�;
�Ǚ$���;���K�      Ǚ$��x �#��:���޿p���ʅ���F�}�
��~����z��$���ս���@2+���ϼPp�����P�]� �*���:�;�8';��:;��C;�H;�}I;�I;s�I;ًI;mgI;�LI; 9I;:+I;""I;�I;-I;�I;$"I;7+I;!9I;�LI;jgI;݋I;q�I;"�I;�}I;H;��C;��:;�8';�;��:�*�P�]�����Pp���ϼ@2+������ս�$���z��~��}�
��F�ʅ��p����޿:��#���x �      3��������㿊�ɿ���ʅ����P�d��<�׾�`��S�H����@��R�a���͡���D��ɻ� �@ح��W�:�;bI-;7|=; CE;��H;�I;��I;v�I;��I;iaI;#HI;�5I;r(I;�I;�I;TI;�I;�I;r(I;�5I;#HI;haI;��I;w�I;��I;�I;��H;!CE;8|=;`I-;�;�W�: ح�� ��ɻ�D�Ρ����R�a��@����S�H��`��<�׾d����P�ʅ�������ɿ�㿳���      ��q�������.蒿��w��F�d��ʰ� ����Yb�)����ѽ�%��D4�ٟ� X�����H���潺���9Hr�:��;�93;'Q@;}vF;�H;�I;��I;��I;�zI;�ZI;CI;�1I;c%I;BI;�I;&I;�I;DI;e%I;�1I;CI;�ZI;�zI;��I;��I;�I;�H;�vF;$Q@;�93;��;<r�:В�9�潺H����� X��؟�D4��%����ѽ)���Yb� ���ʰ�d���F���w�.蒿����q���      ;�}���w�#f���K�q,�}�
�<�׾ �����k���'�fz꽝I���;V�=M�
����iO�lG�qoE����6��:D� ;��$;��8;\�B;��G;/KI;�I;�I;A�I;qI;�SI;�=I;�-I;"I;nI;!I;�I;I;qI;"I;�-I;�=I;�SI;qI;D�I;�I;�I;/KI;��G;\�B;��8;��$;A� ;D��:���soE�jG໬iO�
���<M��;V��I��fz���'���k� ���<�׾}�
�q,���K�#f���w�      H(��$�d��Q������~���`���Yb���'��U�H$��C�m�&����ϼ�/��?��������غP8�9:��:�F;�G.;|=;IE;�\H; �I;y�I;z�I;��I;gI; LI;�7I;)I;qI;uI;uI;(I;tI;uI;rI;)I;�7I;LI;
gI;��I;}�I;v�I;�I;�\H;HE;|=;�G.;�F;H��:X8�9��غ����?���/����ϼ&��C�m�H$���U���'��Yb��`���~�����Q��d���$�      A�׾��Ҿž�j��������z�S�H�)��fz�H$���/v�2+�ݐ�����5��ɻ=4�8(�����:Z��:8o!;P6;lA;��F;s�H;��I;��I;�I;I}I;�\I;]DI;2I;r$I;�I;JI;�I;�I;�I;LI;�I;s$I;	2I;^DI;�\I;N}I;�I;��I;��I;w�H;��F;
lA;P6;9o!;p��:���:H(��94��ɻ��5���ݐ�2+��/v�H$��fz�)��S�H���z������j��ž��Ҿ      �T��f�����z��Yb�'�D��$�����ѽ�I��C�m�2+�������K�K�ﻙ�p�P������9'T�:�/;r�-;g�<;EzD;\H;�mI;��I;��I;��I;�oI;�RI;�<I;,I;�I;I;2I;�I;�I;�I;2I;I;�I;,I;�<I;�RI;�oI;��I;~�I;��I;�mI;]H;KzD;n�<;u�-;�/;/T�:���9D�����p��I�K�������2+�C�m��I����ѽ���$�'�D��Yb���z�f���      �L+�  (���E�������ս�@���%���;V�&��ܐ�����MS�N��'���D� �n8q�:�;d�$;�^7;+�A;f�F;��H;b�I;d�I;��I;߃I;TbI;�HI;5I;'&I;/I;@I;�I;�
I;
I;�
I;�I;@I;0I;'&I;5I;�HI;[bI;�I;��I;b�I;h�I;��H;i�F;1�A;_7;o�$;�;�p�:��n8xD�'��L��MS�����ܐ�&���;V��%���@����ս����E���  (�      ��ս��ѽ<�ƽ1����I�����R�a�D4�<M���ϼ��J�K�O��QG��bf���o���:�B�:�Y;��1;Pl>;�E;�/H;qI;��I;��I;ژI;�rI;�UI;�>I;�-I;b I;�I;�I;�
I;I;2I;I;�
I;�I;�I;b I;�-I;�>I;�UI;sI;ݘI;��I;�I;"qI;�/H;�E;Sl>;��1;�Y;�B�:��:��o�af�NG��N��I�K�����ϼ<M�D4�R�a�����I��1���<�ƽ��ѽ      j��ҷ��%0v�s�a�#�G�@2+���ן�	����/����5��)��df��ج��g:3�:
�;I-;g;;�NC;SG;�I;ɶI;�I;��I;	�I;
cI;~II;�5I;n&I;�I;5I;�I;�I;QI;[I;PI;�I;�I;7I;�I;u&I;�5I;�II;cI;�I;��I; �I;̶I;�I;SG;OC;g;;I-;�;?�:�g:�ج�_f�'�����5��/��	���؟���?2+�$�G�s�a�&0v�ҷ��      
��'�T5���������ϼ͡��X���iO�?���ɻ��p��D���o���g:�_�:AG;p*;p9;��A;�uF;�H;��I;��I;��I;H�I;�pI;3TI;N>I;-I;�I;{I;�I;VI;�I;�I;�I;�I;�I;VI;�I;zI;�I;!-I;T>I;:TI;�pI;D�I;��I;��I;ĔI;"�H;�uF;��A;u9;l*;GG;�_�:�g:��o��D⺙�p��ɻ?���iO�X��͡����ϼ������T5�&�      L�����3���?����N��Pp��D����hG�����64�L�����n8��:;�:GG;�(;��7;Z�@;��E;MQH;mI;��I;��I;��I;#}I;�^I;�FI;�3I;�$I;[I;�I;�	I;I;�I;��H;P�H;��H;�I;I;�	I;�I;aI;�$I;�3I;�FI;�^I;!}I;��I;��I;��I;mI;RQH;��E;_�@;��7;�(;HG;A�:��:��n8B���34�����hG໇���D�Pp��N��@���4������      �iO���K��o@���.���������ɻH��poE���غ0(�����9�p�:�B�:�;l*;��7;�P@;�\E;�H;�II;�I;g�I;�I;V�I;<hI;�NI;b:I;9*I;xI;�I;�I;I;I;2�H;a�H;��H;^�H;/�H;I;I;�I;�I;~I;:*I;f:I;�NI;:hI;_�I;�I;f�I;��I;�II;�H;�\E;�P@;��7;l*;
�;�B�:�p�:���9�'����غjoE�H���ɻ���������.��o@�ߔK�      ��ͻLɻ�����d�����@�]�� ��潺���p8�9���:'T�:�;�Y;I-;u9;Z�@;�\E;��G;05I;��I;D�I;ڵI;S�I;apI;�UI;S@I;2/I;{!I;�I;?I;�I;�I;!�H;��H;�H;��H;�H;��H;�H;�I;�I;DI;�I;}!I;9/I;V@I;�UI;ipI;X�I;ֵI;J�I;��I;75I;��G;�\E;`�@;s9;I-;�Y;�;/T�:���:h8�9����潺� �G�]�����d������Lɻ      ���.��si�X�غd����*�@׭����9<��:>��:h��:�/;g�$;��1;g;;��A;��E;�H;25I;8�I;��I;L�I;��I;�vI;L[I;^EI;�3I;2%I;�I;�I;P	I;�I;|�H;a�H;'�H;��H;n�H;��H;$�H;`�H;�H;�I;T	I;�I;�I;9%I;�3I;\EI;U[I;�vI;��I;P�I;��I;<�I;75I;�H;��E;��A;g;;��1;i�$;�/;n��:B��:@��:Ȓ�9�׭���*�V���r�غ�i�5��      @(m8���80_u9p��9P�9:
��:�W�:Dr�:>� ;�F;8o!;q�-;�^7;Pl>;�NC;�uF;NQH;�II;��I;��I;��I;��I;|zI;�_I;=II;I7I;a(I;^I;�I;I;�I;* I;r�H;��H;�H;��H;t�H;��H;�H;��H;s�H;' I;�I;!I;�I;dI;a(I;I7I;CII;_I;xzI;��I;��I;��I;��I;�II;QQH;�uF;OC;Ol>;�^7;r�-;?o!;�F;=� ;<r�:�W�:��:��9:���9�_u9`��8      Vo�:���:YK�:�Y�:B��:�;�;��;��$;�G.;P6;i�<;+�A;�E;SG; �H;mI;��I;H�I;O�I;��I;�{I;vaI;�KI;�9I;�*I;�I;�I;�I;%I;� I;��H;��H;k�H;��H;�H;��H;�H;��H;k�H;��H;��H;� I;(I;�I;�I;�I;�*I;�9I;�KI;paI;�{I;��I;P�I;J�I;��I;mI;!�H;SG;�E;-�A;m�<;P6;�G.;��$;��;�;�;v��:�Y�:CK�:z��:      n�;z�;];8X;�n!;�8';jI-;�93;��8;|=;lA;MzD;h�F;�/H;�I;ǔI;��I;j�I;ٵI;��I;|zI;qaI;vLI;!;I;`,I;0 I;I;�I;:I;�I;v�H;��H;e�H;m�H;
�H;U�H;"�H;O�H;�H;p�H;g�H;��H;z�H;�I;9I;�I;I;1 I;e,I;;I;rLI;vaI;~zI;��I;ݵI;h�I;��I;ȔI;�I;�/H;i�F;PzD;lA;|=;��8;�93;hI-;�8';�n!;:X;];`�;      R�1;��1;�73;�25;}�7;��:;.|=;#Q@;U�B;HE;��F;ZH;��H;"qI;ɶI;��I;��I;�I;R�I;�vI;}_I;�KI;;I;�,I;� I;I;�I;I;qI;��H;q�H;n�H;!�H;��H;n�H;��H;��H;��H;m�H;��H;#�H;m�H;x�H;��H;qI;I;�I;I;� I;�,I;;I;�KI;}_I;�vI;Q�I;�I;��I;��I;ʶI;qI;��H;]H;��F;HE;X�B;(Q@;-|=;��:;��7;�25;�73;��1;      ��?;�@;�@;�A;��B;�C;'CE;~vF;��G;�\H;z�H;�mI;b�I;�I; �I;��I;��I;a�I;opI;Y[I;III;�9I;e,I;� I;nI;^I;�I;�I;f�H;��H;��H;-�H;U�H;��H;��H;^�H;4�H;X�H;��H;��H;U�H;(�H;��H;��H;f�H;�I;�I;`I;rI;� I;e,I;�9I;III;V[I;opI;_�I;��I;��I;!�I;�I;c�I;�mI;{�H;�\H;��G;}vF;&CE;��C;��B;�A;�@;�@;      �uF;x�F;��F;X!G;@�G;H;��H; �H;2KI;%�I;��I;��I;c�I;��I;��I;K�I;(}I;>hI;�UI;\EI;N7I;�*I;. I;I;\I;�I;EI;��H;��H;��H;$�H;>�H;��H;]�H;��H;�H;��H;�H;��H;^�H;��H;;�H;'�H;��H;��H;��H;BI;�I;`I;I;- I;�*I;N7I;\EI;�UI;;hI;*}I;L�I;��I;��I;c�I;��I;��I;$�I;2KI;�H;��H;�H;W�G;j!G;��F;y�F;      u I;*I;BI;J7I;�YI;�}I;�I;�I;�I;v�I;��I;~�I;��I;ݘI;�I;�pI;�^I;�NI;W@I;�3I;k(I;�I;!I;�I;�I;BI;��H;"�H;��H;2�H;"�H;i�H;�H;�H;��H;�H;��H;�H;�H;�H;�H;f�H;#�H;2�H;��H;#�H;��H;HI;�I;�I;!I;�I;i(I;�3I;V@I;�NI;�^I;�pI;�I;טI;��I;~�I;��I;u�I;�I;�I;�I;�}I;�YI;C7I;@I;I;      e�I;�I;��I;y�I;�I;�I;��I;��I;�I;��I;�I;��I;��I;sI;
cI;5TI;�FI;_:I;4/I;4%I;dI;�I;�I;I;�I;��H;�H;��H;B�H;�H;W�H;��H;��H;�H;[�H;�H;��H;��H;Z�H;�H;��H;��H;Z�H;!�H;B�H;��H;�H;��H;�I;I;�I;�I;bI;4%I;4/I;\:I;�FI;7TI;
cI;sI;߃I;��I;�I;�I;�I;��I;��I;�I;%�I;}�I;��I;ڿI;      ��I;��I;L�I;T�I;N�I;s�I;y�I;��I;=�I;��I;M}I;�oI;VbI;�UI;�II;T>I;�3I;<*I;�!I;�I;�I;�I;6I;pI;b�H;��H;��H;@�H;/�H;U�H;��H;��H;��H;��H;|�H;5�H;.�H;1�H;z�H;��H;��H;��H;��H;U�H;/�H;C�H;��H;��H;g�H;mI;9I;�I;�I;�I;�!I;:*I;�3I;T>I;�II;�UI;UbI;�oI;P}I;��I;>�I;��I;y�I;j�I;W�I;X�I;K�I;��I;      ��I;��I;a�I;M�I;��I;֋I;��I;�zI;qI;gI;�\I;�RI;�HI;�>I;�5I;-I;�$I;vI;�I;�I;"I; I;�I;��H;��H;��H;/�H;!�H;X�H;��H;��H;��H;��H;�H;��H;|�H;]�H;y�H;��H;�H;��H;��H;��H;��H;X�H;%�H;/�H;��H;��H;��H;�I;%I;I;�I;�I;tI;�$I;!-I;�5I;�>I;�HI;�RI;�\I;gI;qI;�zI;��I;ًI;��I;Y�I;_�I;��I;      VvI;�uI;�sI;�pI;�lI;kgI;haI;�ZI;�SI;LI;bDI;�<I;5I;�-I;x&I;�I;fI;�I;DI;X	I;�I;� I;s�H;r�H;��H;!�H;!�H;[�H;��H;��H;��H;��H;��H;Z�H;�H;��H;��H;��H;�H;^�H;��H;��H;��H;��H;��H;[�H;"�H;&�H;��H;r�H;z�H;� I;�I;S	I;FI;�I;fI;�I;x&I;�-I;5I;�<I;dDI;
LI;�SI;�ZI;paI;cgI;�lI;�pI;�sI;�uI;      �WI;/WI;�UI;�SI;gPI;�LI; HI;CI;�=I;�7I;	2I;,I;+&I;i I;�I;~I;�I;�I;�I;�I;1 I;��H;��H;h�H;*�H;3�H;c�H;��H;��H;��H;��H;��H;B�H;��H;|�H;A�H;K�H;A�H;{�H;��H;H�H;��H;��H;��H;��H;��H;c�H;7�H;.�H;e�H;��H;��H;- I;�I;�I;�I;�I;�I;�I;i I;)&I;,I;2I;�7I;�=I;CI;)HI;�LI;pPI;�SI;�UI;/WI;      �AI;tAI;E@I;�>I;<I;9I;�5I;�1I;�-I;	)I;u$I;�I;2I;�I;:I;�I;�	I;I;�I;��H;}�H;��H;a�H;�H;U�H;��H;�H;��H;��H;��H;��H;B�H;��H;\�H;�H;��H;��H;��H;�H;_�H;��H;H�H;��H;��H;��H;��H;�H;��H;Y�H;�H;g�H;��H;w�H;�H;�I;I;�	I;�I;<I;�I;2I;�I;v$I;	)I;�-I;�1I;�5I;9I;<I;�>I;O@I;tAI;      �1I;�1I;�0I;q/I;�-I;-+I;r(I;j%I;	"I;zI;�I;I;GI;�I;�I;]I;I;I;&�H;g�H;��H;j�H;i�H;��H;��H;T�H;�H;�H;��H;�H;U�H;��H;]�H;��H;��H;��H;�H;��H;��H;��H;`�H;��H;U�H;�H;��H;��H;�H;V�H;��H;��H;p�H;h�H;��H;^�H;#�H;I;I;[I;�I;�I;EI;I;�I;xI;"I;e%I;y(I;)+I;�-I;v/I;�0I;�1I;      �'I;�'I;�&I;�%I;$I;"I;�I;LI;tI;�I;TI;@I;�I;�
I;�I;�I;�I;2�H;��H;+�H;�H;��H;�H;b�H;��H;��H;z�H;[�H;~�H;��H;�H;{�H;�H;��H;�H;\�H;W�H;\�H;}�H;��H;�H;�H;�H;��H;y�H;U�H;z�H;��H;��H;b�H;�H;��H;�H;$�H;��H;3�H;�I;�I;�I;�
I;�I;=I;XI;�I;rI;JI;�I;"I;$I;�%I;�&I;�'I;      �!I;�!I;!I;" I;�I;�I;�I;�I;I;|I;�I;�I;�
I;I;TI;�I;��H;^�H;�H;��H;��H;�H;L�H;��H;W�H;�H;�H; �H;8�H;}�H;��H;A�H;��H;��H;a�H;*�H;-�H;-�H;\�H;��H;��H;F�H;��H;x�H;4�H;��H;�H;�H;T�H;��H;P�H;�H;��H;��H;�H;_�H;��H;�I;TI;I;�
I;�I;�I;|I;I;�I;�I;�I;�I;# I;!I;�!I;      �I;�I;AI;.I;�I;#I;WI;*I;�I;+I;�I;�I;
I;;I;dI;�I;Z�H;��H;��H;v�H;��H;��H;�H;��H;.�H;��H;��H;��H;1�H;^�H;��H;J�H;��H;z�H;X�H;(�H;�H;*�H;T�H;{�H;��H;M�H;��H;Y�H;,�H;��H;��H;��H;,�H;��H;"�H;��H;z�H;o�H;��H;��H;W�H;�I;bI;=I;	
I;�I;�I;)I;�I;)I;\I;#I;�I;3I;>I;�I;      �!I;�!I;!I; I;�I;�I;�I;�I;I;{I;�I;�I;�
I;I;SI;�I;��H;\�H;�H;��H;��H;�H;L�H;��H;W�H;�H;�H; �H;:�H;|�H;��H;D�H;��H;��H;a�H;(�H;-�H;+�H;[�H;��H;��H;F�H;��H;v�H;4�H;��H;�H;�H;T�H;��H;O�H;�H;��H;��H;�H;_�H;��H;�I;TI;I;�
I;�I;�I;yI;I;�I;�I;�I;�I;' I;!I;�!I;      �'I;�'I;�&I;�%I;$I;"I;�I;NI;rI;I;SI;?I;�I;�
I;�I;�I;�I;2�H;��H;)�H;�H;��H;�H;`�H;��H;��H;z�H;Z�H;~�H;��H;�H;{�H;�H;��H;~�H;\�H;U�H;\�H;}�H;��H;�H;|�H;�H;��H;y�H;T�H;z�H;��H;��H;`�H;�H;��H;�H;"�H;��H;3�H;�I;�I;�I;�
I;�I;?I;XI;I;rI;PI;�I;"I;$I;�%I;�&I;�'I;      �1I;�1I;�0I;u/I;�-I;2+I;r(I;l%I;	"I;wI;�I;I;EI;�I;�I;[I;I;I;%�H;d�H;��H;k�H;i�H;��H;��H;T�H;�H;�H; �H;�H;U�H;��H;]�H;��H;��H;��H;~�H;��H;��H;��H;]�H;��H;U�H;�H;��H;��H;�H;W�H;��H;��H;o�H;h�H;��H;`�H;%�H;I;I;]I;�I;�I;EI;I;�I;wI;"I;i%I;|(I;/+I;�-I;v/I;�0I;�1I;      �AI;{AI;H@I;>I;<I;9I;�5I;�1I;�-I;)I;r$I;�I;0I;�I;<I;�I;�	I;I;�I;��H;~�H;��H;a�H;�H;Y�H;��H;�H;��H;��H;��H;��H;D�H;��H;]�H;�H;��H;��H;��H;�H;\�H;��H;E�H;��H;��H;��H;��H;�H;��H;U�H;�H;g�H;��H;u�H;��H;�I;I;�	I;�I;<I;�I;4I;�I;w$I;)I;�-I;�1I;�5I;9I;<I;�>I;T@I;vAI;      �WI;3WI;�UI;�SI;gPI;�LI;&HI;CI;�=I;�7I;2I;,I;)&I;h I;�I;I;�I;�I;�I;�I;4 I;��H;��H;g�H;.�H;4�H;c�H;��H;��H;��H;��H;��H;E�H;��H;~�H;?�H;J�H;C�H;z�H;��H;E�H;��H;��H;��H;��H;��H;a�H;4�H;*�H;`�H;��H;��H;, I;�I;�I;�I;�I;I;�I;i I;,&I;,I;2I;�7I;�=I;CI;'HI;�LI;hPI;�SI;�UI;-WI;      NvI;�uI;�sI;�pI;�lI;jgI;iaI;�ZI;�SI;LI;aDI;�<I;5I;�-I;w&I;�I;fI;�I;DI;T	I;�I;� I;t�H;r�H;��H;�H;!�H;[�H;��H;��H;��H;��H;��H;\�H;�H;��H;��H;��H;	�H;]�H;��H;��H;��H;��H;��H;W�H;�H;#�H;��H;p�H;{�H;� I;�I;T	I;GI;�I;hI;�I;x&I;�-I;5I;�<I;dDI;LI;�SI;�ZI;paI;ggI;�lI;�pI;�sI;�uI;      ��I;��I;Y�I;Y�I;��I;�I;��I;�zI;qI;gI;�\I;�RI;�HI;�>I;�5I;-I;�$I;wI;�I;�I;%I;$I;�I;��H;��H;��H;1�H;#�H;[�H;��H;��H;��H;��H;�H;��H;y�H;\�H;{�H;��H;�H;��H;��H;��H;��H;T�H;!�H;.�H;��H;��H;��H;�I;"I;I;�I;�I;tI;�$I; -I;�5I;�>I;�HI;�RI;�\I;gI;qI;�zI;��I;ӋI;��I;`�I;d�I;��I;      ��I;��I;[�I;K�I;@�I;x�I;v�I;��I;B�I;��I;J}I;�oI;TbI;�UI;�II;T>I;�3I;?*I;~!I;�I;�I;�I;4I;qI;f�H;��H;��H;B�H;2�H;T�H;��H;��H;��H;��H;|�H;3�H;-�H;3�H;z�H;��H;��H;��H;��H;T�H;)�H;?�H;��H;��H;c�H;jI;:I;�I;�I;�I;�!I;:*I;�3I;V>I;�II;�UI;UbI;�oI;N}I;��I;>�I;��I;}�I;q�I;O�I;M�I;[�I;��I;      p�I;ؿI;��I;z�I;�I;*�I;��I;��I;�I;�I;�I;��I;߃I;sI;cI;7TI;�FI;`:I;3/I;2%I;eI;�I;�I;I;�I;��H;�H;��H;G�H;�H;X�H;��H;��H;�H;^�H; �H;��H; �H;[�H;�H;��H;��H;[�H;�H;@�H;��H;�H;��H;�I;I;�I;�I;aI;4%I;6/I;\:I;�FI;7TI;cI;sI;߃I;��I;�I;��I;�I;��I;��I;�I;$�I;}�I;��I;ؿI;      c I;-I;?I;V7I;�YI;�}I;�I;�I;�I;v�I;��I;��I;��I;ژI;�I;�pI;�^I;�NI;V@I;�3I;l(I;�I;I;�I;�I;AI;��H;#�H;��H;1�H;"�H;j�H;�H;�H;��H;�H;��H;�H;�H;�H;�H;l�H;#�H;1�H;��H;!�H;��H;GI;�I;�I;$I;�I;g(I;�3I;W@I;�NI;�^I;�pI;�I;٘I;��I;|�I;��I;u�I;�I;�I;�I;�}I;�YI;X7I;?I;I;      �uF;u�F;��F;V!G;D�G;H;��H;!�H;0KI;"�I;��I;��I;d�I;��I; �I;L�I;'}I;AhI;�UI;[EI;P7I;�*I;* I;I;^I;�I;DI;��H;��H;��H;'�H;@�H;��H;^�H;��H;�H;��H;�H;��H;]�H;��H;@�H;(�H;��H;��H;��H;EI;�I;]I;I;. I;�*I;N7I;^EI;�UI;:hI;*}I;M�I;�I;��I;`�I;��I;��I;%�I;,KI;�H;��H;�H;P�G;\!G;��F;j�F;      ��?;�@;�@;�A;��B;�C;#CE;zvF;��G;�\H;w�H;�mI;b�I;�I;$�I;��I;��I;c�I;ppI;W[I;JII;�9I;e,I;� I;tI;YI;�I;�I;k�H;��H;��H;1�H;U�H;��H;��H;[�H;3�H;[�H;��H;��H;V�H;.�H;��H;��H;f�H;�I;�I;]I;nI;� I;h,I;�9I;III;Y[I;rpI;\�I;��I;��I;!�I;�I;b�I;�mI;w�H;�\H;��G;|vF;'CE;��C;��B;�A;�@;�@;      3�1;��1;�73;�25;x�7;��:;.|=;%Q@;[�B;DE;��F;_H;��H;qI;̶I;��I;��I;�I;R�I;�vI;�_I;�KI;;I;�,I;� I;I;�I;I;uI;��H;t�H;t�H;$�H;��H;p�H;��H;��H;��H;k�H;��H;&�H;o�H;w�H;��H;qI;I;�I;I;� I;�,I;;I;�KI;_I;�vI;S�I;�I;��I;��I;ɶI;qI;��H;ZH;��F;GE;U�B;!Q@;1|=;��:;��7;�25;�73;��1;      d�;v�;�\;DX;�n!;�8';dI-;�93;��8;|=;lA;PzD;f�F;�/H;�I;ʔI;��I;m�I;ڵI;��I;~zI;vaI;sLI;!;I;g,I;* I;I;�I;@I;�I;x�H;�H;g�H;m�H;�H;U�H;%�H;S�H;�H;l�H;e�H;�H;{�H;�I;9I;�I;!I;. I;a,I;;I;uLI;taI;~zI;��I;ݵI;d�I;��I;ǔI;�I;�/H;i�F;LzD;lA;|=;��8;�93;dI-;�8';�n!;FX;�\;d�;      Vo�:���:AK�:�Y�:F��: �;�;��;��$;�G.;P6;p�<;-�A;�E;SG;$�H;mI;��I;G�I;P�I;��I;�{I;taI;�KI;�9I;�*I;�I;�I;�I;%I;� I;��H;��H;k�H;��H;�H;��H;�H;��H;j�H;��H;��H;� I;(I;�I;�I;�I;�*I;�9I;�KI;taI;�{I;��I;P�I;H�I;~�I;mI;!�H;SG;�E;-�A;k�<;P6;�G.;��$;��;�;�;p��:�Y�:=K�:r��:      �%m8���8 `u9���9P�9:��:�W�:Br�:D� ;�F;;o!;s�-;�^7;Pl>;OC;�uF;QQH;�II;��I;��I;��I;��I;{zI;�_I;DII;G7I;^(I;bI;�I;I;�I;- I;u�H;��H;�H;��H;u�H;��H; �H;��H;s�H;* I;�I;I;�I;bI;d(I;I7I;?II;�_I;zzI;��I;��I;��I;��I;�II;QQH;�uF;OC;Pl>;�^7;r�-;<o!;�F;@� ;Jr�:�W�:��:��9:���9�`u9���8      |��*��zi�V�غh�����*��׭���9L��:B��:n��:�/;h�$;��1;g;;��A;��E;�H;25I;;�I;��I;Q�I;��I;�vI;U[I;[EI;�3I;6%I;�I;�I;T	I;�I;�H;b�H;'�H;��H;p�H;��H;$�H;^�H;}�H;�I;T	I;�I;�I;5%I;�3I;\EI;O[I;�vI;��I;O�I;��I;9�I;35I;�H;��E;��A;g;;��1;h�$;�/;p��:<��:@��:Ȓ�9`׭��*�V���l�غ|i�1��      ��ͻLɻ�����d�����@�]�� ��潺���h8�9���:/T�:�;�Y;I-;w9;]�@;�\E;��G;35I;��I;J�I;ܵI;S�I;kpI;�UI;T@I;4/I;!I;�I;CI;�I;�I;"�H;��H;�H;��H;�H;��H;�H;�I;�I;DI;�I;{!I;4/I;T@I;�UI;dpI;X�I;ڵI;G�I;��I;55I;��G;�\E;\�@;r9;I-;�Y;�;-T�:���:h8�9����潺� �B�]�����d������Iɻ      �iO�ޔK��o@���.���������ɻ�G��loE���غ(�����9�p�:�B�:�;p*;��7;�P@;�\E;�H;�II;��I;k�I;�I;_�I;<hI;�NI;c:I;<*I;xI;�I;�I;I;I;0�H;a�H;��H;c�H;-�H;I;I;�I;�I;zI;9*I;c:I;�NI;;hI;W�I;�I;h�I;��I;�II;�H;�\E;�P@;��7;n*;
�;�B�:�p�:���9 (����غjoE� H���ɻ���������.��o@�ޔK�      L�����2���>����N��Pp��D����hG�����54�>�����n8��:E�:KG;�(;��7;Z�@;��E;RQH;mI;��I;��I;��I;$}I;�^I;�FI;�3I;�$I;aI;�I;�	I;I;�I;��H;S�H;��H;�I;I;�	I;�I;_I;�$I;�3I;�FI;�^I;!}I;��I;��I;��I;mI;KQH;��E;Z�@;��7;�(;GG;A�:��:@�n8D���34�����gG໇���D�Pp��N��@���4������      
��'�T5���������ϼ͡��X���iO�?���ɻ��p��D���o���g:�_�:CG;p*;r9;��A;�uF;$�H;ǔI;��I;��I;H�I;�pI;3TI;T>I;-I;�I;I;�I;]I;�I;�I;�I;�I;�I;TI;�I;zI;�I;-I;Q>I;5TI;�pI;D�I;��I;��I;ƔI;!�H;�uF;��A;o9;l*;CG;�_�:�g:��o��D⺛�p��ɻ?���iO�X��Ρ����ϼ������U5�'�      k��ҷ��&0v�r�a�#�G�?2+���ן�	����/����5��'��^f��ج���g:?�:
�;I-;g;;OC;SG;�I;ͶI;!�I; �I;�I;cI;�II;�5I;t&I;�I;7I;�I;�I;NI;[I;PI;�I;�I;7I;�I;p&I;�5I;�II;cI;�I;��I;�I;̶I;�I;SG;�NC;g;;I-;�;?�:�g:�ج�af�(�����5��/��	���؟���?2+�$�G�s�a�&0v�ҷ��      ��ս��ѽ=�ƽ1����I�����R�a�D4�<M���ϼ��I�K�N��NG��[f�p�o���:�B�:�Y;��1;Vl>;�E;�/H;#qI;�I;��I;ژI; sI;�UI;�>I;�-I;e I;�I;�I;�
I;I;2I;I;�
I;�I;�I;` I;�-I;�>I;�UI;sI;ژI;��I;��I;#qI;�/H;�E;Kl>;��1;�Y;�B�:��:��o�bf�NG��O��J�K�����ϼ<M�D4�R�a�����I��1���<�ƽ��ѽ      �L+�  (���E�������ս�@���%���;V�&��ܐ�����~MS�M��$��vD�@�n8q�:�;k�$;_7;/�A;l�F; �H;i�I;c�I;��I;��I;[bI;�HI;5I;)&I;2I;BI;�I;�
I;
I;�
I;�I;@I;0I;%&I;5I;�HI;XbI;��I;��I;`�I;a�I;��H;k�F;+�A;�^7;l�$;�;�p�:@�n8~D�&��M��MS�����ܐ�&���;V��%���@����ս����E���  (�      �T��f�����z��Yb�'�D��$�����ѽ�I��C�m�2+�������I�K�ﻖ�p�J������9/T�:�/;y�-;k�<;LzD;cH;�mI;��I;|�I;��I;�oI;�RI;�<I;,I;�I;I;2I;�I;�I;�I;/I;I;�I;,I;�<I;�RI;�oI;��I;z�I;��I;�mI;]H;MzD;g�<;l�-;�/;'T�:���9J�����p��J�K�������2+�C�m��I����ѽ���$�'�D��Yb���z�f���      A�׾��Ҿž�j��������z�S�H�)��fz�H$���/v�2+�ܐ�����5��ɻ:4�H(�����:h��:?o!;P6;lA;��F;z�H;��I;��I;�I;L}I;�\I;aDI;2I;u$I;�I;II;�I;�I;�I;II;�I;s$I;2I;`DI;�\I;L}I;�I;��I;��I;q�H;��F;lA;P6;4o!;h��:���:P(��94��ɻ��5���ݐ�2+��/v�H$��fz�)��S�H���z������j��ž��Ҿ      H(��$�d��P������~���`���Yb���'��U�H$��C�m�&����ϼ�/��>��������غX8�9D��:�F;�G.;|=;LE;�\H; �I;v�I;y�I;��I;	gI;LI;�7I;)I;tI;rI;tI;)I;tI;tI;qI;)I;�7I;LI;gI;��I;|�I;u�I;�I;�\H;KE;|=;�G.;�F;D��:H8�9��غ����?���/����ϼ&��C�m�H$���U���'��Yb��`���~�����Q��d���$�      ;�}���w�#f���K�q,�}�
�<�׾ �����k���'�fz꽝I���;V�<M�	����iO�jG�soE����@��:H� ;��$;��8;_�B;�G;/KI;�I;�I;D�I;qI;�SI;�=I;�-I;	"I;mI;I;�I;I;nI;	"I;�-I;�=I;�SI;	qI;D�I;�I;�I;0KI;��G;`�B;��8;��$;>� ;@��:���soE�jG໬iO�
���<M��;V��I��fz���'���k� ���<�׾}�
�q,���K�#f���w�      ��q�������.蒿��w��F�d��ʰ� ����Yb�)����ѽ�%��D4�؟�X�����H���潺В�9Pr�:��;�93;+Q@;�vF;�H;	�I;��I;��I;�zI;�ZI;CI;�1I;f%I;CI;�I;%I;�I;DI;e%I;�1I;CI;�ZI;�zI;��I;��I;�I;�H;|vF;(Q@;�93;��;:r�:В�9�潺H����� X��ٟ�D4��%����ѽ)���Yb� ���ʰ�d���F���w�.蒿����q���      3��������㿊�ɿ���ʅ����P�d��<�׾�`��S�H����@��R�a���͡���D��ɻ� ��׭��W�:�;dI-;;|=;!CE;��H;�I;��I;w�I;��I;laI;#HI;�5I;u(I;�I;�I;UI;�I;�I;r(I;�5I;%HI;iaI;��I;v�I;��I;�I;��H;CE;;|=;dI-;�;�W�:�׭�� ��ɻ�D�Ρ����R�a��@����S�H��`��<�׾d����P�ʅ�������ɿ�㿳���      Ǚ$��x �#��:���޿p���ʅ���F�}�
��~����z��$���ս���@2+���ϼPp�����N�]��*���:�;�8';��:;��C;�H;�}I;�I;t�I;ۋI;ogI;�LI;9I;:+I;!"I;�I;-I;�I;""I;9+I; 9I;�LI;kgI;ڋI;s�I;"�I;�}I;H;��C;��:;�8';�;
��:�*�R�]�����Pp���ϼ@2+������ս�$���z��~��}�
��F�ʅ��p����޿:��#���x �      J�Q���K���;�Ǚ$��;
��޿�����w�q,���澝���'�D������I��#�G�����N��������T�����9:\��:�n!;��7;��B;J�G;�YI;+�I;\�I;��I;�lI;vPI;<I;�-I;$I;�I;�I;�I;$I;�-I;<I;uPI;�lI;��I;\�I;.�I;�YI;S�G;��B;��7;�n!;V��:x�9:P����������N�����$�G��I������'�D��������q,���w�����޿�;
�Ǚ$���;���K�      T����{���d��F�Ǚ$�:����ɿ.蒿��K�Q���j���Yb�E�1���s�a����?�����.��d��l�غ��9�Y�:.X;�25;!�A;X!G;I7I;t�I;D�I;S�I;�pI;�SI;�>I;}/I;�%I;& I;3I;# I;�%I;y/I;�>I;�SI;�pI;W�I;F�I;w�I;I7I;b!G; �A;�25;*X;�Y�:���9l�غ�d����.�>������s�a�1���E��Yb��j��Q����K�.蒿��ɿ:��Ǚ$��F���d��{�      ����#P�������d���;�#���㿳���#f�d��ž��z���=�ƽ&0v�T5�2����o@�����}i��`u9=K�:];�73;"�@;��F;II;��I;R�I;V�I;�sI;�UI;B@I;�0I;�&I;!I;4I;!I;�&I;�0I;C@I;�UI;�sI;Z�I;P�I;��I;GI;��F;!�@;�73;];7K�:``u9yi������o@�2���T5�&0v�=�ƽ����z�žd��#f�������#����;���d����#P��      �,��a��#P���{���K��x �����q�����w��$���Ҿg���  (���ѽҷ��(�����K�Fɻ*�����8v��:z�;��1;�@;k�F;!I;߿I;�I;��I;�uI;(WI;iAI;�1I;�'I;�!I;�I;�!I;�'I;�1I;jAI;*WI;�uI;��I;�I;�I;!I;x�F;�@;��1;t�;p��:���8)��Hɻ�K����(�ҷ����ѽ  (�g�����Ҿ�$���w�q��������x ���K��{�#P��a��      ඕ�S���Ѭ��-�_���7�{�}߿����,b��V�.l¾Gx�c.���Ž��t�*��f����?�N��)��`�x9���:P�;��2;3@@;`fF;9�H;��I;S�I;!|I;�[I;�CI;2I;�%I;_I;�I;4I;�I;^I;�%I;	2I;�CI;�[I;&|I;R�I;��I;<�H;mfF;1@@;��2;F�;���:�x9&��N����?�f��*����t���Žc.�Gx�.l¾�V��,b����}߿{���7�-�_�Ѭ��S���      S���E���$}��+Y��3�����$ڿ&��Ľ\����(���s��3�5����p�d�U���<<�:������`��9I��:ϻ;R%3;Ep@;�yF;��H;��I;�I;�{I;O[I;RCI;�1I;U%I;!I;[I;I;WI;#I;T%I;�1I;SCI;K[I;�{I;�I;��I;��H;�yF;Dp@;L%3;Ȼ;=��:8��9����;���<<�U��c��p�5����3��s�(�����Ľ\�&���$ڿ����3��+Y�$}�E���      Ѭ��$}�>tf��lG�ע%��p�.�ʿZ����>M����V�����d�Ȥ�̷�.�d��
��I���1�h���d�ຠ��9���:;�U4;��@;ӱF;4�H;܎I;��I;�yI;�YI;<BI;�0I;�$I;�I;�I;�I;�I;�I;�$I;�0I;<BI;�YI;�yI;��I;ގI;1�H;ܱF;��@;�U4;;~��:���9`��i����1��I���
�/�d�̷�ɤ���d�V�������>M�Z���.�ʿ�p�ע%��lG�>tf�$}�      -�_��+Y��lG�f.�{���꿱���M䂿��5���󾌰��O�N�V��S��!�Q����}���i!��g��p�d	:U
�:��;]16;��A;;G;I;9�I;x�I;nvI;LWI;n@I;o/I;�#I;�I;I;�I;	I;�I;�#I;n/I;n@I;HWI;qvI;x�I;6�I;�I;BG;��A;Y16;��;O
�:P	:j񳺎g��i!�}������!�Q�S��V��O�N���������5�M䂿�������{�f.��lG��+Y�      ��7��3�ע%�{��<����ſ
���½\�<����Ͼ����`�3��轻z��}�9�`�Ἓ���z��7}��dt��^:Y+�:��#;��8;��B;sG;q%I;��I;�I;
rI;TI;�=I;t-I;"I;MI;�I;~I;�I;NI;"I;t-I;�=I;TI;rI;�I;��I;n%I;sG;��B;��8;��#;W+�:��^:�dt��7}��z����`��}�9��z����`�3�������Ͼ<��½\�
�����ſ�<��{�ע%��3�      {�����p������ſ%���Ps���1�1r���d���d�}I�ΈŽ��}�`*�KC�� �^��B�~�D�G์ �:��;n);7;;'D;1�G;WHI;��I;��I;�lI;�OI;�:I;+I; I;�I;}I;/I;yI;�I; I;+I;�:I;�OI;�lI;��I;��I;QHI;:�G;'D;7;;l);��;~ �:Gเ�D��B� �^�KC��`*���}�ΈŽ}I��d��d��1r����1��Ps�%����ſ��꿃p����      }߿�$ڿ.�ʿ����
����Ps�PX:����&l¾�ǆ���7����85���Q�����t���75�l�������8�ɼ:��;��.;��=;�EE;�YH;�hI;$�I;��I;(fI;KI;&7I;H(I;�I;�I;�I;{I;�I;�I;�I;H(I;%7I;KI;,fI;��I;$�I;�hI;�YH;�EE;��=;��.;��;�ɼ:��8���m���75��t������Q�85�������7��ǆ�&l¾���PX:��Ps�
�������.�ʿ�$ڿ      ���&��Z���M䂿½\���1�����J˾青�E�N�x��I������V�'�d�Ҽ��|��z��n��Px����&:�P�:��;�W4;Ϡ@;"gF;`�H;�I; �I;2�I;_I;�EI;3I;$%I;GI;�I;�I;�I;�I;�I;GI;#%I;3I;�EI;#_I;2�I;"�I;�I;c�H;%gF;ˠ@;�W4;��;�P�:��&:Px���n���z���|�d�ҼV�'����I���x��E�N�青��J˾�����1�½\�M䂿Z���&��      �,b�Ľ\��>M���5�<��1r��&l¾青�"&W��3�8Sؽ�z��ZG����|I����?���̻��-��
����:��;��&;|9;�C;�dG;KI;A�I;Q�I;RvI;}WI;*@I;�.I;�!I;�I;[I;�I;�I;�I;[I;�I;�!I;�.I;*@I;�WI;SvI;T�I;?�I;KI;�dG;�C;|9;��&;��;��:�
����-���̻��?�|I�����ZG��z��8Sؽ�3�"&W�青�&l¾1r��<����5��>M�Ľ\�      �V������������Ͼ�d���ǆ�E�N��3��c�[����\�3��*C���o���	�숻Z𳺀��9��:�h;O�/;5�=;FE;�2H;�WI;��I;��I;�kI;�OI;":I;�)I;'I;�I;�I;�I;|I;�I;�I;�I;'I;�)I;$:I;�OI;�kI;��I;��I;�WI;�2H;EE;:�=;R�/;h;��:���9\� 숻��	��o�)C��3����\�[���cཱ3�E�N��ǆ��d����Ͼ���������      .l¾(��V������������d���7�x��8Sؽ[���d�D*�dkּ.\����'�,���R�P~��j�:�Z;Σ#;:=7;'�A;�F;V�H;o�I;�I;��I;�`I;�GI;�3I;(%I;uI;�I;UI;N
I;M	I;O
I;XI;�I;wI;'%I;�3I;�GI;�`I;��I;�I;l�I;X�H;�F;+�A;==7;У#;�Z;v�:`~���R�,����'�-\��dkּD*��d�[��8Sؽx����7��d���������V���(��      Gx��s���d�O�N�`�3�}I����H����z����\�C*��ݼJ���0<<��ڻ�V�\dt��&:���:7C;�</;OD=;҈D;��G;�8I;ǘI;��I;tI;'VI;\?I;�-I;e I;�I;\I;�
I;�I;I;�I;�
I;^I;�I;d I;�-I;a?I;/VI;tI;��I;ŘI;�8I;��G;׈D;SD=;�</;DC;���:�&:Ldt��V��ڻ0<<�J����ݼC*���\��z��H������|I�`�3�O�N���d��s�      c.��3�Ȥ�V����ΈŽ85�����ZG�3��dkּI���yC��>�o6}������x9^��:	;)�&;�;8;��A;��F;��H;0yI;��I;��I;1fI;�KI;K7I;|'I;�I;�I;ZI;I;�I;�I;�I;I;ZI;�I;�I;�'I;S7I;�KI;4fI;��I;��I;7yI;��H;��F;��A;�;8;5�&;	;X��:��x9���m6}��>�yC�I���ckּ3��ZG����85��ΈŽ��V��Ȥ��3�      ��Ž5���̷�S���z����}��Q�V�'����)C��-\��0<<��>n��N����&��:&��:�;�'3;��>;�E;cH;^<I;˗I;��I;�vI;�XI;�AI;u/I;�!I;�I;�I;T	I;eI;%I;uI;%I;cI;U	I;�I;�I;�!I;/I;�AI;�XI;�vI;��I;җI;^<I;iH;�E;��>;�'3;�;&��:4��:��L�ຆn���>�0<<�,\��)C�����V�'��Q���}��z��S��̷�5���      ��t��p�.�d�!�Q�}�9�_*����c�Ҽ{I���o���'��ڻp6}�R���9���:Lm�:��;��.;<;�oC;<7G;��H;ҁI;ӜI;҅I;"fI;<LI;�7I;�'I;�I;tI;OI;JI;�I;� I;Q I;� I;�I;KI;PI;uI;�I;�'I;�7I;ELI;"fI;ЅI;ٜI;ӁI;��H;@7G;�oC;<;��.;��;Xm�:��:�9�H��m6}�
�ڻ��'��o�{I��c�Ҽ���_*�~�9�!�Q�/�d��p�      (��c��
����_��KC���t����|���?���	�+���V�$���@���:��:�h;�+;��9;��A;wfF;V�H;q_I;��I;��I;sI;�VI;r@I;�.I;� I;TI;I;�I;kI;P I;�H;�H;~�H;M I;kI;�I;I;[I;� I;�.I;y@I;�VI;�rI;��I;��I;t_I;Z�H;|fF;��A;��9;�+;�h;��:��:��$����V�*����	���?���|��t��JC��`������
�b�      d��T���I��}������ �^��75��z���̻�눻�R�Xdt���x9.��:Tm�:�h;Y�*;ٍ8;��@;ۼE;5(H;d8I;��I;�I;E~I;�`I;�HI;�5I;[&I;tI;2I;�	I;�I;� I;��H;X�H;��H;T�H;��H;� I;�I;�	I;8I;xI;]&I;�5I;�HI;�`I;N~I;�I;��I;h8I;:(H;�E;��@;Ս8;^�*;�h;^m�:6��:��x9@dt��R��눻��̻�z��75��^����~����I��R��      ��?��<<��1��h!��z��B�g���n����-�T�P~���&:P��: ��:��;�+;э8;;�@;�]E;c�G;BI;�I;N�I;5�I;giI;7PI;<I;�+I;�I;nI;OI;)I;qI;��H;��H;R�H;��H;O�H;��H;��H;pI;)I;VI;uI;�I;�+I;<I;4PI;oiI;5�I;L�I;�I;GI;k�G;�]E;:�@;׍8;�+;��;&��:V��:�&:(~��N𳺊�-��n��h���B黶z��h!��1��<<�      N��@��h����g���7}�p�D����>x���
�����9|�:|��:	;�;��.;��9;��@;�]E;f�G;9I;�I;�I;J�I;�pI;VI;�AI;z0I;�"I;�I;�I;�I;�I;��H;^�H;w�H;a�H;��H;^�H;t�H;]�H;��H;�I;�I;�I;�I;�"I;|0I;�AI;�VI;�pI;G�I;�I;�I;?I;j�G;�]E;��@;��9;��.;�;	;���:��:���9�
��Bx�����v�D��7}��g��h���?��      )������P��P񳺴dt��Fเ�8��&:��:��:�Z;>C;.�&;�'3;<;��A;߼E;j�G;:I;U|I;��I;��I;{uI;o[I;FI;�4I;(&I;�I;II;�	I;�I;9�H;��H;6�H;t�H;~�H;�H;x�H;q�H;5�H;��H;7�H;�I;�	I;II;�I;)&I;�4I;	FI;r[I;zuI;��I;ǜI;Y|I;@I;h�G;�E;��A;<;�'3;/�&;EC;�Z;��:��:��&:@�8�F๘dt�j�f��Ǝ��      P�x9Ж�9ث�9<	:��^:� �:�ɼ:�P�:��;�h;Σ#;�</;�;8;��>;�oC;{fF;6(H;II;�I;��I;��I;�wI;m^I;8II;�7I;)I;I;�I;�I;GI;J I;I�H;S�H;:�H;��H;��H;��H;��H;��H;9�H;S�H;E�H;P I;LI;�I;�I;I;)I;�7I;8II;j^I;�wI;��I;��I;�I;II;9(H;|fF;�oC;��>;�;8;�</;ԣ#;�h;��;�P�:�ɼ:| �:�^:H	:0��9�9      ���:c��:���:i
�:I+�:��;��;��;��&;P�/;==7;MD=;��A;�E;=7G;Z�H;g8I;�I;�I;��I;�wI;�_I;�JI;�9I;�*I;�I;2I;9I;I;9I;��H;��H;�H;<�H;��H;�H;��H;�H;��H;=�H;�H;��H;�H;<I;I;<I;2I;�I;�*I;�9I;�JI;�_I;�wI;��I;	�I;�I;l8I;[�H;@7G;�E;��A;SD=;@=7;O�/;��&;��;��;��;+�:W
�:���:O��:      b�;̻;;��;��#;t);��.;�W4;"|9;9�=;.�A;وD;��F;nH;��H;w_I;��I;R�I;J�I;}uI;m^I;�JI;$:I; ,I;5 I;~I;MI;�I;!I;��H;��H;4�H;�H;k�H;c�H;��H;U�H;��H;c�H;n�H;�H;3�H;�H;��H;I;�I;MI;�I;: I;,I;!:I;�JI;q^I;~uI;N�I;N�I;I;x_I;��H;kH;��F;ۈD;4�A;6�=;!|9;�W4;��.;p);��#;��;;��;      ��2;X%3;�U4;S16;��8;7;;��=;ˠ@;�C;EE;�F;��G;��H;^<I;сI;��I;�I;6�I;�pI;m[I;6II;�9I;,I;� I;I;I;QI;�I;H�H;d�H;\�H;*�H;:�H;��H;��H;a�H;�H;[�H;��H;��H;;�H;(�H;a�H;d�H;G�H;�I;OI;I;I;� I;,I;�9I;6II;k[I;�pI;2�I;�I;��I;ҁI;]<I;��H;��G;�F;FE;�C;Р@;��=;7;;��8;U16;�U4;Q%3;      Q@@;Ep@;��@;��A;��B;3D;�EE;%gF;�dG;�2H;Z�H;�8I;2yI;՗I;ۜI;��I;R~I;siI;�VI;FI;�7I;�*I;; I;#I;ZI;�I;=I;��H;��H;��H;�H;"�H;��H;o�H;��H;%�H;��H;�H;��H;r�H;��H;�H; �H;��H;��H;��H;9I;�I;^I;!I;: I;�*I;�7I;FI;�VI;qiI;U~I;��I;ۜI;ԗI;3yI;�8I;^�H;�2H;�dG;#gF;�EE;)D;��B;��A;��@;Cp@;      \fF;�yF;ӱF;5G;�rG;>�G;�YH;l�H;KI;�WI;q�I;ΘI;��I;��I;҅I;sI;�`I;8PI;�AI;�4I;)I;�I;~I;!I;�I;PI;��H;��H;��H;T�H;-�H;h�H;�H;-�H;t�H;�H;�H;�H;q�H;-�H;�H;c�H;0�H;U�H;��H; �H;��H;VI;�I;I;|I;�I;	)I;�4I;�AI;4PI;�`I;sI;҅I;��I;��I;̘I;y�I;�WI;NI;k�H;�YH;3�G;sG;GG;ӱF;�yF;      G�H;��H;,�H; I;d%I;THI;�hI;�I;A�I;��I;�I;��I;�I;�vI;fI;�VI;�HI;<I;~0I;,&I;I;1I;NI;WI;9I;��H;�H;��H;h�H;2�H;l�H;��H;��H;�H;j�H;�H;�H;�H;h�H;	�H;��H;��H;o�H;2�H;f�H;��H;��H;��H;>I;SI;OI;5I;I;)&I;~0I;<I;�HI;�VI;fI;�vI;�I;��I;�I;��I;?�I;�I;�hI;NHI;y%I;�I;+�H;��H;      ��I; �I;׎I;=�I;��I;��I;+�I;�I;S�I;��I;��I;tI;0fI;�XI;<LI;v@I;�5I;�+I;�"I;�I;�I;6I;�I;�I;��H;��H;��H;^�H;E�H;\�H;��H;��H;��H;��H;��H;B�H;'�H;>�H;��H; �H;��H;��H;��H;^�H;E�H;a�H;��H;��H;��H;�I;�I;9I;�I;�I;�"I;�+I;�5I;w@I;>LI;�XI;0fI;tI;��I;��I;S�I;�I;+�I;��I;��I;@�I;ՎI;�I;      Q�I;ޛI;��I;��I;ڔI;��I;��I;7�I;LvI;�kI;�`I;/VI;�KI;�AI;�7I;�.I;b&I;�I;�I;LI;�I;zI;I;G�H;��H;��H;_�H;E�H;_�H;��H;��H;��H;��H;&�H;��H;��H;O�H;�H;��H;'�H;��H;��H;��H;��H;_�H;H�H;_�H;��H;��H;D�H; I;{I;�I;II;�I;�I;b&I;�.I;�7I;�AI;�KI;/VI;�`I;�kI;MvI;5�I;��I;��I;�I;��I;��I;ٛI;      !|I;�{I;�yI;hvI;rI;�lI;)fI;#_I;�WI;�OI;�GI;g?I;R7I;�/I;�'I;� I;{I;kI;�I;�	I;NI;4I;��H;b�H;��H;J�H;/�H;^�H;��H;��H;��H;��H;��H;��H;�H;��H;��H;��H;�H;��H;��H;��H;��H;��H;��H;a�H;-�H;Q�H;��H;`�H;��H;9I;JI;�	I;�I;kI;{I;� I;�'I;}/I;R7I;d?I;�GI;�OI;WI;_I;,fI;�lI;rI;qvI;�yI;�{I;      �[I;a[I;�YI;RWI;TI;�OI;KI;�EI;0@I;):I;�3I;�-I;�'I;�!I;�I;\I;=I;TI;�I;�I;V I;��H;��H;]�H;�H;)�H;l�H;��H;��H;��H;~�H;��H;V�H;��H;x�H;\�H;U�H;Y�H;u�H;��H;Z�H;��H;��H;��H;��H;��H;m�H;/�H; �H;]�H;�H;�H;S I;�I;�I;TI;=I;]I;�I;�!I;�'I;�-I;�3I;):I;0@I;�EI;%KI;�OI;TI;UWI;�YI;a[I;      �CI;VCI;7BI;b@I;�=I;�:I;"7I;
3I;�.I;�)I;'%I;k I;�I;�I;wI;I;
I;,I;�I;>�H;P�H;��H;0�H;&�H;�H;[�H;��H;��H;��H;��H;��H;D�H;��H;N�H;�H;��H;��H;��H;�H;Q�H;��H;B�H;��H;��H;��H;��H;��H;a�H;#�H;!�H;6�H;��H;L�H;:�H;�I;/I;
I;I;zI;�I;�I;h I;.%I;�)I;�.I;3I;,7I;�:I;�=I;k@I;?BI;VCI;      2I;�1I;�0I;n/I;p-I;+I;A(I; %I;�!I;!I;wI;�I;�I;�I;PI;�I;�I;tI;��H;��H;_�H;�H;�H;6�H;��H;�H;��H;��H;��H;��H;S�H;��H;3�H;��H;��H;~�H;o�H;�H;��H;��H;5�H;��H;S�H;��H;��H;��H;��H;�H;��H;7�H;	�H;�H;X�H;��H;��H;tI;�I;�I;SI;�I;�I;�I;{I;!I;�!I;%I;E(I;+I;v-I;m/I;�0I;�1I;      �%I;P%I;�$I;�#I;"I; I;�I;II;�I;�I;�I;eI;aI;\	I;OI;oI;� I;��H;c�H;<�H;A�H;<�H;g�H;��H;k�H;#�H;�H; �H;'�H;��H;��H;Q�H;��H;��H;^�H;8�H;&�H;8�H;\�H;��H;��H;R�H;��H;��H;#�H;��H;�H;(�H;l�H;��H;m�H;<�H;=�H;5�H;a�H;��H;� I;oI;OI;[	I;`I;dI;�I;�I;�I;GI;�I; I;"I;�#I;�$I;\%I;      QI;6I;�I;�I;VI;�I;�I;�I;]I;�I;aI;�
I;I;oI;�I;T I;��H;��H;x�H;x�H;��H;��H;]�H;��H;��H;f�H;b�H;��H;��H;�H;n�H;�H;��H;\�H;�H;�H;�H;�H;�H;^�H;��H;�H;p�H;
�H;��H;��H;c�H;i�H;��H;��H;b�H;��H;��H;q�H;w�H;��H;��H;V I;�I;mI;I;�
I;cI;�I;]I;�I;�I;�I;TI;�I;�I;8I;      �I;]I;�I;	I;�I;sI;�I;�I;�I;�I;T
I;I;�I;*I;� I;~�H;X�H;N�H;b�H;~�H;��H;�H;��H;O�H;�H;�H;�H;?�H;��H;��H;X�H;��H;��H;9�H;	�H;��H;��H;��H;�H;=�H;��H;��H;V�H;��H;��H;<�H;�H;�H;�H;P�H;��H;�H;��H;x�H;a�H;Q�H;[�H;��H;� I;*I;�I; I;X
I;�I;�I;�I;�I;uI;�I;
I;�I;kI;      9I;�I;�I;�I;uI;%I;{I;�I;�I;{I;W	I;I;�I;~I;X I;�H;��H;��H;��H;!�H;��H;��H;Q�H;��H;��H;�H;�H;*�H;V�H;��H;N�H;��H;p�H;!�H;�H;��H;��H;��H;�H;#�H;s�H;��H;N�H;��H;O�H;&�H;�H;	�H;��H;��H;T�H;��H;��H;�H;��H;��H;��H;�H;Z I;I;�I;I;Z	I;{I;�I;�I;�I;%I;sI;�I;�I;
I;      �I;`I;�I;I;�I;vI;�I;�I;�I;�I;R
I;I;�I;*I;� I;~�H;X�H;N�H;b�H;~�H;��H;�H;��H;O�H;�H;�H;�H;?�H;��H;��H;V�H;��H;��H;9�H;�H;��H;��H;��H;�H;<�H;��H;��H;U�H;��H;��H;;�H;�H;�H;�H;O�H;��H;
�H;��H;x�H;a�H;Q�H;Z�H;��H;� I;(I;�I; I;V
I;�I;�I;�I;�I;uI;�I;I;�I;gI;      II;9I;�I;�I;VI;�I;�I;�I;\I;�I;_I;�
I;I;lI;�I;S I;��H;��H;x�H;x�H;��H;��H;]�H;��H;��H;d�H;c�H;��H;��H;�H;n�H;�H;��H;\�H;�H;�H;�H;�H;�H;\�H;��H;�H;m�H;�H;��H;��H;c�H;i�H;��H;��H;`�H;��H;��H;q�H;w�H;��H;��H;V I;�I;mI;I;�
I;bI;�I;\I;�I;�I;�I;VI;�I;�I;;I;      �%I;Q%I;�$I;�#I;"I; I;�I;LI;�I;�I;�I;dI;`I;[	I;OI;nI;� I;��H;c�H;;�H;B�H;=�H;g�H;��H;o�H;%�H;�H;�H;*�H;��H;��H;R�H;��H;��H;_�H;6�H;&�H;9�H;[�H;��H;��H;O�H;��H;}�H;"�H;��H;�H;&�H;l�H;��H;k�H;;�H;:�H;6�H;c�H;��H;� I;qI;QI;\	I;`I;dI;�I;�I;�I;KI;�I; I;"I;�#I;�$I;S%I;      2I;�1I;�0I;k/I;o-I;+I;?(I;$%I;�!I;I;tI;�I;�I;�I;SI;�I;�I;tI;��H;��H;_�H;�H;�H;7�H;��H;�H;��H;��H;��H; �H;S�H;��H;3�H;��H;��H;�H;o�H;�H;��H;��H;2�H;��H;R�H;��H;��H;��H;��H;�H;��H;3�H;	�H;�H;U�H;��H;��H;sI;�I;�I;SI;�I;�I;�I;xI; I;�!I; %I;H(I;+I;s-I;r/I;�0I;�1I;      �CI;ZCI;(BI;b@I;�=I;�:I;)7I;3I;�.I;�)I;+%I;k I;�I;�I;wI;I;
I;/I;�I;=�H;S�H;��H;2�H;$�H;#�H;^�H;��H;��H;��H;��H;��H;D�H;��H;N�H;�H;��H;��H;��H;�H;O�H;��H;D�H;��H;��H;��H;��H;��H;^�H;�H;�H;7�H;��H;J�H;:�H;�I;,I;
I;I;xI;�I;�I;k I;.%I;�)I;�.I;3I;)7I;�:I;�=I;n@I;/BI;UCI;      �[I;a[I;�YI;NWI;TI;�OI;KI;�EI;-@I;':I;�3I;�-I;�'I;�!I;�I;\I;=I;VI;�I;�I;W I;�H;��H;]�H; �H;)�H;j�H;��H;��H;��H;��H;��H;Y�H;��H;z�H;Y�H;T�H;\�H;u�H;��H;Z�H;��H;��H;��H;��H;��H;j�H;,�H;�H;Z�H;�H;�H;P I;�I;�I;SI;?I;\I;�I;�!I;�'I;�-I;�3I;(:I;0@I;�EI;#KI;�OI;TI;WWI;�YI;c[I;      )|I;�{I;�yI;rvI;�qI;�lI;(fI;&_I;�WI;�OI;�GI;d?I;O7I;}/I;�'I;� I;zI;nI;�I;�	I;PI;8I;��H;`�H;��H;J�H;/�H;_�H;��H;��H;��H;��H;��H;��H;�H;��H;��H;��H;�H;��H;��H;��H;��H;��H;��H;^�H;-�H;N�H;��H;]�H;��H;8I;JI;�	I;�I;iI;zI;� I;�'I;/I;P7I;a?I;�GI;�OI;}WI;#_I;,fI;�lI;rI;yvI;�yI;�{I;      Z�I;ܛI;��I;��I;̔I;��I;��I;5�I;RvI;�kI;�`I;.VI;�KI;�AI;�7I;�.I;`&I;�I;�I;II;�I;{I;I;G�H;��H;��H;_�H;G�H;c�H;��H;��H;��H;��H;'�H;��H;��H;P�H;��H;��H;&�H;��H;��H;��H;��H;\�H;D�H;a�H;��H;��H;A�H;!I;|I;�I;II;�I;�I;`&I;�.I;�7I;�AI;�KI;+VI;�`I;�kI;OvI;7�I;��I;��I;ܔI;��I;��I;ԛI;      ��I;�I;ȎI;=�I;��I;��I;-�I;&�I;Q�I;��I;��I;tI;0fI;�XI;?LI;w@I;�5I;�+I;�"I;�I;�I;9I;�I;�I;��H;��H;��H;^�H;K�H;\�H;��H;��H;��H;��H;��H;?�H;)�H;?�H;��H; �H;��H;��H;��H;^�H;D�H;\�H;��H;��H;��H;�I;�I;8I;�I;�I;�"I;�+I;�5I;w@I;?LI;�XI;0fI;tI;��I;��I;P�I;�I;-�I;��I;��I;@�I;ӎI;�I;      9�H;��H;*�H;I;q%I;WHI;�hI;�I;A�I;��I;�I;��I;�I;�vI;fI;�VI;�HI;<I;}0I;(&I;I;5I;MI;ZI;;I;��H; �H;��H;j�H;2�H;m�H;��H;��H;�H;l�H;�H;�H;�H;h�H;	�H;��H;��H;p�H;3�H;f�H;��H;�H;��H;;I;SI;RI;4I;I;+&I;�0I;<I;�HI;�VI;fI;�vI;��I;��I;�I;��I;?�I;�I;�hI;QHI;x%I;I;+�H;��H;      TfF;�yF;ڱF;6G;sG;E�G;�YH;n�H;MI;�WI;r�I;ϘI;��I;��I;ԅI;sI;�`I;:PI;�AI;�4I;)I;�I;|I;!I;�I;PI;��H;�H;��H;T�H;0�H;i�H;�H;-�H;u�H;�H;�H;�H;p�H;,�H;�H;h�H;3�H;U�H;��H;��H;��H;RI;�I;I;I;�I;)I;�4I;�AI;5PI;�`I;sI;ՅI;��I;��I;ʘI;u�I;�WI;FI;e�H;�YH;3�G;sG;9G;��F;�yF;      N@@;@p@;��@;��A;��B;5D;�EE;"gF;�dG;�2H;Z�H;�8I;0yI;їI;ݜI;��I;S~I;viI;�VI;FI;�7I;�*I;: I;#I;`I;�I;9I;��H;��H;��H;�H;%�H;��H;p�H;��H;"�H;��H;"�H;��H;p�H;��H;#�H;!�H;��H;��H;��H;=I;�I;\I;I;< I;�*I;�7I;FI;�VI;oiI;S~I;��I;ܜI;їI;2yI;�8I;Z�H;�2H;�dG;#gF;�EE;'D;��B;��A;~�@;Ap@;      ��2;>%3;�U4;a16;��8;'7;;��=;͠@;�C;CE;�F;��G;��H;[<I;ӁI;��I;�I;6�I;�pI;m[I;9II;�9I;,I;� I;I;I;OI;�I;K�H;c�H;`�H;.�H;;�H;��H;��H;]�H;�H;`�H;��H;��H;=�H;-�H;c�H;d�H;G�H;�I;SI;I;I;� I;,I;�9I;8II;m[I;�pI;1�I;�I;��I;сI;[<I;��H;��G;�F;CE;�C;Ƞ@;��=;7;;��8;u16;�U4;)%3;      T�;ɻ;;�;��#;p);��.;�W4;(|9;:�=;+�A;ۈD;��F;mH;��H;y_I;��I;R�I;J�I;}uI;p^I;�JI; :I; ,I;; I;{I;KI;�I;%I;��H;�H;9�H;�H;m�H;d�H;��H;W�H;��H;`�H;j�H;�H;7�H;�H;��H;I;�I;QI;|I;7 I;,I;":I;�JI;p^I;~uI;N�I;K�I;I;x_I;��H;jH;��F;وD;.�A;9�=;$|9;�W4;��.;p);��#;�;;��;      z��:]��:���:[
�:K+�:��;��;��;��&;O�/;?=7;VD=;��A;�E;A7G;]�H;h8I;�I;�I;��I;�wI;�_I;�JI;�9I;�*I;�I;2I;=I;�I;9I;�H;��H;�H;<�H;��H;�H;��H;�H;��H;;�H;�H;��H;�H;<I;I;<I;6I;�I;�*I;�9I;�JI;�_I;�wI;��I;�I;�I;h8I;Z�H;@7G;�E;��A;QD=;@=7;M�/;��&;��;��;z�;y+�:C
�:���:G��:      ��x9x��9@��9P	:��^:� �:�ɼ:�P�:��;~h;ѣ#;�</;�;8;��>;�oC;~fF;9(H;II;�I;��I;��I;�wI;k^I;8II;�7I;)I;I;�I;�I;GI;O I;L�H;T�H;=�H;��H;��H;��H;��H;��H;9�H;T�H;I�H;P I;JI;�I;�I;	I;)I;�7I;8II;k^I;�wI;��I;��I;�I;EI;:(H;~fF;�oC;��>;�;8;�</;ӣ#;�h;��;�P�:�ɼ:� �:$�^:T	:���9 ��9      ������Z��L��dt��F�`�8��&: ��:��:�Z;BC;/�&;�'3;<;��A;�E;j�G;<I;X|I;ŜI;��I;{uI;o[I;FI;~4I;%&I;�I;LI;�	I;�I;;�H;��H;8�H;t�H;z�H;�H;|�H;q�H;4�H;��H;:�H;�I;�	I;II;�I;+&I;�4I;FI;r[I;}uI;��I;ÜI;X|I;=I;h�G;�E;��A;<;�'3;/�&;?C;�Z;��:��:��&:@�8G๘dt�b�^�຺���      N��@��h����g���7}�o�D����>x��h
�����9|�:���:	;�;��.;��9;��@;�]E;g�G;=I;�I;�I;J�I;�pI;�VI;�AI;z0I;�"I;�I;�I;�I;�I;��H;`�H;w�H;a�H;��H;a�H;t�H;]�H;��H;�I;�I;�I;�I;�"I;|0I;�AI;�VI;�pI;H�I;�I;�I;=I;g�G;�]E;��@;��9;��.;�;	;���:|�:���9x
��8x�����r�D��7}��g��k���=��      ��?��<<��1��h!��z��B�f���n����-�R�0~���&:R��:"��:��;�+;Ս8;;�@;�]E;h�G;FI;�I;Q�I;5�I;oiI;7PI;<I;�+I;�I;nI;TI;.I;sI;��H;��H;Q�H;��H;T�H;��H;��H;sI;+I;TI;oI;�I;�+I;<I;4PI;jiI;5�I;N�I;�I;CI;h�G;�]E;9�@;ҍ8;�+;��;"��:R��:�&:(~��R𳺋�-��n��f���B黶z��h!�
�1��<<�      d��T���I��}�������^��75��z���̻�눻�R�<dt���x90��:`m�:�h;^�*;؍8;��@;�E;:(H;h8I;��I;�I;Q~I;�`I;�HI;�5I;_&I;uI;8I;�	I;�I;� I;��H;W�H;��H;W�H;��H;� I;�I;�	I;6I;tI;]&I;�5I;�HI;�`I;H~I;�I;��I;g8I;3(H;�E;��@;Ս8;\�*;�h;Zm�:4��:��x9Ddt��R��눻��̻�z��75��^����}����I��S��      (��c��
����_��JC���t����|���?���	�*���V�"�������:��:�h;�+;��9;��A;~fF;[�H;w_I;��I;��I;sI;�VI;s@I;�.I;� I;YI;I;�I;nI;Q I;~�H;�H;�H;M I;jI;�I;I;VI;� I;�.I;u@I;�VI;�rI;��I;��I;u_I;X�H;tfF;��A;��9;�+;�h;��:��:��$����V�+����	���?���|��t��JC��`������
�c�      ��t��p�/�d� �Q�}�9�_*����c�Ҽ{I���o���'�
�ڻm6}�F��`9���:Tm�:��;��.;<;�oC;@7G;��H;ՁI;ٜI;҅I;fI;>LI;�7I;�'I;�I;wI;PI;MI;�I;� I;Q I;� I;�I;KI;OI;tI;�I;�'I;�7I;?LI;fI;хI;ҜI;ӁI;��H;?7G;�oC;<;��.;��;Xm�:��:�9�H��o6}��ڻ��'��o�{I��c�Ҽ���_*�~�9�!�Q�/�d��p�      ��Ž5���̷�R���z����}��Q�U�'����)C��,\��/<<��>n��>�຀�.��:(��:�;�'3;��>;�E;jH;d<I;ԗI;��I;�vI;�XI;�AI;y/I;�!I;�I;�I;T	I;cI;#I;uI;&I;aI;U	I;�I;�I;�!I;|/I;�AI;�XI;�vI;��I;ʗI;a<I;kH;�E;��>;�'3;�;&��:0��:��H�ຆn���>�0<<�,\��)C�����U�'��Q���}��z��S��̷�5���      c.��3�Ȥ�V����ΈŽ85�����ZG�3��ckּI���yC��>�h6}������x9\��:
	;0�&;�;8;��A;��F;��H;7yI;��I;�I;0fI;�KI;P7I;�'I;�I;�I;]I;I;�I;�I;�I;I;ZI;�I;�I;�'I;O7I;�KI;1fI;�I;��I;0yI;��H;��F;��A;�;8;3�&;	;V��:��x9���l6}��>�yC�I���dkּ3��ZG����85��ΈŽ��V��Ȥ��3�      Gx��s���d�O�N�`�3�|I����H����z����\�C*��ݼI���0<<�
�ڻ�V�Pdt��&:���:?C;�</;QD=;ڈD;��G;�8I;ȘI;��I;tI;+VI;]?I;�-I;e I;�I;`I;�
I;�I;I;�I;�
I;]I;�I;d I;�-I;^?I;,VI;tI;��I;ǘI;�8I;��G;وD;OD=;�</;AC;|��:�&:Xdt��V��ڻ0<<�J����ݼC*���\��z��H������|I�`�3�O�N���d��s�      .l¾(��V������������d���7�x��8Sؽ[���d�C*�dkּ-\����'�,���R�h~��r�:�Z;գ#;==7;-�A;�F;[�H;q�I;�I;��I;�`I;�GI;�3I;*%I;wI;�I;WI;O
I;N	I;O
I;WI;�I;wI;'%I;�3I;�GI;�`I;��I;�I;o�I;T�H;�F;+�A;9=7;ɣ#;�Z;j�:`~���R�,����'�-\��dkּD*��d�[��8Sؽx����7��d���������V���(��      �V������������Ͼ�d���ǆ�E�N��3��c�[����\�3��)C���o���	��눻\𳺠��9��:�h;R�/;:�=;JE;�2H;�WI;��I;��I;�kI;�OI;':I;�)I;'I;�I;�I;�I;|I;�I;�I;�I;'I;�)I;%:I;�OI;�kI;��I;��I;�WI;�2H;FE;<�=;O�/;}h;��:x��9\� 숻��	��o�)C��3����\�[���cཱ3�E�N��ǆ��d����Ͼ���������      �,b�Ľ\��>M���5�<��1r��&l¾青�"&W��3�8Sؽ�z��ZG����|I����?���̻��-��
����:��;��&;|9;�C;�dG;KI;@�I;P�I;SvI;WI;.@I;�.I;�!I;�I;XI;�I;�I;�I;YI;�I;�!I;�.I;,@I;}WI;RvI;Q�I;?�I;NI;�dG;�C;|9;��&;��;��:�
����-���̻��?�|I�����ZG��z��8Sؽ�3�"&W�青�&l¾1r��<����5��>M�Ľ\�      ���&��Z���M䂿½\���1�����J˾青�E�N�x��I������V�'�d�Ҽ��|��z��n��Jx����&:�P�:��;�W4;Ҡ@;(gF;`�H;�I;�I;1�I;_I;�EI;	3I;$%I;GI;�I;�I;�I;�I;�I;GI;$%I;3I;�EI;!_I;1�I; �I;�I;c�H;"gF;Р@;�W4;��;�P�:��&:Rx���n���z���|�d�ҼV�'����I���x��E�N�青��J˾�����1�½\�M䂿Z���&��      }߿�$ڿ.�ʿ����
����Ps�PX:����&l¾�ǆ���7����85���Q�����t���75�l�������8�ɼ:��;��.;��=;�EE;�YH;�hI;#�I;��I;)fI;KI;&7I;I(I;�I;�I;�I;zI;�I;�I;�I;H(I;&7I;KI;+fI;��I;&�I;�hI;�YH;�EE;��=;��.;��;�ɼ:��8���l���75��t������Q�85�������7��ǆ�&l¾���PX:��Ps�
�������.�ʿ�$ڿ      {�����p������ſ%���Ps���1�1r���d���d�}I�ΈŽ��}�_*�KC���^��B�}�D��F๐ �:��;p);7;;)D;1�G;UHI;��I;��I;�lI;�OI;�:I;+I; I;�I;|I;/I;|I;�I; I;+I;�:I;�OI;�lI;��I;��I;THI;:�G;'D;7;;n);��;� �:Gเ�D��B��^�KC��`*���}�ΈŽ}I��d��d��1r����1��Ps�%����ſ��꿃p����      ��7��3�ע%�{��<����ſ
���½\�<����Ͼ����`�3��轻z��}�9�_�Ἓ���z��7}��dt��^:_+�:��#;��8;��B;	sG;o%I;��I;�I;	rI;TI;�=I;s-I;"I;HI;�I;}I;�I;KI;"I;s-I;�=I;TI;rI;�I;��I;r%I;sG;��B;��8;��#;]+�:��^:�dt��7}��z����`��}�9��z����`�3�������Ͼ<��½\�
�����ſ�<��{�ע%��3�      -�_��+Y��lG�f.�{���꿱���M䂿��5���󾌰��O�N�V��S��!�Q����}���i!��g��h�l	:W
�:��;]16;��A;8G;�I;8�I;x�I;lvI;NWI;l@I;m/I;�#I;�I;I;�I;
I;�I;�#I;o/I;o@I;KWI;rvI;x�I;9�I; I;CG;��A;\16;��;Q
�:P	:j񳺎g��i!�}������!�Q�S��V��O�N���������5�M䂿�������{�f.��lG��+Y�      Ѭ��$}�>tf��lG�ע%��p�/�ʿZ����>M����V�����d�ɤ�̷�/�d��
��I���1�h���^�ຠ��9���:;�U4;��@;ұF;2�H;ݎI;��I;�yI;�YI;<BI;�0I;�$I;�I;�I;�I;�I;�I;�$I;�0I;<BI;�YI;�yI;��I;��I;4�H;ܱF;��@;�U4;;~��:���9Z��i����1��I���
�/�d�̷�ɤ���d�V�������>M�Z���/�ʿ�p�ע%��lG�>tf�$}�      S���E���$}��+Y��3�����$ڿ&��Ľ\����(���s��3�5����p�c�U���<<�9������p��9I��:ϻ;R%3;Ep@;�yF;��H;��I;�I;�{I;O[I;RCI;�1I;U%I;#I;ZI;I;WI;#I;U%I;�1I;SCI;K[I;�{I;�I;��I;��H;�yF;Dp@;N%3;Ȼ;=��:8��9����<���<<�U��c��p�5����3��s�(�����Ľ\�&���$ڿ����3��+Y�$}�F���      �Aq���i���U�G:�@�����;���v���{A�d5�� ��~^Z�����A���]�����d��K",��5����Ѻ ��9���:�;^Y4;H�@;LVF;��H;�GI;�bI;OI;!:I;�)I;$I;�I;�I;�I;�I;�I;�I;�I;"I;�)I;:I;$OI;�bI;�GI;��H;XVF;H�@;XY4;�;���: ��9��Ѻ�5��K",��d������]��A�����~^Z�� ��d5�{A�v���;�������@�G:���U���i�      ��i���b�Z�O�.5�2i�������������q<�����e��`
V�GE	�!���IY�j9�E�����(��R��
�ȺX�:Q��:�;A�4;>�@;hF;��H;II;|bI;�NI;�9I;�)I;�I;_I;�I;dI;^I;`I;�I;_I;�I;�)I;�9I;�NI;|bI;II;��H;'hF;>�@;<�4;ڔ;I��:@�:�Ⱥ�R����(�E���j9��IY�!��GE	�`
V��e������q<������������2i�.5�Z�O���b�      ��U�Z�O�H-?�.�'���M�ῴ欿`�{�fa/���뾝���I����d���ZN�\5������=H�d ��l���|�":��:}�;��5;�`A;��F;L�H;MI;�aI;�MI;�8I;�(I;FI;�I;=I;I;I;I;=I;�I;FI;�(I;�8I;�MI;�aI;MI;L�H;��F;�`A;��5;s�;��:h�":d���g ��=H�����\5���ZN�d������I�������fa/�`�{��欿M����.�'�H-?�Z�O�      G:�.5�.�'��������jȿ���k$_���W�Ҿܕ���6�����*���`=�>�漮)��JG�(6�����$�Q:��:�/";
�7;^&B;��F;��H;�RI;�`I;zKI;7I;�'I;AI;I;�I;uI;t
I;oI;�I;I;AI;�'I;7I;KI;�`I;�RI;��H;��F;]&B;�7;�/";��:�Q:���)6��JG��)��>���`=��*������6�ܕ��W�Ҿ��k$_����jȿ�������.�'�.5�      @�2i�������I�ѿk��� ���q<��:��a����q����Wн罅���'�Ub̼�zl��.��N�X�h����:��;ю&;ȫ9;#C;<MG;��H;9YI;�^I;�HI;�4I;�%I;�I;I;�I;�
I;�	I;�
I;�I;
I;�I;�%I;�4I;�HI;�^I;:YI;��H;CMG;!C;«9;ˎ&;��;��:`��Q�X��.���zl�Ub̼��'�罅��Wн����q��a���:��q<� ��k���I�ѿ������2i�      �������M��jȿk���������O���z]׾{����I�����A��>�d�n�~֮�RH��jλP�$��(�q��:FN;��+;�<;�3D;��G;�I;�^I;l[I;�DI;"2I;�#I;II;�I;bI;�	I;�I;�	I;aI;�I;GI;�#I;!2I;�DI;l[I;�^I;�I;��G;�3D;�<;��+;FN;c��:�(�S�$��jλRH�֮�n�>�d��A������I�{���z]׾����O�����k���jȿM�Ῡ��      ;��������欿��� ����O��x����� ���l���"��ܽ���`=����w���k"�-R��Dۺ���9�?�:_L;��0;��>;�ME;K#H;�%I;�aI;�VI;�@I;�.I;B!I;DI;I;I;SI;�I;PI;I;I;AI;?!I;�.I;�@I; WI;�aI;�%I;P#H;�ME;��>;}�0;[L;|?�:���9Fۺ.R���k"�w������`=����ܽ��"��l�� ����뾁x���O� ������欿����      v�������`�{�k$_��q<�������}��w��	�6�����!���h����ⷾ�� d��.���^e�I[���Z:`��:�, ;��5;�A;�VF;��H;�@I;pbI;�QI;�;I;>+I;qI;I;:I;�	I;�I;2I;�I;�	I;<I;I;mI;=+I;�;I;�QI;ubI;�@I;��H;�VF;�A;��5;�, ;T��:��Z:I[��^e�~.��� d�ⷾ�����h�!������	�6�w���}��������q<�k$_�`�{�����      {A��q<�fa/����:�z]׾� ��w��>�DE	�����ڽ����3�_�꼚���",��W��a��@Q�w��:�M
;�f);��:;'@C;�?G;R�H;KTI;�_I;)KI;�6I;O'I;kI;�I;AI;�I;tI;�I;qI;�I;AI;�I;jI;P'I;�6I;,KI;�_I;GTI;R�H;�?G;%@C;��:;�f);�M
;���: Q�d���W��",�����^�꼘�3�ڽ������DE	�>�w��� ��z]׾�:���fa/��q<�      d5�������W�Ҿ�a��{����l�	�6�DE	���Ƚk���aG����f֮��W����q�k�2���c,:���:��;��1;?�>;@E;"�G;I;)_I;CZI;7DI;�1I;2#I;HI;I;
I;I;�I;%I;�I;I;
I; I;CI;3#I;�1I;:DI;GZI;&_I;I;&�G;=E;B�>;��1;��;���:�c,:6��m�k�����W�e֮�����aG�k����ȽDE	�	�6��l�{����a��W�Ҿ������      � ���e�����ܕ����q��I���"���������k���ZN�[�"¼P�y��$��Q���� � hX���:0;%�&;�w8;n B;��F;ԐH;W@I;�aI;lRI;=I;,I;�I;�I;^I;�I;:I; I;hI;!I;:I;�I;^I;�I;�I;,I;=I;pRI;�aI;T@I;ؐH;��F;q B;�w8;#�&;#0;��: pX��� ��Q���$�P�y�"¼[��ZN�k������������"��I���q�ܕ������e��      ~^Z�`
V��I��6�������ܽ!��ڽ���aG�[�
�ȼ�)��}�(�j��NG5������Z:�:S;'1;��=;��D;/�G;��H;�XI;^I;II;�5I;�&I;�I;�I;�
I;�I;NI;d I;��H;d I;NI;�I;�
I;�I;�I;�&I;�5I;�II;^I;�XI;��H;/�G;��D;��=;'1;S;�:��Z:���KG5�j��|�(��)��
�ȼ[��aG�ڽ��!���ܽ������6��I�`
V�      ���GE	��������Wн�A�����h���3����!¼�)��2x/��һv�X�v#����9L��:�>;,f);g`9;^&B;��F;g}H;�6I;PaI;�UI;a@I;�.I;� I;HI;)I;�I;OI;S I;��H;��H;��H;Q I;OI;�I;'I;MI;!I;�.I;d@I;�UI;NaI;�6I;i}H;��F;a&B;e`9;7f);�>;F��:��9p#��s�X��һ2x/��)��!¼�����3��h��󑽢A���Wн��콺��GE	�      �A��!��c���*��潅�?�d��`=����^��e֮�O�y�~�(��һ�]e�򄮺@�f9���:6�;D1";�4;�m?;�E;��G;e�H;�WI;�^I;KI;r7I;�'I;�I;%I;�
I;&I;I;n�H;��H;<�H;��H;m�H;I;#I;�
I;)I;�I;�'I;v7I;KI;|^I;�WI;g�H;��G;�E;�m?; �4;H1";4�;���:`�f9ꄮ��]e��һ|�(�N�y�e֮�]�꼗���`=�>�d�罅��*��c��!��      �]��IY��ZN��`=���'�n����᷾������W��$�k��y�X�􄮺�9v��:W��:o�;��0;��<;Q�C; G;��H;�?I;%aI;�TI;>@I;/I;W!I;�I;I;{I;�I;��H;~�H;�H;��H;�H;}�H;��H;�I;xI;I;�I;[!I;/I;A@I;�TI;,aI;�?I;��H;%G;R�C;��<;��0;i�;_��:v��:9ꄮ�u�X�h���$��W�����᷾����m���'��`=��ZN��IY�      ���j9�[5��<��Ub̼~֮�v��� d�",�����Q��RG5�|#��`�f9t��:��:�;��-;��:;�KB;8VF;KH;�I;�\I;\I;�HI;6I;'I;I;�I;
I;CI;��H;��H;��H;[�H;��H;Z�H;��H;��H;��H;BI;
I;�I;I;"'I;6I;�HI;#\I;�\I;�I;KH;<VF;�KB;��:;��-;�;��:|��:`�f9|#��KG5��Q�����",�� d�v��}֮�Vb̼=��\5��i9�      �d��D��������)���zl�RH��k"�y.���W��i�k��� ������9���:c��:�;�-;̫9;BaA;��E;%�G;t�H;�RI;`I;�OI;�<I;�,I;�I;/I;I;{I;UI;��H;��H;��H;��H;c�H;��H;��H;��H;��H;UI;I;I;1I;�I;�,I;�<I;�OI;`I;�RI;y�H;(�G;��E;GaA;ȫ9;�-;�;g��:���:��9����� �g�k��W��z.���k"�RH��zl��)������B���      D",���(�<H�FG��.���jλ(R���^e�a��.�� hX�x�Z:<��:2�;l�;��-;«9;wA;�cE;�G;��H;NGI;�`I;�UI;8BI;�1I;�#I;�I;�I;�I;�I;��H;I�H;��H;�H;�H;��H;�H;
�H;��H;G�H;�H;�I;�I;�I;�I;�#I;�1I;>BI;�UI;�`I;SGI;��H;"�G;�cE;uA;ɫ9;��-;m�;2�;B��:��Z: LX�&��Y���^e�(R���jλ�.��HG�:H���(�      �5���R��f ��'6��R�X�B�$�2ۺ�H[��
Q��c,:��:�:�>;D1";��0;��:;BaA;�cE;��G;r�H;�=I;+`I;nYI;�FI;�5I;�'I;�I;�I;�
I;�I;��H;�H;�H;��H;��H;��H;>�H;��H;~�H;��H;�H;�H;��H;�I;�
I;�I;�I;�'I;�5I;�FI;mYI;.`I;�=I;w�H;��G;�cE;HaA;��:;��0;E1";�>;�:��:�c,:�
Q��H[�6ۺH�$�P�X�*6��f ���R��      ��Ѻ�ȺX������t���(���9��Z:��:���:#0;S;0f);�4;��<;�KB;��E;$�G;u�H;\:I;O_I;[I; JI;9I;�*I;�I;�I;�I;\I;I;��H;��H;�H;1�H;��H;9�H;��H;3�H;��H;/�H;�H;��H;��H;I;\I;I;�I;�I;�*I;9I;!JI;�[I;S_I;_:I;y�H;!�G;��E;�KB;��<;�4;3f);S;%0;���:���:��Z:�9@(�X�����l���$�Ⱥ      ��9�:�":��Q:��:i��:v?�:Z��:�M
;��;#�&;'1;b`9;�m?;P�C;>VF;%�G;��H;�=I;N_I;\I;�KI;;I;�,I;� I;�I;�I;�I;HI;��H;5�H;x�H;5�H;��H;��H;��H;��H;��H;��H;��H;2�H;r�H;9�H;��H;FI;�I;�I;�I;� I;�,I;;I;�KI;\I;O_I;�=I;��H;(�G;@VF;T�C;�m?;e`9;
'1;'�&;��;�M
;T��:�?�:]��:��: �Q:@�": �:      ���:q��:��:��:��;FN;ZL;�, ;�f);��1;�w8;��=;]&B;�E;%G;KH;y�H;UGI;/`I;�[I;�KI;�;I;�-I;0"I;-I;I;	I;cI;��H;��H;��H;j�H;y�H;�H;F�H;��H;e�H;��H;C�H;�H;y�H;h�H;��H;��H;��H;dI;	I;I;1I;/"I;�-I;�;I;�KI;�[I;1`I;RGI;{�H;KH;%G;�E;_&B;��=;�w8;��1;�f);�, ;aL;@N;��;��:��:]��:      1�;��;s�;�/";��&;��+;��0;��5;��:;D�>;v B;��D;��F;��G;��H;�I;SI;�`I;nYI;!JI;;I;�-I;�"I;I;�I;�	I;)I;H�H;q�H;X�H;��H;��H;��H;��H;��H;��H;a�H;��H;��H;��H;��H;��H;��H;X�H;m�H;L�H;)I;�	I;�I;�I;�"I;�-I;;I;!JI;qYI;�`I;SI;�I;��H;��G;��F;��D;} B;A�>;��:;��5;��0;��+;ю&;�/";q�;̔;      ZY4;G�4;��5;�7;��9;�<;��>;�A;@C;=E;��F;,�G;c}H;g�H;�?I;�\I;`I;�UI;�FI; 9I;�,I;("I;�I;#I;X
I;�I;��H;��H;��H;��H;��H;��H;��H;��H;��H;��H;g�H;��H;��H;��H;��H;��H;��H;��H;��H;��H;��H;�I;]
I;!I;�I;,"I;�,I;�8I;�FI;�UI;`I;�\I;�?I;e�H;c}H;1�G;��F;=E;$@C;�A;��>;�<;ū9;�7;��5;=�4;      f�@;?�@;�`A;U&B;C;4D;�ME;�VF;�?G;&�G;ڐH;��H;�6I;�WI;,aI;)\I;�OI;EBI;�5I;�*I;� I;1I;�I;c
I;�I; I;.�H;��H;"�H;��H;��H;��H;L�H;{�H;��H;��H;f�H;��H;��H;|�H;I�H;��H;�H;��H;�H;��H;,�H; I;�I;b
I;�I;5I;� I;�*I;�5I;ABI;�OI;+\I;-aI;�WI;�6I;��H;ܐH;&�G;�?G;�VF;�ME;�3D;'C;[&B;�`A;>�@;      JVF;-hF;��F;��F;0MG;��G;N#H;��H;O�H;I;Y@I;�XI;RaI;�^I;�TI;�HI;�<I;�1I;�'I;�I;�I;I;�	I;�I; I;<�H;�H;Y�H;��H;��H;y�H;I�H;?�H;z�H;�H;��H;}�H;��H;�H;{�H;?�H;G�H;z�H;��H;��H;Y�H;�H;B�H; I;�I;�	I;I;�I;�I;�'I;�1I;�<I;�HI;�TI;�^I;RaI;�XI;a@I;I;R�H;��H;P#H;��G;GMG;��F;��F;*hF;      ��H;��H;G�H;��H;��H;�I;�%I;�@I;HTI;'_I;�aI;^I;�UI;KI;>@I;6I;�,I;�#I;�I;�I;�I;	I;*I;��H;*�H;�H;G�H;�H;,�H;o�H;(�H;�H;6�H;��H;8�H;��H;��H;��H;5�H;��H;9�H;�H;)�H;o�H;)�H;�H;D�H;�H;0�H;��H;,I;	I;�I;�I;�I;�#I;�,I;6I;>@I;KI;�UI;^I;�aI;$_I;GTI;�@I;�%I;�I;��H;��H;G�H;��H;      �GI;II;MI;�RI;*YI;�^I;�aI;pbI;�_I;EZI;pRI;�II;`@I;v7I;/I;'I;�I;�I;�I;�I;�I;^I;B�H;��H;��H;Q�H;�H;�H;z�H;(�H;�H;�H;d�H;��H;u�H;@�H;4�H;;�H;t�H;��H;g�H;	�H;�H;&�H;z�H;�H;�H;X�H;��H;��H;E�H;aI;�I;�I;�I;�I;�I;#'I;/I;x7I;^@I;�II;tRI;JZI;�_I;pbI;�aI;w^I;6YI;�RI;MI;II;      �bI;ubI;�aI;�`I;�^I;l[I;WI;�QI;"KI;7DI;=I;�5I;�.I;�'I;Z!I;I;5I;�I;�
I;`I;NI;��H;k�H;��H;�H;��H;%�H;|�H;�H;��H;��H;:�H;��H;*�H;��H;��H;��H;��H;��H;-�H;��H;8�H;��H;��H;�H;|�H;$�H;��H;�H;��H;n�H;��H;MI;\I;�
I;�I;6I;I;\!I;�'I;�.I;�5I;=I;9DI;&KI;�QI;WI;d[I;�^I;�`I;�aI;qbI;      OI;�NI;�MI;rKI;�HI;�DI;�@I;�;I;�6I;�1I;,I;�&I;!I;�I;�I;�I;I;�I;�I;I;��H;��H;T�H;��H;��H;��H;k�H;)�H;��H;��H;%�H;}�H;��H;��H;C�H; �H;�H;�H;A�H;��H;��H;}�H;&�H;��H;��H;(�H;i�H;��H;��H;��H;X�H;��H;��H;I;�I;�I;I;�I;�I;�I;!I;�&I;,I;�1I;�6I;�;I;�@I;�DI;�HI;zKI;�MI;�NI;      :I;�9I;�8I;#7I;�4I;!2I;�.I;G+I;R'I;9#I;�I;�I;QI;/I;I; 
I;�I;�I;��H;��H;?�H;��H;��H;��H;��H;u�H;&�H;�H;��H;*�H;��H;��H;[�H;�H;��H;��H;��H;��H;��H;�H;_�H;��H;��H;)�H;��H;�H;&�H;z�H;��H;��H;��H;��H;<�H;��H;��H;�I;�I;$
I;I;.I;RI;�I;�I;:#I;V'I;D+I;�.I;2I;�4I;&7I;�8I;�9I;      �)I;�)I;�(I;�'I;�%I;�#I;<!I;qI;kI;HI;�I;�I;+I;�
I;{I;HI;[I;��H;�H;��H;�H;i�H;��H;��H;��H;@�H;	�H;�H;;�H;�H;��H;u�H;��H;��H;v�H;M�H;8�H;M�H;q�H;��H;��H;w�H;��H;}�H;7�H;�H;�H;E�H;��H;��H;��H;l�H;{�H;��H;�H;��H;\I;II;}I;�
I;+I;�I;�I;II;kI;pI;F!I;�#I;�%I;�'I;�(I;�)I;      %I;�I;MI;AI;�I;;I;=I;I;�I;�I;_I;�
I;�I;(I;�I;  I;��H;K�H;#�H;�H;@�H;|�H;��H;��H;I�H;9�H;6�H;i�H;��H;��H;X�H;��H;��H;T�H;�H;�H;�H; �H;�H;W�H;��H;��H;X�H;��H;��H;h�H;8�H;<�H;N�H;��H;��H;{�H;<�H;�H;#�H;L�H;��H; I;�I;(I;�I;�
I;aI;�I;�I;I;AI;5I;�I;>I;TI;�I;      vI;ZI;�I;I;I;�I;I;<I;>I;
I;�I;�I;VI;$I;��H;��H;��H;��H;��H;5�H;��H;�H;��H;��H;u�H;q�H;��H;��H;,�H;��H;�H;��H;W�H;�H;��H;��H;��H;��H;��H;�H;X�H;��H;�H;��H;(�H;��H;��H;w�H;x�H;��H;��H;�H;��H;.�H;��H;��H;��H;��H;��H;#I;SI;�I;�I;
I;?I;9I;I;�I;	I;I;�I;eI;      �I;�I;@I;�I;�I;WI;I;�	I;�I;I;AI;[I;] I;x�H;��H;��H;��H;�H;��H;��H;��H;C�H;��H;��H;��H;��H;1�H;r�H;��H;F�H;��H;w�H;�H;��H;��H;��H;��H;��H;��H;��H;�H;x�H;��H;@�H;��H;q�H;4�H;�H;��H;��H;��H;B�H;��H;��H;��H;�H;��H;��H;��H;w�H;] I;XI;CI;I;�I;�	I;I;XI;�I;�I;@I;�I;      ~I;dI;I;qI;�
I;�	I;TI;�I;mI;�I;%I;h I;��H;��H;�H;X�H;��H;�H;��H;9�H;��H;��H;��H;z�H;��H;��H;��H;>�H;��H;$�H;��H;Q�H;�H;��H;��H;|�H;z�H;~�H;��H;��H;�H;Q�H;��H;�H;��H;=�H;��H;��H;��H;z�H;��H;��H;��H;3�H;��H;�H;��H;\�H;�H;��H;��H;e I;'I;�I;pI;�I;^I;�	I;�
I;oI; I;rI;      �I;WI;I;r
I;�	I;�I;�I;3I;�I;"I;pI;��H;�H;E�H;��H;��H;k�H;��H;A�H;��H;��H;h�H;^�H;_�H;e�H;r�H;��H;9�H;��H;$�H;��H;9�H;�H;��H;��H;v�H;��H;v�H;��H;��H;�H;<�H;��H;�H;��H;4�H;��H;w�H;c�H;]�H;a�H;e�H;��H;��H;A�H;��H;k�H;��H;��H;C�H;�H;��H;sI;"I;�I;3I;�I;�I;�	I;w
I;I;dI;      ~I;eI; I;nI;�
I;�	I;SI;�I;mI;�I;$I;i I;��H;��H;�H;X�H;��H;�H;��H;9�H;��H;��H;��H;z�H;��H;��H;��H;@�H;��H;"�H;��H;Q�H;�H;��H;��H;|�H;z�H;~�H;��H;��H;�H;Q�H;��H;�H;��H;:�H;��H;��H;��H;x�H;��H;��H;��H;3�H;��H;�H;��H;[�H;�H;��H;��H;e I;(I;�I;pI;�I;ZI;�	I;�
I;rI;I;lI;      �I;�I;;I;�I;�I;TI;I;�	I;�I;I;>I;YI;[ I;w�H;��H;��H;��H;�H;��H;��H;��H;D�H;��H;��H;��H;��H;3�H;t�H;��H;D�H;��H;w�H;�H;��H;��H;��H;��H;��H;��H;��H;�H;w�H;��H;?�H;��H;n�H;3�H;�H;��H;��H;��H;C�H;��H;��H;��H;�H;��H;��H;��H;w�H;] I;YI;CI;I;�I;�	I;I;TI;�I;�I;AI;�I;      vI;[I;�I;I;I;�I;I;?I;?I;	
I;�I;�I;SI;#I;��H;��H;��H;��H;��H;4�H;��H;�H;��H;��H;z�H;t�H;��H;��H;/�H;��H;�H;��H;W�H;�H;��H;��H;��H;��H;��H;�H;X�H;��H;�H;��H;(�H;��H;��H;v�H;u�H;��H;��H;�H;��H;/�H;��H;��H;��H;��H;��H;#I;SI;�I;�I;
I;?I;=I;I;�I;
I;I;�I;\I;      "I;�I;PI;?I;�I;=I;;I;I;�I;�I;\I;�
I;�I;(I;�I;  I;��H;K�H;!�H;�H;B�H;|�H;��H;��H;N�H;6�H;8�H;k�H;��H;��H;V�H;��H;��H;T�H;�H;�H;�H;�H;�H;U�H;��H;��H;X�H;��H;��H;e�H;6�H;9�H;I�H;��H;��H;y�H;6�H;�H;!�H;I�H;��H; I;�I;(I;�I;�
I;aI;�I;�I;I;BI;9I;�I;EI;XI;�I;      �)I;�)I;�(I;�'I;�%I;�#I;C!I;mI;hI;FI;�I;�I;+I;�
I;|I;FI;[I;��H;
�H;��H;��H;l�H;��H;��H;��H;A�H;�H;�H;>�H;}�H;��H;u�H;��H;��H;x�H;I�H;8�H;M�H;q�H;��H;��H;u�H;��H;|�H;7�H;�H;	�H;B�H;��H;��H;��H;j�H;y�H;��H;
�H;��H;\I;II;}I;�
I;,I;�I;�I;HI;jI;mI;D!I;�#I;�%I;�'I;�(I;�)I;      :I;�9I;�8I;!7I;�4I; 2I;�.I;H+I;P'I;6#I;�I;�I;QI;.I;I;!
I;�I;�I;��H;��H;@�H;��H;��H;��H;��H;s�H;%�H;�H;��H;)�H;��H;��H;\�H;�H;��H;��H;��H;��H;��H;�H;]�H;��H;��H;&�H;��H;�H;(�H;w�H;��H;��H;��H;��H;9�H;��H;��H;�I;�I; 
I;I;/I;QI;�I;�I;6#I;S'I;H+I;�.I;2I;�4I;*7I;�8I;�9I;      &OI;�NI;�MI;KI;|HI;�DI;�@I;�;I;�6I;�1I;,I;�&I;!I;�I;�I;�I;I;�I;�I;I;��H;��H;S�H;��H;��H;��H;k�H;(�H;�H; �H;&�H;��H;��H;��H;D�H;�H;�H; �H;A�H;��H;��H;��H;%�H;��H;��H;&�H;l�H;��H;��H;��H;Z�H;��H;��H;I;�I;�I;I;�I;�I;�I;!I;�&I;,I;�1I;�6I;�;I;�@I;�DI;�HI;�KI;�MI;�NI;      �bI;rbI;�aI;�`I;~^I;q[I; WI;�QI;*KI;5DI;=I;�5I;�.I;�'I;\!I;I;4I;�I;�
I;]I;OI;��H;j�H;��H;�H;��H;$�H;|�H;"�H;��H;��H;<�H;��H;*�H;��H;��H;��H;��H;��H;*�H;��H;;�H;��H;��H;�H;y�H;%�H;��H;�H;��H;o�H;��H;KI;\I;�
I;�I;4I;I;\!I;�'I;�.I;�5I;=I;5DI;$KI;�QI;WI;j[I;�^I;�`I;�aI;kbI;      �GI;II;MI;�RI;'YI;�^I;�aI;wbI;�_I;EZI;oRI;�II;^@I;u7I;/I;"'I;�I;�I;�I;�I;�I;aI;B�H;��H;��H;O�H;�H;�H;~�H;&�H;�H;�H;e�H;��H;v�H;=�H;6�H;@�H;r�H;��H;g�H;�H;�H;&�H;y�H;�H;�H;T�H;��H;��H;H�H;`I;�I;�I;�I;�I;�I;"'I;/I;t7I;^@I;�II;qRI;HZI;�_I;pbI;�aI;}^I;5YI;�RI;MI;II;      ��H;��H;D�H;��H;��H;�I;�%I;�@I;JTI;&_I;�aI;!^I;�UI;KI;>@I;6I;�,I;�#I;�I;�I;�I;	I;&I;��H;.�H;�H;F�H;�H;/�H;o�H;(�H;�H;8�H;��H;:�H;��H;��H;��H;5�H;��H;8�H;�H;)�H;o�H;)�H;�H;H�H;�H;-�H;��H;.I;	I;�I;�I;�I;�#I;�,I;	6I;?@I;KI;�UI;^I;�aI;#_I;ETI;�@I;�%I;�I;��H;��H;E�H;��H;      @VF;(hF;��F;��F;7MG;��G;M#H;��H;P�H;I;Z@I;�XI;SaI;�^I;�TI;�HI;�<I;�1I;�'I;�I;�I;I;�	I;�I; I;;�H;�H;]�H;��H;��H;y�H;K�H;=�H;z�H;	�H;��H;~�H;��H;�H;z�H;?�H;K�H;}�H;��H;��H;Y�H;�H;>�H; I;�I;�	I;I;�I;�I;�'I;�1I;�<I;�HI;�TI;�^I;RaI;�XI;]@I;I;I�H;��H;M#H;��G;@MG;��F;��F;hF;      d�@;:�@;�`A;[&B;C;4D;�ME;�VF;�?G;%�G;ڐH;��H;�6I;�WI;0aI;+\I;�OI;EBI;�5I;�*I;� I;5I;�I;c
I;�I; I;.�H;��H;$�H;��H;��H;��H;I�H;z�H;��H;��H;h�H;��H;��H;|�H;K�H;��H;�H;��H; �H;��H;.�H; I;�I;_
I;�I;4I;� I;�*I;�5I;?BI;�OI;+\I;.aI;�WI;�6I;��H;ڐH;%�G;�?G;�VF;�ME;�3D;#C;[&B;�`A;;�@;      5Y4;.�4;��5;�7;��9;�<;��>;�A;%@C;:E;��F;/�G;c}H;d�H;�?I;�\I;`I;�UI;�FI;�8I;�,I;)"I;�I;#I;]
I;�I;��H;��H;��H;��H;��H;��H;��H;��H;��H;��H;j�H;��H;��H;��H;��H;��H;��H;��H;��H;��H;��H;�I;Y
I;!I;�I;)"I;�,I;9I;�FI;�UI;`I;�\I;�?I;d�H;c}H;,�G;��F;<E;@C;�A;��>;�<;ɫ9;%�7;��5;�4;      �;ٔ;e�;�/";��&;��+;��0;��5;��:;D�>;r B;��D;��F;��G;��H;�I;SI;�`I;nYI;!JI;;I;�-I;�"I; I;�I;�	I;)I;L�H;r�H;V�H;��H;��H;��H;��H;��H;��H;d�H;��H;��H;��H;��H;��H;��H;Z�H;n�H;I�H;-I;�	I;�I;�I;�"I;�-I;;I;#JI;rYI;�`I;SI;�I;��H;��G;��F;��D;u B;B�>;��:;��5;��0;��+;��&;�/";f�;Ŕ;      ���:k��:��:��:��;LN;_L;�, ;�f);��1;�w8;��=;_&B;�E;'G;KH;y�H;UGI;.`I;�[I;�KI;�;I;�-I;/"I;3I;I;	I;eI;��H;��H;��H;m�H;y�H;�H;D�H;��H;g�H;��H;B�H;�H;y�H;l�H;��H;��H;��H;cI;	I;I;.I;0"I;�-I;�;I;�KI;�[I;1`I;QGI;y�H;KH;%G;�E;^&B;��=;�w8;��1;�f);�, ;[L;6N;��;��:��:W��:      ���9d�:L�":�Q:��:q��:|?�:^��:�M
;��;$�&;'1;c`9;�m?;U�C;@VF;(�G;��H;�=I;O_I;\I;�KI;;I;�,I;� I;�I;�I;�I;HI;��H;6�H;{�H;5�H;��H;��H;��H;��H;��H;��H;��H;5�H;y�H;9�H;��H;FI;�I;�I;�I;� I;�,I;;I;�KI;\I;Q_I;�=I;��H;(�G;@VF;U�C;�m?;e`9;'1;'�&;��;�M
;`��:�?�:i��:��:�Q:��":$�:      ��Ѻ�Ⱥd������|��0(��9��Z:���:���:%0;S;2f);�4;��<;�KB;��E;"�G;u�H;_:I;S_I;�[I; JI;9I;�*I;�I;�I; I;_I;I;��H;��H;�H;2�H;��H;4�H;��H;7�H;��H;.�H;�H;��H;��H;I;]I;�I;�I;�I;�*I;9I;!JI;�[I;R_I;_:I;w�H; �G;��E;�KB;��<;�4;2f);S;%0;���:���:��Z:ؓ�9�(�X�����f����Ⱥ      �5���R��f ��$6��W�X�B�$�6ۺ�H[�@
Q��c,:��:�:�>;C1";��0;��:;EaA;�cE;��G;v�H;�=I;/`I;pYI;�FI;�5I;�'I;�I;�I;�
I;�I;��H;�H;�H;��H;�H;��H;>�H;��H;}�H;��H;�H;�H;��H;�I;�
I;�I;�I;�'I;�5I;�FI;pYI;,`I;�=I;w�H;��G;�cE;EaA;��:;��0;E1";�>;�:��:�c,:�
Q��H[�6ۺE�$�T�X�$6��h ���R��      H",���(�>H�FG��.���jλ&R���^e�\��,�� XX���Z:@��:2�;p�;��-;ȫ9;uA;�cE; �G;��H;SGI;�`I;�UI;>BI;�1I;�#I;�I;�I;�I;�I;��H;H�H;��H;�H;�H;��H;�H;	�H;��H;I�H;��H;�I;�I;�I;�I;�#I;�1I;8BI;�UI;�`I;RGI;��H;"�G;�cE;uA;ƫ9;��-;p�;2�;<��:��Z: XX�,��]���^e�(R���jλ�.��HG�@H���(�      �d��D��������)���zl�RH��k"�y.���W��g�k��� ������9���:k��:�;�-;ʫ9;DaA;��E;)�G;y�H;�RI;`I;�OI;�<I;�,I;�I;2I;I;I;UI;��H;��H;��H;��H;d�H;��H;��H;��H;��H;UI;I;I;1I;�I;�,I;�<I;�OI;`I;�RI;v�H;#�G;��E;DaA;ȫ9;�-;�;g��:���:��9����� �i�k��W��y.���k"�RH��zl��)������C���      ���i9�\5��;��Ub̼~֮�v��� d�",�����Q��JG5�|#��`�f9~��:��:�;��-;��:;�KB;@VF;KH;�I;�\I;#\I;�HI;6I;'I;I;�I;
I;EI;��H;��H;��H;Z�H;��H;Z�H;��H;��H;��H;CI;
I;�I;I;'I;6I;�HI;\I;�\I;�I;KH;8VF;�KB;��:;��-;�;��:x��:`�f9|#��OG5��Q�����",�� d�w��~֮�Vb̼<��]5��j9�      �]��IY��ZN��`=���'�m����෾������W��$�h��u�X�섮�P9x��:_��:m�;��0;��<;W�C;%G;��H;�?I;*aI;�TI;<@I;/I;[!I;�I;I;|I;�I;��H;��H;�H;��H;�H;}�H;��H;�I;yI;I;�I;\!I;/I;<@I;�TI;%aI;�?I;��H;#G;M�C;��<;��0;i�;c��:t��:�9ꄮ�w�X�i���$��W�����᷾����m���'��`=��ZN��IY�      �A��!��d���*��潅�>�d��`=����^��e֮�N�y�|�(��һ�]e�℮���f9���:4�;E1";�4;�m?;�E;��G;j�H;�WI;�^I;KI;r7I;�'I;�I;+I;�
I;$I;I;p�H;��H;>�H;��H;m�H;I;$I;�
I;'I;�I;�'I;t7I;
KI;}^I;�WI;h�H;��G;�E;�m?;�4;A1";2�;���:`�f9섮��]e��һ|�(�N�y�e֮�^�꼗���`=�>�d�罅��*��c��!��      ���GE	��������Wн�A�����h���3���� ¼�)��1x/��һo�X�n#����9L��:�>;3f);l`9;a&B;��F;j}H;�6I;RaI;�UI;b@I;�.I;!I;MI;+I;�I;SI;T I;��H;��H;��H;S I;PI;�I;(I;JI;!I;�.I;a@I;�UI;NaI;�6I;g}H;��F;^&B;b`9;6f);�>;B��:��9t#��s�X��һ2x/��)��!¼�����3��h��󑽢A���Wн��콺��GE	�      ~^Z�`
V��I��6�������ܽ!��ڽ���aG�[�
�ȼ�)��|�(�f��JG5������Z:�:S;'1;��=;��D;2�G;��H;�XI;^I;II;�5I;�&I;�I;�I;�
I;�I;OI;b I;��H;d I;NI;�I;�
I;�I;�I;�&I;�5I;II;^I;�XI;��H;1�G;��D;��=;'1;S;�:��Z:���NG5�h��}�(��)��
�ȼ[��aG�ڽ��!���ܽ������6��I�`
V�      � ���e�����ܕ����q��I���"���������k���ZN�[�!¼P�y��$��Q���� � pX���:0;+�&;�w8;s B;��F;ڐH;Z@I;�aI;pRI;=I;,I;�I;�I;_I;�I;7I;!I;hI;!I;7I;�I;_I;�I;�I;,I;=I;pRI;�aI;V@I;ԐH;��F;s B;�w8;�&;0;��: pX��� ��Q���$�P�y�"¼[��ZN�k������������"��I���q�ܕ������e��      d5�������W�Ҿ�a��{����l�	�6�DE	���Ƚk���aG����f֮��W����m�k�6���c,:���:�;��1;B�>;CE;&�G;I;&_I;DZI;:DI;�1I;6#I;FI;I;	
I;I;�I;"I;�I;I;
I;I;EI;4#I;�1I;9DI;DZI;$_I;I;"�G;@E;E�>;��1;�;���:�c,:6��m�k�����W�f֮�����aG�k����ȽDE	�	�6��l�{����a��W�Ҿ������      {A��q<�fa/����:�z]׾� ��w��>�DE	�����ڽ����3�^�꼙���",��W��c�� Q���:�M
;�f);��:;'@C;�?G;R�H;HTI;�_I;,KI;�6I;S'I;jI;�I;AI;�I;qI;�I;pI;�I;?I;�I;jI;R'I;�6I;,KI;�_I;HTI;S�H;�?G;*@C;��:;�f);�M
;���: Q�c���W��",�����^�꼙�3�ڽ������DE	�>�w��� ��z]׾�:���fa/��q<�      v�������`�{�k$_��q<�������}��w��	�6�����!���h����ⷾ�� d�~.���^e��H[���Z:h��:�, ;��5;�A;�VF;��H;�@I;rbI;�QI;�;I;A+I;qI;I;<I;�	I;�I;0I;�I;�	I;:I;I;nI;A+I;�;I;�QI;sbI;�@I;��H;�VF;�A;��5;�, ;R��:��Z:I[��^e�~.��� d�ⷾ�����h�!������	�6�w���}��������q<�k$_�`�{�����      ;��������欿��� ����O��x����� ���l���"��ܽ���`=����w���k"�-R��@ۺГ�9�?�:^L;��0;��>;�ME;H#H;�%I;�aI;WI;�@I;�.I;B!I;BI;I;I;PI;�I;OI;I;I;BI;@!I;�.I;�@I;WI;�aI;�%I;Q#H;�ME;��>;��0;[L;z?�:Г�9Jۺ.R���k"�w������`=����ܽ��"��l�� ����뾁x���O� ������欿����      �������M��jȿk���������O���z]׾{����I�����A��>�d�n�~֮�RH��jλO�$��(�q��:FN;��+;�<;�3D;��G;�I;�^I;n[I;�DI;'2I;�#I;GI;�I;aI;�	I;�I;�	I;aI;�I;GI;�#I;"2I;�DI;n[I;�^I;�I;��G;�3D;�<;��+;BN;e��:�(�T�$��jλRH�֮�n�>�d��A������I�{���z]׾����O�����k���jȿL�Ῡ��      @�2i�������I�ѿk��� ���q<��:��a����q����Wн罅���'�Ub̼�zl��.��M�X�`����:��;Ύ&;ƫ9;&C;8MG;��H;9YI;�^I;�HI;�4I;�%I;�I;I;�I;�
I;�	I;�
I;�I;I;�I;�%I;�4I;�HI;�^I;<YI;��H;CMG;$C;ƫ9;ˎ&;��;��:`��Q�X��.���zl�Ub̼��'�罅��Wн����q��a���:��q<� ��k���I�ѿ������2i�      G:�.5�.�'��������jȿ���k$_���W�Ҿܕ���6�����*���`=�>�漮)��JG�&6�����(�Q:��:�/";�7;^&B;��F;��H;�RI;�`I;zKI;7I;�'I;?I;I;�I;tI;u
I;qI;�I;I;BI;�'I;7I;�KI;�`I;�RI;��H;��F;^&B;	�7;�/";��:�Q:���)6��IG��)��=���`=��*������6�ܕ��W�Ҿ��k$_����jȿ�������.�'�.5�      ��U�Z�O�H-?�.�'���M�ῴ欿`�{�fa/���뾝���I����d���ZN�\5������=H�d ��j�����":��:{�;��5;�`A;��F;L�H;MI;�aI;�MI;�8I;�(I;DI;�I;;I;
I;I;I;=I;�I;FI;�(I;�8I;�MI;�aI;MI;N�H;��F;�`A;��5;t�;��:h�":`���g ��=H�����\5���ZN�d������I�������fa/�`�{��欿M����.�'�H-?�Z�O�      ��i���b�Z�O�.5�2i�������������q<�����e��`
V�GE	�!���IY�j9�E�����(��R���ȺX�:Q��:�;A�4;>�@;hF;��H;II;|bI;�NI;�9I;�)I;�I;_I;�I;bI;`I;^I;�I;_I;�I;�)I;�9I;�NI;|bI;II;��H;*hF;>�@;?�4;ڔ;I��:@�:�Ⱥ�R����(�E���j9��IY�!��GE	�`
V��e������q<������������2i�.5�Z�O���b�      �>���8���*�O������˿p��E�b�C\�4m־^��R�:��J�)��E�B�=��������1/��T����>:it�:p ;�J6;�DA;]IF;�NH;��H;�!I;�I;�I;�I;UI;�I;P I;��H;�H;��H;M I;�I;SI;�I;�I;�I;�!I;��H;�NH;gIF;�DA;�J6;p ;at�:ԑ>:R���2/���������=��E�B�)���J�R�:�^��4m־C\�E�b�p���˿����O���*���8�      ��8��4��g&�6��<����<ƿ񲗿�>]����P�Ѿ�p���*7����%W��LR?� }�r8�������؅����G:s �:�!;�6;�kA;hYF;�TH;G�H;�!I;�I;�I;nI;/I;�I;A I;��H;��H;��H;A I;�I;-I;nI;�I;�I;�!I;I�H;�TH;pYF;�kA;�6;�!;k �:|�G:҅�������r8�� }�LR?�%W�����*7��p��P�Ѿ����>]�񲗿�<ƿ<���6���g&��4�      ��*��g&��#�t�U[�pL�������M�r5��>ľ����,��D�蒐��5�2�ݼ���q
��x�(uk���b:+l�:�#;Ɨ7;V�A;��F;�dH;�I;&"I;�I;II;I;�I;�I;��H;`�H;��H;Y�H;��H;�I;�I;I;DI;�I;&"I;�I;�dH;��F;S�A;��7;�#;l�:��b:uk��x��q
���2�ݼ�5�蒐��DὪ�,����>ľr5���M����pL��U[�t��#��g&�      O�6��t����˿@1��6�y�Î6��z �����1�l�+��ͽ$�����&���˼@�k�$�����X� � �v��:8�;�&;�9;k�B;��F;�}H;�	I;5"I;I;�I;I;[I;)I;��H;�H;h�H;�H;��H;)I;VI;}I;�I; I;5"I;�	I;�}H;��F;j�B;z9;�&;4�;l��:�� ���X�$���@�k���˼��&�$����ͽ+�1�l������z �Î6�6�y�@1���˿���t�6��      ����<���U[忶˿�T���{�R�����E۾ӗ����M���	������j��3�d����O�;�׻��/�`��?��:� 
;�*;P;;�jC;�'G;؛H;�I;�!I;�I;{I;�
I;�I;�I;(�H;��H;��H;��H;(�H;�I;�I;�
I;vI;�I;�!I;�I;؛H;�'G;�jC;L;;�*;� 
;1��:H����/�<�׻��O�d���3���j������	���M�ӗ���E۾���{�R���T���˿U[�<���      �˿�<ƿpL��@1����>]���)��$��ֳ���{���,�r��'��Q`I��J���,���3/� ,��� ��,69�4�:Ԅ;�o.;.=;?aD;��G;V�H;�I;!I;BI;-I;�	I;�I;� I;��H;��H;H�H;��H;��H;� I;�I;�	I;*I;FI;!I;�I;Q�H;��G;=aD;.=;�o.;΄;�4�: -69� �,���3/��,���J��Q`I�'��q�齤�,���{�ֳ��$����)��>]��@1��pL���<ƿ      p��񲗿���6�y�{�R���)�nv��>ľ^���I�Xl����������&�ԮҼ�}�1B�̮�����t�!:�*�:$z;[3;Kj?;r\E;��G;��H;LI;�I;nI;�I;[I;�I;��H;��H;I�H;��H;F�H;��H;��H;�I;WI;�I;tI;�I;KI;��H;��G;s\E;Ij?;Y3; z;�*�:��!:���ή��1B��}�ԮҼ��&��������Xl��I�^���>ľnv���)�{�R�6�y����񲗿      E�b��>]���M�Î6�����$���>ľ"q��y�Z�+�Q9ݽ!W����L����"F���G��׻;�@o�|Ȋ:�i;P$;��7;W�A;�IF;CH;��H;� I;GI;ZI;�I;I;�I;��H;��H;y�H;��H;x�H;��H;��H;�I;
I;�I;^I;EI;� I;��H;CH;�IF;Q�A;��7;P$;zi;�Ȋ:Ho�;��׻�G�"F�������L�!W��Q9ݽ+�y�Z�"q���>ľ�$�����Î6���M��>]�      C\����r5��z ��E۾ֳ�^��y�Z�L?#����A����j�&��Dϼ�����̵���lۺ`9�9`4�:A�;G�,;W�;;�C;G; �H;�I;�!I;�I;(I;	I;wI;(I;��H;��H;��H;�H;��H;��H;��H;&I;vI;I;+I;�I;�!I;�I;"�H;�G;�C;X�;;H�,;:�;l4�:X9�9�lۺ˵�������Dϼ%����j��A�����L?#�y�Z�^��ֳ��E۾�z �r5����      4m־P�Ѿ�>ľ����ӗ����{��I�+�����V���{�?�/�%���,��@=�D�һq�@�H� ���k:��:�a;��3;	j?;R2E;��G;B�H;I;P I;�I;�I;	I;�I;��H;��H;��H;��H;<�H;��H;��H;��H;��H;�I; 	I;�I;�I;Q I;I;A�H;��G;P2E;j?;��3;�a;��:��k:T� �n�@�D�һ@=��,��%��?�/��{��V�����+��I���{�ӗ�������>ľP�Ѿ      ^���p����1�l���M���,�Xl�Q9ݽ�A���{���5��J��
;���T[�"?�����dP�� P�9��:��;*;�9;4kB;��F;WNH;W�H; I;iI;�I;I;�I;%I;H�H;��H;��H;��H;M�H;��H;��H;��H;G�H;"I;�I;I;�I;lI;�I;V�H;ZNH;��F;7kB;�9;
*;��;��:�O�9\P������"?��T[�	;���J����5��{��A��Q9ݽXl���,���M�1�l����p��      Q�:��*7���,�+���	�q�齂���!W����j�?�/��J���I���k�m�.��h��`���Ȋ:'o�:�;Cr3; �>;�D;O�G;%�H;�I;!I;�I;hI;c
I;�I;B I;��H;|�H;��H;��H;D�H;��H;��H;�H;��H;B I;�I;i
I;oI;�I;!I;�I;(�H;O�G;	�D;�>;Cr3;�;/o�:�Ȋ:0��h��.��l��k��I���J��?�/���j�!W������q�齂�	�+���,��*7�      �J�����D��ͽ���'�������L�%��%��	;���k����nI����/��/��>:��:�B;<�,;��:;�B;ixF;v<H;��H;�I;tI;�I;I;�I;�I;p�H;Z�H;�H;R�H;��H;Q�H;��H;R�H;�H;W�H;n�H;�I;�I;!I;�I;sI;�I;��H;v<H;kxF;�B;��:;H�,;�B;��:$�>:�/���/�lI������k�	;��%��%����L����'������ͽ�D����      (��%W��蒐�$�����j�R`I���&����Dϼ�,���T[�n�oI��h;��nk�h:�4�:�;�&;��6;�!@;2E;��G;��H;�I;� I;3I;�I;�
I;I;S I;��H;��H;��H;D�H;x�H;*�H;x�H;C�H;��H;��H;��H;W I;#I;�
I;�I;2I;� I;�I;��H;��G;2E;�!@;��6;�&;�;�4�:h:�nk�d;�mI��l��T[��,��Cϼ�����&�Q`I���j�$���蒐�$W��      D�B�MR?��5���&��3��J��ԮҼ F����?=�!?�.����/��nk�ȭ�9׳:��;!;93;��=;��C;��F;�cH;��H;lI;�I;�I;I;�I;�I;"�H;��H;u�H;b�H;$�H;g�H;�H;g�H;#�H;d�H;u�H;��H;%�H;�I;�I;I;�I;�I;qI;��H;�cH; �F;��C;��=;?3;!;��;׳:ȭ�9�nk���/�.�� ?�?=���!F��ԮҼ�J���3���&��5�MR?�      :���|�1�ݼ��˼d���,���}��G����D�һ����k���/�d:׳:�;Mb;��0;m<;�B;�IF;KH; �H;�I;L I;�I;I;9
I;�I; I;�H;8�H;��H;�H;�H;^�H;�H;]�H;�H;	�H;��H;6�H;�H; I;�I;=
I;I;�I;S I;�I;�H;OH;�IF;��B;q<;��0;Pb;�;&׳:h:�/�f������C�һ����G��}��,��d����˼1�ݼ�|�      ����p8����A�k���O��3/�/B�
�׻ȵ��i�@�TP��H��$�>:�4�:��;Sb;�/;;;�A;d�E;��G;ѭH;�
I;D I;�I;�I;�I;�I;�I;h�H;�H;��H;{�H;��H;��H;R�H;�H;N�H;��H;��H;z�H;��H; �H;l�H;�I;�I;�I;�I;�I;G I;�
I;խH;��G;o�E; �A;;;��/;Sb;��;�4�:$�>:(��NP��g�@�ǵ��
�׻0B��3/���O�B�k���o8��      ������q
����6�׻�+��Ȯ��;��lۺ<� �P�9�Ȋ:��:�;!;��0;	;;��A;�pE;M�G;��H;��H;�I;I;.I; I;�I;SI;��H;%�H;Z�H;��H; �H;��H;��H;I�H;�H;F�H;��H;��H;��H;��H;^�H;*�H;��H;VI;�I;�I;5I;I;�I;��H;��H;T�G;�pE;��A;;;��0;!;�;��:�Ȋ:8P�90� ��lۺ;�ʮ���+��2�׻ ����q
���      &/��&����x���X���/�� �
���o칈9�9��k:��:!o�:�B;�&;=3;n<;�A;�pE;@tG;�|H;�H;I;OI;#I;�I;K
I;�I;1 I;-�H;�H;��H;`�H;��H;��H;��H;[�H;F�H;X�H;��H;��H;��H;]�H;��H;�H;-�H;5 I;�I;H
I;�I;&I;NI;	I;�H;�|H;CtG;�pE;!�A;n<;A3;�&;�B;)o�:��:��k:�9�9o����� ���/���X��x�&���      N���䅍��tk��� ����0-69��!:zȊ:l4�:��:��;�;C�,;��6;��=;��B;m�E;W�G;�|H;t�H;VI;�I;_I;9I;�I;I;hI;'�H;��H;�H;��H;��H;��H;��H;��H;q�H;V�H;k�H;��H;��H;��H;��H;��H;�H;��H;-�H;fI;I;�I;:I;_I;�I;[I;u�H;�|H;S�G;o�E;��B;��=;��6;G�,;�;��;��:n4�:�Ȋ:��!:p-69H��� �uk�􅍺      T�>:@�G:h�b:`��:��:�4�:�*�:|i;;�;�a;
*;<r3;��:;�!@;��C;�IF;��G;��H;
�H;SI;�I;I;I;�I;�I;9I;��H;m�H;��H;Z�H;,�H;��H;|�H;��H;��H;��H;d�H;��H;��H;��H;z�H;��H;0�H;^�H;��H;n�H;��H;9I;�I;�I;I;!I; I;VI;�H;��H;��G;�IF;��C;�!@;��:;Br3;*;�a;9�;zi;�*�:�4�:5��:f��:��b:H�G:      at�:� �:Al�:E�;� 
;҄;z; P$;K�,;��3;�9;��>;�B;2E;�F;OH;խH;��H;
I;�I;"I;\I;I;�I;�I;��H;�H;0�H;��H;y�H;��H;��H;r�H;��H;�H;��H;��H;��H;�H;��H;r�H;��H;��H;|�H;��H;1�H; �H;��H;�I;�I;I;^I;%I;�I;
I;��H;٭H;PH;�F;2E;�B;�>;�9;��3;K�,;P$;&z;΄;� 
;<�;-l�:{ �:      $p ;�!;�#;�&;�*;�o.;c3;��7;\�;;j?;;kB;	�D;kxF;��G;�cH;�H;�
I;�I;QI;aI;I;I;�I;:I;�H;o�H;o�H;�H;��H;��H;��H;d�H;t�H;��H;8�H;�H;��H;��H;6�H;��H;t�H;c�H;��H;��H;��H;�H;n�H;r�H;�H;7I;�I;I;I;bI;RI;�I;�
I;
�H;�cH;��G;nxF;�D;BkB;j?;_�;;��7;b3;�o.;�*;�&;�#;�!;      �J6;�6;��7;z9;A;;.=;Ej?;S�A;�C;P2E;��F;J�G;r<H;�H;��H;�I;E I;I;%I;6I;�I;�I;3I;-�H;��H;��H;A�H;�H; �H;��H;h�H;U�H;v�H;�H;��H;T�H;,�H;O�H;��H;�H;v�H;T�H;m�H;��H;�H;�H;?�H;��H;��H;-�H;3I;�I;�I;6I;&I;I;J I;�I;��H;�H;r<H;O�G;��F;R2E;�C;[�A;Ej?;.=;P;;z9;��7;�6;       EA;�kA;M�A;d�B;�jC;MaD;{\E;�IF;�G;��G;`NH;+�H;��H;�I;tI;X I;�I;9I;�I;�I;�I;�I;�H;��H;��H;]�H;�H;0�H;��H;y�H;N�H;f�H;��H;B�H;��H;��H;��H;��H;��H;C�H;��H;b�H;R�H;{�H;��H;0�H;�H;`�H;��H;��H;�H;�I;�I;�I;�I;7I;�I;[ I;uI;�I;��H;0�H;aNH;��G;�G;�IF;{\E;CaD;�jC;j�B;O�A;�kA;      ZIF;sYF;��F;��F;t'G;��G;��G;CH;�H;E�H;W�H;�I;�I;� I;�I;�I;�I; I;J
I;I;=I;��H;n�H;��H;\�H;8�H;C�H;��H;{�H;]�H;G�H;��H;�H;}�H;7�H;�H;�H;�H;4�H;}�H;�H;��H;I�H;\�H;{�H;��H;A�H;>�H;`�H;��H;o�H;��H;?I;I;M
I;�I;�I;�I;�I;� I;�I;�I;_�H;F�H;"�H;CH;��G;��G;�'G;��F;��F;rYF;      �NH;�TH;�dH;�}H;̛H;S�H;��H;��H;�I;I;  I;!I;oI;0I;�I;I;�I;�I;�I;jI;�H;��H;o�H;F�H;�H;@�H;��H;�H;M�H;M�H;��H;��H;V�H;��H;��H;��H;x�H;��H;��H;��H;W�H;��H;��H;N�H;J�H;�H;��H;G�H;�H;D�H;p�H;�H;�H;iI;�I;�I;�I;I;�I;/I;pI;!I; I;I;�I;��H;��H;O�H;�H;�}H;�dH;yTH;      ��H;J�H;�I;�	I;�I;�I;UI;� I;�!I;U I;lI;�I;�I;�I;�I;<
I;�I;RI;3 I;(�H;n�H;,�H;�H;�H;)�H;��H;|�H;]�H;C�H;u�H;��H;3�H;��H;r�H;2�H;�H;��H;��H;2�H;u�H;��H;2�H;��H;u�H;B�H;]�H;{�H;��H;/�H;�H;	�H;0�H;q�H;*�H;3 I;RI;�I;@
I;I;�I;�I;�I;pI;W I;�!I;� I;UI;�I;�I;�	I;�I;?�H;      �!I;�!I;#"I;D"I;�!I;!I;�I;GI;�I;�I;�I;mI; I;�
I;�I;�I;�I;��H;1�H;��H;��H;��H;��H; �H;��H;r�H;D�H;F�H;��H;��H;!�H;��H;?�H;��H;��H;��H;��H;��H;��H;��H;D�H;��H;%�H;��H;��H;D�H;C�H;v�H;��H;�H;��H;��H;��H;��H;3�H;��H;�I;�I;�I;�
I; I;mI;�I;�I;�I;GI;�I;!I;�!I;I"I;"I;�!I;      �I;�I;�I;I;�I;<I;mI;[I;'I;�I;I;k
I;�I;!I;�I; I;o�H;"�H;�H;!�H;a�H;v�H;��H;��H;t�H;Q�H;I�H;v�H;��H;�H;��H;=�H;��H;��H;a�H;B�H;1�H;@�H;^�H;��H;��H;<�H;��H;�H;��H;v�H;F�H;Y�H;{�H;��H;��H;x�H;^�H;�H;�H;"�H;p�H; I;�I;I;�I;i
I;I;�I;)I;ZI;qI;<I;�I;I;�I;�I;      �I;�I;NI;�I;tI;*I;�I;�I;I;	I;�I;�I;�I;] I;)�H;�H;%�H;^�H;��H;��H;6�H;��H;��H;j�H;M�H;C�H;��H;��H;(�H;��H;�H;��H;m�H;2�H;�H;��H;��H;��H;�H;6�H;p�H;��H;�H;��H;#�H;��H;��H;J�H;R�H;j�H;��H;��H;3�H;��H;��H;^�H;(�H;�H;+�H;] I;�I;�I;�I;	I;I;�I;�I;"I;�I;�I;LI;�I;      �I;rI;I;qI;�
I;�	I;XI;I;{I;�I;"I;F I;r�H;��H;��H;<�H;��H;��H;e�H;��H;��H;��H;a�H;R�H;c�H;��H;��H;3�H;��H;?�H;��H;N�H;�H;��H;��H;��H;��H;��H;��H;��H;�H;L�H;��H;<�H;��H;2�H;��H;��H;h�H;N�H;h�H;��H;��H;��H;d�H;��H;��H;=�H;��H;��H;r�H;E I;)I;�I;wI;I;aI;�	I;�
I;yI;I;pI;      WI;6I;�I;XI;�I;�I;�I;I;I;��H;J�H;��H;\�H;��H;w�H;��H;��H;�H;��H;��H;��H;v�H;t�H;t�H;��H;�H;U�H;��H;F�H;��H;j�H;�H;��H;��H;��H;e�H;`�H;g�H;��H;��H;��H;�H;i�H;��H;C�H;��H;W�H;�H;��H;v�H;z�H;u�H;��H;��H;��H;�H;��H;��H;w�H;��H;]�H;��H;M�H;��H;!I;|I;�I;�I;�I;UI;�I;3I;      �I;�I;�I;I;�I;� I;��H;��H;��H;��H;��H;��H; �H;��H;i�H;�H;��H;��H;��H;��H;��H;��H;��H;�H;>�H;x�H;��H;u�H;��H;��H;.�H;��H;��H;g�H;Q�H;B�H;5�H;B�H;Q�H;h�H;��H;��H;/�H;��H;��H;r�H;��H;{�H;?�H;�H;��H;��H;��H;��H;��H;��H;��H;�H;f�H;��H;�H;��H;��H;��H;��H;��H; I;� I;�I;I;�I;�I;      E I;Q I; I;��H;0�H;z�H;��H;��H;��H;��H;��H;��H;Z�H;K�H;+�H;�H;��H;��H;��H;��H; �H;�H;5�H;��H;��H;,�H;��H;2�H;��H;e�H;��H;��H;��H;P�H;.�H;�H;%�H;"�H;,�H;Q�H;��H;��H;��H;^�H;��H;/�H;��H;0�H;��H;��H;9�H;�H;��H;��H;��H;��H;��H;
�H;(�H;J�H;Z�H;��H;��H;��H;��H;��H;��H;{�H;0�H;��H; I;S I;      ��H;��H;X�H;�H;��H;��H;L�H;y�H;��H;��H;��H;��H;��H;z�H;g�H;\�H;T�H;C�H;[�H;o�H;��H;��H;��H;F�H;��H;�H;��H;�H;��H;G�H;��H;��H;k�H;C�H;%�H;�H;
�H;�H; �H;H�H;n�H;��H;��H;B�H;��H;��H;��H;�H;��H;F�H; �H;��H;��H;j�H;Z�H;I�H;U�H;^�H;g�H;{�H;��H;��H;��H;��H;��H;x�H;V�H;��H;��H;�H;T�H;��H;      �H;��H;��H;h�H;��H;>�H;��H;��H;�H;9�H;V�H;L�H;V�H;2�H; �H;�H;�H;�H;I�H;\�H;p�H;��H;��H;%�H;��H;��H;t�H;��H;��H;6�H;��H;��H;b�H;3�H;%�H;�H;�H;�H;"�H;4�H;g�H;��H;��H;1�H;��H;��H;w�H;�H;��H;#�H;��H;��H;i�H;W�H;I�H;�H;�H;"�H; �H;1�H;V�H;I�H;X�H;9�H;�H;��H;��H;>�H;��H;l�H;��H;��H;      ��H;��H;R�H;�H;��H;��H;L�H;x�H;��H;��H;��H;��H;��H;{�H;g�H;\�H;T�H;C�H;[�H;o�H;��H;��H;��H;F�H;��H;�H;��H;�H;��H;F�H;��H;��H;l�H;E�H;%�H;�H;�H;�H;�H;F�H;n�H;��H;��H;@�H;��H;��H;��H;�H;��H;E�H; �H;��H;��H;j�H;Z�H;G�H;T�H;^�H;g�H;x�H;��H;��H;��H;��H;��H;{�H;S�H;��H;��H;�H;V�H;��H;      : I;S I;��H;��H;2�H;w�H;��H;��H;��H;��H;��H;��H;\�H;J�H;*�H;�H;��H;��H;��H;��H;�H;�H;5�H;��H;��H;,�H;��H;2�H;��H;c�H;��H;��H;��H;P�H;-�H; �H;#�H;"�H;,�H;Q�H;��H;��H;��H;^�H;��H;,�H;��H;0�H;��H;��H;9�H;�H;��H;��H;��H;��H;��H;
�H;'�H;J�H;Y�H;��H;��H;��H;��H;��H;��H;x�H;6�H;��H; I;T I;      �I;�I;�I; I;�I;� I;��H;��H;��H;��H;��H;��H;�H;��H;g�H;�H;��H;��H;��H;��H;��H;��H;��H;�H;A�H;y�H;��H;u�H;��H;��H;.�H;��H;��H;g�H;T�H;A�H;5�H;B�H;P�H;h�H;��H;��H;.�H;��H;��H;q�H;��H;{�H;?�H; �H;��H;��H;��H;��H;��H;��H;��H;�H;g�H;��H;�H;��H;��H;��H;��H;��H; I;� I;�I;!I;�I;�I;      VI;:I;�I;UI;�I;�I;�I;�I; I;��H;G�H;��H;\�H;��H;y�H;��H;��H;�H;��H;��H;��H;v�H;q�H;v�H;��H;�H;V�H;��H;H�H;��H;h�H;�H;��H;��H;��H;g�H;`�H;g�H;��H;��H;��H;�H;i�H;��H;@�H;��H;V�H;�H;��H;q�H;z�H;t�H;��H;��H;��H;�H;��H;��H;v�H;��H;^�H;��H;K�H;��H;!I;�I;�I;�I;�I;[I;�I;6I;      rI;pI;I;rI;�
I;�	I;^I;
I;tI;�I;%I;H I;r�H;��H;��H;<�H;��H;��H;d�H;��H;��H;��H;d�H;R�H;h�H;��H;��H;4�H;��H;=�H;��H;L�H;�H;��H;��H;��H;��H;��H;��H;��H;�H;M�H;��H;<�H;��H;/�H;��H;��H;c�H;J�H;g�H;��H;��H;��H;b�H;��H;��H;<�H;��H;��H;t�H;F I;%I;�I;wI;	I;^I;�	I;�
I;yI;I;kI;      �I;�I;II;�I;zI;)I;�I;�I;
I;	I;�I;�I;�I;] I;)�H;�H;'�H;^�H;��H;��H;7�H;��H;��H;k�H;Q�H;C�H;��H;��H;)�H;��H;�H;��H;o�H;4�H;�H;��H;��H;��H;�H;6�H;o�H;��H;�H;��H;"�H;��H;��H;G�H;M�H;e�H;��H;��H;2�H;��H;��H;^�H;(�H;�H;+�H;] I;�I;�I;�I;	I;I; I;�I;%I;�I;�I;PI;�I;      �I;�I;�I;I;�I;HI;nI;aI;)I;�I;I;j
I;�I;I;�I; I;m�H;#�H;�H;�H;b�H;y�H;��H;��H;y�H;R�H;I�H;v�H;��H;�H;��H;=�H;��H;��H;c�H;@�H;1�H;C�H;_�H;��H;��H;?�H;��H;�H;��H;u�H;I�H;X�H;v�H;��H;��H;x�H;\�H;�H;�H;!�H;m�H; I;�I; I;�I;i
I;I;�I;(I;]I;rI;:I;�I;$I;�I;�I;      �!I;�!I;0"I;?"I;�!I;!I;�I;GI;�I;�I;�I;mI;I;�
I;�I;�I;�I;��H;0�H;��H;��H;��H;��H;�H;��H;q�H;D�H;F�H;��H;��H;"�H;��H;@�H;��H;��H;��H;��H;��H;��H;��H;A�H;��H;#�H;��H;��H;B�H;F�H;u�H;��H;�H;��H;��H;��H;��H;3�H;��H;�I;�I;�I;�
I;I;jI;�I;�I;�I;HI;�I;!I;�!I;?"I;0"I;�!I;      ��H;?�H;xI;�	I;�I;�I;VI;� I;�!I;U I;kI;�I;�I;�I;I;<
I;�I;UI;0 I;'�H;p�H;.�H;�H;�H;/�H;��H;{�H;]�H;F�H;s�H;��H;3�H;��H;r�H;5�H;�H;��H;�H;2�H;t�H;��H;3�H;��H;u�H;B�H;[�H;|�H;��H;)�H;�H;�H;-�H;m�H;(�H;3 I;NI;�I;<
I;I;�I;�I;�I;oI;W I;�!I;� I;VI;�I;�I;�	I;�I;?�H;      �NH;�TH;�dH;�}H;ۛH;V�H;��H;��H;�I;I;  I;!I;mI;/I;�I;I;�I;�I;�I;hI;�H;�H;k�H;H�H;�H;@�H;��H;��H;N�H;M�H;��H;��H;U�H;��H;��H;��H;x�H;��H;��H;��H;V�H;��H;��H;M�H;J�H;}�H;��H;F�H;�H;C�H;s�H;�H;�H;jI;�I;�I;�I;I;�I;.I;mI;!I;  I;I;�I;��H;��H;Q�H;�H;�}H;�dH;�TH;      PIF;oYF;��F;��F;{'G;ǈG;��G;CH;"�H;C�H;]�H;�I;�I;� I;�I;�I;�I;I;K
I;I;@I;��H;k�H;��H;_�H;7�H;C�H;��H;�H;\�H;I�H;��H;�H;�H;7�H;�H;
�H;�H;4�H;}�H;�H;��H;J�H;\�H;x�H;��H;F�H;:�H;]�H;��H;q�H;��H;=I;I;M
I;�I;�I;�I;�I;� I;�I;�I;^�H;F�H;�H;CH;��G;��G;�'G;��F;��F;bYF;      �DA;�kA;J�A;h�B;�jC;QaD;{\E;�IF;�G;��G;`NH;/�H;��H;�I;vI;Z I;�I;:I;�I;�I;�I;�I;�H;��H;��H;Y�H;�H;2�H;��H;y�H;O�H;h�H;��H;B�H;��H;��H;��H;��H;��H;E�H;��H;h�H;T�H;{�H;��H;/�H;�H;_�H;��H;��H;�H;�I;�I;�I;�I;6I;�I;[ I;xI;�I;��H;,�H;]NH;��G;�G;�IF;}\E;CaD;�jC;h�B;H�A;�kA;      �J6;��6;��7;�9;;;;.=;Ij?;V�A; �C;M2E;��F;O�G;r<H;|�H;��H;�I;G I;I;#I;5I;�I;�I;2I;/�H;��H;��H;?�H;�H;!�H;��H;k�H;X�H;w�H;�H;��H;S�H;-�H;T�H;��H;�H;z�H;X�H;n�H;��H;�H;�H;C�H;��H;��H;-�H;4I;�I;�I;6I;&I;I;H I;�I;��H;~�H;q<H;L�G;��F;P2E;�C;P�A;Hj?;.=;S;;�9;��7;�6;      p ;�!;�#;�&;�*;�o.;_3;��7;b�;;j?;8kB;�D;kxF;��G;�cH;
�H;�
I;�I;QI;aI;I;I;�I;9I;�H;j�H;n�H;�H;��H;��H;��H;h�H;t�H;��H;;�H;�H;��H;�H;5�H;��H;u�H;h�H;��H;��H;��H;�H;s�H;o�H;�H;7I;�I;I;I;bI;SI;�I;�
I;�H;�cH;��G;mxF;�D;8kB;j?;_�;;��7;_3;�o.;�*;�&;�#;�!;      Yt�:� �:!l�:>�;� 
;ڄ;$z;P$;K�,;��3;�9;�>;�B;2E;�F;PH;խH;��H;I;�I;$I;]I;I;�I;�I;��H;�H;3�H;��H;y�H;��H;��H;r�H;��H;�H;��H;��H;��H;�H;��H;v�H;��H;��H;}�H;��H;0�H;�H;��H;�I;�I;I;]I;%I;�I;
I;��H;׭H;PH;�F;2E;�B; �>;	�9;��3;K�,;P$; z;;� 
;0�;'l�:{ �:      (�>:��G:��b:p��:#��:�4�:�*�:~i;>�;�a;*;Br3;��:;�!@;��C;�IF;��G;��H;
�H;VI;�I;!I;I;�I;�I;6I;��H;n�H;��H;Z�H;-�H;��H;}�H;��H;��H;��H;f�H;��H;��H;��H;~�H;��H;2�H;^�H;��H;n�H;��H;7I;�I;�I;I;I;�I;WI;�H;��H;��G;�IF;��C;�!@;��:;?r3;*;�a;:�;�i;�*�:�4�:G��:n��:��b:T�G:      (���څ��uk��� �����-69��!:�Ȋ:v4�:��:��;�;D�,;��6;��=;��B;n�E;V�G;�|H;u�H;ZI;�I;_I;7I;�I;I;eI;*�H;��H;�H;��H;��H;��H;��H;��H;m�H;W�H;n�H;��H;��H;��H;��H;��H;�H;��H;*�H;jI;I;�I;:I;cI;�I;XI;u�H;�|H;S�G;o�E;��B;��=;��6;D�,;�;��;��:l4�:�Ȋ:��!: -698��ܙ �uk�䅍�      %/��&����x���X���/�� ���� o치9�9��k:��:)o�:�B;�&;C3;r<;�A;�pE;@tG;�|H;�H;	I;QI;#I;�I;J
I;�I;3 I;.�H;�H;��H;a�H;��H;��H;��H;X�H;F�H;Z�H;��H;��H;��H;b�H;��H;�H;-�H;3 I;�I;H
I;�I;&I;QI;I;�H;�|H;@tG;�pE;�A;n<;A3;�&;�B;)o�:��:��k:�9�9�n����� ���/���X�!�x�$���      ������q
����4�׻�+��Ȯ���;��lۺ8� � P�9�Ȋ:��:�;!;��0;;;��A;�pE;S�G;��H;��H;�I;I;3I;�I;�I;UI;��H;%�H;^�H;��H;�H;��H;��H;I�H;�H;J�H;��H;��H; �H;��H;^�H;&�H;��H;VI;�I;�I;.I;I;�I;��H;��H;T�G;�pE;��A;;;��0;!;�;��:�Ȋ:(P�9<� ��lۺ�;�ɮ���+��4�׻����q
���      ����p8����?�k���O��3/�/B�	�׻ȵ��g�@�RP����$�>:�4�:��;Vb;��/;;;�A;k�E;��G;ԭH;�
I;G I;�I;�I;�I;�I;�I;h�H; �H;��H;}�H;��H;��H;R�H;�H;R�H;��H;��H;{�H;��H;!�H;i�H;�I;�I;�I;�I;�I;E I;�
I;ѭH;��G;n�E;�A;;;��/;Tb;��;�4�:(�>:0��NP��i�@�Ƶ��
�׻0B��3/���O�A�k���p8��      :���|�1�ݼ��˼d���,���}��G����D�һ����e���/�d:(׳:�;Ob;��0;n<;��B;�IF;OH;�H;�I;S I;�I;I;9
I;�I; I;�H;;�H;��H;�H;�H;]�H;�H;]�H;�H;�H;��H;9�H;�H; I;�I;:
I;I;�I;M I;�I;�H;NH;�IF;��B;m<;��0;Rb;�;&׳:h:�/�i������D�һ����G��}��,��d����˼3�ݼ�|�      E�B�LR?��5���&��3��J��ԮҼ F����?=�!?�.����/��nk���9"׳:��;!;=3;��=;��C;�F;�cH;��H;rI;�I;�I;I;�I;�I;'�H;��H;v�H;f�H;$�H;g�H;�H;h�H;!�H;d�H;v�H;��H;%�H;�I;�I;I;�I;�I;lI;��H;�cH; �F;��C;��=;93;!;��;׳:���9�nk���/�.��!?�@=���!F��ԮҼ�J���3���&��5�MR?�      (��%W��蒐�$�����j�Q`I���&����Cϼ�,���T[�l�mI��d;��nk�x:�4�:�;�&;��6;�!@;2E;��G;��H;�I;� I;2I;�I;�
I;I;X I;��H;��H;��H;C�H;w�H;*�H;z�H;?�H;��H;��H;��H;V I;I;�
I;�I;/I;� I;�I;��H;��G;2E;�!@;��6;�&;�;�4�:h:�nk�e;�nI��l��T[��,��Cϼ�����&�Q`I���j�$���蒐�%W��      �J�����D��ͽ���'�������L�%��%��	;���k����lI����/��/� �>:��:�B;D�,;��:;�B;pxF;y<H;��H;�I;qI;�I;!I;�I;�I;r�H;\�H;�H;R�H;��H;Q�H;��H;P�H;�H;Z�H;p�H;�I;�I; I;�I;qI;�I;��H;u<H;pxF;�B;��:;G�,;�B;��: �>:�/���/�mI������k�	;��%��%����L����'������ͽ�D����      Q�:��*7���,�+���	�q�齂��� W����j�?�/��J���I���k�l�.��e��H���Ȋ:-o�:�;Jr3;�>;	�D;Q�G;+�H;�I;!I;�I;lI;c
I;�I;B I;��H;�H;��H;��H;E�H;��H;��H;~�H;��H;B I;�I;g
I;mI;�I;!I;�I;$�H;P�G;�D;��>;=r3;�;#o�:�Ȋ:H��i��.��m��k��I���J��?�/���j�!W������q�齂�	�+���,��*7�      ^���p����1�l���M���,�Xl�Q9ݽ�A���{���5��J��	;���T[�!?�����bP���O�9��:��;*;�9;9kB;��F;ZNH;Z�H;  I;kI;�I;I;�I;%I;H�H;��H;��H;��H;O�H;��H;��H;��H;H�H;"I;�I;I;�I;lI;�I;W�H;WNH;��F;8kB;�9;*;��;��:�O�9\P������"?��T[�
;���J����5��{��A��Q9ݽXl���,���M�1�l����p��      4m־P�Ѿ�>ľ����ӗ����{��I�+�����V���{�>�/�%���,��?=�C�һm�@�T� ���k:��:�a;��3;j?;T2E;��G;C�H;I;Q I;�I;�I;	I;�I;��H;��H;��H;��H;=�H;��H;��H;��H;��H;�I;	I;�I;�I;R I;I;B�H;��G;Q2E;j?;��3;�a;��:��k:T� �n�@�D�һ@=��,��&��?�/��{��V�����+��I���{�ӗ�������>ľP�Ѿ      C\����r5��z ��E۾ֳ�^��y�Z�L?#����A����j�%��Dϼ�����˵���lۺp9�9l4�:B�;G�,;X�;; �C;�G;"�H;�I;�!I;�I;(I;I;wI;(I;��H;��H;��H;	�H;��H;��H;��H;&I;xI;	I;)I;�I;�!I;�I;#�H;�G; �C;X�;;F�,;:�;l4�:X9�9�lۺ̵�������Dϼ%����j��A�����L?#�y�Z�^��ֳ��E۾�z �r5����      E�b��>]���M�Î6�����$���>ľ"q��y�Z�+�Q9ݽ!W����L����!F���G��׻;�0o칄Ȋ:�i;P$;��7;X�A;�IF;CH;��H;� I;GI;ZI;�I;I;�I;��H;��H;v�H;��H;v�H;��H;��H;�I;I;�I;`I;GI;� I;��H;	CH;�IF;T�A;��7;P$;xi;�Ȋ:Ho�;��׻�G�"F�������L�!W��Q9ݽ+�y�Z�"q���>ľ�$�����Î6���M��>]�      p��񲗿���6�y�{�R���)�nv��>ľ^���I�Xl����������&�ԮҼ�}�0B�ή�������!:�*�:$z;Y3;Kj?;t\E;��G;��H;LI;�I;pI;�I;[I;�I;��H;��H;F�H;��H;F�H;��H;��H;�I;]I;�I;tI;�I;LI;��H;��G;r\E;Kj?;\3; z;�*�:��!:���ή��0B��}�ծҼ��&��������Xl��I�^���>ľnv���)�{�R�6�y����񲗿      �˿�<ƿpL��@1����>]���)��$��ֳ���{���,�q��'��Q`I��J���,���3/�,��� �0-69�4�:҄;�o.;.=;@aD;��G;S�H;�I;!I;EI;1I;�	I;�I;� I;��H;��H;H�H;��H;��H;� I;�I;�	I;-I;HI;!I;�I;T�H;��G;?aD;.=;�o.;΄;�4�: -69� �,���3/��,���J��Q`I�'��q�齤�,���{�ֳ��$����)��>]��@1��pL���<ƿ      ����<���U[忶˿�T���{�R�����E۾ӗ����M���	������j��3�d����O�<�׻��/�P��?��:� 
;�*;P;;�jC;~'G;؛H;�I;�!I;�I;{I;�
I;�I;�I;#�H;��H;��H;��H;&�H;�I;�I;�
I;xI;�I;�!I;�I;ۛH;�'G;�jC;P;;�*;� 
;1��:8����/�<�׻��O�d���3���j������	���M�ӗ���E۾���{�R���T���˿U[�<���      O�6��t����˿@1��6�y�Î6��z �����1�l�+��ͽ$�����&���˼@�k�$�����X��� �z��:7�;�&;}9;m�B;��F;�}H;�	I;5"I;I;�I;I;XI;)I;��H;�H;h�H;�H;��H;'I;YI;�I;�I;$I;6"I;�	I;�}H;��F;j�B;~9;�&;5�;n��:�� ���X�#���@�k���˼��&�$����ͽ+�1�l������z �Î6�6�y�@1���˿���t�6��      ��*��g&��#�t�U[�pL�������M�r5��>ľ����,��D�蒐��5�2�ݼ���q
��x� uk���b:%l�:�#;ɗ7;W�A;��F;�dH;�I;&"I;�I;KI;I;�I;�I;��H;]�H;��H;Y�H;��H;�I;�I;I;GI;�I;&"I;�I;�dH;��F;T�A;×7;�#;l�:��b:uk��x��q
���2�ݼ�5�蒐��DὪ�,����>ľr5���M����pL��U[�t��#��g&�      ��8��4��g&�6��<����<ƿ񲗿�>]����P�Ѿ�p���*7����%W��LR?� }�r8�������օ����G:s �:�!;�6;�kA;fYF;�TH;G�H;�!I;�I;�I;nI;/I;�I;A I;��H;��H;��H;A I;�I;-I;oI;�I;�I;�!I;J�H;�TH;rYF;�kA;�6;�!;k �:|�G:Ѕ�� �����r8�� }�LR?�%W�����*7��p��P�Ѿ����>]�񲗿�<ƿ<���6���g&��4�      ��$������꿯�ſ�ޞ�%3s��2�=����� j���yHͽŸ����'�B<ͼq�n�e���AQ^��-.�p��:mW;_S%;ho8;��A;DF;�H;~�H;��H;��H;%�H;�H;(�H;��H;��H;��H;�H;��H;��H;��H;&�H;�H;"�H;��H;��H;~�H;�H;DF;��A;bo8;VS%;gW;h��:�-.�CQ^�e���r�n�B<ͼ��'�Ÿ��yHͽ�� j���=����2�%3s��ޞ���ſ������$�      $�������忇�����cm�V�-�����Qh��Vde�"-�תɽ�v��(�$���ɼ{mj�8���X�$���ņ:gx;�%;4�8;FB;"RF;�H;�H;�H;��H;I�H;�H;�H;|�H;��H;��H;�H;��H;��H;{�H;�H;�H;E�H;��H;�H;�H;�H;*RF;CB;.�8;�%;ax;�ņ: ��X�8���{mj���ɼ(�$��v��תɽ"-�Vde�Qh������V�-�cm��������忝����      ����������ԿLw�����:�\�"����k��Y0X�����;����w����������]� ���F�����ɒ:��;�';��9;�oB;�zF;�!H;u�H;��H;�H;s�H;�H;!�H;��H;��H;��H;��H;��H;��H;��H;�H;�H;o�H;�H;��H;t�H;�!H;�zF;�oB;��9;��';��;�ɒ:����F�!�黬�]����������w��;�����Z0X�k�����"�:�\����Lw���Կ��𿝏�      ������Կp���ޞ�_F�h�C�-E�"�;�I��D���"��f�c�|��֯���J��ѻѢ)��K���:
�
;�M*;n�:;�C;ʸF;�8H;/�H;M�H;\�H;��H;�H;!�H;��H;��H;��H;��H;��H;��H;��H;�H;�H;��H;b�H;K�H;+�H;�8H;иF;�C;j�:;�M*;�
;��:�K�Ӣ)��ѻ��J��֯�|�f�c�"����D��I��"�;-E�h�C�_F��ޞ�p���Կ��      ��ſ���Lw���ޞ�����>�W�5�%�����hɰ��|x�g{+�ұ����J��  �ζ��Z�1�(���+� 
9��:��;�-;��<;^�C;�G;�TH;'�H;��H;��H;��H;0�H;�H;j�H;��H;{�H;��H;v�H;��H;h�H;�H;,�H;��H;��H;��H;&�H;�TH;�G;[�C;��<;۷-;��;��:@ 
9"+�)���[�1�϶���  ��J���ұ�g{+��|x�hɰ�����5�%�>�W������ޞ�Lw�����      �ޞ�������_F�>�W�W�-���?Kɾ�G����O����ƽƸ��΄-���ۼㄼ64�ǐ�϶�]:��:;|�1;�c>;E�D;y\G;0sH;z�H;8�H;G�H; �H;N�H;�H;L�H;o�H;c�H;��H;^�H;n�H;I�H;�H;M�H;��H;K�H;5�H;x�H;-sH;\G;B�D;�c>;x�1;|;��:]:϶�ǐ�64�ㄼ��ۼ΄-�Ƹ��ƽ�����O��G��?Kɾ��W�-�>�W�_F�������      %3s�cm�:�\�h�C�5�%����TҾj��
 j��C(����^P����[�|������Y�;��eX�l�<���k:6��:�� ;ԟ5;2R@;8uE;ѲG;�H;#�H;��H;��H;$�H;J�H;�H;E�H;R�H;=�H;q�H;:�H;P�H;E�H;
�H;G�H; �H;��H;��H; �H;�H;ղG;6uE;0R@;ҟ5;�� ;$��: �k:p�<�fX�;����Y����|���[�^P����콪C(�
 j�j���TҾ��5�%�h�C�:�\�cm�      �2�U�-�"�-E�����?Kɾj����s�8�5���v㻽�v��	z0��;��+���*����26�@BS�GM�:O�	;p�(;�9;�/B;JDF;"H;��H;_�H;��H;��H;N�H;g�H;��H;�H;�H;!�H;=�H;�H;"�H;�H;��H;d�H;M�H;��H;��H;]�H;��H;#H;JDF;�/B;�9;p�(;F�	;MM�:@BS�26�����*��+���;�	z0��v��v㻽��8�5���s�j��?Kɾ����-E�"�U�-�      =����������"�;hɰ��G��	 j�7�5��	�ΪɽY����J�s���沼��]�����	x�V	��n:���:�v;��/;d-=;��C;�F;�HH;��H;�H;��H;�H;~�H;j�H;��H;��H;��H;��H;	�H;��H;��H;��H;��H;j�H;~�H;�H;��H;�H;|�H;�HH;�F;��C;g-=;��/;�v;���:n:^	���	x������]��沼s���J�Y���Ϫɽ�	�7�5�
 j��G��hɰ�"�;��徶���      ��Qh��k���I���|x���O��C(���Ϫɽ����QDX�I��'<ͼ	ㄼ�X!��s���W��uK���:�y;��#;�H6;R@;�PE;h�G;\�H;��H;
�H;��H;��H;��H;X�H;��H;��H;��H;��H;��H;��H;��H;��H;��H;T�H;��H;��H;��H;�H;��H;[�H;k�G;�PE;R@;�H6;��#;�y;��: vK��W��s���X!�	ㄼ'<ͼI��RDX�����Ϊɽ���C(���O��|x��I��k��Ph��       j�Vde�Z0X�D�f{+�������v㻽Y���RDX������ۼ˾����;�H>ۻ#X�x�y��>":���:��;��-;��;;��B;mzF;�H;`�H;Z�H;��H;��H;��H;��H;Q�H;��H;~�H;u�H;��H;_�H;��H;w�H;��H;��H;M�H;��H;��H;��H;�H;X�H;]�H;�H;kzF;��B;��;;��-;��;���:�>":h�y�"X�H>ۻ��;�˾����ۼ���RDX�Y���v㻽��콂��g{+�D�Z0X�Vde�      ��"-������ѱ�ƽ^P���v���J�H����ۼ��d�J������+���rѺ�'
9�M�:��;p $;��5;��?;\�D;@\G;�eH;��H;��H;��H;��H; �H;��H;6�H;V�H;=�H;6�H;H�H;�H;H�H;6�H;@�H;T�H;3�H;��H;�H;��H;��H;��H;��H;�eH;>\G;b�D;��?;��5;z $;��;�M�: (
9�rѺ�+������d�J�����ۼI���J��v��^P��ƽұ轄����"-�      yHͽ֪ɽ�;��"����Ƹ����[�	z0�s��&<ͼ˾��d�J�����j���*���ਂ:4b�:6�;��/;}L<;�C;mF;m�G;ۡH;��H;��H;��H;�H;2�H;��H;�H;�H;��H;��H;��H;��H;��H;��H;��H;�H;�H;��H;9�H; �H;��H;��H;��H;ߡH;m�G;mF;�C;~L<;��/;;�;,b�:訂:��*��j�����c�J�˾��'<ͼs��	z0���[�Ƹ����"���;��֪ɽ      ĸ���v����w�f�c��J�΄-�|��;缅沼ㄼ��;������j���5�����>Q:.��:Li;�M*;d�8;d�@;�PE;�uG;iH;��H;��H;��H;��H;��H;W�H;��H;��H;��H;��H;��H;��H;��H;��H;��H;��H;��H;��H;��H;_�H;��H;�H;��H;��H;��H;iH;�uG;�PE;d�@;l�8;�M*;Ki;8��:�>Q:x�깧5��j��������;�ㄼ�沼�;�|�΄-��J�g�c���w��v��      ��'�(�$����|��  ���ۼ����+����]��X!�F>ۻ�+���*������>:���:��; �%;Ο5;v�>;�(D;��F;R!H;�H;)�H;��H;��H;��H;��H;M�H;��H;��H;m�H;p�H;M�H;8�H;S�H;6�H;L�H;s�H;m�H;��H;��H;T�H;��H;��H;��H;��H;-�H;�H;U!H;��F;�(D;~�>;ҟ5;�%;��;���:��>:x��*��+��D>ۻ�X!���]��+�������ۼ�  �|����(�$�      @<ͼ�ɼ�����֯�ζ��ㄼ��Y��*�����s��X��rѺ���>Q:���:��
;1�#;O�3;qc=;�#C;DF;��G;�H;��H;��H;�H;��H;5�H;��H;G�H;p�H;G�H;�H;4�H;��H;��H;��H;��H;��H;4�H;�H;D�H;t�H;L�H;�H;:�H;��H;�H;��H;��H;�H;��G;DF;�#C;tc=;K�3;3�#;��
;���:�>Q:���rѺX��s������*���Y�ㄼ϶���֯�����~�ɼ      m�n�xmj���]���J�Z�1�54�6������	x��W�P�y��'
9ꨂ:8��:��;6�#;:�2;�<;KpB; �E;��G;�eH;��H;�H;��H;��H;��H;��H;�H;*�H;�H;��H;��H;��H;��H;��H;��H;��H;��H;��H;��H;��H;�H;.�H;�H;��H;��H;��H;��H;�H;��H;�eH;��G;�E;NpB;�<;;�2;6�#;��;<��:訂:P(
9D�y��W��	x����8��44�Z�1���J���]�vmj�      X���4��� ���ѻ#���ǐ�]X�,6�Z	���uK��>":�M�:&b�:Hi;�%;H�3;߆<;*0B;��E;R\G;�HH;!�H;v�H;>�H;��H;�H;�H;��H;��H;��H;��H;��H;��H;E�H;8�H;8�H;�H;7�H;7�H;F�H;��H;��H;��H;�H;��H;��H;�H;�H;��H;<�H;v�H;$�H;�HH;Y\G;��E;(0B;�<;I�3; �%;Ii;*b�:�M�:�>":�uK�L	��,6�bX�ǐ�����ѻ��4���      .Q^�X��F�Ϣ)�%+��ζ�H�<�@AS� n:��:���:��;8�;�M*;ҟ5;tc=;KpB;��E;�JG;,8H;I�H;d�H;��H;�H;b�H;��H;r�H;��H;��H;��H;v�H;]�H;8�H;��H;��H;��H;��H;��H;��H;��H;7�H;Z�H;y�H;��H;��H;��H;p�H;��H;g�H;�H;��H;h�H;N�H;28H;�JG;��E;OpB;sc=;ԟ5;�M*;;�;��;���:��:4n: AS�T�<��ζ�"+�آ)��F�X�       ..�H����깰~K��
9,]:,�k:AM�:���:�y;��;v $;��/;j�8;��>;�#C;�E;]\G;08H;��H;��H;��H;l�H;�H;e�H;1�H;��H;��H;��H;e�H;�H;��H;��H;��H;�H;x�H;]�H;r�H;|�H;��H;��H;��H;�H;d�H;��H;��H;��H;.�H;k�H;�H;j�H;��H;��H;��H;38H;Y\G;�E;�#C;��>;j�8;��/;~ $;��;�y;���:QM�: �k:@]:P 
9�K����h��      ���:�ņ:�ɒ:��:��:��:$��:I�	;�v;��#;��-;��5;yL<;c�@;�(D;DF;��G;�HH;K�H;��H;��H;'�H;��H;=�H;��H;l�H;��H;��H;A�H;�H;��H;��H;V�H;H�H;�H;�H;�H;	�H;�H;H�H;S�H;��H;��H;�H;A�H;��H;��H;l�H;��H;;�H;��H;+�H;��H;��H;N�H;�HH;��G;DF;�(D;a�@;}L<;��5;·-;��#;�v;H�	;0��:��:��:��:�ɒ:�ņ:      jW;ux;��;�
;��;�;�� ;n�(;��/;�H6;��;;��?;�C;�PE;��F;��G;�eH;'�H;h�H;��H;,�H;��H;�H;��H;?�H;b�H;k�H;J�H;��H;��H;��H;/�H;��H;��H;��H;��H;��H;��H;��H;��H;��H;)�H;��H;��H;��H;L�H;g�H;e�H;C�H;��H;�H;��H;/�H; �H;j�H;%�H;�eH;��G;��F;�PE;�C;��?;��;;�H6;��/;t�(;�� ;z;��;�
;��;jx;      vS%;�%;��';�M*;׷-;��1;ޟ5;��9;k-=;R@;��B;b�D;mF;�uG;X!H;�H;��H;{�H;��H;j�H;��H;�H;��H;H�H;`�H;W�H;�H;��H;��H;{�H;	�H;��H;��H;��H;n�H;Y�H;:�H;T�H;m�H;��H;��H;��H;�H;y�H;��H;��H;�H;Z�H;d�H;F�H;��H;�H;��H;l�H;��H;y�H;��H;�H;Y!H;�uG;mF;f�D;��B;R@;n-=;��9;ܟ5;��1;�-;�M*;��';��%;      bo8;8�8;��9;j�:;z�<;�c>;.R@;�/B;��C;�PE;izF;=\G;l�G;iH;�H;��H;�H;B�H;
�H;�H;;�H;��H;C�H;S�H;I�H;)�H;��H;��H;S�H;��H;��H;��H;F�H;�H;�H;�H;��H;	�H;�H;�H;D�H;��H;��H;��H;P�H;��H;��H;-�H;M�H;Q�H;B�H;��H;>�H;�H;
�H;?�H;�H;��H;�H;iH;l�G;A\G;pzF;�PE;��C;�/B;0R@;�c>;��<;i�:;��9;.�8;      ��A;CB;�oB;�C;S�C;S�D;@uE;JDF;�F;l�G;�H;�eH;ߡH;��H;0�H;��H;��H;��H;n�H;q�H;�H;E�H;d�H;S�H;�H;��H;��H;Y�H;��H;��H;`�H;2�H;��H;��H;��H;��H;��H;��H;��H;��H;��H;.�H;d�H;��H;��H;Y�H;��H;��H;�H;Q�H;e�H;H�H;�H;o�H;q�H;��H;��H;��H;4�H;��H;�H;�eH;�H;n�G;�F;KDF;@uE;I�D;d�C;�C;�oB;CB;      DF;,RF;�zF;ŸF;�G;�\G;ԲG;,H;�HH;`�H;`�H;��H;��H;��H;��H;�H;��H;�H;��H;.�H;o�H;a�H;V�H;0�H;��H;t�H;H�H;��H;��H;T�H;�H;��H;��H;��H;f�H;U�H;b�H;P�H;c�H;��H;��H;��H;	�H;T�H;��H;��H;E�H;y�H;��H;.�H;W�H;d�H;r�H;0�H;��H;�H;��H;�H;��H;��H;��H;��H;h�H;b�H;�HH;,H;ղG;x\G;�G;иF;�zF;*RF;      �H;H;�!H;�8H;�TH;-sH;"�H;��H;|�H;��H;X�H;��H;��H;��H;��H;��H;��H;�H;u�H;��H;��H;h�H;�H;��H;��H;D�H;��H;x�H;<�H;�H;��H;��H;U�H;8�H;!�H; �H;�H;��H;�H;9�H;W�H;��H;��H;�H;7�H;w�H;��H;L�H;��H;��H;�H;l�H;��H;��H;v�H;�H;��H;��H;��H;��H;��H;��H;[�H;��H;{�H;��H;�H;'sH;�TH;�8H;�!H;�H;      ��H;	�H;q�H;5�H;�H;{�H;+�H;]�H;�H;�H;�H;��H;��H; �H;��H;8�H;��H;��H;��H;��H;��H;F�H;��H;��H;P�H;��H;t�H;J�H;��H;��H;h�H;=�H;�H;��H;��H;��H;��H;��H;��H;��H;�H;;�H;h�H;��H;��H;H�H;r�H;��H;V�H;��H;��H;J�H;��H;��H;��H;��H;��H;;�H;��H;�H;��H;��H;�H;�H;�H;`�H;.�H;o�H;(�H;6�H;q�H;��H;      ��H;�H;��H;\�H;��H;5�H;��H;��H;��H;��H;��H;��H;�H;��H;��H;�H; �H;��H;��H;��H;H�H;��H;��H;R�H;��H;��H;3�H;��H;��H;a�H;*�H;��H;��H;��H;��H;��H;v�H;��H;��H;��H;��H;��H;-�H;_�H;��H;��H;2�H;��H;��H;O�H;��H;��H;H�H;��H;��H;��H;!�H;�H;��H;��H;�H;��H;��H;��H;��H;��H;��H;0�H;��H;_�H;��H;�H;      ��H;��H;�H;S�H;��H;A�H;��H;��H;�H;��H;��H;�H;5�H;_�H;N�H;I�H;/�H;��H;��H;e�H;�H;��H;u�H;��H;��H;H�H;�H;��H;a�H;#�H;��H;��H;��H;��H;`�H;E�H;7�H;B�H;]�H;��H;��H;��H;��H; �H;_�H;��H;��H;O�H;��H;��H;y�H;��H;�H;d�H;��H;��H;2�H;M�H;N�H;\�H;8�H;�H;��H;��H;�H;��H;��H;C�H;��H;X�H;�H;��H;      '�H;^�H;z�H;��H;��H;��H;$�H;T�H;��H;��H;��H;��H;��H;��H;��H;v�H;!�H;��H;z�H;%�H;��H;��H;�H;��H;_�H;�H;��H;j�H;/�H;��H;��H;}�H;o�H;8�H;�H; �H;�H;�H;�H;;�H;s�H;}�H;��H;��H;+�H;i�H;��H;�H;c�H;��H;�H;��H;��H;"�H;|�H;��H;$�H;z�H;��H;��H;��H;��H;��H;��H;��H;S�H;.�H;��H;��H;��H;z�H;]�H;      �H;�H;�H;�H;$�H;D�H;G�H;g�H;m�H;U�H;N�H;9�H;�H;��H;��H;J�H;��H;��H;`�H;��H;��H;/�H;��H;��H;/�H;��H;�H;=�H;��H;��H;v�H;[�H;:�H;�H;��H;��H;��H;��H;��H;�H;?�H;Z�H;u�H;��H;��H;=�H;��H;��H;2�H;��H;��H;2�H;��H;��H;a�H;��H;��H;M�H;��H;��H;�H;7�H;T�H;X�H;m�H;g�H;O�H;F�H;2�H;�H; �H;�H;      /�H;#�H;(�H;�H;�H;�H;�H;��H;��H;��H;��H;Y�H;�H;��H;o�H;�H;��H;��H;<�H;��H;`�H;�H;��H;F�H;��H;��H;U�H;�H;��H;��H;l�H;<�H;��H;��H;��H;��H;��H;��H;��H;��H;��H;>�H;k�H;��H;��H;�H;U�H;��H;��H;F�H;��H;�H;\�H;��H;<�H;��H;��H;!�H;o�H;��H;�H;Y�H;��H;��H;��H;��H;
�H;��H;�H;�H;0�H;"�H;      {�H;u�H;��H;x�H;d�H;>�H;D�H;�H;��H;��H;��H;D�H;�H;��H;w�H;9�H;��H;H�H;��H;��H;P�H;��H;~�H;�H;��H;��H;2�H;��H;��H;��H;3�H;
�H;��H;��H;��H;��H;��H;��H;��H;��H;��H;�H;3�H;}�H;��H;��H;5�H;��H;��H;�H;��H;��H;L�H;��H;��H;J�H;��H;9�H;v�H;��H;�H;C�H;��H;��H;��H;�H;I�H;;�H;k�H;y�H;��H;�H;      ��H;��H;��H;��H;��H;a�H;U�H;#�H;��H;��H;~�H;A�H;�H;��H;S�H;��H;��H;8�H;��H;��H;�H;��H;j�H;�H;��H;\�H;�H;��H;��H;b�H;�H;��H;��H;��H;��H;��H;��H;��H;��H;��H;��H;��H;�H;[�H;��H;��H;�H;_�H;��H;�H;p�H;��H;�H;|�H;��H;;�H;��H;��H;S�H;��H;�H;A�H;��H;��H;��H;%�H;Z�H;c�H;��H;��H;��H;��H;      ��H;��H;��H;��H;h�H;V�H;A�H;�H;��H;��H;��H;M�H;��H;��H;6�H;��H;��H;5�H;��H;v�H;�H;��H;Q�H;�H;��H;I�H;��H;��H;��H;I�H;�H;��H;��H;��H;��H;��H;��H;��H;��H;��H;��H;��H;�H;C�H;��H;��H;��H;L�H;��H;�H;X�H;��H;�H;r�H;��H;:�H;��H;��H;6�H;��H;��H;K�H;��H;��H;��H;!�H;I�H;W�H;m�H;��H;��H;��H;      �H;�H;
�H;��H;��H;��H;t�H;=�H;	�H;��H;g�H;%�H;��H;��H;Z�H;��H;��H;�H;��H;e�H;�H;��H;:�H;��H;��H;[�H;�H;��H;|�H;?�H;�H;��H;��H;��H;��H;��H;{�H;��H;��H;��H;��H;��H;�H;:�H;u�H;��H;�H;^�H;��H;��H;?�H;��H;	�H;a�H;��H;�H;��H;��H;X�H;��H;��H;$�H;j�H;��H;�H;>�H;{�H;��H;��H;��H;
�H;�H;      ��H;��H;��H;��H;j�H;Y�H;@�H;�H;��H;��H;��H;M�H;��H;��H;6�H;��H;��H;5�H;��H;v�H;�H;��H;Q�H;�H;��H;I�H;��H;��H;��H;H�H;�H;��H;��H;��H;��H;��H;��H;��H;��H;��H;��H;��H;�H;B�H;��H;��H;��H;M�H;��H;�H;V�H;��H;�H;r�H;��H;:�H;��H;��H;6�H;��H;��H;J�H;��H;��H;��H;"�H;E�H;V�H;m�H;��H;��H;��H;      ��H;��H;��H;��H;��H;^�H;U�H;%�H;��H;��H;|�H;A�H;�H;��H;T�H;��H;��H;:�H;��H;��H;"�H;��H;j�H;�H;��H;\�H;�H;��H;��H;a�H;�H;��H;��H;��H;��H;��H;��H;��H;��H;��H;��H;��H;�H;[�H;��H;��H;�H;a�H;��H;�H;p�H;��H;�H;|�H;��H;;�H;��H;��H;P�H;��H;�H;C�H;~�H;��H;��H;)�H;\�H;^�H;��H;��H;��H;��H;      |�H;u�H;�H;|�H;e�H;A�H;B�H;�H;��H;��H;��H;C�H;�H;��H;w�H;9�H;��H;J�H;��H;��H;P�H;��H;~�H;�H;��H;��H;5�H;��H;��H;��H;3�H;�H;��H;��H;��H;��H;��H;��H;��H;��H;��H;
�H;1�H;~�H;��H;��H;4�H;��H;��H;�H;��H;��H;I�H;��H;��H;I�H;��H;;�H;w�H;��H;�H;C�H;��H;��H;��H;�H;K�H;>�H;m�H;|�H;��H;v�H;      -�H;)�H;*�H;�H;�H;�H;�H;��H;��H;��H;��H;[�H;�H;��H;p�H; �H;��H;��H;?�H;��H;a�H;�H;��H;F�H;��H;��H;T�H;�H;��H;��H;k�H;;�H;��H;��H;��H;��H;��H;��H;��H;��H;��H;>�H;k�H;��H;��H;�H;T�H;��H;��H;C�H;��H;�H;Y�H;��H;>�H;��H;��H; �H;m�H;��H;�H;X�H;��H;��H;��H;��H;�H;�H;�H;"�H;3�H;#�H;      �H;�H;�H;	�H;"�H;N�H;M�H;d�H;j�H;U�H;Q�H;9�H;�H;��H;��H;M�H;��H;��H;`�H;��H;��H;2�H;��H;��H;2�H;��H;�H;?�H;��H;��H;u�H;X�H;;�H;�H;��H;��H;��H;��H;��H;�H;<�H;Z�H;s�H;��H;��H;;�H;~�H;��H;/�H;��H;��H;2�H;��H;��H;`�H;��H;��H;J�H;��H;��H;�H;9�H;Q�H;U�H;j�H;d�H;O�H;C�H;%�H;�H;�H;�H;      �H;[�H;v�H;��H;��H;��H;&�H;T�H;�H;��H;��H;��H;��H;��H;��H;x�H;$�H;��H;|�H;#�H;��H;��H;	�H;��H;c�H;�H;��H;j�H;1�H;��H;��H;~�H;p�H;:�H;�H;�H;�H; �H;�H;;�H;r�H;~�H;��H;��H;*�H;i�H;��H;�H;_�H;��H;�H;��H;��H;"�H;|�H;��H;$�H;w�H;��H;��H;��H;��H;��H;��H;��H;U�H;*�H;��H;��H;��H;|�H;Z�H;      ��H;��H;	�H;^�H;��H;M�H;��H;��H;�H;��H;��H;�H;6�H;^�H;Q�H;J�H;1�H;��H;��H;g�H;�H;��H;t�H;��H;��H;H�H;�H;��H;b�H;$�H;��H;��H;��H;��H;`�H;C�H;7�H;E�H;]�H;��H;��H;��H;��H;!�H;^�H;��H;�H;N�H;��H;��H;|�H;��H;�H;b�H;��H;��H;/�H;J�H;P�H;\�H;5�H;�H;��H;��H;�H;��H;��H;?�H;��H;c�H;�H;��H;      ��H;�H;	�H;X�H;��H;:�H;��H;��H;��H;��H;��H;��H;�H;��H;��H;�H;�H;��H;��H;��H;J�H;��H;��H;S�H;��H;��H;2�H;��H;��H;_�H;*�H;��H;��H;��H;��H;��H;v�H;��H;��H;��H;��H;��H;+�H;a�H;��H;��H;5�H;��H;��H;K�H;��H;��H;E�H;��H;��H;��H;�H;�H;��H;��H;�H;��H;��H;��H;��H;��H;��H;3�H;��H;V�H;�H;
�H;      ��H;��H;c�H;5�H;�H;��H;-�H;f�H;�H;�H;�H;��H;��H; �H;��H;;�H;��H;��H;��H;��H;��H;I�H;��H;��H;W�H;��H;r�H;H�H;��H;��H;h�H;=�H;�H;��H;��H;��H;��H;��H;��H;��H;�H;=�H;i�H;��H;��H;G�H;u�H;��H;R�H;��H;��H;I�H;��H;��H;��H;��H;��H;:�H;��H; �H;��H;��H;�H;�H;�H;`�H;+�H;t�H;$�H;5�H;m�H;��H;      �H;H;�!H;�8H;�TH;1sH;"�H;��H;~�H;��H;Z�H;��H;��H;��H;��H;��H;��H;"�H;u�H;��H;��H;k�H;�H;��H;��H;D�H;��H;x�H;<�H;�H;��H;��H;T�H;8�H;#�H;��H;�H;��H;�H;9�H;U�H;��H;��H;�H;7�H;w�H;��H;K�H;��H;��H;�H;k�H;��H;��H;u�H;�H;��H;��H;��H;��H;��H;��H;X�H;��H;{�H;��H;$�H;,sH;�TH;�8H;�!H;�H;      DF;)RF;�zF;ŸF;�G;�\G;ѲG;.H;�HH;_�H;e�H;��H;��H;��H;��H;�H;��H;�H;��H;.�H;r�H;b�H;T�H;0�H;��H;r�H;E�H;��H;��H;T�H;�H;��H;��H;��H;h�H;Q�H;e�H;T�H;c�H;��H;��H;��H;�H;T�H;��H;��H;I�H;v�H;��H;-�H;X�H;b�H;o�H;.�H;��H;�H;��H;�H;��H;��H;��H;��H;d�H;`�H;�HH;&H;ϲG;x\G;�G;ŸF;vzF;RF;      ��A;?B;�oB;�C;V�C;V�D;@uE;KDF;�F;n�G;�H;�eH;ߡH;��H;4�H;��H;��H;��H;p�H;n�H;�H;H�H;b�H;S�H;�H;��H;��H;Y�H;��H;��H;b�H;3�H;��H;��H;��H;��H;��H;��H;��H;��H;��H;3�H;f�H;��H;��H;V�H;��H;��H;�H;P�H;g�H;H�H;�H;o�H;r�H;��H;��H;��H;4�H;��H;�H;�eH;�H;n�G;�F;KDF;?uE;I�D;^�C;�C;�oB;?B;      >o8;�8;��9;u�:;t�<;�c>;2R@;�/B;��C;�PE;mzF;A\G;l�G;iH;�H;��H;�H;C�H;�H;�H;>�H;��H;A�H;S�H;M�H;&�H;��H;��H;U�H;��H;��H;��H;F�H;�H;�H;�H;��H;�H;�H;�H;H�H;��H;��H;��H;R�H;��H;��H;*�H;J�H;Q�H;C�H;��H;>�H;�H;�H;>�H;�H;��H;�H;iH;k�G;>\G;lzF;�PE;��C;�/B;1R@;�c>;��<;��:;��9;�8;      _S%;��%;�';�M*;ӷ-;|�1;؟5;��9;r-=;R@;��B;f�D;mF;�uG;[!H;�H;��H;}�H;��H;j�H;��H;�H;��H;H�H;d�H;S�H;�H;��H;��H;x�H;�H;��H;��H;��H;p�H;Y�H;=�H;Y�H;m�H;�H;��H;��H;�H;|�H;��H;��H;�H;W�H;a�H;E�H;��H;�H;��H;l�H;��H;y�H;��H;�H;[!H;�uG;mF;b�D;��B;
R@;n-=;��9;؟5;|�1;Է-;�M*;�';��%;      fW;ux;��;�
;��;�;�� ;t�(;��/;�H6;��;;��?;�C;�PE;��F;��G;�eH;'�H;g�H; �H;.�H;��H;�H;��H;E�H;^�H;i�H;L�H;��H;��H;��H;0�H;��H;��H;��H;��H;��H;��H;��H;��H; �H;2�H;��H;��H;��H;J�H;l�H;d�H;A�H;��H;�H;��H;.�H;�H;j�H;%�H;�eH;��G;��F;�PE;�C;��?;��;;�H6;��/;t�(;�� ;n;��;�
;��;kx;      ���:�ņ:�ɒ:��:��:���:0��:L�	;�v;��#;��-;��5;zL<;a�@;�(D;DF;��G;�HH;K�H;��H;��H;+�H;��H;=�H;��H;i�H;��H;��H;B�H;�H;��H;��H;U�H;K�H;�H;�H;�H;�H;�H;H�H;V�H;��H;��H;�H;A�H;��H;��H;k�H;��H;=�H;��H;(�H;��H;��H;M�H;�HH;��G;DF;�(D;a�@;}L<;��5;·-;��#;�v;M�	;2��:��:��:��:�ɒ:�ņ:      �-.�4�����p~K��
9H]:,�k:]M�:���:�y;��;~ $;��/;h�8;��>;�#C;�E;\\G;08H;��H;��H; �H;j�H;�H;k�H;.�H;��H;��H;��H;a�H;�H;��H;��H;��H;�H;t�H;`�H;u�H;|�H;��H;��H;��H;"�H;e�H;��H;��H;��H;0�H;g�H;�H;m�H;��H;��H;��H;28H;Y\G;�E;�#C;��>;h�8;��/;z $;��;�y;���:OM�:�k: ]:` 
9@K����@��      -Q^�X��F�̢)�)+��ζ�T�<��@S�4n:��:���:��;9�;�M*;֟5;uc=;MpB;��E;�JG;08H;N�H;g�H;��H;�H;i�H;��H;p�H;��H;��H;��H;w�H;]�H;8�H;��H;��H;��H;��H;��H;��H;��H;8�H;^�H;z�H;��H;��H;��H;s�H;��H;c�H;
�H;��H;e�H;M�H;28H;�JG;��E;MpB;sc=;ԟ5;�M*;8�;��;���:��:,n:@@S�X�<��ζ�&+�̢)��F�X�      `���.���"���ѻ"���ǐ�[X�%6�N	���uK��>":�M�:,b�:Ii;!�%;K�3;�<;)0B;��E;X\G;�HH;$�H;z�H;>�H;��H;�H;�H;��H;��H;��H;��H;��H;��H;H�H;8�H;7�H;�H;:�H;5�H;H�H;��H;��H;��H;��H;��H;��H;�H;�H;��H;<�H;y�H;!�H;�HH;Y\G;��E;(0B;��<;I�3; �%;Ii;&b�:�M�:�>":�uK�L	��)6�^X�ǐ�!����ѻ&��1���      m�n�xmj���]���J�Y�1�44�8������	x��W�L�y�`(
9ꨂ:<��:��;9�#;<�2;�<;KpB;�E;��G;�eH;��H;�H;��H;��H;��H;��H;�H;*�H;�H;��H;��H;��H;��H;��H;��H;��H;��H;��H;��H;��H;�H;-�H;�H;��H;��H;��H;��H;�H;��H;�eH;��G;�E;KpB;�<;;�2;8�#;��;<��:ꨂ:0(
9D�y��W��	x����9��44�[�1���J���]�wmj�      ?<ͼ�ɼ�����֯�ζ��ㄼ��Y��*�����s��X��rѺ���>Q:���:��
;2�#;K�3;sc=;�#C;	DF;��G;�H;��H;��H;�H;��H;5�H;�H;G�H;t�H;I�H;�H;9�H;��H;��H;��H;��H;��H;5�H;�H;I�H;t�H;J�H; �H;8�H;��H;�H;��H;��H;��H;��G;DF;�#C;qc=;H�3;3�#;��
;���:�>Q:���rѺX��s������*���Y�ㄼ϶���֯������ɼ      ��'�(�$����|��  ���ۼ����+����]��X!�F>ۻ�+��~*�x����>:���:��;�%;П5;|�>;�(D;��F;\!H;�H;-�H;��H;��H;��H;��H;N�H;��H;��H;m�H;t�H;M�H;5�H;S�H;6�H;L�H;t�H;l�H;��H;��H;P�H;��H;��H;��H;��H;*�H;�H;X!H;��F;(D;~�>;Ο5;�%;��;���:��>:x�깁*��+��F>ۻ�X!���]��+�������ۼ�  �|����(�$�      Ÿ���v����w�f�c��J�΄-�|��;缅沼ㄼ��;������j���5�H�� ?Q:8��:Ki;�M*;h�8;j�@;�PE;�uG;iH;��H;��H;��H; �H;��H;Z�H;��H;��H;��H;��H;��H;��H;��H;��H;��H;��H;��H;��H;��H;^�H;��H; �H;��H;��H;��H;iH;�uG;�PE;`�@;j�8;�M*;Ki;8��:�>Q:x�깧5��j��������;�ㄼ�沼�;�|�΄-��J�f�c���w��v��      yHͽ֪ɽ�;��"����Ƹ����[�	z0�s��&<ͼʾ��c�J�����j��z*���訂:0b�:8�;��/;�L<;�C;mF;r�G;�H;��H;��H;��H; �H;5�H;��H;�H;�H;�H;��H;��H;��H;��H;��H;��H;�H;�H;��H;9�H; �H;��H;��H;��H;ۡH;m�G;mF;�C;wL<;��/;5�;,b�:訂:��~*��j�����d�J�˾��'<ͼs��	z0���[�Ƹ����"���;��֪ɽ      ��"-������ұ�ƽ^P���v���J�H����ۼ��d�J������+���rѺ(
9�M�:��;x $;��5;��?;d�D;C\G;�eH;��H;��H;��H;��H; �H;��H;5�H;Y�H;@�H;6�H;F�H;�H;H�H;5�H;?�H;V�H;5�H;��H;�H;��H;��H;��H;��H;�eH;A\G;d�D;��?;��5;z $;��;�M�:(
9�rѺ�+������d�J�����ۼH���J��v��^P��ƽұ轄����"-�       j�Vde�Z0X�D�f{+�������v㻽Y���RDX������ۼ˾����;�F>ۻ X�l�y��>":���:��;ķ-;��;;��B;mzF;�H;a�H;Z�H;�H;��H;��H;��H;Q�H;��H;��H;t�H;��H;`�H;��H;t�H;�H;��H;N�H;��H;��H;��H;�H;X�H;^�H;�H;mzF;��B;�;;��-;��;���:�>":h�y�#X�H>ۻ��;�˾����ۼ���RDX�Y���v㻽��콂��g{+�D�Z0X�Vde�      ��Ph��k���I���|x���O��C(���Ϫɽ����QDX�H��'<ͼ	ㄼ�X!��s���W��uK���:�y;�#;�H6;R@;�PE;l�G;]�H;��H;
�H;��H;��H;��H;V�H;��H;��H;��H;��H;��H;��H;��H;��H;��H;U�H;��H;��H;��H;�H;��H;\�H;h�G;�PE;R@;�H6;��#;�y;��:�uK��W��s���X!�	ㄼ'<ͼI��QDX�����Ϫɽ���C(���O��|x��I��k��Ph��      =����������"�;hɰ��G��	 j�8�5��	�ΪɽY����J�s���沼��]�����	x�\	�� n:���:�v;��/;g-=;��C;�F;�HH;~�H;��H;��H;�H;��H;j�H;��H;��H;��H;��H;
�H;��H;��H;��H;��H;k�H;~�H;�H;��H;�H;�H;�HH;�F;��C;h-=;��/;�v;���:n:Z	���	x������]��沼s���J�Y���Ϊɽ�	�8�5�
 j��G��hɰ�"�;��徶���      �2�U�-�"�-E�����?Kɾj����s�8�5���v㻽�v��	z0��;��+���*����66��AS�IM�:P�	;p�(;�9;�/B;MDF; H;��H;]�H;��H;��H;P�H;g�H;��H;�H;�H;�H;=�H;�H;!�H;�H;��H;f�H;N�H;��H;��H;_�H;��H;%H;HDF;�/B;�9;p�(;H�	;MM�:�BS�26�����*��+���;�	z0��v��v㻽��8�5���s�j��?Kɾ����-E�"�U�-�      %3s�cm�:�\�h�C�5�%����TҾj��
 j��C(����^P����[�|������Y�:��fX�l�<� �k:6��:�� ;ԟ5;2R@;8uE;ѲG;�H; �H;��H;��H;&�H;J�H;�H;E�H;O�H;:�H;q�H;9�H;P�H;D�H;
�H;J�H;#�H;��H;��H;#�H;�H;ֲG;5uE;2R@;֟5;�� ;(��:�k:t�<�fX�:����Y����|���[�^P����콪C(�
 j�j���TҾ��5�%�h�C�:�\�cm�      �ޞ�������_F�>�W�W�-���?Kɾ�G����O����ƽƸ��΄-���ۼㄼ54�ǐ�϶�$]:���:};|�1;�c>;E�D;x\G;.sH;z�H;8�H;J�H;�H;Q�H;�H;L�H;n�H;`�H;��H;`�H;m�H;K�H;�H;Q�H;��H;M�H;:�H;}�H;1sH;�\G;D�D;�c>;z�1;z;��: ]:
϶�ǐ�64�ㄼ��ۼ΄-�Ƹ��ƽ�����O��G��?Kɾ��W�-�>�W�_F�������      ��ſ���Lw���ޞ�����>�W�5�%�����hɰ��|x�g{+�ұ����J��  �ζ��Z�1�)���+�@ 
9��:��;߷-;��<;^�C;�G;�TH;&�H;��H;��H;��H;/�H;�H;k�H;��H;y�H;��H;u�H;��H;g�H;�H;/�H;��H;��H;��H;*�H;�TH;�G;[�C;��<;ܷ-;��;��:@ 
9"+�(���[�1�ζ���  ��J���ұ�g{+��|x�hɰ�����5�%�>�W������ޞ�Lw�����      ������Կp���ޞ�_F�h�C�-E�"�;�I��D���"��f�c�|��֯���J��ѻϢ)��K�!��:�
;�M*;m�:;�C;ȸF;�8H;.�H;K�H;[�H;��H;�H;�H;��H;��H;��H;��H;��H;��H;��H;!�H;�H;��H;c�H;N�H;/�H;�8H;ѸF;�C;m�:;�M*;�
;��:�K�Ӣ)��ѻ��J��֯�|�f�c�"����D��I��"�;-E�h�C�`F��ޞ�p���Կ��      ����������ԿLw�����:�\�"����k��Z0X�����;����w����������]�!���F�����ɒ:��; �';��9;�oB;�zF;�!H;u�H;��H;�H;u�H;�H;�H;��H;��H;��H;��H;��H;��H;��H;�H;�H;p�H;�H;��H;x�H;�!H;�zF;�oB;��9;��';��;�ɒ:����F� �黬�]����������w��;�����Z0X�k�����"�:�\����Lw���Կ��𿝏�      $�������忇�����cm�V�-�����Qh��Vde�"-�תɽ�v��(�$���ɼ{mj�9���	X� ���ņ:gx;	�%;4�8;FB; RF;�H;�H;�H;��H;I�H;�H;�H;|�H;��H;��H;�H;��H;��H;{�H;�H;�H;E�H;��H;�H;�H; H;-RF;CB;0�8;�%;cx;�ņ:��X�8���|mj���ɼ(�$��v��תɽ"-�Vde�Qh������V�-�cm��������忝����      dܿ3�ֿ�aǿ=^��/���Yo���7����iþ�(���-=��` �A���_�0]�/p����I�R�ѻ��)���R���:0�
;�*;"�:;��B;�HF;+�G;�lH;��H;y�H;@�H;��H;��H;O�H;�H;�H;��H;	�H;}�H;O�H;��H;��H;<�H;��H;��H;�lH;+�G;IF;��B;�:;�*;,�
;��:`�R���)�R�ѻ��I�/p��0]��_�A���` ��-=��(���iþ����7�Yo�/���=^���aǿ3�ֿ      2�ֿCpѿ�¿������_Xi�Е3��
�UD��Fl��@�9��.���R�� \� �ex��0�E��ͻ�$�@ �ݍ�:>�;K�*;6�:;�B;�TF;��G;,nH;��H;·H;m�H;��H;��H;^�H;��H;!�H;��H;�H;��H;[�H;��H;��H;g�H;ɷH;��H;)nH;��G;�TF;�B;1�:;D�*;;�;э�:0 ��$��ͻ0�E�ex�� � \��R���.��@�9�Fl��VD���
�Е3�_Xi��������¿Cpѿ      �aǿ�¿����������"Y��f'�����7o���.}��k/����%ڟ�!<Q�-#�ע��(;�/���7�� h7���:�;r,;��;;�C;�vF;�G;�rH; �H;��H;�H;��H;��H;��H;��H;P�H;��H;G�H;��H;��H;��H;��H;�H;��H;�H;�rH;�G;wF;�C;��;;k,;�;��: d7�;��0����(;�ע�-#�!<Q�%ڟ�����k/��.}�7o�������f'��"Y�����������¿      =^������k���Yo���@�)�$�޾����8ce�0����ڽ󻒽 g@������R���O*�IG�����pC^9,��:;[d.;��<;��C;��F;��G;�yH;��H;�H;"�H;��H;n�H;��H;��H;��H;�H;�H;��H;��H;k�H;��H;�H;!�H;��H;�yH;��G;��F;��C;��<;Sd.; ;$��:�C^9���IG���O*��R������ g@�󻒽��ڽ0��9ce�����$�޾)���@�Yo�k�������      /����������Yo��!J�K�#��\��VD������zPH�����b��C��� +���ټ(����쿐����\�:$��:E�;�Y1;	>;�0D;}�F;bH;F�H;ƨH;�H;\�H;��H;�H;e�H;M�H;��H;b�H;��H;L�H;e�H;�H;��H;W�H;�H;ĨH;E�H;dH;��F;�0D;>;�Y1;C�;��:l�:������(����ټ� +� C���b�����zPH�����VD���\��K�#��!J�Yo��������      Yo�_Xi��"Y���@�K�#��
��о�A���i���(�~��vr���_��5��ɺ�p�`��<��f�d�`�\�L�X:�P�:�`;ȱ4;��?;��D;w8G;n0H;��H;n�H;u�H;�H;��H;��H;��H;��H;�H;��H;�H;��H;��H;��H;��H;�H;{�H;m�H;��H;m0H;|8G;��D;��?;±4;�`;�P�:T�X:l�\�f�d��<��q�`��ɺ��5��_�vr��~����(��i��A���о�
�K�#���@��"Y�_Xi�      ��7�Е3��f'�)��\���о�����.}��-=�{
���Ľ[��+:��������� �7�"GĻ$� O�����:�{;�D&;�+8;JA;�E;��G;~LH;�H;y�H;5�H;��H;�H;��H;��H;�H;��H;�H;��H;�H;��H;��H; �H;��H;;�H;x�H;�H;zLH;��G;�E;JA;�+8;�D&;�{;ÿ�: O��ă$�"GĻ�7���������+:�[����Ľ{
��-=��.}������о�\��)��f'�Е3�      ���
�����$�޾VD���A���.}�(�D�ht���ڽ�!��\����[�ļ�
v�<��ʿ���Iɺ�R�9���:(;�-;��;;��B;hIF;��G;fH;��H;�H;.�H;��H;i�H;��H;^�H;��H;��H;j�H;��H;��H;`�H;��H;d�H;��H;5�H;�H;��H;fH;��G;iIF;��B;��;;�-;(;���:�R�9�Iɺʿ��<���
v�[�ļ���\��!����ڽht�(�D��.}��A��VD��$�޾�����
�      �iþUD��7o�����������i��-=�ht� ���R��hys�z +����y񗼔(;�*�ѻ�s@���!�4j:�P�:��;�D3;1�>;FD;��F;�	H;;|H;��H;t�H;6�H;��H;��H;��H;�H;0�H;r�H;��H;o�H;2�H;�H;��H;��H;��H;;�H;t�H;��H;;|H;�	H;��F;FD;3�>;�D3;��;�P�:4j:��!��s@�+�ѻ�(;�y����z +�hys��R�� ��ht��-=��i���������7o��UD��      �(��Fl���.}�8ce�zPH���(�{
���ڽ�R�� �{�C�6�� �-p��_�`�ͨ��,��JIҺ@L^9���:٣;�~(;-�8;�IA;|E;jG;�=H;C�H;֬H;�H;_�H;(�H;m�H;��H;��H;��H;��H;M�H;��H;��H;��H;��H;j�H;(�H;f�H; �H;֬H;B�H;�=H;jG;|E;�IA;/�8;�~(;ߣ;���: L^9JIҺ�,��ͨ�_�`�-p��� �C�6� �{��R����ڽ{
���(�zPH�8ce��.}�Fl��      �-=�@�9��k/�0�����~��Ľ�!��hys�C�6�$#��ɺ��vz����A^��i�$��~�<�r:���:��;�Y1;�H=;&xC;'wF;�G;�eH;J�H;��H;��H;��H;Q�H;��H;��H;��H;e�H;z�H;��H;|�H;g�H;��H;��H;��H;P�H;��H;��H;��H;I�H;�eH;�G;$wF;)xC;�H=;�Y1;��;��:<�r:�~�i�$�A^������vz��ɺ�$#�C�6�hys��!����Ľ~���0���k/�@�9�      �` ��.�����ڽ�b��vr��[��\�z +�� ��ɺ�@��O*�Hͻ�5R�ǅ���:(��:��;�);�t8;b�@;U*E;m8G;>$H;<�H;E�H;��H;"�H;��H;n�H;b�H;�H;O�H;��H;��H;!�H;��H;��H;R�H;��H;`�H;n�H;��H;)�H;�H;>�H;<�H;?$H;j8G;Z*E;d�@;�t8;�);��;(��:̜:ǅ��5R�Fͻ�O*�?��ɺ�� �y +�\�[��vr���b����ڽ��.��      A���R��%ڟ�󻒽C���_�+:�������-p���vz��O*��4ֻk�0����09*�:
1;M� ;�D3;E�=;��C;�kF;��G;�\H;��H;O�H;�H;;�H;��H;w�H;��H;��H;	�H;��H;W�H;��H;U�H;��H;
�H;��H;��H;z�H;��H;>�H;�H;K�H;��H;�\H;��G;�kF;��C;D�=;�D3;R� ;1;4�: �09,���k��4ֻ�O*��vz�,p����輤��+:��_� C��󻒽%ڟ��R��      �_� \�!<Q� g@� +��5�����Z�ļy�]�`����Hͻk�Iɺ �6�<�:�P�:(�;�d.;C�:;!�A;'|E;vNG;C'H;��H;ƥH;]�H;��H;#�H;J�H;Z�H;4�H;��H;��H;�H;��H;��H;��H;�H;��H;��H;2�H;]�H;T�H;*�H;��H;[�H;åH; �H;C'H;{NG;*|E; �A;L�:;�d.;%�;�P�:<�: �6��Hɺk�Fͻ���]�`�x�Z�ļ�����5�� +�g@�!<Q�\�      /]� �-#�������ټ�ɺ������
v��(;�ͨ�?^���5R�2��� �6����:���:�;&�*;�+8;!@;V�D;`�F;��G;�eH;~�H;��H;��H;��H;��H;��H; �H;u�H;��H;d�H;{�H;,�H;Y�H;+�H;z�H;e�H;��H;p�H;#�H;��H;��H;��H;��H;��H;��H;�eH;��G;c�F;X�D;�!@;�+8; �*;��;���:���: �6�.����5R�=^��ͨ��(;��
v������ɺ���ټ����-#� �      ,p��dx��ע��R��(��q�`���7�:��*�ѻ�,��e�$�ǅ��09<�:���:�;�~(;�Z6;��>;ȨC;�HF;٠G;�DH;F�H;��H;��H;�H;)�H;�H;��H;��H;��H;��H;�H;��H;��H;��H;��H;��H;�H;��H;��H;��H;��H;�H;,�H;�H;��H;��H;F�H;�DH;ܠG;�HF;ϨC;��>;�Z6;�~(;�;���:<�:��09ǅ�b�$��,��(�ѻ:�� �7�n�`�)���R��ע�cx��      �I�.�E��(;��O*����<��GĻƿ���s@�:IҺ�~���:6�:�P�:��;�~(;	�5;�>;6C;-�E;wcG;8$H;�{H;7�H;�H;��H;��H;;�H;��H;�H;W�H;��H;P�H;��H;A�H;��H;��H;��H;?�H;��H;M�H;��H;Z�H;!�H;��H;;�H;��H;��H;�H;8�H;�{H;;$H;zcG;5�E;6C;�>;�5;�~(;��;�P�:6�:М:x~�6IҺ�s@�ſ�� GĻ�<�����O*��(;�,�E�      F�ѻ�ͻ.���DG��运�d�d���$��Iɺ��!��L^9H�r:��:1;&�;"�*;�Z6;�>;;�B;��E;�8G;�	H;�mH;�H;F�H;��H;b�H;��H;��H;H�H;��H;��H;x�H;��H;��H;��H;	�H;#�H;�H;��H;��H;��H;t�H;��H;�H;H�H;��H;��H;`�H;��H;G�H;�H; nH;�	H;�8G;��E;8�B;�>;�Z6;$�*;&�;1;$��:`�r:�L^9ą!��Iɺ��$�_�d�俐�FG��+����ͻ      m�)�+�$�:��������4�\��N�� S�94j:���:��:~�;R� ;�d.;�+8;��>;6C;��E;�)G;��G;dH;~�H;��H;\�H;��H;3�H;��H;��H;��H;��H;��H;J�H;}�H;b�H;��H;9�H;L�H;6�H;��H;`�H;z�H;F�H;��H;��H;��H;��H;��H;3�H;��H;_�H;��H;��H;dH;��G;�)G;��E;:C;��>;�+8;�d.;U� ;��;��:���:$4j: S�9�N��D�\����"���9��+�$�      ��R�� � ]7��D^9T�:X�X:׿�:���:�P�:�;��;�);�D3;J�:;�!@;ϨC;4�E;�8G;��G;�`H;l�H;�H;�H;x�H;8�H;0�H;L�H;^�H;��H;��H;��H;�H;��H;��H;/�H;o�H;e�H;j�H;-�H;��H;��H;	�H;��H;��H;��H;`�H;J�H;0�H;>�H;y�H;�H;�H;r�H;�`H;��G;�8G;4�E;ШC;�!@;I�:;�D3;�);��;�;�P�:���:Ͽ�:t�X:l�:�C^9 e7�P �      ��:���:��:��:��:�P�:�{;(;��;�~(;�Y1;�t8;B�=;�A;V�D;�HF;wcG;�	H;dH;k�H;E�H;ӶH;0�H;��H;��H;:�H;H�H;��H;#�H;��H;~�H;��H;U�H;��H;H�H;��H;��H;��H;I�H;��H;T�H;��H;��H;��H; �H;��H;D�H;9�H;��H;��H;.�H;ֶH;L�H;o�H;dH;�	H;zcG;�HF;Y�D;�A;E�=;�t8;�Y1;�~(;��;(;�{;�P�:��:��:��:���:      ,�
;I�;��;;A�;�`;�D&;�-;�D3;2�8;I=;b�@;��C;+|E;c�F;ߠG;>$H;nH;��H;�H;ֶH;��H;6�H;�H;d�H;��H;��H;r�H;i�H;�H; �H;��H;��H;!�H;g�H;��H;��H;��H;c�H;�H;��H;��H; �H;�H;g�H;s�H;��H;��H;j�H;�H;3�H;��H;ܶH;�H;��H;nH;A$H;ߠG;h�F;*|E;��C;i�@;I=;0�8;�D3;�-;�D&;�`;X�;
;�;<�;      �*;I�*;k,;jd.;�Y1;ӱ4;�+8;��;;:�>;�IA;0xC;\*E;�kF;�NG;��G;�DH;�{H;�H;��H;�H;/�H;5�H;��H;��H;��H;[�H;�H;��H;��H;��H;��H;p�H;��H;;�H;��H;��H;��H;��H;��H;=�H;��H;j�H;��H;��H;��H;��H;�H;_�H;��H;��H;��H;:�H;5�H;�H;��H;�H;�{H;�DH;��G;�NG;�kF;a*E;4xC;�IA;<�>;��;;�+8;α4;�Y1;hd.;k,;3�*;      �:;;�:;�;;��<;�>;��?;JA;��B;FD;|E;$wF;j8G;��G;E'H;�eH;K�H;:�H;L�H;_�H;u�H;��H;�H;��H;��H;�H;��H;��H;2�H;u�H;p�H;�H;��H;�H;\�H;}�H;��H;��H;��H;|�H;^�H;�H;��H;�H;o�H;r�H;4�H;��H;��H;�H;��H;��H;�H;��H;v�H;_�H;I�H;<�H;M�H;�eH;E'H;��G;m8G;+wF;|E;FD;��B;JA;��?;>;��<;��;;/�:;      ңB;�B;�C;��C;�0D;��D;��E;iIF;��F;jG;#�G;D$H;�\H;�H;��H;��H;$�H;��H;��H;C�H;��H;j�H;��H;�H;��H;o�H;��H;B�H;(�H;��H;��H;��H;-�H;q�H;��H;��H;��H;��H;��H;t�H;,�H;��H;��H;��H;'�H;C�H;��H;s�H;��H;�H;��H;p�H;��H;B�H;��H;��H;)�H;��H;��H;�H;�\H;I$H;$�G;jG;��F;iIF;��E;��D;�0D;��C;�C;�B;      �HF;�TF;wF;�F;s�F;8G;��G;��G;�	H;�=H;�eH;B�H;��H;ͥH;��H;��H;��H;e�H;3�H;/�H;=�H;��H;[�H;��H;m�H;��H; �H;�H;��H;C�H;��H;"�H;3�H;q�H;��H;��H;��H;��H;��H;q�H;4�H;�H;��H;C�H;��H;	�H;�H;��H;q�H;��H;\�H;��H;@�H;0�H;6�H;d�H;��H;��H;��H;ʥH;��H;C�H;fH;�=H;�	H;��G;��G;t8G;��F;��F;wF;�TF;      ;�G;��G;�G;��G;YH;m0H;�LH;fH;7|H;B�H;I�H;>�H;I�H;]�H;��H;�H;��H;��H;��H;L�H;L�H;��H;�H;��H;��H;�H;��H;��H;N�H;��H;��H;/�H;L�H;t�H;��H;��H;��H;��H;��H;v�H;R�H;/�H;��H;��H;M�H;��H;��H;&�H;��H;��H;�H;��H;P�H;L�H;��H;��H;��H;�H;��H;Z�H;K�H;B�H;L�H;A�H;7|H;fH;�LH;f0H;pH;��G;�G;��G;      �lH;,nH;�rH;�yH;:�H;��H;�H;��H;��H;۬H;��H;��H;��H;��H;��H;*�H;=�H;��H;��H;^�H;��H;o�H;��H;4�H;>�H;�H;��H;3�H;��H;��H;�H;;�H;^�H;d�H;�H;��H;��H;��H;}�H;g�H;`�H;7�H;�H;��H;��H;2�H;��H;�H;B�H;4�H;��H;s�H;��H;]�H;��H;��H;>�H;/�H;��H;��H;��H;��H;��H;ܬH;��H;��H;��H;��H;H�H;�yH;�rH;nH;      �H;��H;�H;��H;��H;k�H;}�H;�H;j�H;�H;��H;&�H;=�H;(�H;��H;�H;��H;O�H;��H;��H;(�H;f�H;��H;u�H;#�H;��H;F�H;��H;��H;�H;)�H;K�H;`�H;e�H;d�H;o�H;m�H;j�H;c�H;g�H;a�H;H�H;,�H;�H;��H;��H;F�H;��H;'�H;p�H;��H;g�H;(�H;��H;��H;L�H;��H;�H;��H;(�H;;�H;%�H;��H; �H;o�H;�H;|�H;d�H;¨H;��H;�H;��H;      {�H;��H;��H;�H;�H;p�H;4�H;-�H;6�H;`�H;��H;��H;��H;R�H;��H;��H;$�H;�H;��H;��H;��H;�H;��H;m�H;��H;9�H;��H;��H;�H;!�H;>�H;B�H;O�H;d�H;N�H;\�H;q�H;Y�H;I�H;d�H;P�H;@�H;@�H;!�H;�H;��H;��H;A�H;��H;j�H;��H;�H;��H;��H;��H; �H;&�H; �H;��H;O�H;��H;��H;��H;f�H;9�H;.�H;6�H;p�H;�H;�H;��H;��H;      C�H;��H;�H;%�H;U�H; �H;��H;��H;��H;*�H;T�H;v�H;~�H;a�H;&�H;��H;`�H;��H;��H;��H;��H;!�H;��H;�H;��H;��H;��H;
�H;-�H;D�H;U�H;N�H;=�H;@�H;a�H;O�H;/�H;K�H;]�H;A�H;A�H;N�H;V�H;B�H;,�H;	�H;��H;��H;��H;�H;��H;#�H;��H;��H;��H;��H;d�H;��H;&�H;`�H;��H;x�H;W�H;-�H;��H;��H;��H;��H;c�H;#�H;�H;��H;      ��H;��H;��H;��H;��H;��H;�H;g�H;��H;i�H;��H;e�H;��H;;�H;u�H;��H;��H;|�H;O�H;�H;��H;��H;k�H;��H;��H;�H;*�H;;�H;I�H;D�H;H�H;U�H;:�H;9�H;K�H;,�H;%�H;,�H;H�H;:�H;A�H;V�H;H�H;B�H;H�H;9�H;,�H;�H;��H;��H;r�H;��H;��H;�H;O�H;}�H;��H;��H;u�H;9�H;��H;g�H;��H;m�H;��H;i�H;	�H;��H;��H;��H;��H;��H;      ��H;��H;�H;l�H;�H;��H;��H;��H;��H;��H;��H;�H;�H;��H;��H;��H;V�H;�H;��H;��H;_�H;��H;��H;�H;-�H;/�H;N�H;e�H;d�H;S�H;:�H;>�H;D�H;>�H;�H;�H;L�H;�H;�H;@�H;E�H;>�H;9�H;N�H;a�H;c�H;O�H;3�H;0�H;�H;��H;��H;\�H;��H;��H;�H;W�H;��H;��H;��H;�H;�H;��H;��H;��H;��H;��H;��H;�H;g�H;�H;��H;      E�H;W�H;��H;��H;c�H;��H;��H;\�H;�H;��H;��H;Y�H;�H;��H;k�H;�H;��H;�H;d�H;��H;��H;"�H;7�H;W�H;q�H;k�H;o�H;e�H;d�H;e�H;9�H;:�H;>�H;)�H;�H;�H;&�H;�H;�H;)�H;A�H;9�H;9�H;a�H;a�H;a�H;r�H;n�H;t�H;V�H;@�H;!�H;��H;��H;c�H;�H;��H;�H;k�H;��H;�H;V�H;��H;��H;�H;]�H;��H;��H;l�H;��H;��H;b�H;      x�H;��H;��H;��H;W�H;��H;#�H;��H;3�H;��H;o�H;��H;��H;�H;��H;��H;G�H;��H; �H;3�H;N�H;c�H;��H;r�H;��H;��H;��H;}�H;d�H;O�H;W�H;L�H;�H;�H;#�H;�H;��H;�H;!�H;�H;"�H;N�H;V�H;H�H;`�H;y�H;��H;��H;��H;t�H;��H;c�H;I�H;-�H;��H;��H;K�H;��H;��H;�H;��H;��H;r�H;��H;6�H;��H;(�H;��H;W�H;��H;��H;��H;      �H; �H;J�H;~�H;��H;�H;��H;��H;m�H;��H;��H;��H;Z�H;��H;.�H;��H;��H;�H;9�H;m�H;��H;��H;��H;��H;��H;��H;�H;��H;o�H;^�H;I�H;0�H;!�H;�H;�H;�H;�H;�H;�H;"�H;"�H;0�H;H�H;Y�H;k�H;��H;��H;��H;��H;��H;��H;��H;��H;h�H;7�H;	�H;��H;��H;.�H;��H;X�H;��H;��H;��H;o�H;��H;��H;�H;��H;{�H;G�H;+�H;      ��H;��H;��H;�H;[�H;��H;�H;j�H;��H;M�H;��H;+�H;��H;�H;b�H;��H;��H;)�H;O�H;m�H;��H;��H;��H;��H;��H;��H;��H;��H;o�H;x�H;*�H;)�H;P�H;%�H;��H;�H;��H;�H;��H;&�H;S�H;*�H;*�H;r�H;k�H;��H;��H;��H;��H;��H;��H;��H;��H;g�H;O�H;*�H;��H;��H;`�H;�H;��H;*�H;��H;M�H;��H;k�H;!�H;��H;]�H;�H;��H;��H;      �H;!�H;F�H;}�H;��H;	�H;��H;��H;k�H;��H;}�H;��H;Z�H;��H;.�H;��H;��H;�H;9�H;m�H;��H;��H;��H;��H;��H;��H;�H;��H;q�H;]�H;I�H;2�H;"�H;�H;�H;�H;�H;�H;�H;�H;"�H;0�H;H�H;Y�H;k�H;��H;��H;��H;��H;��H;��H;��H;��H;h�H;7�H;	�H;��H;��H;.�H;��H;X�H;��H;��H;��H;n�H;��H;��H;�H;��H;��H;L�H;(�H;      k�H;��H;��H;��H;X�H;��H;#�H;��H;2�H;��H;n�H;��H;��H;�H;��H;��H;G�H;��H; �H;3�H;O�H;e�H;��H;t�H;��H;��H;��H;�H;d�H;N�H;V�H;N�H;!�H;�H;%�H;�H;��H;�H;!�H;�H;"�H;L�H;V�H;H�H;`�H;y�H;��H;��H;��H;r�H;��H;d�H;H�H;-�H;��H;��H;J�H;��H;��H;�H;��H;��H;n�H;��H;3�H;��H;(�H;��H;]�H;��H;��H;��H;      F�H;W�H;��H;��H;e�H;��H;��H;^�H;�H;��H;��H;U�H;�H;��H;l�H;�H;��H;�H;g�H;��H;��H;%�H;:�H;Z�H;u�H;k�H;q�H;d�H;e�H;e�H;9�H;;�H;>�H;)�H;�H;�H;&�H;�H;�H;)�H;@�H;:�H;7�H;a�H;`�H;c�H;q�H;m�H;o�H;S�H;@�H;"�H;��H;��H;d�H;�H;��H;�H;k�H;��H;�H;U�H;��H;��H;�H;`�H;��H;��H;l�H;��H;��H;X�H;      ��H;��H;�H;h�H;�H;��H;��H;��H;��H;��H;��H;�H;�H;��H;��H;��H;V�H;�H;��H;��H;`�H;��H;��H;�H;0�H;-�H;N�H;d�H;g�H;U�H;9�H;=�H;B�H;>�H;�H;�H;L�H;�H;�H;@�H;B�H;@�H;9�H;O�H;^�H;`�H;N�H;2�H;-�H;�H;��H;��H;X�H;��H;��H; �H;V�H;��H;��H;��H;�H;�H;��H;��H;��H;��H;��H;��H;�H;o�H;�H;��H;      y�H;��H;��H;��H;��H;��H;�H;f�H;��H;i�H;��H;e�H;��H;9�H;w�H;��H;��H;}�H;O�H;�H;��H;��H;n�H;��H;��H;�H;*�H;;�H;L�H;D�H;G�H;V�H;;�H;9�H;L�H;,�H;%�H;/�H;H�H;9�H;>�H;U�H;E�H;A�H;G�H;7�H;)�H;�H;��H;��H;t�H;��H;��H;�H;M�H;{�H;��H;��H;u�H;9�H;��H;e�H;��H;j�H;��H;f�H;�H;��H;��H;��H;��H;��H;      7�H;��H;�H;�H;\�H; �H;��H;��H;��H;*�H;U�H;v�H;�H;c�H;'�H;��H;b�H;��H;��H;��H;��H;$�H;��H;�H;��H;��H;��H;	�H;/�H;E�H;U�H;O�H;>�H;A�H;c�H;N�H;/�H;O�H;^�H;A�H;@�H;N�H;S�H;A�H;(�H;�H;��H;��H;��H;�H;��H;#�H;��H;��H;��H;��H;d�H;��H;&�H;`�H;~�H;v�H;T�H;*�H;��H;��H;��H;��H;i�H;)�H;�H;~�H;      ��H;��H;��H;�H;�H;{�H;5�H;4�H;:�H;c�H;��H;��H;��H;Q�H;��H;��H;$�H;�H;��H;��H;��H;�H;��H;m�H;��H;:�H;��H;��H;�H;#�H;@�H;B�H;L�H;d�H;N�H;Z�H;q�H;\�H;I�H;c�H;P�H;B�H;>�H;�H;	�H;��H;��H;?�H;��H;h�H;��H;�H;��H;��H;��H; �H;$�H;��H;��H;Q�H;��H;��H;��H;c�H;6�H;3�H;8�H;k�H;�H;!�H;��H;��H;      ��H;��H;+�H;��H;��H;q�H;{�H;�H;s�H;�H;��H;&�H;=�H;)�H;��H;�H;��H;P�H;��H;��H;+�H;i�H;��H;v�H;'�H;��H;F�H;��H;��H;�H;)�H;L�H;`�H;e�H;d�H;n�H;k�H;m�H;a�H;d�H;`�H;I�H;)�H;�H;��H;��H;F�H;��H;$�H;n�H;��H;i�H;(�H;��H;��H;L�H;��H;�H;��H;&�H;=�H;#�H;��H;�H;p�H;�H;�H;j�H;��H;��H;*�H;��H;      �lH;nH;�rH;�yH;5�H;��H;��H;��H;��H;ܬH;��H;��H;��H;��H;��H;-�H;=�H;��H;��H;]�H;��H;r�H;��H;7�H;C�H;�H;��H;2�H;��H;��H;�H;:�H;]�H;e�H;�H;��H;��H;��H;|�H;e�H;a�H;:�H;�H;��H;��H;/�H;��H;�H;>�H;0�H;��H;r�H;��H;]�H;��H;��H;>�H;-�H;��H;��H;��H;��H;��H;۬H;��H;��H;�H;��H;C�H;�yH;�rH;nH;      .�G;��G;�G;��G;gH;q0H;�LH; fH;:|H;B�H;J�H;B�H;H�H;[�H;��H;�H;��H;��H;��H;J�H;N�H;��H;�H;��H;��H;�H;��H;��H;O�H;��H;��H;2�H;N�H;u�H;��H;��H;��H;��H;��H;u�H;O�H;2�H;��H;��H;J�H;��H;��H;&�H;��H;��H;�H;��H;L�H;O�H;��H;��H;��H;�H;��H;Z�H;I�H;A�H;I�H;A�H;7|H;"fH;�LH;j0H;oH;��G;�G;��G;      �HF;�TF;wF;�F;|�F;�8G;��G;��G;�	H;�=H;fH;F�H;��H;˥H;��H;��H;��H;h�H;3�H;-�H;@�H;��H;X�H;��H;s�H;��H;�H;�H;��H;C�H;��H;#�H;4�H;r�H;��H;��H;��H;��H;��H;q�H;4�H;"�H;��H;D�H;��H;�H;"�H;��H;o�H;��H;\�H;��H;>�H;0�H;6�H;a�H;��H;��H;��H;ǥH;��H;B�H;fH;�=H;�	H;��G;��G;t8G;��F;�F;�vF;�TF;      ̣B;�B;�C;��C;�0D;��D;��E;jIF;��F;jG;#�G;I$H;�\H;�H;��H;¨H;%�H;��H;��H;A�H;��H;m�H;��H; �H;��H;m�H;��H;C�H;*�H;��H;��H;��H;,�H;r�H;��H;��H;��H;��H;��H;u�H;-�H;��H;��H;��H;(�H;B�H;��H;s�H;��H;�H;��H;n�H;��H;B�H;��H;��H;(�H;��H;��H;�H;�\H;E$H;!�G;jG;��F;hIF;��E;��D;�0D;��C;�C;�B;      ��:;!�:;x�;;�<;�>;ŧ?;JA;��B;FD;|E;'wF;n8G;��G;B'H;�eH;M�H;:�H;M�H;]�H;u�H;��H;�H;��H;��H;�H;��H;��H;4�H;u�H;m�H;�H;��H;�H;\�H;}�H;��H;��H;��H;{�H;]�H;�H;��H;�H;s�H;w�H;4�H;��H;��H;�H;��H;��H;�H;��H;y�H;`�H;J�H;<�H;M�H;�eH;C'H;��G;k8G;'wF;|E;FD;��B;JA;��?;>;�<;v�;;�:;      �*;>�*;^,;qd.;�Y1;ʱ4;�+8;��;;?�>;�IA;*xC;^*E;�kF;�NG;��G;�DH;�{H;�H;��H;�H;0�H;6�H;��H;��H;��H;Z�H;�H;��H;��H;��H;��H;p�H;��H;;�H;��H;��H;��H;��H;��H;:�H;��H;r�H;��H;��H;��H;��H;�H;^�H;��H;��H;��H;7�H;3�H;�H;��H;�H;�{H;�DH;��G;NG;�kF;\*E;-xC;�IA;<�>;��;;�+8;ȱ4;�Y1;rd.;`,;(�*;      (�
;I�;��;;D�;�`;�D&;�-;�D3;-�8;I=;i�@;��C;)|E;e�F;�G;>$H;nH;��H;�H;ڶH;��H;3�H;�H;m�H;��H;��H;u�H;i�H;�H;�H;��H;��H;!�H;d�H;��H;��H;��H;a�H;�H;��H;��H;$�H;
�H;j�H;u�H;��H;��H;g�H;�H;6�H;��H;ڶH;�H;��H;nH;?$H;�G;g�F;*|E;��C;d�@;I=;,�8;�D3;�-;�D&;�`;X�;�;�;@�;      ��:鍨:��:&��:
��:�P�:�{;(;��;�~(;�Y1;�t8;E�=;�A;[�D;�HF;ycG;�	H;dH;l�H;H�H;ֶH;.�H;��H;��H;7�H;E�H;��H;#�H;��H;~�H;��H;T�H;��H;I�H;��H;��H;��H;H�H;��H;U�H;��H;��H;��H;!�H;��H;I�H;9�H;��H;��H;/�H;նH;K�H;o�H;dH;�	H;zcG;�HF;Y�D;�A;E�=;�t8;�Y1;�~(;��;(;�{;�P�:,��: ��:��:Ǎ�:      P�R�p � d7��D^9\�:|�X:ۿ�:���:�P�:�;��;�);�D3;I�:;�!@;ҨC;4�E;�8G;��G;�`H;r�H;�H;�H;y�H;?�H;/�H;I�H;^�H;��H;��H;��H;�H;��H;��H;0�H;k�H;e�H;m�H;-�H;��H;��H;�H;��H;��H;��H;^�H;L�H;/�H;:�H;|�H;�H;�H;q�H;�`H;��G;�8G;7�E;ҨC;�!@;G�:;�D3;�);��;ߣ;�P�:���:Ͽ�:T�X:p�:D^9 a7�� �      l�)�*�$�<�����$���,�\��N�� S�9$4j:���:��:��;T� ;�d.;�+8;��>;7C;��E;�)G;��G;dH;��H;��H;]�H;��H;2�H;��H;��H;��H;��H;��H;I�H;}�H;b�H; �H;7�H;L�H;7�H;��H;b�H;}�H;J�H;��H;��H;��H;��H;��H;2�H;��H;_�H;��H;�H;dH;��G;�)G;��E;7C;��>;�+8;�d.;R� ;��;��:���:$4j:8S�9�N��@�\� ������B��&�$�      M�ѻ�ͻ2���CG��翐�Z�d���$��Iɺ̅!��L^9L�r:$��:1;$�;&�*;�Z6;�>;9�B;��E;�8G;�	H; nH;�H;G�H;��H;b�H;��H;��H;I�H;��H;��H;y�H;��H;��H;��H;�H;#�H;	�H;��H;��H;��H;y�H;��H;�H;K�H;��H;��H;a�H;��H;F�H;�H;�mH;�	H;�8G;��E;8�B;�>;�Z6;&�*;$�;1;"��:X�r:PL^9̅!��Iɺ��$�b�d�翐�EG��6����ͻ      �I�-�E��(;��O*����<�� GĻſ���s@�6IҺ�~�М:6�:�P�:��;�~(;�5;�>;6C;1�E;{cG;:$H;�{H;8�H;�H;��H;��H;9�H;��H;�H;[�H;��H;P�H;��H;C�H;��H;��H;��H;?�H;��H;M�H;��H;]�H;!�H;��H;;�H;��H;��H;�H;7�H;�{H;8$H;vcG;5�E;6C;�>;�5;�~(;��;�P�:6�:̜:�~�:IҺ�s@�ƿ��!GĻ�<�����O*��(;�,�E�      ,p��dx��ע��R��(��n�`���7�:��*�ѻ�,��d�$�ǅ��096�:���:�;�~(;�Z6;��>;ΨC;�HF;ޠG;�DH;I�H;��H;��H;�H;)�H;�H;��H;��H;��H;��H;�H;��H;��H;��H;��H;��H;�H;��H;��H;��H;��H;�H;,�H;�H;��H;��H;F�H;�DH;۠G;�HF;ϨC;~�>;�Z6;�~(;�;���:<�:�09ǅ�c�$��,��*�ѻ:�� �7�n�`�)���R��ע�dx��      /]� �.#�������ټ�ɺ������
v��(;�̨�>^���5R�,��� �6����:���:��;#�*;�+8;�!@;\�D;d�F;��G;�eH;��H;��H;��H;��H;��H;��H;$�H;u�H;��H;g�H;}�H;)�H;Y�H;+�H;z�H;h�H;��H;s�H;#�H;��H;��H;��H;��H;��H;�H;�eH;��G;d�F;T�D;�!@;�+8; �*;��;���:���: �6�0����5R�>^��ͨ��(;��
v������ɺ���ټ����.#� �      �_�\�!<Q� g@�� +��5�����Z�ļx�^�`����Dͻk��Hɺ �6�D�:�P�:&�;�d.;G�:;'�A;*|E;~NG;F'H;�H;ȥH;]�H;��H;*�H;N�H;^�H;6�H;��H;��H;�H;��H;��H;��H;�H;��H;��H;4�H;\�H;Q�H;)�H;��H;[�H;ĥH;��H;F'H;�NG;&|E;�A;L�:;�d.;%�;�P�:<�: �6��Hɺk�Fͻ���^�`�x�Y�ļ�����5�� +� g@�!<Q�\�      A���R��%ڟ�󻒽C���_�+:�������,p���vz��O*��4ֻk�$��� �090�:1;Q� ;�D3;K�=;��C;�kF;��G;�\H;��H;L�H; �H;@�H;��H;{�H;��H;��H;�H;��H;U�H;��H;W�H;��H;�H;��H;��H;z�H;��H;@�H; �H;K�H;��H;�\H;��G;�kF;��C;B�=;�D3;N� ;1;.�:�09,���k��4ֻ�O*��vz�-p����輤��+:��_� C��󻒽%ڟ��R��      �` ��.�����ڽ�b��vr��[��\�z +�� ��ɺ�?��O*�Fͻ�5R�ǅ�Ĝ:"��:��;�);�t8;f�@;^*E;n8G;B$H;@�H;A�H;�H;%�H;��H;r�H;b�H;�H;R�H;��H;��H;$�H;��H;��H;R�H;�H;b�H;o�H;��H;(�H;�H;@�H;>�H;>$H;m8G;_*E;c�@;�t8;�);��;"��:Ĝ:ǅ��5R�Fͻ�O*�?��ɺ�� �z +�\�[��vr���b����ڽ��.��      �-=�@�9��k/�0�����~��Ľ�!��hys�C�6�$#��ɺ��vz����>^��g�$��~�<�r:���:��;�Y1;�H=;-xC;(wF;�G;�eH;H�H;��H;��H;��H;T�H;��H;��H;��H;e�H;|�H;��H;|�H;e�H;��H;��H;��H;Q�H;��H;��H;��H;H�H;�eH;�G;'wF;+xC;�H=;�Y1;��;���:8�r:�~�i�$�A^������vz��ɺ�$#�C�6�hys��!����Ľ~���0���k/�@�9�      �(��Fl���.}�8ce�zPH���(�{
���ڽ�R�� �{�C�6�� �-p��^�`�̨��,��BIҺ L^9���:ޣ;�~(;-�8;�IA;|E;jG;�=H;B�H;֬H; �H;b�H;)�H;l�H;��H;��H;��H;��H;O�H;��H;��H;��H;��H;j�H;)�H;d�H;!�H;֬H;B�H;�=H;jG;|E;�IA;,�8;�~(;ޣ;���:L^9DIҺ�,��ͨ�^�`�-p��� �C�6� �{��R����ڽ{
���(�zPH�8ce��.}�Fl��      �iþVD��7o�����������i��-=�ht� ���R��hys�z +����y񗼔(;�*�ѻ�s@��!�4j:�P�:��;�D3;5�>;FD;��F;�	H;;|H;��H;v�H;7�H;��H;��H;��H;�H;/�H;n�H;��H;n�H;0�H;�H;��H;��H;��H;9�H;v�H;��H;<|H;�	H;��F;FD;5�>;�D3;��;�P�:�3j:�!��s@�*�ѻ�(;�y����z +�hys��R�� ��ht��-=��i���������7o��UD��      ���
�����$�޾VD���A���.}�(�D�ht���ڽ�!��\����[�ļ�
v�<��ʿ���IɺS�9���:(;�-;��;;��B;iIF;��G;fH;��H;�H;.�H;��H;i�H;��H;^�H;��H;��H;j�H;��H;��H;\�H;��H;f�H;��H;5�H;�H;��H;fH;��G;fIF;��B;��;;�-;(;���:�R�9�Iɺʿ��<���
v�[�ļ���\��!����ڽht�(�D��.}��A��VD��$�޾�����
�      ��7�Е3��f'�)��\���о�����.}��-=�{
���Ľ[��+:��������� �7� GĻŃ$�O�����:�{;�D&;�+8;JA;�E;��G;zLH;�H;y�H;5�H;��H;�H;��H;��H;�H;��H;�H;��H;�H;��H;��H;�H;��H;;�H;y�H;�H;}LH;��G;�E;JA;�+8;�D&;�{;ɿ�: O��Ń$�!GĻ�7���������+:�[����Ľ{
��-=��.}������о�\��)��f'�Е3�      Yo�_Xi��"Y���@�K�#��
��о�A���i���(�~��vr���_��5��ɺ�p�`��<��h�d�`�\�X�X:�P�:�`;ȱ4;��?;��D;t8G;k0H;��H;n�H;x�H;�H;��H;��H;��H;��H;�H;��H;�H;��H;��H;��H;��H;�H;{�H;p�H;��H;p0H;|8G;��D;��?;ȱ4;�`;�P�:`�X:l�\�h�d��<��p�`��ɺ��5��_�vr��~����(��i��A���о�
�K�#���@��"Y�_Xi�      /����������Yo��!J�K�#��\��VD������zPH�����b��C��� +���ټ(��������l�:&��:E�;�Y1;	>;�0D;z�F;aH;E�H;ŨH;�H;\�H;��H;�H;f�H;H�H;��H;`�H;��H;I�H;b�H;�H;��H;Z�H;�H;ƨH;F�H;hH;��F;�0D;	>;�Y1;D�;��:p�:���쿐���(����ټ� +� C���b�����zPH�����VD���\��K�#��!J�Yo��������      =^������k���Yo���@�)�$�޾����9ce�0����ڽ󻒽 g@������R���O*�IG������C^9.��:;Zd.;��<;��C;�F;��G;�yH;��H;�H;#�H;��H;l�H;��H;��H;��H;�H;��H;��H;��H;n�H;��H; �H;$�H;��H;�yH;��G;��F;��C;��<;Vd.;�;$��: D^9���HG���O*��R������ g@�󻒽��ڽ0��8ce�����$�޾)���@�Yo�k�������      �aǿ�¿����������"Y��f'�����7o���.}��k/����%ڟ�!<Q�-#�ע��(;�0���7�� g7���:�;q,;��;;�C;�vF;�G;�rH;�H;��H;�H;��H;��H;��H;��H;M�H;��H;I�H;��H;��H;��H;��H;�H;��H; �H;�rH;�G;wF;�C;��;;k,;�;��: a7�:��/����(;�ע�-#�!<Q�%ڟ�����k/��.}�7o�������f'��"Y�����������¿      3�ֿCpѿ�¿������_Xi�Е3��
�UD��Fl��@�9��.���R�� \� �ex��0�E��ͻ�$�@ �ߍ�:?�;K�*;6�:;�B;�TF;��G;,nH;��H;·H;m�H;��H;��H;]�H;��H; �H;��H;�H;��H;]�H;��H;��H;g�H;ɷH;��H;)nH;��G;�TF;�B;2�:;D�*;9�;э�: ��$��ͻ1�E�ex�� � \��R���.��@�9�Fl��VD���
�Е3�_Xi��������¿Cpѿ      �?��|h��=v��� ��7�X��O/�/y�@�;ఖ��+X����ѽ����_n;�[�������B(�ښ��V��`�e9�:�;�Y.;V�<;iWC;�ZF;��G;0H;7jH;:�H;H�H;��H;+�H;��H;[�H;��H;��H;��H;V�H;��H;(�H;�H;C�H;B�H;4jH;0H;��G;�ZF;bWC;Q�<;�Y.;�;�:��e9Z��ښ���B(�����\��_n;������ѽ���+X�ఖ�@�;/y��O/�7�X�� ��=v��|h��      |h��/���a�����y�VvS�pM+��v�9ɾ�����T� ]�\ν����x\8�����x��%�N���t��P�9s-�:j�;��.; �<;�nC;�dF;�G;�1H;�jH;��H;��H;͵H;k�H;��H;g�H;��H;��H;��H;g�H;��H;i�H;˵H;��H;��H;�jH;�1H;�G;�dF;�nC;�<;��.;d�;g-�:h�9x��M���%��x�����x\8�����\ν ]��T�����9ɾ�v�pM+�VvS���y�a���/���      =v��b���W ��`�h�6E�W��i���|㼾}���nH�ӈ�y�ý�Ȅ��s/��o��#�����$J��(кH	�9Xg�:�l;$0;!]=;ܲC;ڀF;r�G;6H;mH;(�H;��H;��H; �H;A�H;��H;
�H;��H; �H;��H;@�H;��H;�H;��H;/�H; mH;6H;r�G;�F;زC;]=;0;�l;Pg�:h	�90к$J������#���o��s/��Ȅ�y�ýӈ��nH�}��|㼾i���W��6E�`�h�W ��a���      � ����y�`�h���N��O/����B�߾B���*|��6�p}�䳽iSt�<�!�orμAF{��_��X��Γ��<:.��:�Z;�2;�O>;oD;)�F;{�G;=H;�pH;��H;I�H;ͷH;��H;��H;_�H;~�H;a�H;w�H;_�H;��H;��H;̷H;D�H;��H;�pH;=H;{�G;1�F;jD;�O>;�2;�Z;"��:T:ғ���X���_�AF{�orμ<�!�iSt�䳽p}��6��*|�B��B�߾����O/���N�`�h���y�      7�X�VvS�6E��O/��S�GW����������LS\��� ���9����Y�z��Ѓ����]�����$�b���Y�8�Y:��:f`;9�4;�?;9�D;��F;�G;FH;GuH;ēH;��H;��H;�H;��H; �H;�H;��H;�H; �H;��H;�H;��H;��H;ƓH;FuH;FH;�G;��F;8�D;�?;1�4;``;��:@�Y:��Y�%�b�������]�Ѓ��{���Y�9����彑� �LS\���������GW���S��O/�6E�VvS�      �O/�pM+�W�����GW��9ɾA���Mw�� :�i��w�ý�L��\n;�]���sv���E<��˻��-�0��dy�:�^;�%;~�7;v�@;5E;�"G;�G;8PH;�zH;��H;Z�H;|�H;��H;��H;�H;��H;��H;��H;�H;��H;��H;|�H;T�H;H;�zH;8PH;�G;�"G;5E;r�@;|�7;�%;�^;hy�:@����-��˻�E<�sv��]���[n;��L��w�ýi��� :��Mw�A��9ɾGW�����X��pM+�      /y��v�i���B�߾����A��?����nH���CὝu����d�/O�irμI"�����	�����`r89X;�:a�;�+;Q|:;y7B;��E;�aG;rH;�ZH;e�H;,�H;��H;�H;J�H;G�H;�H;��H;u�H;��H;�H;G�H;F�H;�H;��H;0�H;c�H;�ZH;qH;bG;��E;v7B;O|:;�+;Z�;\;�:Pr89���	�����I"��irμ0O���d��u��C����nH�?���A������B�߾i����v�      @�;9ɾ|㼾B�������Mw��nH�����Z�䳽˕��q\8�n#������^N�M���b� Ix�<5:ۮ�:1�;��0;]=;@�C;�[F;ӞG;�)H;�eH;s�H;&�H;=�H;��H;�H;��H;+�H;��H;n�H;��H;-�H;��H;�H;��H;;�H;+�H;s�H;�eH;�)H;؞G;�[F;:�C;]=;��0;)�;��:85:Ix�
�b�M��^N�����n#��q\8�ʕ��䳽�Z񽰯��nH��Mw�����B��|㼾9ɾ      ఖ�����}���*|�LS\�� :����Z�l$�������K�v���Oļ����������B&����A/�:�^;��#;�G6;5�?;��D;E�F;��G;@H;�pH;��H;u�H;�H;N�H;3�H;n�H;r�H;��H;z�H;��H;r�H;m�H;-�H;L�H;�H;z�H;ޏH;�pH;@H;��G;H�F;��D;8�?;�G6;��#;�^;C/�:0��C&������������Oļv���K�����k$���Z���� :�LS\��*|�}������      �+X��T��nH��6��� �i��C�䳽�����mR����ټ�����E<��?ݻ8d\������ :�d�:��;'�,;y�:;U7B;��E;mLG;,H;ZSH;�{H;}�H;�H;�H;@�H;V�H;�H;��H;��H;��H;��H;��H;�H;Q�H;:�H;�H;�H;�H;�{H;YSH;+H;oLG;��E;V7B;y�:;"�,;��;�d�:� :����7d\��?ݻ�E<�����ټ����mR�����䳽C�i���� ��6��nH��T�      �� ]�ӈ�p}���w�ý�u��ʕ���K�����o�jv���&R���V^����� �>����:[B;7";f�4;��>;;D;��F;�G;�)H;fdH;r�H;	�H;a�H;(�H;/�H;��H;��H;�H;�H;��H;�H;�H;��H;~�H;*�H;(�H;f�H;�H;q�H;ddH;�)H;�G;��F;=D;��>;b�4;>";]B;���: �>����V^�����&R�iv���o�����K�ʕ���u��w�ý��p}�ӈ� ]�       �ѽ\νy�ý䳽9����L����d�q\8�v��ټhv����Y��_����?���[���Y:U��:Im;�r-;
�:;l�A;(oE;�"G;J�G;WGH;�sH;�H;��H;�H;%�H;�H;��H;v�H;~�H;'�H;��H;'�H;~�H;{�H;��H;�H;&�H;�H;��H;�H;�sH;WGH;K�G;�"G;,oE;l�A;�:;�r-;Im;U��:��Y:�[�=������_���Y�hv��ټu��q\8���d��L��:���䳽y�ý\ν      ���������Ȅ�jSt��Y�\n;�/O�m#���Oļ�����&R��_������N3��Y��3:��:ӯ;�?&;�G6;}X?;�D;"xF;��G;*!H;�^H;��H;�H;ĭH;>�H;��H;��H;��H;	�H;��H;P�H;�H;P�H;��H;	�H;��H;��H;�H;E�H;ɭH;�H;��H;�^H;0!H;��G;$xF;�D;}X?;�G6;�?&;ϯ;�:�3:��Y��N3������_��&R������Oļm#��/O�[n;��Y�jSt��Ȅ�����      ]n;�x\8��s/�<�!�y��_���hrμ��������E<�������N3�XHx���9��:�^;Q ;)2;]�<;�B;��E;!5G; �G;'FH;vqH;��H;>�H;��H;F�H;��H;��H;��H;��H;�H;n�H;�H;n�H;�H;��H;��H;��H;��H;P�H;��H;A�H;��H;uqH;+FH; �G;'5G;��E;�B;e�<;*2;N ;�^;��:��9HHx��N3�������E<��������irμ]���z��=�!��s/�w\8�      Z������o�orμЃ��rv��I"��^N�����?ݻT^��D���Y���9��:Ѧ�:��;N�.;z|:;�>A;��D; �F;��G;�)H;aH;	�H;t�H;ڬH;-�H;�H;/�H;W�H;��H;�H;O�H;��H;��H;��H;N�H;�H;��H;S�H;2�H;�H;2�H;�H;t�H;�H;aH;�)H;��G;#�F;��D;�>A;||:;J�.;��;Ѧ�:��:��9�Y�?��S^���?ݻ���^N�I"��qv��҃��orμ�o����      �����x���#��?F{���]��E<����I�뻨���6d\�z���[��3:��:Ӧ�:v[;_�,;��8;!@;�0D;o[F;{G;�
H;;PH;vH;ڐH;6�H;��H;�H;]�H;q�H;��H;��H;t�H;o�H;��H;��H;��H;m�H;t�H;��H;��H;t�H;c�H;#�H;��H;6�H;֐H;vH;;PH;�
H;{G;p[F;�0D;!@;��8;d�,;v[;٦�:��:�3:�[�v��3d\�����H�뻢���E<���]�@F{��#���x��      �B(�%�����_������˻	���b�;&����� |>���Y:�:�^;��;e�,;`8;a�?;��C;iF;�FG;?�G;�?H;kH;�H;��H;�H;L�H;��H;b�H;k�H;�H;u�H;��H;��H;~�H;��H;z�H;��H;��H;r�H;�H;o�H;f�H;��H;M�H;�H;��H;��H;kH;�?H;B�G;�FG;qF;��C;X�?;`8;e�,;��;�^;�:��Y: t>�����:&��b�	���˻�����_���� %�      ̚��I���$J���X���b���-�����Hx����� :���:G��:̯;N ;J�.;��8;U�?;��C;��E;'#G;��G;�1H;�aH;@�H;j�H;m�H;��H;��H;S�H;�H;(�H;0�H;��H;�H;��H;5�H;��H;2�H;�H;�H;��H;,�H;,�H;�H;U�H;��H;��H;j�H;o�H;>�H;�aH;�1H;��G;.#G;��E;��C;X�?;��8;K�.;N ;ί;Q��:	��:!:����Hx������-��b��X�� J��I���      *�����.кȓ����Y�����r89P5:I/�:�d�:dB;Em;�?&;,2;~|:;!@;��C;��E;oG;��G;K(H;�ZH;`zH;/�H;ǤH;��H;Z�H;��H;��H;U�H;��H;��H;D�H;&�H;D�H;��H;v�H;��H;A�H;&�H;A�H;��H;��H;Z�H;��H;��H;Y�H;��H;ͤH;0�H;]zH;�ZH;O(H;��G;rG;��E;��C;!@;|:;,2;�?&;Im;fB;�d�:O/�:X5:�r89�����Y�ޓ��.к���      0�e9(�9�	�9�:$�Y:py�:t;�:ۮ�:�^;��;>";�r-;�G6;e�<;�>A;�0D;sF;5#G;��G;�$H;RWH;�vH;i�H;4�H;5�H;n�H;�H;��H;q�H;0�H;��H;x�H;��H;"�H;�H;��H;��H;��H;�H;!�H;��H;t�H;��H;.�H;n�H;��H;�H;l�H;;�H;5�H;f�H;�vH;WWH;�$H;��G;1#G;sF;�0D;�>A;b�<;�G6;�r-;D";��;�^;��:p;�:|y�:@�Y:<:P	�9��9      Z�:S-�: g�:��:��:�^;Z�;)�;��#;&�,;f�4;�:;~X?;�B;��D;s[F;�FG;��G;O(H;MWH;\uH;~�H;�H;�H;�H;��H;��H;��H;��H;��H;��H;��H;��H;��H;��H;S�H;M�H;L�H;��H;��H;��H;��H;��H;��H;��H;��H;��H;��H;�H;�H;�H;��H;buH;SWH;Q(H;��G;�FG;s[F;��D;�B;X?;�:;i�4;&�,;��#;'�;`�;�^;��:��:6g�:K-�:      �;t�;�l;�Z;``;�%;�+;��0;�G6;}�:;��>;l�A;�D;��E;'�F;{G;F�G;�1H;�ZH;�vH;��H;?�H;��H;øH;|�H;H�H;��H;��H;��H;��H;3�H;4�H;��H;��H;e�H;��H;��H;��H;b�H;��H;��H;.�H;4�H;��H;��H;��H;��H;J�H;�H;¸H;��H;A�H;��H;�vH;�ZH;�1H;G�G;{G;*�F;��E;�D;q�A;��>;z�:;�G6;��0;�+;�%;v`;�Z;�l;g�;      �Y.;��.;0;�2;,�4;��7;`|:;&]=;?�?;]7B;ED;/oE;'xF;25G;��G;�
H;�?H;�aH;azH;d�H;�H;��H;?�H;��H;[�H;��H;��H;��H;�H;��H;��H;X�H;R�H;A�H;��H;�H;@�H;�H;��H;B�H;N�H;R�H;��H;��H;�H;��H;��H;��H;_�H;��H;>�H;��H;�H;i�H;dzH;�aH;�?H;�
H;��G;05G;+xF;4oE;KD;\7B;B�?;&]=;_|:;��7;<�4;�2;0;��.;      P�<;$�<;]=;�O>;�?;{�@;y7B;=�C;�D;��E;��F;�"G;��G;�G;�)H;>PH;!kH;H�H;0�H;1�H;�H;��H;��H;.�H;)�H;,�H;>�H;��H;�H;5�H;��H;	�H;�H;��H;?�H;{�H;��H;t�H;=�H;��H;�H;�H;��H;3�H;�H;��H;:�H;.�H;,�H;.�H;��H;¸H;�H;2�H;0�H;A�H;!kH;BPH;�)H;�G;��G;�"G;��F;��E;��D;G�C;{7B;j�@;�?;�O>;]=;�<;      �WC;�nC;ӲC;iD;4�D;&5E;��E;�[F;K�F;rLG;��G;P�G;0!H;2FH;aH;vH;��H;y�H;ԤH;?�H;�H;�H;_�H;2�H;��H;��H;:�H;��H;��H;��H;��H;��H;��H;1�H;��H;��H;��H;��H;��H;4�H;��H;��H;��H;��H;��H;��H;6�H;��H;��H;2�H;a�H;��H;�H;>�H;פH;u�H;��H;vH;aH;2FH;4!H;W�G;��G;tLG;N�F;�[F;��E;5E;@�D;hD;ղC;�nC;      �ZF;�dF;݀F;'�F;��F;�"G;bG;��G;��G;2H;�)H;^GH;�^H;qH;�H;ݐH;��H;p�H;��H;k�H;��H;F�H;��H;.�H;��H;�H;��H;��H;h�H;��H;��H;��H;�H;t�H;��H;�H;�H;�H;��H;t�H; �H;��H;��H;��H;e�H;��H;��H;!�H; �H;.�H;��H;J�H;��H;l�H;��H;l�H;��H;ސH;�H;|qH;�^H;^GH;�)H;3H;��G;��G;bG;�"G;��F;-�F;�F;�dF;      �G;�G;p�G;}�G;�G;�G;{H;�)H; @H;\SH;fdH;�sH;��H;��H;r�H;8�H;�H;��H;]�H;�H;��H;��H;��H;A�H;7�H;��H;��H;8�H;{�H;��H;]�H;��H;o�H;��H;�H;5�H;O�H;/�H;��H;��H;q�H;��H;]�H;��H;z�H;8�H;�H;��H;9�H;?�H;��H;��H;��H;�H;]�H;��H;�H;<�H;u�H;��H;��H;�sH;hdH;YSH;�?H;�)H;xH;�G;�G;o�G;n�G;ܪG;      0H;�1H;6H;=H;�EH;:PH;�ZH;�eH;�pH;�{H;q�H;�H;�H;C�H;۬H;��H;M�H;��H;��H;��H;��H;��H;��H;��H;��H;��H;8�H;r�H;Z�H;F�H;��H;a�H;��H;�H;@�H;V�H;A�H;R�H;@�H;�H;��H;^�H;��H;F�H;Y�H;r�H;5�H;��H;��H;��H;��H;��H;��H;��H;��H;��H;O�H;��H;ݬH;C�H;�H;�H;u�H;�{H;�pH;�eH;�ZH;0PH;FH;=H;6H;�1H;      /jH;�jH;mH;�pH;5uH;�zH;i�H;p�H;׏H;|�H;�H;��H;ǭH;��H;0�H;#�H;��H;Z�H;��H;t�H;��H;��H;�H;�H;��H;a�H;r�H;\�H;O�H;��H;L�H;��H;��H;0�H;`�H;g�H;X�H;c�H;]�H;2�H;��H;��H;N�H;��H;O�H;Z�H;q�H;a�H;��H;�H;�H;��H;��H;o�H;��H;W�H;��H;&�H;0�H;��H;ǭH;��H;�H;�H;׏H;p�H;i�H;�zH;DuH;�pH;mH;�jH;      ;�H;��H;2�H;��H;ēH;��H;,�H;$�H;w�H;�H;c�H;�H;A�H;N�H;�H;`�H;i�H;�H;T�H;0�H;��H;��H;��H;0�H;��H;��H;��H;F�H;��H;B�H;��H;��H;,�H;Y�H;d�H;z�H;��H;x�H;b�H;X�H;/�H;��H;��H;@�H;��H;I�H;}�H;��H;��H;.�H;��H;��H;��H;-�H;T�H;�H;i�H;c�H;�H;L�H;A�H;�H;e�H;�H;w�H;$�H;.�H;��H;œH;��H;5�H;��H;      O�H;��H;��H;K�H;��H;V�H;��H;=�H;�H;�H;-�H;,�H;�H;��H;6�H;x�H;v�H;2�H;��H;��H;��H;6�H;��H;��H;��H;��H;X�H;��H;N�H;��H;��H;"�H;V�H;i�H;��H;��H;{�H;~�H;�H;j�H;\�H;"�H;��H;��H;M�H;��H;X�H;��H;��H;��H;��H;7�H;��H;��H;��H;0�H;y�H;z�H;5�H;��H;�H;/�H;/�H;�H;�H;>�H;��H;L�H;��H;H�H;��H;��H;      ��H;ԵH;~�H;��H;{�H;n�H;�H;��H;O�H;=�H;-�H;�H;��H;��H;Z�H;��H;�H;6�H;��H;~�H;��H;4�H;T�H;�H;��H;��H;��H;b�H;��H;��H;�H;:�H;`�H;��H;��H;��H;��H;��H;��H;��H;g�H;:�H;�H;��H;��H;a�H;��H;��H;��H;�H;Y�H;6�H;��H;{�H;��H;7�H;�H;��H;Z�H;��H;��H;�H;2�H;@�H;O�H;��H;��H;r�H;��H;·H;��H;ҵH;      .�H;r�H;�H;��H;�H;��H;F�H;�H;'�H;R�H;��H;��H;��H;��H;��H;��H;z�H;��H;K�H;��H;��H;��H;N�H; �H;��H;�H;l�H;��H;��H;2�H;U�H;d�H;w�H;��H;��H;��H;��H;��H;��H;��H;z�H;d�H;T�H;+�H;��H;��H;p�H;�H;��H;�H;S�H;��H;��H;��H;K�H;��H;��H;��H;��H;��H;��H;��H;��H;U�H;,�H;�H;I�H;z�H;�H;��H;�H;q�H;      ��H;��H;A�H;��H;��H;��H;H�H;��H;m�H;�H;��H;��H;�H;��H;�H;{�H;��H;�H;*�H;)�H;��H;��H;;�H;��H;+�H;m�H;��H;�H;,�H;Y�H;b�H;��H;��H;��H;��H;��H;��H;��H;��H;��H;��H;��H;b�H;V�H;+�H;�H;��H;o�H;.�H;��H;C�H;��H;��H;"�H;'�H;�H;��H;{�H;�H;��H;�H;�H;��H;�H;q�H;��H;L�H;��H;��H;��H;G�H;��H;      S�H;u�H;��H;_�H;+�H;��H;�H;+�H;t�H;��H;$�H;��H;��H;�H;Y�H;u�H;��H;��H;G�H;	�H;��H;b�H;��H;4�H;��H;��H;��H;?�H;`�H;f�H;z�H;��H;��H;��H;��H;��H;��H;��H;��H;��H;��H;��H;x�H;`�H;Y�H;:�H;��H;��H;��H;4�H;��H;a�H;��H;�H;C�H;��H;��H;u�H;V�H;�H;��H;��H;'�H;��H;z�H;.�H;�H;�H;+�H;a�H;��H;v�H;      ��H;��H;�H;w�H;�H;��H;��H;��H;��H;��H;�H;.�H;T�H;t�H;��H;��H;��H;5�H;��H;��H;T�H;��H;�H;l�H;��H;�H;.�H;T�H;g�H;~�H;|�H;��H;��H;��H;��H;��H;��H;��H;��H;��H;��H;��H;{�H;x�H;d�H;R�H;2�H;�H;��H;m�H;�H;��H;Q�H;��H;��H;6�H;��H;��H;��H;r�H;U�H;.�H;�H;��H;��H;��H;��H;��H;�H;s�H; �H;��H;      ��H;��H;��H;^�H;��H;��H;y�H;l�H;{�H;��H;��H;��H;�H;�H;��H;��H;��H;��H;{�H;��H;V�H;��H;?�H;��H;��H;�H;K�H;G�H;[�H;��H;u�H;��H;��H;��H;��H;��H;��H;��H;��H;��H;��H;��H;u�H;��H;V�H;D�H;O�H;�H;��H;��H;F�H;��H;Q�H;��H;y�H;��H;��H;��H;��H;�H;�H;��H;��H;��H;~�H;p�H;�H;��H;��H;_�H;��H;��H;      ��H;��H;��H;v�H;�H;��H;��H;��H;��H;��H;�H;.�H;T�H;t�H;��H;��H;�H;3�H;��H;��H;W�H;��H;�H;l�H;��H;�H;.�H;U�H;i�H;|�H;|�H;��H;��H;��H;��H;��H;��H;��H;��H;��H;��H;��H;{�H;w�H;d�H;Q�H;/�H;�H;��H;l�H;�H;��H;Q�H;��H;��H;6�H;��H;��H;��H;q�H;S�H;,�H;�H;��H;��H;��H;��H;��H;�H;w�H;�H;��H;      F�H;w�H;��H;X�H;,�H;��H;�H;.�H;t�H;��H;#�H;��H;��H;�H;[�H;u�H;��H;��H;G�H;
�H;��H;d�H;��H;4�H;��H;��H;��H;@�H;_�H;d�H;x�H;��H;��H;��H;��H;��H;��H;��H;��H;��H;��H;��H;x�H;_�H;\�H;:�H;��H;��H;��H;2�H;��H;b�H;��H;�H;C�H;��H;��H;u�H;U�H;�H;��H;��H;$�H;��H;u�H;5�H;�H;��H;2�H;\�H;��H;y�H;      ��H;��H;>�H;��H;��H;��H;E�H;��H;n�H;�H;��H;}�H;�H;��H;�H;{�H;��H;�H;*�H;(�H;��H;��H;>�H;��H;.�H;o�H;��H;�H;0�H;Y�H;c�H;��H;��H;��H;��H;��H;��H;��H;��H;��H;��H;��H;`�H;V�H;(�H;�H;��H;q�H;-�H;��H;C�H;��H;��H;"�H;(�H;�H;��H;{�H;�H;��H;�H;}�H;��H;�H;n�H;��H;N�H;��H;��H;��H;G�H;��H;      ,�H;u�H;�H;��H;�H;��H;C�H;�H;)�H;U�H;��H;��H;��H;��H;��H;��H;}�H;��H;I�H;��H;��H;��H;O�H;�H;��H;�H;m�H;��H;��H;2�H;T�H;b�H;u�H;��H;��H;��H;��H;��H;��H;��H;u�H;d�H;T�H;,�H;��H;��H;m�H;�H;��H;��H;U�H;��H;��H;��H;G�H;��H;z�H;��H;��H;��H;��H;��H;��H;T�H;*�H;�H;L�H;��H;�H;��H;�H;p�H;      q�H;еH;r�H;��H;z�H;}�H;��H;��H;N�H;=�H;.�H;�H;��H;��H;]�H;��H;�H;7�H;��H;~�H;��H;8�H;V�H;�H;��H;��H;��H;b�H;��H;��H;�H;:�H;c�H;�H;��H;��H;��H;��H;��H;�H;c�H;9�H;�H;��H;��H;^�H;��H;��H;��H;��H;[�H;5�H;��H;x�H;��H;4�H;�H;��H;X�H;��H;��H;�H;.�H;=�H;P�H;��H;��H;q�H;{�H;ķH;x�H;ʵH;      A�H;��H;��H;E�H;��H;V�H;��H;>�H;�H;�H;,�H;/�H;�H;��H;7�H;z�H;w�H;0�H;��H;��H;��H;9�H;��H;��H;��H;��H;X�H;��H;S�H;��H;��H;"�H;X�H;i�H;��H;�H;{�H;�H;~�H;i�H;[�H;"�H;��H;��H;J�H;��H;Z�H;��H;��H;��H;��H;7�H;��H;��H;��H;0�H;z�H;z�H;6�H;��H;�H;-�H;,�H;�H;�H;B�H;��H;S�H;��H;O�H;��H;��H;      C�H;��H;+�H;��H;��H;H;-�H;*�H;z�H;�H;c�H;�H;B�H;M�H;�H;b�H;g�H;�H;T�H;0�H;��H;��H;��H;1�H;��H;��H;��H;I�H;��H;C�H;��H;��H;)�H;X�H;c�H;w�H;��H;x�H;`�H;X�H;.�H;��H;��H;?�H;��H;C�H;��H;��H;��H;*�H;��H;��H;��H;-�H;U�H;�H;i�H;`�H;�H;M�H;A�H;�H;e�H;�H;w�H;(�H;.�H;��H;œH;��H;3�H;��H;      ;jH;�jH;,mH;�pH;/uH;{H;h�H;p�H;ݏH;{�H;�H;��H;ɭH;��H;2�H;&�H;��H;\�H;��H;q�H;��H;��H;�H;�H;��H;^�H;r�H;Z�H;S�H;��H;M�H;��H;��H;/�H;]�H;d�H;V�H;d�H;\�H;/�H;��H;��H;M�H;��H;L�H;Y�H;r�H;c�H;��H;�H;�H;��H;��H;q�H;��H;W�H;��H;'�H;2�H;��H;ǭH;��H;�H;{�H;ۏH;v�H;l�H;�zH;=uH;�pH;*mH;�jH;      0H;�1H;6H;=H;�EH;DPH;�ZH;�eH;�pH;�{H;t�H;�H;�H;C�H;ެH;��H;M�H;��H;��H;��H;��H;��H;��H;��H;��H;��H;5�H;r�H;]�H;F�H;��H;b�H;��H;�H;?�H;R�H;A�H;T�H;=�H;	�H;��H;_�H;��H;F�H;Z�H;r�H;6�H;��H;��H;��H;��H;��H;��H;��H;��H;��H;O�H;��H;ެH;A�H;�H;�H;u�H;�{H;�pH;�eH;�ZH;3PH;FH;=H;6H;�1H;      �G;��G;j�G;��G;�G;�G;{H;�)H;@H;ZSH;gdH;�sH;��H;��H;t�H;;�H;�H;��H;\�H;�H;��H;��H;��H;E�H;:�H;��H;�H;9�H;|�H;��H;[�H;��H;m�H;��H;�H;0�H;O�H;0�H;��H;��H;p�H;��H;]�H;��H;z�H;8�H;��H;��H;6�H;<�H;��H;��H;��H;�H;^�H;��H;�H;<�H;u�H;��H;��H;�sH;fdH;YSH;�?H;�)H;|H;	�G;�G;��G;n�G;�G;      �ZF;�dF;�F;%�F;��F;�"G;�aG;�G;��G;0H;�)H;_GH;�^H;}qH;�H;ߐH;��H;q�H;��H;i�H;��H;H�H;��H;1�H;��H;�H;��H;��H;h�H;��H;��H;��H;�H;s�H;��H;�H;�H;�H;��H;s�H;�H;��H;��H;��H;c�H;��H;��H;�H;��H;,�H;��H;H�H;��H;l�H;��H;l�H;��H;ߐH;�H;{qH;�^H;\GH;�)H;2H;��G;ܞG;�aG;�"G;��F;%�F;̀F;�dF;      �WC;�nC;βC;fD;7�D;(5E;��E;�[F;N�F;rLG;��G;R�G;0!H;1FH;aH;vH;��H;x�H;֤H;>�H;�H;��H;_�H;4�H;��H;��H;6�H;��H;��H;��H;��H;��H;��H;/�H;��H;��H;��H;��H;��H;1�H;��H;��H;��H;��H;��H;��H;:�H;��H;��H;/�H;a�H;��H;�H;A�H;ؤH;u�H;��H;vH;aH;0FH;1!H;R�G;��G;tLG;I�F;�[F;��E;5E;<�D;hD;ϲC;�nC;      -�<;�<;]=;�O>;؁?;�@;|7B;A�C;��D;��E;��F;�"G;��G;�G;�)H;APH; kH;G�H;/�H;1�H;�H;��H;��H;1�H;-�H;)�H;>�H;��H;�H;1�H;��H;
�H;�H;��H;=�H;x�H;��H;z�H;<�H;��H;�H;�H;��H;5�H;�H;��H;?�H;-�H;*�H;.�H;��H;��H;�H;5�H;3�H;C�H;"kH;APH;�)H;�G;��G;�"G;��F;��E;��D;=�C;y7B;t�@;�?;�O>;]=;��<;      �Y.;��.;0;�2;*�4;��7;X|:;&]=;C�?;\7B;BD;2oE;'xF;/5G;��G;�
H;�?H;�aH;azH;f�H;
�H;��H;>�H;��H;a�H;��H;��H;��H;�H;��H;��H;X�H;O�H;A�H;��H;�H;C�H;�H;��H;?�H;R�H;Y�H;��H;��H;�H;��H;��H;��H;\�H;��H;>�H;��H;�H;j�H;dzH;�aH;�?H;�
H;��G;.5G;)xF;/oE;DD;\7B;C�?;)]=;Y|:;��7;*�4;�2;0;��.;      �;t�;�l;�Z;b`;�%;�+;��0;�G6;y�:;��>;q�A;�D;��E;)�F;{G;D�G;�1H;�ZH;�vH;��H;@�H;��H;øH;��H;G�H;��H;��H;��H;��H;3�H;2�H;��H;��H;b�H;��H;��H;��H;b�H;��H;��H;4�H;9�H;��H;��H;��H;��H;J�H;~�H;ŸH;��H;A�H;��H;�vH;�ZH;�1H;F�G;{G;)�F;��E;�D;p�A;��>;z�:;�G6;��0;�+;�%;x`;�Z;�l;j�;      B�:�-�:Bg�:&��:��:�^;^�;,�;��#;#�,;g�4;�:;~X?;�B;��D;u[F;�FG;��G;N(H;PWH;]uH;��H;
�H;�H;�H;��H;��H;��H;��H;��H;��H;��H;��H;��H;��H;O�H;O�H;P�H;��H;��H;��H;��H;��H;��H;��H;��H;��H;��H;�H;�H;�H;��H;`uH;UWH;Q(H;��G;�FG;s[F;��D;�B;~X?;�:;j�4;$�,;��#;.�;`�;�^;��: ��:\g�:[-�:      `�e9P�9X	�9�:0�Y:|y�:|;�:��:�^;��;C";�r-;�G6;b�<;�>A;�0D;qF;3#G;��G;�$H;VWH;�vH;i�H;5�H;<�H;l�H;�H;��H;r�H;*�H;��H;x�H;��H;$�H;�H;��H;��H;��H;�H; �H;��H;x�H;��H;0�H;q�H;��H;�H;n�H;7�H;8�H;i�H;�vH;VWH;�$H;��G;1#G;tF;�0D;�>A;d�<;�G6;�r-;D";��;�^;��:p;�:jy�:H�Y:\:h	�9(�9      *�����0к����Y�����r89X5:O/�:�d�:dB;Im;�?&;)2;�|:;!@;��C;��E;oG;��G;Q(H;�ZH;czH;0�H;ΤH;��H;Z�H;��H;��H;T�H;��H;��H;B�H;&�H;F�H;��H;v�H;��H;D�H;$�H;B�H;��H;��H;X�H;��H;��H;\�H;��H;ɤH;3�H;czH;�ZH;O(H;��G;pG;��E;��C;!@;�|:;)2;�?&;Hm;dB;�d�:O/�:d5:�r89�����Y�ȓ��:к���      Ԛ��D���'J���X���b���-�����Hx����!:��:U��:ѯ;M ;N�.;��8;W�?;��C;��E;-#G;��G;�1H;�aH;A�H;q�H;l�H;��H;��H;V�H;�H;*�H;/�H;��H;�H;��H;3�H;��H;5�H;~�H;�H;��H;0�H;-�H;�H;V�H;��H;��H;j�H;k�H;A�H;�aH;�1H;��G;0#G;��E;��C;W�?;��8;N�.;K ;˯;O��:��:� :����Hx������-��b��X��+J��D���      �B(�%�����_������˻	����b�<&����� |>���Y:
�:�^;��;h�,;
`8;\�?;��C;pF;�FG;C�G;�?H; kH;��H;��H;�H;J�H;��H;`�H;n�H;�H;u�H;��H;��H;}�H;��H;}�H;��H;��H;s�H;�H;p�H;d�H;��H;L�H;�H;��H;�H;kH;�?H;?�G;�FG;qF;��C;[�?;`8;e�,;��;�^;�:��Y: |>�����8&��b�	���˻�����_���� %�      �����x���#��>F{���]��E<����H�뻨���5d\�v�뺨[��3:��:ݦ�:z[;a�,;��8;!@;�0D;v[F;{G;�
H;=PH;vH;ېH;5�H;��H;#�H;_�H;t�H;��H;��H;v�H;q�H;��H;��H;��H;m�H;s�H;��H;��H;t�H;b�H;#�H;��H;4�H;֐H;vH;:PH;�
H;{G;l[F;�0D;!@;��8;b�,;t[;צ�:��:�3:�[�x��5d\�����I�뻣���E<���]�?F{��#���x��      Z������o�nrμЃ��rv��I"��^N�����?ݻT^��?����Y���9��:צ�:��;K�.;||:;�>A;��D;&�F;��G;�)H;aH;�H;t�H;ݬH;2�H;�H;3�H;W�H;��H;�H;O�H;��H;��H;��H;O�H;�H;��H;V�H;2�H;�H;3�H;ݬH;q�H;�H;aH;�)H;��G;%�F;��D;�>A;{|:;G�.;��;Ϧ�:��:��9�Y�@��T^���?ݻ���^N�I"��rv��҃��prμ�o����      ^n;�w\8��s/�<�!�y��]���hrμ��������E<�������N3�DHx���9��:�^;M ;)2;b�<;��B;��E;)5G;�G;.FH;|qH;��H;?�H;��H;J�H;��H;��H;��H;��H;�H;m�H;�H;p�H;�H;��H;��H;��H;��H;N�H;��H;A�H;��H;uqH;)FH;�G;.5G;��E;�B;e�<;&2;M ;�^;��:��9HHx��N3�������E<��������irμ^���z��<�!��s/�w\8�      ���������Ȅ�jSt��Y�\n;�/O�m#���Oļ�����&R��_������N3�ЅY��3: �:ѯ;�?&;�G6;�X?;�D;*xF;��G;1!H;�^H;��H;�H;˭H;A�H;�H;��H;��H;�H;��H;Q�H;�H;Q�H;��H;�H;��H;��H;�H;C�H;ʭH;�H;��H;�^H;,!H;��G;*xF;�D;xX?;�G6;�?&;̯; �:�3:܅Y��N3������_��&R������Oļm#��/O�[n;��Y�jSt��Ȅ�����       �ѽ\νy�ý䳽9����L����d�q\8�v��ټhv����Y��_����;���[���Y:K��:Im;�r-;�:;n�A;2oE;�"G;N�G;YGH;�sH;�H;��H;�H;)�H;�H;��H;{�H;�H;'�H;��H;)�H;~�H;y�H;��H;�H;&�H;�H;��H;�H;�sH;UGH;I�G;�"G;2oE;l�A;�:;�r-;Fm;K��:��Y:�[�=������_���Y�hv��ټv��q\8���d��L��:���䳽y�ý\ν      �� ]�ӈ�p}���w�ý�u��ʕ���K�����o�iv���&R���T^��~�� �>����:[B;:";j�4;��>;DD;��F;�G;�)H;fdH;q�H;�H;b�H;*�H;.�H;��H;��H;�H;�H;��H;�H;�H;��H;��H;+�H;(�H;f�H;�H;q�H;ddH;�)H;�G;��F;BD;��>;_�4;:";ZB;���: �>����V^�����&R�iv���o�����K�ʕ���u��w�ý��p}�ӈ� ]�      �+X��T��nH��6��� �i��C�䳽�����mR����ټ�����E<��?ݻ6d\������ :�d�:��;*�,;y�:;\7B;��E;qLG;/H;ZSH;�{H;��H;�H;�H;?�H;V�H;�H;��H;��H;��H;��H;��H;�H;R�H;<�H;�H;�H;��H;�{H;YSH;,H;mLG;��E;Z7B;v�:;�,;��;�d�:� :����8d\��?ݻ�E<�����ټ����mR�����䳽C�i���� ��6��nH��T�      ఖ�����}���*|�LS\�� :����Z�l$�������K�v���Oļ����������A&� ��C/�:�^;��#;�G6;9�?;��D;K�F;��G;@H;�pH;��H;w�H;�H;N�H;1�H;n�H;q�H;��H;{�H;��H;q�H;m�H;-�H;N�H;�H;z�H;��H;�pH;@H;��G;H�F;��D;;�?;�G6;��#;�^;?/�: ��A&������������Oļv���K�����k$���Z���� :�LS\��*|�}������      @�;9ɾ|㼾B�������Mw��nH�����Z�䳽ʕ��q\8�n#������^N�L���b�Ix�D5:߮�:1�;��0;]=;?�C;�[F;՞G;�)H;�eH;s�H;$�H;>�H;��H;�H;��H;*�H;��H;n�H;��H;+�H;��H;�H;��H;=�H;+�H;v�H;�eH;�)H;֞G;�[F;=�C;]=;��0;)�;��:85:Ix��b�M��^N�����n#��q\8�ʕ��䳽�Z񽰯��nH��Mw�����B��|㼾9ɾ      /y��v�i���B�߾����A��?����nH���CὝu����d�/O�irμI"�����	�����Pr89\;�:a�;�+;Q|:;x7B;��E;�aG;pH;�ZH;f�H;-�H;��H;�H;I�H;G�H;�H;��H;u�H;��H;�H;E�H;F�H;�H;��H;3�H;h�H;�ZH;tH;bG;��E;y7B;T|:;�+;Z�;b;�:0r89���	�����I"��irμ0O���d��u��C����nH�?���A������B�߾j����v�      �O/�pM+�X�����GW��9ɾA���Mw�� :�i��w�ý�L��[n;�]���sv���E<��˻��-�(��hy�:�^;�%;~�7;v�@;5E;�"G;	�G;7PH;�zH;��H;[�H;}�H;��H;��H;�H;��H;��H;��H;�H;��H;��H;}�H;W�H;ėH; {H;:PH;�G;�"G;5E;u�@;��7;�%;�^;ny�:@����-��˻�E<�sv��]���\n;��L��w�ýi��� :��Mw�A��9ɾGW�����X��pM+�      7�X�VvS�6E��O/��S�GW����������LS\��� ���9����Y�z��Ѓ����]�����&�b���Y�@�Y:��:f`;6�4;�?;<�D;��F;�G;FH;GuH;H;��H;��H;�H;��H;�H;�H;��H;�H;�H;��H;�H;��H;��H;˓H;HuH;FH;�G;��F;9�D;�?;3�4;b`;��:H�Y:��Y�#�b�������]�Ѓ��z���Y�9����彑� �LS\���������GW���S��O/�6E�VvS�      � ����y�`�h���N��O/����B�߾B���*|��6�p}�䳽iSt�<�!�orμAF{��_��X��̓��H:.��:�Z;�2;�O>;oD;&�F;y�G;=H;�pH;��H;K�H;ͷH;��H;��H;_�H;|�H;b�H;y�H;\�H;��H;��H;ϷH;H�H;��H;�pH;=H;}�G;1�F;jD;�O>;�2;�Z;&��:\:ғ���X���_�AF{�orμ<�!�iSt�䳽p}��6��*|�B��B�߾����O/���N�`�h���y�      =v��b���W ��`�h�6E�W��j���|㼾}���nH�ӈ�y�ý�Ȅ��s/��o��#�����$J��*кP	�9\g�:�l;"0;!]=;ݲC;ـF;q�G;6H; mH;(�H;��H;��H;��H;@�H;��H;�H;��H;�H;��H;>�H;��H;�H;��H;/�H; mH;6H;t�G;�F;زC;]=;0;�l;Pg�:p	�90к$J������#���o��s/��Ȅ�y�ýӈ��nH�}��|㼾j���W��6E�`�h�W ��b���      |h��/���b�����y�VvS�pM+��v�9ɾ�����T� ]�\ν����x\8�����x��%�N���r��`�9w-�:j�;��.; �<;�nC;�dF;�G;�1H;�jH;��H;��H;εH;k�H;��H;h�H;��H;��H;��H;e�H;��H;i�H;͵H;��H;��H;�jH;�1H;�G;�dF;�nC;�<;��.;d�;g-�:p�9z��M���%��x�����x\8�����\ν ]��T�����9ɾ�v�pM+�VvS���y�b���/���      EEb�`]��N��7����s� ���˾��(�j��!,�o���L��Cm�+��8,˼��x�\���1�����T�:t�:�;�1;9,>;g�C;VwF;�G;q H;�>H;�hH;-�H;D�H;�H;��H;��H;�H;o�H;�H;��H;��H;�H;A�H;)�H;�hH;�>H;n H;�G;awF;c�C;4,>;
�1;�;l�:\�:����1��\����x�7,˼+��Cm�L��o����!,�(�j�����˾s� �����7��N�`]�      `]�d�W��TI�v3��D�������Ǿv����f�7)�$��r;���Fi��k���Ǽ�[t�N�	�+Ȅ�X��̠:��:��;,J2;TZ>;*	D;>F;=�G;�H;�?H;xiH;ňH;��H;T�H;�H;��H;8�H;��H;1�H;��H;�H;Q�H;��H;��H;~iH;�?H;�H;=�G;HF;%	D;QZ>;$J2;��;��:Ԡ:X��*Ȅ�N�	��[t���Ǽ�k��Fi�r;��$��7)��f�v�����Ǿ�����D�v3��TI�d�W�      �N��TI���;�/�'�l��쾀���x󐾳Z��K ��s�@����&^���"����g����Шu�� ���2<:��:�
;9g3;��>;XBD;x�F;�G;lH;BH;^kH;/�H;��H;�H;��H;E�H;��H;%�H;��H;C�H;��H;�H;��H;(�H;ekH;BH;kH;�G;��F;UBD;��>;2g3;�
;��:�2<:� ��Ѩu������g��"����&^�A����s潥K ��Z�x󐾀�����l�/�'���;��TI�      �7�v3�/�'����s� ��{Ծ ���H���y�F�����ӽ���^�L�Jv��뮼QT����PV���=�X)i:v��:�z ;�$5;��?;�D;��F;�G;uH;fFH;unH;d�H;N�H;N�H;��H;�H;4�H;��H;.�H;�H;��H;K�H;K�H;]�H;znH;eFH;pH;�G;��F;�D;��?;w$5;�z ;r��:`)i:��=��PV���QT��뮼Jv�^�L�����ӽ���y�F�H��� ����{Ծs� ����/�'�v3�      ����D�l�s� �V�ݾj���V͓��f��>/�����'���섽O�6�~t�w��^�:�(Tʻ}.�8۷�<t�:�;��$;�Y7;S�@;�	E;��F;+�G;�H;
LH;�rH;��H;��H; �H;��H;�H;'�H;��H;"�H;�H;��H;��H;��H;��H;�rH;LH;�H;-�G;��F;�	E;O�@;Y7;��$;�;Dt�:H۷�~.�(Tʻ^�:�w��t�O�6��섽�'������>/��f�V͓�j���V�ݾs� �l��D�      s� ��������{Ծj���v���Z�x��SC��^��޽?���x�e�'��C�Ѽ$G������R������ݤ8Ç�:�Y;G�);��9;��A;��E;G;�G;A!H;SH;�wH;L�H;\�H;�H;��H;N�H;Y�H;��H;S�H;L�H;��H;�H;\�H;G�H;�wH;
SH;@!H;�G;�G;��E;��A;��9;C�);�Y;Ň�:�ݤ8����R�����$G��C�Ѽ(��x�e�?����޽�^��SC�Z�x�v���j����{Ծ�쾠���      ��˾��Ǿ���� ���V͓�Z�x���J��K �m���������?����뮼+�[����3|��W����:;�:�';a/;=g<;�C;DF;�NG;��G;
-H;=[H;�}H;��H;��H;��H;��H;��H;��H;��H;��H;��H;��H;��H;��H;��H;�}H;=[H;-H;��G;�NG;FF;�C;;g<;^/;�';=�:|�:�W��3|����*�[��뮼���?������m����K ���J�Y�x�V͓� ���������Ǿ      ��v���x�H����f��SC��K �nn����Ž����Z��k�}ռ-X��ay-�,���r.����P�:�+�:~�;4;�>;�D;�wF;��G;��G;�9H;)dH;V�H;��H;5�H;K�H;��H;��H;.�H;H�H;+�H;��H;��H;G�H;0�H;}�H;[�H;)dH;�9H;��G;�G;�wF;�D;�>;4;w�;�+�:�P�:���s.�,���`y-�-X��}ռ�k��Z������Žnn���K ��SC��f�H���x�v���      (�j��f��Z�y�F��>/��^�m�����ŽF ���Fi��Q+�{t�nT��n�W�����1��,ȺX�9uP�:�Y;��(;��8;�A;�E;��F;8�G;sH;�FH;�mH;m�H;��H;�H;K�H;��H;b�H;��H;��H;��H;b�H;��H;D�H;�H;��H;q�H;�mH;�FH;rH;6�G;��F;�E;�A;��8;}�(;�Y;qP�: X�9,Ⱥ�1�����m�W�nT��{t�Q+��Fi�F ����Žm����^��>/�y�F��Z��f�      �!,�7)��K ��������޽������Fi��0����鷼��x�����.��S�(� ���*i:t��:$�;��0;6�<;nC;��E;�<G;��G;�$H;;TH;�wH;ʒH;�H;$�H;[�H;�H;g�H;t�H;Q�H;q�H;f�H;�H;U�H;�H;�H;̒H;�wH;;TH;�$H;��G;�<G;��E;oC;8�<;��0;)�;t��:�*i:���S�(��.�������x�鷼����0��Fi�������޽�������K �7)�      o���$��s��ӽ�'��?������
�Z��Q+�����"��G����0���׻˕b�>W���X�9ҡ�:`;|*';�Y7;�#@;�D;��F;�G;��G;8H;�aH;΁H;6�H;|�H;K�H;n�H;y�H;X�H;%�H;�H;&�H;Z�H;y�H;i�H;F�H;z�H;<�H;сH;�aH;8H;��G;�G;ݖF;�D;�#@;�Y7;�*';`;ʡ�:�X�9>W��ʕb���׻��0�G���"������Q+�
�Z����?����'���ӽ�s�$��      K��s;��@�������섽x�e��?��k�{t�鷼G���e7���� Ȅ�t0�@�t�u�:�+�:l;j1;A�<;H�B;��E;�G;��G;0H;RJH;4oH;ӋH;��H;�H;n�H;��H;��H;j�H;��H;��H;��H;j�H;��H;��H;j�H;�H;��H;ًH;4oH;PJH;/H;��G;�G;�E;K�B;A�<;v1;l;�+�:u�:@�t�r0��Ǆ���껃e7�G��鷼{t��k��?�w�e��섽���A���r;��      Cm��Fi��&^�_�L�O�6�(����}ռnT����x���0����������ط��n`:|�:�;�*;�8;��@;�D;A�F;�}G;x�G;i1H;�[H;E|H;��H;��H;Y�H;��H;��H;^�H;h�H;��H;E�H;��H;g�H;^�H;��H;��H;]�H;��H;��H;E|H;�[H;h1H;}�G;�}G;D�F;�D;��@;#�8;�*;�;��:�n`:�ط��������껾�0���x�mT��}ռ��'��P�6�_�L��&^��Fi�      *���k��Jv�|t�D�Ѽ�뮼,X��m�W������׻Ȅ���(���4<:Q��:�Y;�t%;�$5;�Z>;�`C;��E;
*G;@�G;�H;�GH;FlH;ǈH;ӞH;��H;��H;p�H;��H;��H;J�H;F�H;�H;E�H;H�H;��H;��H;k�H;��H;��H;ܞH;ʈH;ElH;�GH;�H;@�G;*G;��E;�`C;�Z>;�$5;�t%;�Y;M��:�4<:�����Ǆ���׻���l�W�,X���뮼C�Ѽ~t�Jv���k�      6,˼��Ǽ�"���뮼w��$G��*�[�_y-�����.��Ǖb�~0��ط��4<:�L�:�\;n�!;�J2;�g<;,0B;CE;	�F;#�G;��G;^4H;u\H;�{H;~�H;v�H;/�H;��H;�H;i�H;$�H;%�H;��H;��H;��H;%�H;&�H;h�H;�H;��H;6�H;|�H;��H;�{H;r\H;b4H;��G;$�G;�F;CE;40B;�g<;�J2;t�!;�\;�L�: 5<:�ط�t0�ĕb��.�����_y-�*�[�#G��w���뮼�"����Ǽ      ��x��[t���g�OT�_�:�������)����1��R�(�8W�� �t��n`:S��:�\; { ;��0;O;;�<A;��D;�wF;�cG;*�G;�!H;�MH;VoH;J�H;Z�H;��H;e�H;9�H;��H;/�H;D�H;��H;m�H;��H;k�H;��H;D�H;,�H;��H;<�H;k�H;��H;]�H;H�H;RoH;�MH;�!H;+�G;�cG;�wF;��D;�<A;K;;��0; { ;�\;S��:�n`:@�t�4W��P�(��1��(���������a�:�PT���g��[t�      Y��L�	������%Tʻ�R��3|�m.�"Ⱥ���Y�9u�:��:�Y;r�!;��0;ԕ:;��@;�BD;c2F;V8G;��G;�H;?@H;�cH;��H;K�H;�H;�H;!�H;d�H;��H;��H;B�H;��H;��H;Z�H;��H;��H;C�H;��H;��H;i�H;%�H;�H;�H;H�H;��H;�cH;@@H;�H;��G;X8G;i2F;�BD;��@;ו:;��0;v�!;�Y;��:u�:(Y�9���Ⱥl.�3|��R��(Tʻ�����J�	�      �1��'Ȅ�Ѩu��PV�q.�����W��X��X�9+i:ԡ�:�+�:�;�t%;�J2;H;;��@;\D;�F; G;T�G;dH;U5H;UZH;xH;�H;��H;�H;�H;-�H;?�H;��H;�H;��H;�H;3�H;��H;0�H;�H;��H;��H;��H;C�H;4�H;�H;�H;��H;�H;xH;TZH;S5H;gH;W�G;G;�F;YD;��@;F;;�J2;�t%;�;�+�:ࡼ:+i:HX�9H��W�����m.��PV�ʨu�&Ȅ�      䥥�8X��� ����=�H۷� ߤ8��:�P�:yP�:z��:$`;h;�*;�$5;�g<;�<A;�BD;�F;�G;S�G;=�G;v-H;�RH;+qH;��H;��H;S�H;�H;�H;��H;��H;��H;'�H;��H;t�H;k�H;��H;h�H;q�H;��H;$�H;��H;��H;��H;
�H;�H;N�H;��H;��H;.qH;�RH;y-H;A�G;X�G;�G;�F;�BD;�<A;�g<;�$5;�*;l;)`;z��:P�:�P�:��:�ޤ88۷���=�� ��8X��      @�:��:�2<:�)i:4t�:ɇ�:W�:�+�:�Y;)�;�*';s1;#�8;�Z>;70B;��D;i2F;G;Y�G;��G;U)H;ZNH;IlH;�H;6�H;U�H;p�H;�H;Z�H;��H;�H; �H;�H;0�H;��H;��H;��H;��H;��H;0�H;�H;��H;�H;��H;X�H;�H;n�H;T�H;;�H; �H;FlH;\NH;[)H;��G;\�G;	G;i2F;��D;80B;�Z>;#�8;w1;�*';+�;�Y;�+�:Q�:ׇ�:@t�:D)i:�2<:��:      ��:���:���:Z��:�;�Y;�';w�;��(;��0;�Y7;=�<;��@;�`C;CE;�wF;X8G;a�G;A�G;R)H;�LH;�iH;	�H;.�H;w�H;��H;��H;7�H;��H;��H;��H;/�H;��H;r�H;��H;~�H;��H;w�H;��H;q�H;��H;(�H;��H;��H;��H;7�H;��H;��H;{�H;.�H;�H;�iH;�LH;U)H;C�G;[�G;Z8G;�wF;CE;�`C;��@;A�<;�Y7;��0;~�(;u�;�';�Y;�;Z��:���:���:      �;��;;�z ;��$;D�);^/;
4;��8;<�<; $@;H�B;�D;��E;�F;�cG;��G;lH;{-H;\NH;�iH;�H;��H;��H;��H;��H;x�H;w�H;�H;��H;J�H;�H;�H;��H;��H;G�H;��H;A�H;��H;��H;�H;�H;K�H;��H;�H;v�H;t�H;��H;��H;��H;��H;�H;�iH;^NH;{-H;jH;��G;�cG;�F;��E;!�D;N�B;$@;8�<;��8;4;d/;>�);��$;�z ;�
;��;      )�1;*J2;2g3;�$5;{Y7;��9;Mg<;�>;�A;vC;�D;�E;H�F;*G;(�G;1�G;�H;^5H;�RH;ElH;�H;��H;��H;��H;\�H;<�H;2�H;	�H;��H;��H;a�H;��H;^�H;��H;��H;�H;L�H;�H;��H;��H;]�H;��H;d�H;�H;��H;�H;/�H;>�H;a�H;��H;��H;��H;�H;HlH;�RH;X5H;�H;1�G;*�G;*G;I�F;�E;�D;tC;�A;�>;Kg<;��9;�Y7;�$5;1g3;J2;      3,>;]Z>;��>;��?;H�@;��A;�C;�D;�E;��E;��F;�G;�}G;D�G;��G;�!H;B@H;\ZH;-qH;�H;+�H;~�H;��H;�H;��H;��H;�H;��H;��H;��H;<�H;�H;��H;{�H;@�H;��H;��H;��H;=�H;{�H;�H;�H;?�H;��H;��H;��H;�H;��H;��H;�H;��H;��H;.�H;�H;-qH;XZH;C@H;�!H;��G;B�G;�}G;�G;�F;��E;�E;�D;�C;��A;S�@;��?;��>;SZ>;      ��C;$	D;QBD;�D;�	E;��E;QF;�wF;��F;�<G;��G;��G;}�G;�H;c4H;�MH; dH;xH;��H;@�H;�H;��H;`�H;��H;!�H;��H;��H;O�H;V�H;��H;��H;Z�H;x�H;3�H;��H;>�H;A�H;8�H;��H;4�H;w�H;T�H;��H;��H;S�H;M�H;��H;��H;%�H;��H;a�H;��H;��H;=�H;��H;xH;dH;�MH;f4H;�H;��G;��G;��G;�<G;��F;�wF;RF;��E;�	E;��D;SBD;%	D;      OwF;EF;{�F;��F;��F;�G;�NG;�G;8�G;��G;��G;6H;l1H;�GH;v\H;YoH;��H;�H;��H;S�H;��H;��H;8�H;��H;��H;?�H;�H;�H;��H;y�H;�H;H�H;(�H;��H;g�H;��H;��H;��H;e�H;��H;)�H;C�H;�H;y�H;��H;�H;
�H;C�H;��H;��H;;�H;��H;��H;S�H;��H;�H;��H;ZoH;v\H;�GH;n1H;9H;��G;��G;9�G;�G;�NG;G;��F;��F;�F;DF;      �G;?�G;ߔG;�G;"�G;
�G;��G;��G;mH;�$H;8H;NJH;�[H;FlH;�{H;J�H;L�H; �H;S�H;p�H;��H;v�H;2�H;�H;��H;�H;��H;X�H;>�H;��H;'�H;�H;��H;}�H;��H;��H;	�H;��H;��H;��H;��H;�H;(�H;��H;=�H;W�H;��H;�H;��H;�H;4�H;z�H;��H;p�H;S�H;��H;O�H;N�H;�{H;ElH;�[H;RJH;8H;�$H;mH;��G;��G;�G;9�G;ݣG;ߔG;,�G;      m H;�H;gH;yH;�H;A!H;-H;�9H;�FH;ATH;�aH;9oH;C|H;̈H;~�H;Z�H;�H;�H;�H; �H;7�H;s�H;�H;��H;I�H;
�H;W�H;O�H;��H;��H;��H;��H;n�H;��H;�H;W�H;\�H;T�H;�H;��H;o�H;��H;��H;��H;��H;N�H;S�H;�H;M�H;��H;�H;u�H;9�H;�H;�H;�H;�H;^�H;~�H;̈H;C|H;:oH;�aH;ATH;�FH;�9H;-H;7!H;�H;vH;hH;�H;      �>H;z?H;BH;sFH;�KH;
SH;A[H;%dH;�mH;�wH;ҁH;ًH;��H;؞H;y�H;��H;�H;�H;�H;\�H;��H;�H;��H;��H;P�H;~�H;9�H;��H;�H;��H;��H;b�H;��H;/�H;i�H;��H;��H;��H;h�H;1�H;��H;`�H;��H;��H;�H;��H;6�H;�H;R�H;��H;��H;�H;��H;X�H;�H;�H;!�H;��H;{�H;֞H;��H;׋H;ԁH;�wH;�mH;%dH;A[H;SH;LH;sFH;BH;?H;      �hH;piH;hkH;mnH;�rH;�wH;�}H;S�H;n�H;̒H;:�H;��H;��H;��H;2�H;e�H;'�H;0�H;��H;��H;��H;��H;z�H;��H;��H;o�H;��H;��H;��H;��H;h�H;��H;�H;t�H;��H;��H;��H;��H;��H;v�H;�H;��H;i�H;��H;��H;��H;��H;t�H;��H;��H;�H;��H;��H;��H;��H;-�H;'�H;i�H;3�H;��H;��H;��H;<�H;ϒH;n�H;W�H;�}H;�wH;�rH;pnH;jkH;oiH;      3�H;׈H;3�H;d�H;��H;H�H;��H;��H;��H;�H;��H;�H;a�H;��H;��H;?�H;n�H;G�H;��H;�H;��H;J�H;^�H;:�H;��H;�H;'�H;��H;��H;n�H;��H;'�H;~�H;��H;��H;��H;��H;��H;��H;��H;��H;'�H;��H;l�H;��H;��H;%�H;	�H;��H;:�H;d�H;K�H;��H;�H;��H;D�H;q�H;@�H;��H;��H;c�H;�H;��H;�H;��H;��H;��H;@�H;��H;a�H;5�H;׈H;      A�H;��H;��H;@�H;��H;O�H;��H;2�H;�H;!�H;K�H;r�H;��H;w�H;�H;��H;��H;��H;��H;�H;2�H;�H;��H;�H;W�H;@�H;�H;��H;a�H;��H;!�H;t�H;��H;��H;��H;��H;�H;��H;��H;��H;��H;t�H;!�H;��H;`�H;��H; �H;C�H;Z�H;�H;��H;�H;0�H;�H;��H;��H;��H;��H;�H;t�H;��H;r�H;Q�H;$�H;�H;6�H;��H;R�H;��H;C�H;��H;��H;      �H;]�H;�H;J�H;�H;�H;��H;B�H;@�H;X�H;o�H;��H;��H;��H;l�H;3�H;��H;�H;+�H;
�H;��H;!�H;[�H;}�H;x�H;#�H;��H;u�H;��H;�H;}�H;��H;��H;��H;�H;�H;��H;�H;�H;��H;��H;��H;}�H;�H;��H;p�H;��H;&�H;{�H;}�H;a�H;!�H;��H;�H;+�H;�H;��H;6�H;l�H;��H;��H;��H;r�H;[�H;D�H;D�H;��H;�H;�H;D�H;�H;]�H;      �H;�H;��H;��H;��H;��H;��H;��H;��H;�H;��H;��H;h�H;��H;+�H;K�H;I�H;�H;��H;6�H;v�H;��H;��H;p�H;/�H;��H;y�H;��H;-�H;w�H;��H;��H;��H;��H;(�H;2�H;�H;0�H;'�H;��H;��H;��H;��H;s�H;+�H;��H;z�H;��H;3�H;p�H;��H;��H;r�H;/�H;��H;�H;L�H;I�H;+�H;��H;g�H;��H;��H;�H;��H;��H;��H;��H;��H;��H;��H;�H;      ��H;��H;L�H;�H;�H;@�H;��H;�H;d�H;n�H;b�H;u�H;u�H;U�H;.�H;��H;��H;�H;u�H;��H;��H;��H;|�H;0�H;��H;]�H;��H;�H;h�H;��H;��H;��H;�H;)�H;�H;'�H;F�H;(�H;	�H;)�H;�H;��H;��H;��H;e�H;�H;��H;`�H;��H;2�H;��H;��H;��H;��H;q�H;�H;��H;��H;-�H;T�H;v�H;x�H;g�H;q�H;i�H;��H;��H;B�H;�H;�H;M�H;��H;      �H;3�H;��H;-�H;�H;I�H;��H;,�H;��H;z�H;-�H;��H;��H;L�H;��H;n�H;��H;2�H;m�H;��H;��H;D�H;��H;��H;5�H;��H;��H;X�H;��H;��H;��H;��H;�H;5�H;)�H;�H;2�H;�H;'�H;6�H;�H;��H;��H;��H;��H;W�H;��H;��H;8�H;��H;�H;A�H;{�H;��H;j�H;3�H;��H;o�H;��H;M�H;��H;��H;2�H;}�H;��H;0�H;��H;L�H;!�H;'�H;��H;A�H;      q�H;��H;:�H;��H;��H;��H;��H;E�H;��H;R�H;�H;��H;P�H;�H;��H;��H;c�H;��H;��H;��H;��H;��H;H�H;��H;>�H;��H;�H;c�H;��H;��H;��H;�H;��H;�H;F�H;0�H; �H;/�H;C�H;�H;�H;�H;��H;��H;��H;_�H;	�H;��H;A�H;��H;O�H;��H;��H;��H;��H;��H;c�H;�H;��H;�H;R�H;��H;�H;U�H;��H;I�H;��H;��H;��H;��H;:�H;��H;      �H;5�H;��H;+�H;�H;O�H;��H;,�H;��H;z�H;,�H;��H;��H;M�H;��H;n�H;��H;2�H;m�H;��H;��H;F�H;��H;��H;5�H;��H;��H;X�H;��H;��H;��H;��H;�H;5�H;,�H;�H;2�H;�H;'�H;5�H;�H;��H;��H;��H;��H;T�H;��H;��H;7�H;��H;�H;@�H;{�H;��H;j�H;3�H;��H;o�H;��H;J�H;��H;��H;2�H;z�H;��H;0�H;��H;L�H;"�H;.�H;��H;<�H;      ��H;��H;F�H;�H;�H;>�H;��H;��H;d�H;n�H;b�H;u�H;s�H;T�H;.�H;��H;��H;�H;u�H;��H;��H;��H;|�H;2�H;��H;[�H;��H;�H;i�H;��H;��H;��H;�H;(�H;�H;(�H;F�H;(�H;	�H;)�H;�H;��H;��H;��H;e�H;	�H;��H;`�H;��H;0�H;��H;��H;��H;��H;q�H;�H;��H;��H;,�H;R�H;v�H;x�H;d�H;n�H;e�H;��H;��H;>�H;�H;	�H;L�H;��H;      �H;�H;��H;��H;��H;��H;��H;��H;��H;�H;��H;��H;e�H;��H;-�H;I�H;L�H;�H;��H;5�H;x�H;��H;��H;r�H;2�H;��H;y�H;��H;/�H;w�H;��H;��H;��H;��H;)�H;0�H;�H;0�H;%�H;��H;��H;��H;��H;s�H;(�H;��H;z�H;��H;0�H;k�H;��H;��H;n�H;/�H;��H;�H;J�H;K�H;+�H;��H;e�H;��H;��H;�H;��H;��H;��H;��H; �H;��H;��H;�H;      �H;a�H;�H;G�H;��H;�H;��H;G�H;A�H;Z�H;o�H;��H;��H;��H;o�H;6�H;��H;�H;,�H;�H;��H;"�H;Z�H;~�H;{�H;"�H;��H;s�H;��H;!�H;}�H;��H;��H;��H;�H;	�H;��H;�H;�H;��H;��H;��H;{�H;�H;��H;n�H;��H;%�H;x�H;z�H;b�H;�H;��H;�H;+�H;�H;��H;4�H;l�H;��H;��H;��H;o�H;X�H;D�H;G�H;��H;�H;�H;M�H;�H;[�H;      4�H;��H;��H;A�H;��H;^�H;��H;3�H;�H;!�H;M�H;r�H;��H;u�H;�H;��H;��H;��H;��H;�H;6�H;�H;��H;�H;Z�H;A�H;��H;��H;e�H;��H;!�H;s�H;��H;��H;��H;��H;�H;��H;��H;��H;��H;s�H;�H;��H;^�H;��H;��H;D�H;W�H;�H;��H;�H;-�H;�H;��H;��H;��H;��H;�H;t�H;��H;r�H;K�H;"�H;�H;5�H;��H;S�H;��H;C�H;��H;��H;      &�H;ֈH;3�H;`�H;��H;I�H;��H;��H;��H;�H;��H;�H;a�H;��H;��H;@�H;p�H;G�H;��H;�H;��H;N�H;a�H;<�H;��H;�H;$�H;��H;��H;o�H;��H;(�H;�H;��H;��H;��H;��H;��H;��H;��H;��H;'�H;��H;k�H;��H;��H;$�H;�H;��H;6�H;e�H;K�H;��H;�H;��H;D�H;r�H;@�H;��H;��H;a�H;�H;��H;�H;��H;��H;��H;G�H;��H;i�H;9�H;ԈH;      �hH;siH;akH;wnH;�rH;�wH;�}H;Z�H;q�H;ϒH;:�H;��H;��H;��H;3�H;g�H;'�H;0�H;��H;��H;��H;��H;{�H;��H;��H;o�H;��H;��H;��H;��H;i�H;��H;�H;t�H;��H;��H;��H;��H;��H;t�H;�H;��H;h�H;��H;��H;��H;��H;v�H;��H;��H;��H;��H;��H;��H;��H;-�H;'�H;h�H;2�H;��H;��H;��H;<�H;ϒH;n�H;Z�H;�}H;�wH;�rH;{nH;kkH;oiH;      �>H;z?H;!BH;pFH;�KH;SH;>[H;%dH;�mH;�wH;сH;ًH;��H;ٞH;|�H;��H;�H;�H;�H;Z�H;��H;�H;��H;��H;U�H;{�H;4�H;��H;�H;��H;��H;d�H;��H;.�H;h�H;��H;��H;��H;f�H;.�H;��H;a�H;��H;��H;�H;��H;7�H;��H;O�H;��H;��H;�H;��H;Z�H;�H;�H;�H;��H;{�H;֞H;��H;֋H;ҁH;�wH;�mH;*dH;B[H;
SH;LH;mFH; BH;y?H;      y H;�H;]H;wH;�H;L!H;-H;�9H;�FH;ATH;�aH;9oH;E|H;̈H;��H;^�H;�H;�H;�H;�H;:�H;w�H;�H;��H;O�H;�H;S�H;N�H;��H;��H;��H;��H;l�H;��H;�H;T�H;\�H;U�H;�H;��H;o�H;��H;��H;��H;��H;K�H;U�H;�H;I�H;��H;	�H;u�H;7�H;�H;�H;�H;�H;]�H;��H;ʈH;C|H;9oH;�aH;ATH;�FH;�9H;-H;<!H;�H;vH;gH;�H;      �G;I�G;۔G;��G;1�G;�G;��G;��G;oH;�$H;8H;RJH;�[H;FlH;�{H;M�H;O�H;�H;T�H;n�H;��H;z�H;0�H;#�H;��H;�H;��H;W�H;@�H;��H;'�H;�H;��H;~�H;��H;��H;�H;��H;��H;~�H;��H;�H;(�H;��H;=�H;W�H;��H;�H;��H;�H;4�H;x�H;��H;r�H;T�H;��H;O�H;N�H;�{H;ElH;�[H;QJH;8H;�$H;lH;��G;��G;
�G;8�G;�G;ޔG;4�G;      CwF;DF;��F;��F;��F;�G;�NG;�G;;�G;��G;��G;9H;n1H;�GH;w\H;\oH;��H;�H;��H;S�H;��H;��H;8�H;��H;��H;>�H;�H;�H;��H;x�H;	�H;G�H;&�H;��H;e�H;��H;��H;��H;b�H;��H;&�H;G�H;�H;y�H;��H;�H;�H;C�H;��H;��H;;�H;��H;��H;T�H;��H;�H;��H;\oH;z\H;�GH;l1H;6H;��G;��G;2�G;�G;�NG;�G;��F;��F;m�F;6F;      ��C;#	D;MBD;�D;�	E;��E;RF;�wF;��F;�<G;��G;��G;�G;�H;h4H;�MH;dH;xH;��H;?�H;��H;��H;`�H;��H;%�H;��H;��H;M�H;V�H;��H;��H;Z�H;u�H;3�H;��H;:�H;?�H;:�H;��H;3�H;x�H;Z�H;��H;��H;S�H;L�H;��H;��H;!�H;��H;c�H;��H;��H;?�H;��H;xH;dH;�MH;i4H;�H;��G;��G;�G;�<G;��F;�wF;OF;��E;�	E;��D;MBD;!	D;      ,>;EZ>;��>;��?;A�@;��A;�C;�D;�E;��E;�F;�G;�}G;B�G;��G;�!H;C@H;]ZH;.qH;�H;/�H;��H;��H;��H;��H;��H;�H;��H;��H;��H;=�H;�H;��H;z�H;=�H;��H;��H;��H;;�H;x�H;��H;�H;A�H;��H;��H;��H;�H;��H;��H;�H;��H;��H;/�H;�H;/qH;YZH;E@H;�!H;��G;D�G;�}G;�G;�F;��E;�E;�D;�C;��A;W�@;Ư?;��>;*Z>;      �1;$J2;$g3;�$5;yY7;��9;Gg<;�>;�A;uC;	�D;	�E;G�F;*G;+�G;3�G;�H;^5H;�RH;FlH;�H;��H;��H;��H;a�H;8�H;2�H;�H;��H;{�H;b�H;��H;]�H;��H;��H;�H;N�H;�H;��H;��H;^�H;��H;g�H;��H;��H;	�H;4�H;>�H;]�H;��H;��H;��H;�H;HlH;�RH;X5H;�H;1�G;,�G;*G;H�F;�E;
�D;uC;�A;�>;Fg<;��9;xY7;�$5;&g3;J2;      �;��;�
;�z ;��$;K�);b/;4;��8;8�<;�#@;O�B;�D;��E;�F;�cG;��G;lH;z-H;^NH;�iH;�H;��H;��H;��H;��H;x�H;w�H;�H;��H;J�H;�H;�H;��H;��H;C�H;��H;F�H;��H;��H;�H;�H;N�H;��H;�H;w�H;z�H;��H;��H;��H;��H;�H;�iH;`NH;{-H;jH;��G;�cG;�F;��E;�D;L�B;�#@;8�<;��8;4;[/;3�);��$;�z ;�
;��;      ��:��:��:n��:�;�Y;�';x�;��(;��0;�Y7;@�<;��@;�`C;CE;�wF;X8G;^�G;C�G;U)H;�LH;�iH;	�H;/�H;|�H;��H;��H;7�H;��H;��H;��H;-�H;��H;q�H;��H;z�H;��H;{�H;��H;n�H;��H;,�H;��H;��H;��H;7�H;��H;��H;x�H;0�H;	�H;�iH;�LH;W)H;C�G;[�G;Z8G;�wF;CE;�`C;��@;@�<;�Y7;��0;��(;{�;�';�Y;�;f��:��:���:      ��:̠:�2<:�)i:8t�:Ӈ�:Y�:�+�:�Y;+�;�*';v1;#�8;�Z>;70B;��D;h2F;
G;Y�G;��G;[)H;^NH;IlH; �H;<�H;T�H;n�H;�H;[�H;��H;�H;��H;�H;2�H;��H;��H;��H;��H;��H;.�H;�H; �H;�H;��H;[�H;�H;q�H;W�H;8�H;#�H;IlH;]NH;Y)H;��G;Z�G;	G;j2F;��D;80B;�Z>;#�8;s1;�*';(�;�Y;�+�:Q�:Ç�:Bt�:l)i:�2<:��:      ⥥�4X��� ����=�h۷� ߤ8��:�P�:}P�:z��:$`;n;�*;�$5;�g<;�<A;�BD;�F;�G;X�G;D�G;z-H;�RH;-qH;��H;��H;N�H;�H;�H;��H;��H;��H;'�H;��H;t�H;j�H;��H;j�H;q�H;��H;%�H;��H;��H;��H;�H;�H;S�H;��H;��H;/qH;�RH;y-H;A�G;Y�G;�G;�F;�BD;�<A;�g<;�$5;�*;j;#`;t��:}P�:�P�:��:�ޤ8h۷���=�!��,X��      �1��"Ȅ�֨u��PV�n.�����W��(��@X�9+i:ء�:�+�:�;�t%;�J2;J;;��@;WD;�F;G;Z�G;hH;[5H;VZH;
xH;�H;��H;�H;�H;,�H;A�H;��H;�H; �H;�H;2�H;��H;2�H;�H;��H;�H;��H;D�H;3�H;�H;�H; �H;�H;xH;VZH;Z5H;gH;U�G;G;�F;WD;��@;H;;�J2;�t%;�;�+�:ܡ�:+i:@X�98��W�����q.��PV�ߨu�"Ȅ�      Y��L�	������#Tʻ�R��3|�l.�$Ⱥ���Y�9"u�:��:�Y;v�!;��0;Օ:;��@;�BD;h2F;]8G;��G;�H;@@H;�cH;��H;H�H;�H;�H; �H;g�H;��H;��H;C�H;��H;��H;[�H;��H;��H;B�H;��H;��H;j�H;%�H;�H;�H;K�H;��H;�cH;B@H;�H;��G;V8G;i2F;�BD;��@;Օ:;��0;v�!;�Y;��:u�:Y�9���Ⱥm.�3|��R��)Tʻ�����J�	�      ��x��[t���g�NT�_�:�������(����1��R�(�4W����t��n`:S��:�\;{ ;��0;K;;�<A;��D;�wF;�cG;1�G;�!H;�MH;YoH;G�H;Y�H;��H;e�H;<�H;��H;/�H;G�H;��H;k�H;��H;k�H;��H;D�H;-�H;��H;=�H;i�H;��H;]�H;J�H;UoH;�MH;�!H;1�G;�cG;�wF;��D;�<A;H;;��0;�z ;�\;S��:�n`:��t�6W��R�(��1��(���������a�:�OT���g��[t�      6,˼��Ǽ�"���뮼w��#G��*�[�_y-�����.��ŕb�x0㺰ط��4<:�L�:�\;r�!;�J2;�g<;00B;CE;�F;,�G;��G;b4H;v\H;�{H;~�H;}�H;2�H;��H;�H;i�H;'�H;&�H;��H;��H;��H;&�H;'�H;i�H;�H;��H;3�H;}�H;��H;�{H;r\H;^4H;��G;*�G;�F;CE;30B;�g<;�J2;r�!;�\;�L�:�4<:�ط�x0�Ǖb��.�����^y-�+�[�#G��w���뮼�"����Ǽ      *���k��Jv�|t�C�Ѽ�뮼,X��m�W������׻�Ǆ�����5<:Y��:�Y;�t%;�$5;�Z>;�`C;��E;*G;B�G;�H;�GH;FlH;ʈH;؞H;��H;��H;p�H;��H;��H;M�H;C�H;�H;I�H;H�H;��H;��H;n�H;��H;��H;ٞH;ɈH;ClH;�GH;�H;D�G;*G;��E;�`C;�Z>;�$5;�t%;�Y;Q��:�4<:�����Ǆ���׻���l�W�,X���뮼C�Ѽ~t�Jv���k�      Cm��Fi��&^�_�L�O�6�(����}ռnT����x���0����������ط��n`:��:�;�*; �8; �@;�D;I�F;�}G;�G;k1H;�[H;E|H;��H;��H;\�H;��H;��H;b�H;k�H;��H;G�H;��H;h�H;`�H;��H;��H;\�H;��H;��H;E|H;�[H;g1H;y�G;�}G;I�F;�D;��@;!�8;�*;�;��:�n`:�ط��������껿�0���x�mT��}ռ��(��P�6�_�L��&^��Fi�      K��r;��A�������섽x�e��?��k�{t�鷼G���e7�����Ǆ�p0���t�u�:�+�:j;q1;G�<;K�B;�E;�G;��G;3H;QJH;3oH;׋H;��H;�H;n�H;��H;��H;m�H;��H;��H;��H;j�H;��H;��H;m�H;�H;��H;ًH;3oH;PJH;/H;��G;�G;	�E;I�B;=�<;s1;j;�+�:u�:��t�p0� Ȅ���껄e7�G��鷼{t��k��?�w�e��섽���A���r;��      o���$��s��ӽ�'��?�������Z��Q+�����"��G����0���׻ȕb�:W���X�9̡�:`;�*';�Y7;�#@;	�D;��F;�G;��G;8H;�aH;сH;7�H;~�H;K�H;n�H;|�H;Z�H;(�H;�H;(�H;Z�H;{�H;k�H;H�H;|�H;<�H;ҁH;�aH;8H;��G;�G;�F;	�D;�#@;�Y7;�*';`;ʡ�:�X�9>W��̕b���׻��0�G���"������Q+��Z����?����'���ӽ�s�$��      �!,�7)��K ��������޽������Fi��0����鷼��x�����.��Q�(�����*i:x��:'�;��0;8�<;rC;��E;�<G;��G;�$H;:TH;�wH;˒H;�H;"�H;[�H;�H;g�H;s�H;Q�H;s�H;f�H;�H;X�H;!�H;�H;ΒH;�wH;;TH;�$H;��G;�<G;��E;tC;4�<;��0;)�;r��:�*i:���T�(��.�������x�鷼����0��Fi�������޽�������K �7)�      (�j��f��Z�y�F��>/��^�m�����ŽF ���Fi��Q+�{t�mT��m�W�����1��(Ⱥ�W�9uP�:�Y;��(;��8;�A;�E;��F;8�G;rH;�FH;�mH;n�H;��H;�H;K�H;��H;a�H;��H;��H;��H;a�H;��H;G�H;�H;��H;o�H;�mH;�FH;sH;8�G;��F;�E;�A;��8;}�(;�Y;oP�:�W�9,Ⱥ�1�����m�W�nT��{t�Q+��Fi�F ����Žm����^��>/�y�F��Z��f�      ��v���x�H����f��SC��K �nn����Ž����Z��k�}ռ-X��`y-�,���s.����P�:�+�:��;4;�>;�D;�wF; �G;��G;�9H;'dH;V�H;��H;5�H;K�H;��H;��H;+�H;G�H;+�H;��H;��H;H�H;2�H;��H;]�H;*dH;�9H;��G;�G;�wF;�D;�>;4;x�;�+�:�P�:���p.�-���ay-�-X��}ռ�k��Z������Žnn���K ��SC��f�H���x�v���      ��˾��Ǿ���� ���V͓�Y�x���J��K �m���������?����뮼+�[����3|��W��|�:=�:�';b/;=g<;�C;FF;�NG;��G;-H;=[H;�}H;��H;��H;��H;��H;��H;��H;��H;��H;��H;��H;��H;��H;��H;�}H;@[H;
-H;��G;�NG;DF;�C;Bg<;`/;�';C�:x�:�W��3|����+�[��뮼���?������m����K ���J�Z�x�V͓� ���������Ǿ      s� ��������{Ծj���v���Z�x��SC��^��޽?���x�e�'��C�Ѽ$G������R������ݤ8Ç�:�Y;D�);��9;��A;��E;G;�G;A!H;SH;�wH;N�H;]�H;�H;��H;L�H;V�H;��H;V�H;L�H;��H;�H;]�H;I�H;�wH;SH;C!H;�G;�G;��E;��A;��9;C�);�Y;ɇ�:`ݤ8����R�����$G��C�Ѽ(��x�e�?����޽�^��SC�Z�x�v���j����{Ծ�쾠���      ����D�l�s� �V�ݾj���V͓��f��>/�����'���섽O�6�~t�w��^�:�'Tʻ�.�8۷�@t�:�;��$;�Y7;R�@;�	E;��F;)�G;�H;
LH;�rH;��H;��H;��H;��H;�H;'�H;��H;"�H;�H;��H;��H;��H;��H;�rH;
LH;�H;0�G;��F;�	E;S�@;�Y7;��$;�;Dt�:H۷�}.�(Tʻ^�:�w��t�O�6��섽�'������>/��f�V͓�j���V�ݾs� �l��D�      �7�v3�/�'����s� ��{Ծ ���H���y�F�����ӽ���^�L�Jv��뮼QT����PV���=�\)i:|��:�z ;}$5;��?;�D;��F;�G;uH;fFH;tnH;e�H;N�H;M�H;��H;�H;2�H;��H;.�H;�H;��H;M�H;N�H;b�H;~nH;fFH;sH;�G;��F;�D;��?;{$5;�z ;r��:p)i:��=��PV���QT��뮼Jv�^�L�����ӽ���y�F�H��� ����{Ծs� ����/�'�v3�      �N��TI���;�/�'�l��쾀���x󐾳Z��K ��s�@����&^���"����g����Ѩu�� ���2<:��:�
;8g3;��>;XBD;w�F;�G;nH;BH;`kH;0�H;��H;�H;��H;C�H;��H;$�H;��H;C�H;��H;	�H;��H;,�H;ekH;BH;lH;�G;��F;UBD;��>;4g3;�
;��:�2<:� ��Ҩu������g��"����&^�A����s潥K ��Z�x󐾀�����l�/�'���;��TI�      `]�d�W��TI�v3��D�������Ǿv����f�8)�$��r;���Fi��k���Ǽ�[t�N�	�+Ȅ�X��Ԡ:��:��;,J2;TZ>;*	D;=F;=�G;�H;�?H;xiH;ňH;��H;T�H;�H;��H;7�H;��H;1�H;��H;�H;Q�H;��H;��H;iH;�?H;�H;>�G;IF;$	D;QZ>;$J2;��;��:ܠ: X��*Ȅ�N�	��[t���Ǽ�k��Fi�r;��$��8)��f�v�����Ǿ�����D�v3��TI�d�W�      1�$��� ����#��?��'�þ�*��0Dx���=�����Pν���#'K��c���p�V����E^���S�|w[:���:e;)�4;E`?;�mD;U�F;OvG;�G;@H;dOH;�sH;��H;|�H;��H;�H;U�H;&�H;O�H;�H;��H;{�H;��H;�sH;mOH;=H;�G;QvG;a�F;�mD;A`?;"�4;e;���:�w[:��S�E^����p�V����c�#'K�����Pν�����=�0Dx��*��'�þ?��#������� �      �� ����R��O��/������0��4�s�ր:�g9��ʽ1Z����G��8�
.���5S�����/X�x�D�nBd:�B�: ;��4;ʈ?;�~D;�F;yG;��G;P H;-PH;tH;�H;΢H;ɰH;,�H;r�H;5�H;n�H;,�H;ưH;̢H;�H;tH;3PH;O H;��G;yG;�F;�~D;ǈ?;��4; ;�B�:vBd:|�D��/X���껭5S�
.���8���G�1Z���ʽg9�ր:�4�s��0�����/��O��R�����      ���R��8�
������Yؾ���ޥ����f���0�Z[�N8��ϐ���>�����JȤ��6H�a�ܻrF�����}:��:d";/�5;��?;W�D;��F;�G;��G;2#H;cRH;�uH;I�H;ƣH;x�H;źH;�H;��H;�H;ĺH;v�H;��H;F�H;�uH;iRH;0#H;��G;�G;��F;S�D;��?;&�5;_";��:�}:Ԗ�rF�b�ܻ�6H�IȤ������>�ϐ��N8��Z[���0���f�ޥ������Yؾ����8�
�Q��      #��O������>I�(�þ�R��;���tS��Q"��s������}��0��켈�����6�F�ƻ9}*������:}x;Z%;�l7;ڳ@;��D;��F;��G;��G;�'H;�UH;`xH;Q�H;I�H;��H;��H;��H;z�H;��H;��H;��H;D�H;M�H;XxH;�UH;�'H;��G;��G;��F;��D;ٳ@;�l7;V%;zx;��:���:}*�F�ƻ��6��������0���}�����s��Q"�tS�;����R��(�þ=Iᾣ���O��      ?��/�待Yؾ(�þĪ�|쏾�k�ր:�~�{�ؽ�����c�]y���Ҽ����C� �j�+�� "(7A�:��
;��(;�_9;��A;h\E;o�F;��G;��G;�.H;�ZH;�{H;�H;L�H;S�H;�H;��H;x�H;��H;�H;Q�H;H�H;�H;�{H;�ZH;�.H;��G;��G;u�F;g\E;��A;z_9;��(;��
;I�: (7,��j�C� �������Ҽ]y��c�����{�ؽ~�ր:��k�|쏾Ī�(�þ�Yؾ/��      '�þ��� ����R��|쏾4�s��H�����������ΐ����D��c�����<�f�S,�����P��H�9ɳ�:�;"j-;M�;;u�B;��E;[G;��G;��G;�6H;�`H;Z�H;O�H;ةH;Q�H;��H;U�H;��H;P�H;��H;M�H;ҩH;L�H;V�H;�`H;�6H;��G;��G;bG;��E;p�B;I�;;j-;�;ͳ�:@�9�P�����T,�<�f������c���D�ΐ�������������H�4�s�|쏾�R�� ������      �*���0��ޥ��;����k��H��#%�Z[��Pνt��`�f�2/%���伆���u�=��?ػ�FL���D�h�R:��:4�;42;��=;��C;f0F;FGG;��G;&H;�?H;�gH;��H;.�H;��H;��H;��H;��H;u�H;��H;��H;��H;��H;*�H;��H;�gH;�?H;#H;��G;JGG;f0F;��C;��=;42;/�;��:\�R:��D��FL��?ػt�=��������2/%�`�f�t���PνZ[��#%��H��k�;���ޥ���0��      0Dx�4�s���f�tS�ր:����Z[��7ս�榽��}���;��8�U�����r����:G��	�� ͬ�%��:	�;�}$;Ä6;�?;��D;ƔF;�pG;��G;�H;"JH;AoH;>�H;y�H; �H;9�H;��H;��H;)�H;��H;��H;9�H;��H;s�H;9�H;GoH;$JH;�H;��G;�pG;ǔF;�D;��?;Ä6;�}$;�;!��: ͬ�	��;G�������r�U����8���;���}��榽�7սZ[����׀:�sS���f�4�s�      ��=�ր:���0��Q"�~������Pν�榽@����G�1����Ҽ ��IE:�<�ܻ�D^�����`i:=��:�;8|,;��:;K�A;AiE;��F;�G;�G;�(H;2UH;}wH;q�H;$�H;��H;��H;��H;��H;�H;��H;��H;�H;��H;#�H;o�H;�wH;5UH;�(H;~�G;�G;��F;<iE;K�A;��:;6|,;�;?��:Xi:�����D^�<�ܻHE:� ����Ҽ1����G�?���榽�Pν����~��Q"���0�ր:�      ���g9�Z[��s�z�ؽ���t����}���G������1c��W�V�E,��*����� ����:��:Q ;c�3;�0>;ÚC;�F;�8G;*�G;kH;�7H;�`H;�H;�H;��H;N�H;��H;I�H;��H;�H;��H;I�H;��H;G�H;��H;�H;�H;�`H;�7H;iH;'�G;�8G;�F;ÚC;�0>;_�3;V ;��:��:�������*��E,�V�V�0c��������G���}�t�����{�ؽ�s�Z[�g9�      �Pν�ʽN8���������ΐ��`�f���;�1�����BȤ�3�f�)��Lߵ�Vo5���D�0�-:D��:�>;�+;�_9;�A;c�D; �F;�vG;��G;H;uGH;ZlH;��H;��H;��H;/�H;��H;��H;�H;%�H;�H;��H;��H;*�H;�H;��H;ǈH;`lH;vGH;H;��G;�vG;�F;e�D;�A;�_9;�+;�>;@��:<�-:��D�To5�Kߵ�)��2�f�BȤ����1����;�`�f�ΐ���������N8���ʽ      ���1Z��ϐ����}��c���D�2/%��8���Ҽ0c��2�f�����ƻ/X�\������9�::�;�";��3;=>;?YC;r�E;�G;�G;c�G;�,H;WH;xH;��H;/�H;�H;�H;��H;3�H;G�H;0�H;E�H;3�H;��H;�H;�H;2�H;��H;xH;WH;�,H;`�G;�G;�G;w�E;DYC;=>;��3;�";:�;	�:���9Z���|/X��ƻ���1�f�0c����Ҽ�8�2/%���D��c���}�ϐ��1Z��      #'K���G��>��0�\y��c����T��� ��V�V�(���ƻ�od���º {(7�4�:���:��;�P.;ϡ:;zA;)�D;ƨF;MnG;8�G;�H;�@H;$fH;]�H;.�H;��H;׸H;��H;��H;��H;~�H;9�H;}�H;��H;��H;��H;иH;��H;5�H;c�H;%fH;�@H;�H;<�G;KnG;ǨF;-�D;zA;ڡ:;�P.;��;���:�4�: ~(7|�º�od��ƻ(��V�V� ��S�����伕c�^y��0��>���G�      �c��8���������Ҽ����������r�HE:�D,�Jߵ��/X���º Ǭ�d�}:�:�;H�);#m7;�?;��C;F;U)G;�G;E�G;�)H;�SH;�tH;\�H;|�H;�H;��H;��H;��H;�H;��H;M�H;��H;�H;��H;��H;��H;�H;��H;f�H;�tH;�SH;�)H;I�G;�G;Y)G;F;��C;�?;%m7;E�);�;� �:l�}:�Ƭ���º|/X�Hߵ�E,�GE:���r�����������Ҽ�켶����8�      ��.��JȤ���������;�f�t�=����=�ܻ�*��Qo5�h��� z(7h�}:�n�:*�;�>&;��4;��=;��B;�E;�F;��G;��G;+H;�AH;�eH;<�H;јH;Y�H;ڷH;i�H;!�H;��H;m�H;��H;Q�H;��H;k�H;��H;�H;c�H;ݷH;_�H;ؘH;A�H;�eH;{AH;/H;��G;��G;�F;�E;��B;��=;��4;�>&;)�;�n�:t�}: |(7\���No5��*��9�ܻ���t�=�9�f���������KȤ�.��      j�V��5S��6H���6�C� �T,��?ػ8G���D^������D����9�4�:�:)�;�%;��3;�<;UB;�E;��F;�XG;��G;E H;h0H;LWH;YvH;�H;{�H;��H;��H;��H;o�H;O�H;��H;��H;:�H;��H;��H;N�H;l�H;��H;��H;ñH;�H;�H;[vH;GWH;l0H;D H;��G;�XG;��F;�E;VB;�<;��3;�%;,�; �:�4�:���9��D�����D^�6G���?ػQ,�F� ���6��6H��5S�      ��ﻬ��g�ܻH�ƻf󩻸���FL����������H�-:�:���:�;�>&;��3;Q9<;�A;ذD;>ZF;5G;��G;��G;i!H;,JH;/kH;��H;��H;c�H;��H;��H;��H;��H;��H;��H;f�H;��H;b�H;��H;��H;��H;��H;��H;��H;g�H;��H;��H;*kH;/JH;i!H;��G;��G;5G;EZF;۰D;�A;T9<;��3;�>&;�;���:�:T�-:����������FL����j�L�ƻk�ܻ���      �D^��/X�rF�.}*����P����D��̬�`i:��:J��:5�;��;E�);��4;�<;
�A;#�D;s9F;�G;m�G;C�G;=H;?H;ZaH;}H;|�H;v�H;��H;�H;��H;b�H;�H;�H;��H;(�H;��H;%�H;��H;�H;{�H;]�H;��H;�H;��H;v�H;{�H;}H;\aH;?H;7H;C�G;n�G;�G;t9F; �D;�A;�<;��4;E�);��;7�;V��:��:ti:@̬���D��P����6}*�rF��/X�      @�S���D�Ж�膪� !(7��9��R:-��:C��:��:�>;�";�P.;'m7;��=;VB;ڰD;{9F;G;�G;R�G;�H;�6H;iYH;�uH;�H;�H;��H;��H;��H;�H;��H;�H;8�H;a�H;��H;��H;��H;^�H;6�H;�H;��H; �H;��H;��H;��H;�H;�H;�uH;iYH;�6H;�H;T�G;�G;G;v9F;ްD;SB;��=;'m7;�P.;�";�>;��:I��:/��:��R:p�9 "(7P���Ж���D�      tw[:^Bd:,�}:��:7�:ϳ�:�:	�;�;W ;�+;��3;١:;�?;��B;�E;EZF;�G;�G;o�G;>H;S1H;�SH;`pH;ׇH;H�H;�H;{�H;��H;��H;��H;��H;r�H;"�H;��H;�H;\�H;�H;��H;!�H;p�H;��H;��H;��H;��H;|�H;�H;D�H;ۇH;`pH;�SH;S1H;AH;o�G;�G;�G;EZF;�E;��B;�?;١:;��3;�+;W ;�;�;�:ݳ�:C�:��: �}:"Bd:      &��:�B�:���:lx;��
;�;0�;�}$;6|,;b�3;�_9;7>;zA;��C;�E;�F;5G;u�G;T�G;=H;�/H;�PH;mH;H�H;��H;��H;n�H;��H;��H;�H;\�H;��H;��H;��H;k�H;L�H;��H;D�H;j�H;��H;��H;��H;^�H;�H;��H;��H;i�H;��H;��H;E�H;�lH;�PH;�/H;=H;U�G;q�G;5G;�F;�E;��C;zA;=>;�_9;b�3;2|,;�}$;6�;�;��
;mx;І�:�B�:      e; ;n";f%;��(;!j-;02;��6;��:;�0>;�A;>YC;-�D;
F;�F;�XG;��G;I�G;�H;T1H;�PH;�kH;t�H;{�H;1�H;,�H;׼H;��H;��H;�H;m�H;��H;v�H;p�H;��H;a�H;��H;[�H;��H;p�H;u�H;��H;n�H;�H;��H;��H;ӼH;.�H;5�H;x�H;m�H;�kH;�PH;S1H;�H;F�G;��G;�XG;�F;F;.�D;EYC;�A;�0>;��:;Ȅ6;62;j-;��(;X%;d";  ;      ?�4;��4;%�5;�l7;y_9;T�;;��=;	�?;U�A;ʚC;o�D;x�E;ʨF;_)G;��G;�G;��G;BH;�6H;�SH;�lH;r�H;��H;�H;��H;O�H;#�H;2�H;��H;��H;�H;��H;2�H;��H;��H;b�H;��H;[�H;��H;��H;2�H;��H;�H;�H;��H;3�H;�H;P�H;��H;�H;��H;r�H;mH;�SH;�6H;=H;��G;�G;��G;])G;ͨF;~�E;q�D;ǚC;U�A;	�?;��=;P�;;�_9;�l7;%�5;��4;      B`?;ш?;��?;ӳ@;��A;u�B;��C;�D;8iE;�F;#�F;�G;KnG;�G;��G;F H;i!H;?H;iYH;[pH;E�H;t�H;�H;C�H;��H;%�H;C�H;�H;��H;s�H;S�H;��H;��H;��H;��H;<�H;M�H;5�H;��H;��H;��H;��H;V�H;r�H;��H;�H;?�H;(�H;��H;A�H;�H;w�H;C�H;ZpH;hYH;?H;i!H;H H;��G;�G;KnG;�G;&�F;�F;?iE;��D;��C;e�B;��A;ѳ@;��?;Ȉ?;      �mD;�~D;P�D;��D;a\E;��E;r0F;ǔF;��F;�8G;�vG;�G;>�G;O�G;/H;o0H;5JH;eaH;�uH;��H;��H;5�H;��H;��H;��H;��H;j�H;�H;��H;��H;\�H;A�H;��H;��H;��H;��H;)�H;��H;��H;��H;��H;;�H;_�H;��H;��H;�H;d�H;��H;��H;��H;��H;6�H;��H;ۇH;�uH;baH;6JH;r0H;2H;M�G;@�G;��G;�vG;�8G;��F;ʔF;u0F;��E;m\E;��D;S�D;�~D;      M�F;�F;��F;��F;l�F;dG;PGG;�pG;�G;4�G;��G;i�G;�H;*H;AH;NWH;/kH;}H;�H;A�H;��H;(�H;K�H;%�H;��H;/�H;��H;�H;��H;�H;�H;��H;��H;��H;:�H;��H;��H;��H;7�H;��H;��H;��H;�H;�H;��H;�H;��H;3�H;��H;"�H;L�H;)�H;��H;A�H;�H;}H;0kH;NWH;~AH;*H;�H;j�G;��G;2�G;�G;�pG;QGG;[G;��F;��F;��F;�F;      dvG;yG;
�G;��G;��G;��G;��G;��G;~�G;lH;!H;�,H;�@H;�SH;�eH;[vH;��H;�H;�H;�H;p�H;ӼH;#�H;D�H;g�H;��H;c�H;]�H;��H;��H;^�H;��H;��H;@�H;��H;&�H;#�H;�H;��H;B�H;��H;��H;`�H;��H;��H;\�H;^�H;��H;k�H;@�H;#�H;ԼH;r�H;�H;�H;y�H;��H;]vH;�eH;�SH;�@H;�,H;!H;kH;}�G;��G;��G;��G;˝G;��G;�G; yG;      �G;��G;��G;��G;��G;��G;1H;�H;�(H;�7H;yGH;WH;$fH;�tH;:�H;�H;��H;v�H;��H;v�H;��H;��H;-�H;�H;�H;}�H;]�H;��H;��H;d�H;��H;��H;U�H;��H;O�H;��H;��H;��H;M�H;��H;W�H;��H;��H;e�H;��H;��H;X�H;�H;�H;�H;0�H;��H;��H;v�H;��H;q�H;��H;�H;<�H;�tH;$fH;
WH;|GH;�7H;�(H;�H;3H;��G;��G;��G;��G;��G;      :H;E H;,#H;(H;w.H;�6H;�?H; JH;.UH;�`H;alH;xH;a�H;b�H;֘H;�H;j�H;��H;�H;��H;��H;��H;��H;��H;��H;��H;��H;��H;1�H;��H;��H;O�H;��H;s�H;��H;��H;��H;��H;��H;u�H;��H;I�H;��H;��H;3�H;��H;��H;��H;��H;��H;��H;��H;��H;��H;��H;��H;j�H;��H;֘H;`�H;`�H;xH;blH;�`H;.UH; JH;�?H;6H;�.H; (H;-#H;I H;      cOH;%PH;kRH;�UH;�ZH;�`H;�gH;@oH;�wH;�H;ǈH;��H;3�H;��H;[�H;��H;��H;�H;��H;��H;�H;�H;z�H;n�H;��H;	�H;��H;d�H;��H;��H;I�H;��H;e�H;��H;��H;�H;4�H;�H;��H;��H;g�H;��H;H�H;��H;��H;d�H;��H;�H;��H;k�H;~�H;�H;�H;��H;��H;߾H;��H;��H;Y�H;��H;3�H;��H;ǈH;�H;wH;EoH;�gH;�`H;�ZH;�UH;nRH;"PH;      �sH;-tH;�uH;`xH;�{H;X�H;��H;;�H;s�H;�H;��H;9�H;��H;��H;�H;��H;��H;��H;#�H;��H;a�H;m�H;�H;S�H;\�H;�H;`�H;��H;��H;O�H;��H;k�H;��H;�H;X�H;c�H;[�H;_�H;U�H;�H;��H;h�H;��H;L�H;��H;��H;[�H;�H;a�H;R�H;�H;k�H;^�H;��H;"�H;��H;��H;��H;�H;��H;��H;;�H;��H;�H;t�H;@�H;��H;P�H;�{H;^xH;�uH;.tH;      ��H;�H;F�H;D�H;�H;B�H;4�H;w�H;(�H;��H;��H;�H;۸H;��H;i�H;��H;��H;d�H;��H;��H;��H;��H;��H;��H;@�H;��H;��H;��H;L�H;��H;e�H;��H;�H;Z�H;��H;�H;��H;�H;��H;[�H;�H;��H;d�H;��H;K�H;��H;��H;��H;B�H;��H;��H;��H;��H;��H;��H;f�H;��H;��H;i�H;��H;ڸH;�H;��H;��H;(�H;|�H;:�H;E�H;��H;G�H;O�H;�H;      ��H;ڢH;̣H;D�H;O�H;ЩH;��H;��H;��H;N�H;4�H;�H;��H;��H;$�H;v�H;��H;��H;�H;w�H;��H;w�H;/�H;��H;��H;��H;��H;Z�H;��H;l�H;��H;�H;Q�H;��H;��H;��H;��H;��H;��H;��H;S�H;�H;��H;g�H;��H;Y�H;��H;��H;��H;��H;6�H;w�H;��H;u�H;�H;��H;��H;w�H;%�H;��H;��H;�H;4�H;O�H;��H;��H;��H;ʩH;U�H;B�H;٣H;ڢH;      |�H;°H;x�H;��H;S�H;C�H;��H;;�H;��H;��H;�H;��H;��H;��H;��H;V�H;��H;�H;;�H;&�H;��H;n�H;��H;��H;��H;��H;=�H;��H;p�H;��H;	�H;Z�H;��H;��H;��H;��H;��H;��H;��H;��H;��H;Z�H;	�H;��H;n�H;��H;>�H;��H;��H;��H;��H;p�H;��H;�H;9�H;#�H;��H;V�H;��H;��H;��H;��H;�H;��H;��H;@�H;��H;C�H;[�H;��H;��H;ͰH;      �H;=�H;ѺH;��H;�H;��H;��H;��H;��H;R�H;��H;<�H;��H;�H;t�H;��H;��H;��H;`�H;��H;n�H;��H;��H;��H;��H;2�H;��H;P�H;��H;�H;T�H;��H;��H;��H;��H;��H;��H;��H;��H;��H;��H;��H;Q�H;��H;��H;L�H;��H;3�H;��H;��H;��H;��H;k�H;��H;`�H;��H;��H;��H;t�H;�H;��H;>�H;��H;S�H;��H;��H;��H;��H;�H;��H;ҺH;A�H;      N�H;o�H;�H;��H;��H;E�H; �H;��H;��H;��H;�H;L�H;��H;��H;��H;��H;f�H;%�H;��H;�H;N�H;]�H;Z�H;,�H;��H;��H;"�H;��H;��H;$�H;a�H;��H;��H;��H;��H;��H;��H;��H;��H;��H;��H;��H;_�H;�H;��H;��H;#�H;��H;��H;.�H;a�H;]�H;K�H;�H;��H;)�H;i�H;��H;��H;��H;��H;L�H;�H;��H;��H;��H;�H;I�H;��H;��H;�H;}�H;      +�H;1�H;��H;u�H;r�H;��H;z�H;'�H;�H;�H;5�H;?�H;D�H;[�H;[�H;?�H;��H;��H;��H;b�H;��H;��H;��H;D�H;*�H;��H;�H;��H;��H;=�H;X�H;��H;��H;��H;��H;��H;��H;��H;��H;��H;��H;��H;X�H;8�H;��H;��H;#�H;��H;*�H;F�H;��H;��H;��H;]�H;��H;��H;��H;B�H;[�H;[�H;F�H;>�H;6�H;�H;�H;-�H;��H;��H;t�H;u�H;��H;;�H;      O�H;r�H;�H;��H;��H;K�H;��H;��H;��H;��H;�H;L�H;��H;��H;��H;��H;e�H;%�H;��H;�H;O�H;^�H;Z�H;,�H;��H;��H;"�H;��H;��H;#�H;a�H;��H;��H;��H;��H;��H;��H;��H;��H;��H;��H;��H;_�H;�H;��H;��H;"�H;��H;��H;,�H;a�H;[�H;K�H;�H;��H;)�H;h�H;��H;��H;��H;��H;L�H;�H;��H;��H;��H;�H;I�H;��H;��H;�H;{�H;      ܹH;@�H;ʺH;��H;�H;��H;��H;��H;��H;S�H;��H;<�H;��H;�H;u�H;��H;��H;��H;`�H;��H;p�H;��H;��H;��H;��H;2�H;��H;Q�H;��H;�H;S�H;��H;��H;��H;��H;��H;��H;��H;��H;��H;��H;��H;Q�H;��H;��H;J�H;��H;4�H;��H;��H;��H;��H;j�H;��H;`�H;��H;��H;��H;r�H;�H;��H;?�H;��H;S�H;��H;��H;��H;��H;�H;��H;κH;A�H;      |�H;��H;w�H;��H;S�H;G�H;��H;>�H;��H;��H;�H;��H;��H;��H;��H;V�H;��H;"�H;;�H;#�H;��H;q�H;��H;��H;��H;��H;=�H;��H;r�H;��H;	�H;Z�H;��H;��H;��H;��H;��H;��H;��H;��H;��H;Z�H;�H;��H;l�H;��H;=�H;��H;��H;��H;��H;q�H;��H;!�H;;�H;"�H;��H;X�H;��H;��H;��H;��H; �H;��H;��H;A�H;��H;D�H;Z�H;��H;��H;ðH;      ��H;ݢH;ͣH;B�H;K�H;ҩH;��H;��H;��H;O�H;3�H;�H;��H;��H;'�H;t�H;��H;��H;�H;w�H;��H;w�H;,�H;��H;��H;��H;��H;]�H;��H;l�H;��H;�H;P�H;��H;��H;��H;��H;��H;��H;��H;P�H;�H;��H;g�H;��H;W�H;��H;��H;��H;��H;7�H;v�H;��H;u�H;�H;��H;��H;w�H;%�H;��H;��H;�H;3�H;N�H;��H; �H;��H;ΩH;P�H;I�H;ףH;آH;      ��H;�H;8�H;D�H;�H;P�H;5�H;|�H;&�H;��H;��H;�H;ڸH;��H;i�H;��H;��H;f�H;��H;��H;��H;��H;��H;��H;B�H;��H;��H;��H;P�H;��H;d�H;��H;�H;X�H;��H;��H;��H;��H;��H;Z�H;�H;��H;b�H;��H;K�H;��H;��H;��H;@�H;��H;��H;��H;��H;��H;��H;f�H;��H;��H;i�H;��H;ڸH;�H;��H;��H;+�H;|�H;;�H;F�H;�H;C�H;>�H;�H;      �sH;)tH;�uH;ZxH;�{H;X�H;��H;:�H;s�H;�H;��H;<�H;��H;��H;�H;��H;��H;��H;#�H;��H;c�H;n�H;�H;S�H;b�H;�H;[�H;��H;��H;N�H;��H;i�H;��H;�H;Z�H;b�H;[�H;c�H;W�H;�H;��H;i�H;��H;K�H;��H;��H;]�H;�H;\�H;O�H;�H;n�H;]�H;��H;%�H;��H;��H;��H;�H;��H;��H;<�H;��H;��H;t�H;B�H;��H;V�H;�{H;exH;�uH;*tH;      mOH;)PH;fRH;�UH;�ZH;�`H;�gH;GoH;�wH;�H;ǈH;��H;3�H;��H;[�H;��H;��H;�H;��H;��H;�H;	�H;x�H;l�H;��H;�H;��H;g�H;��H;��H;I�H;��H;d�H;��H;��H;�H;4�H;�H;��H;��H;g�H;��H;H�H;�H;��H;a�H;��H;�H;��H;h�H;��H;�H;�H;��H;��H;�H;��H;��H;[�H;��H;5�H;��H;ɈH;�H;�wH;GoH;�gH;�`H;�ZH;�UH;qRH;#PH;      BH;E H;=#H;�'H;m.H;�6H;�?H; JH;5UH;�`H;`lH;xH;^�H;`�H;טH;�H;g�H;��H;��H;��H;��H;��H;��H;��H;��H;��H;��H;��H;5�H;��H;��H;O�H;��H;s�H;��H;��H;��H;��H;��H;s�H;��H;L�H;��H;��H;.�H;��H;��H;��H;��H;��H;��H;��H;��H;��H;�H;��H;h�H;��H;טH;`�H;a�H;xH;alH;�`H;4UH;%JH;�?H;�6H;|.H;�'H;=#H;B H;      !�G;��G;��G;��G;��G;��G;0H;�H;�(H;�7H;yGH;WH;"fH;�tH;?�H;�H;��H;v�H;��H;u�H;��H;��H;,�H;�H;�H;y�H;Y�H;��H;��H;d�H;��H;��H;U�H;��H;O�H;��H;��H;��H;O�H;��H;W�H;��H;��H;d�H;��H;��H;Y�H;��H;�H;�H;3�H;��H;��H;x�H;��H;s�H;��H;�H;?�H;�tH;$fH;	WH;{GH;�7H;�(H;�H;1H;��G;��G;��G;��G;��G;      PvG;yG;�G;��G;��G;��G;��G;��G;~�G;kH;H;�,H;�@H;�SH;�eH;\vH;��H;��H;�H;�H;p�H;ּH;�H;F�H;j�H;��H;`�H;]�H;��H;��H;^�H;��H;��H;A�H;��H; �H;#�H; �H;��H;A�H;��H;��H;`�H;��H;��H;[�H;`�H;��H;h�H;@�H;&�H;ּH;o�H;�H;�H;|�H;��H;_vH;�eH;�SH;�@H;�,H;H;kH;~�G;��G;��G;��G;ȝG;��G;�G;yG;      @�F;�F;��F;��F;n�F;iG;GGG;�pG;�G;0�G;��G;i�G;�H;*H;�AH;OWH;/kH;}H;�H;A�H;��H;)�H;I�H;%�H;��H;-�H;��H;��H;��H;�H;�H;��H;��H;��H;9�H;��H;��H;��H;7�H;��H;��H;��H;�H;�H;��H;�H;��H;3�H;��H;"�H;N�H;)�H;��H;D�H;�H;}H;2kH;OWH;�AH;*H;�H;i�G;��G;4�G;�G;�pG;IGG;[G;x�F;��F;��F;�F;      �mD;�~D;M�D;��D;a\E;��E;r0F;ƔF;��F;�8G;�vG;�G;;�G;L�G;2H;u0H;6JH;haH;�uH;݇H;��H;8�H;��H;��H;��H;��H;g�H;�H;��H;��H;^�H;A�H;��H;��H;��H;��H;)�H;��H;��H;��H;��H;>�H;a�H;��H;��H;�H;g�H;��H;��H;��H;��H;8�H;��H;��H;�uH;baH;7JH;s0H;4H;M�G;@�G;�G;�vG;�8G;��F;ȔF;p0F;��E;h\E;��D;O�D;�~D;      #`?;��?;��?;߳@;��A;y�B;��C;�D;CiE;�F;&�F;�G;KnG;�G;��G;I H;j!H;?H;iYH;[pH;H�H;w�H;�H;E�H;��H;!�H;@�H;�H;��H;p�H;U�H;��H;��H;��H;��H;9�H;N�H;:�H;��H;��H;��H;��H;W�H;s�H;��H;�H;A�H;(�H;��H;E�H;�H;w�H;F�H;^pH;jYH;?H;l!H;K H;��G;�G;MnG;�G;$�F;�F;>iE;��D;��C;o�B;��A;��@;��?;��?;      /�4;��4;�5;�l7;v_9;O�;;��=;
�?;[�A;ɚC;j�D;{�E;ɨF;])G;��G;�G;��G;EH;�6H;�SH;mH;r�H;��H;
�H;��H;I�H; �H;2�H;��H;}�H;�H;��H;2�H;��H;��H;a�H;��H;_�H;��H;��H;0�H;��H;�H;��H;��H;2�H;#�H;P�H;��H;�H;��H;r�H;mH;�SH;�6H;>H;��G;�G;��G;[)G;ʨF;y�E;j�D;ǚC;V�A;�?;��=;M�;;v_9;�l7;�5;��4;      e; ;b";\%;��(;'j-;82;Ä6;��:;�0>;�A;EYC;.�D;F;�F;�XG;��G;J�G;�H;T1H;�PH;�kH;q�H;z�H;5�H;(�H;ԼH;��H;��H;�H;n�H;��H;u�H;p�H;��H;]�H;��H;^�H;��H;n�H;v�H;��H;r�H;�H;��H;��H;׼H;,�H;4�H;}�H;r�H;�kH;�PH;U1H;�H;F�G;��G;�XG;�F;	F;.�D;DYC;�A;�0>;��:;Ƅ6;02;j-; �(;N%;c"; ;      
��:�B�:ކ�:wx;��
;�;4�;�}$;6|,;a�3;�_9;;>;zA;��C;�E;�F;5G;u�G;W�G;>H;�/H;�PH;mH;H�H;��H;��H;i�H;��H;��H;�H;]�H;��H;��H;��H;j�H;H�H;��H;I�H;j�H;��H;��H;��H;^�H;�H;��H;��H;l�H;��H;��H;I�H;mH;�PH;�/H;?H;W�G;t�G;"5G;�F;�E;��C;zA;:>;�_9;b�3;6|,;�}$;6�;�;��
;rx;���:�B�:      �w[:vBd:�}:��:=�:۳�:�:�;�;W ;�+;��3;١:;�?;��B;�E;FZF;�G;�G;p�G;DH;W1H;�SH;^pH;ۇH;B�H;�H;y�H;��H;��H;��H;��H;s�H;#�H;��H;�H;\�H;�H;��H;�H;p�H;��H;��H;��H;��H;y�H;�H;H�H;هH;dpH;�SH;S1H;?H;p�G;�G;�G;FZF;�E;��B;�?;١:;��3;�+;W ;�;�;�:˳�:E�:��:�}:ZBd:      D�S���D�Ж����� (7��9��R:+��:G��:��:�>;�";�P.;%m7;��=;XB;۰D;y9F;G;�G;X�G;�H;�6H;fYH;�uH;�H;�H;��H; �H;��H;�H;��H;�H;9�H;a�H;��H;��H;��H;^�H;6�H;�H;��H;"�H;��H;��H;��H;�H;�H;�uH;mYH;�6H;�H;T�G;�G; G;w9F;۰D;SB;��=;%m7;�P.;�";�>;��:G��:3��:��R:��9 (7��������D�      E^��/X�rF�.}*����P����D��ˬ�pi:��:J��:7�;��;E�);��4;�<;�A;#�D;v9F;�G;o�G;E�G;>H;?H;^aH;}H;x�H;v�H;��H;�H;��H;b�H;�H;�H;��H;&�H;��H;&�H;��H;�H;�H;`�H;��H;�H;��H;v�H;|�H;}H;ZaH;?H;>H;C�G;m�G;�G;t9F;#�D;�A;�<;��4;D�);��;6�;R��:��:pi: ̬���D��P����4}*�rF��/X�      ��ﻬ��f�ܻE�ƻe󩻸���FL����������H�-:�:���:�;�>&;��3;T9<;�A;۰D;CZF;!5G;��G;��G;i!H;2JH;-kH;��H;��H;j�H;��H;��H;��H;��H;��H;��H;c�H;��H;e�H;��H;��H;��H;��H;��H;��H;g�H;��H;��H;,kH;,JH;j!H;��G;��G;5G;CZF;ڰD;�A;R9<;��3;�>&;�;���:�:H�-:����������FL����k�J�ƻk�ܻ���      j�V��5S��6H���6�D� �R,��?ػ6G���D^������D����9�4�: �:-�;�%;��3;�<;UB;�E;�F;�XG;�G;E H;n0H;NWH;YvH;�H;�H;��H;��H;��H;p�H;T�H;��H;��H;:�H;��H;��H;N�H;m�H;��H;��H;��H;|�H;�H;XvH;HWH;g0H;E H;�G;�XG;��F;�E;SB;�<;��3;�%;*�;�:�4�:���9��D�����D^�6G���?ػR,�F� ���6��6H��5S�      ��.��LȤ���������:�f�t�=����<�ܻ�*��Po5�^��� }(7t�}:�n�:-�;�>&;��4;��=;��B;�E;�F;��G;��G;/H;AH;�eH;?�H;ؘH;[�H;ݷH;f�H;!�H;��H;m�H;��H;Q�H;��H;k�H;��H; �H;c�H;۷H;\�H;ؘH;<�H;�eH;}AH;*H;��G;��G;�F;�E;��B;��=;��4;�>&;'�;�n�:l�}: z(7b���Qo5��*��:�ܻ���u�=�:�f���������KȤ�.��      �c��8���������Ҽ����������r�HE:�E,�Iߵ�}/X���º�Ƭ�t�}:
�:�;E�);$m7;�?;��C;F;[)G;�G;L�G;*H;�SH;�tH;c�H;�H;�H;��H;��H;��H;�H;��H;M�H;��H;�H;��H;��H;��H;�H;��H;c�H;�tH;�SH;�)H;E�G;�G;\)G;F;��C;�?;!m7;D�);�;�:h�}:�Ƭ���º~/X�Jߵ�E,�HE:���r�����������Ҽ�켵����8�      #'K���G��>��0�\y��c����T��� ��V�V�(���ƻ�od�~�º �(7�4�:���:��;�P.;ա:;zA;,�D;̨F;NnG;<�G;�H;�@H;$fH;d�H;0�H;��H;ָH;��H;��H;��H;~�H;9�H;~�H;��H;��H;��H;ԸH;��H;2�H;c�H;!fH;�@H;�H;8�G;MnG;ʨF;*�D;	zA;ء:;�P.;��;���:�4�: (7��º�od��ƻ(��V�V� ��T�����伕c�^y��0��>���G�      ���1Z��ϐ����}��c���D�2/%��8���Ҽ0c��1�f�����ƻ~/X�V������9�:6�;�";��3;B>;AYC;y�E;�G;�G;f�G;�,H;WH;xH;��H;4�H;�H;�H;��H;3�H;E�H;1�H;G�H;0�H;��H;�H;�H;1�H;��H;xH;WH;�,H;`�G;�G;�G;y�E;?YC;8>;��3;�";7�;�:���9X���/X��ƻ���2�f�0c����Ҽ�8�2/%���D��c���}�ϐ��0Z��      �Pν�ʽN8���������ΐ��`�f���;�1�����BȤ�2�f�(��Lߵ�Ro5���D�0�-:B��:�>;�+;�_9;�A;h�D; �F;�vG;��G;H;xGH;`lH;H;��H;��H;/�H;��H;��H;�H;'�H;�H;��H;��H;,�H;��H;��H;ňH;`lH;uGH;H;��G;�vG;!�F;h�D;�A;�_9;�+;�>;>��:4�-:��D�Vo5�Lߵ�)��3�f�BȤ����1����;�a�f�ΐ���������N8���ʽ      ���g9�Z[��s�z�ؽ���t����}���G�����0c��V�V�E,��*����������:��:T ;f�3;�0>;ǚC;�F;�8G;-�G;kH;�7H;�`H;
�H;�H;��H;N�H;��H;I�H;��H;�H;��H;H�H;��H;K�H;��H;�H;�H;�`H;�7H;iH;)�G;�8G;�F;ʚC;�0>;[�3;T ;��:��:�������*��E,�W�V�0c���������G���}�t�����{�ؽ�s�Z[�g9�      ��=�ր:���0��Q"�~������Pν�榽@����G�1����Ҽ ��HE:�<�ܻ�D^�����Pi:C��:�;:|,;��:;L�A;?iE;��F;�G;�G;�(H;5UH;|wH;q�H;#�H;��H;��H;��H;��H;�H;��H;��H;��H;��H;$�H;p�H;�wH;5UH;�(H;��G;�G;��F;CiE;O�A;��:;2|,;�;?��:Xi:�����D^�<�ܻHE:� ����Ҽ1����G�@���榽�Pν����~��Q"���0�ր:�      0Dx�4�s���f�sS�ր:����Z[��7ս�榽��}���;��8�U�����r����:G�����ͬ�'��:
�;�}$;Ä6;�?;��D;ʔF;�pG;��G;�H;"JH;@oH;=�H;y�H; �H;:�H;��H;��H;'�H;��H;��H;9�H;��H;u�H;:�H;GoH;"JH;�H;��G;�pG;ȔF;�D;�?;6;�}$;�;��:@ͬ���;G�������r�U����8���;���}��榽�7սZ[����ր:�sS���f�4�s�      �*���0��ޥ��;����k��H��#%�Z[��Pνt��`�f�2/%���伆���t�=��?ػ�FL���D�d�R:��:4�;42;��=;��C;h0F;IGG;��G;#H;�?H;�gH;��H;-�H;��H;��H;��H;��H;u�H;��H;��H;��H;��H;-�H;��H;�gH;�?H;&H;��G;MGG;h0F;��C;��=;22;-�;��:\�R:��D��FL��?ػt�=��������2/%�`�f�t���PνZ[��#%��H��k�;���ޥ���0��      '�þ��� ����R��|쏾5�s��H�����������ΐ����D��c�����;�f�S,�����P��H�9ͳ�:�;"j-;M�;;u�B;��E;\G;��G;��G;�6H;�`H;[�H;O�H;թH;Q�H;��H;R�H;��H;R�H;��H;O�H;թH;O�H;W�H;�`H;�6H;��G;��G;bG;��E;v�B;M�;;j-;�;ѳ�:8�9�P�����S,�;�f������c���D�ΐ�������������H�5�s�|쏾�R�� ������      @��/�待Yؾ(�þĪ�|쏾�k�ր:�~�{�ؽ�����c�]y���Ҽ����C� �i�.��  (7E�:��
;��(;~_9;��A;j\E;l�F;��G;��G;�.H;�ZH;�{H;�H;I�H;S�H;�H;��H;x�H;��H;�H;P�H;H�H;�H;�{H;�ZH;�.H;��G;ÝG;v�F;g\E;��A;~_9;��(;��
;I�: (7+��j�C� �������Ҽ]y��c�����{�ؽ~�ր:��k�|쏾Ī�(�þ�Yؾ/��      #��N������>I�(�þ�R��;���tS��Q"��s������}��0��켈�����6�F�ƻ:}*������:}x;X%;�l7;ڳ@;��D;��F;��G;��G;�'H;�UH;`xH;N�H;F�H;��H;��H;��H;{�H;��H;��H;��H;F�H;N�H;]xH;�UH;�'H;��G;��G;��F;��D;ܳ@;�l7;V%;zx;��:���8}*�F�ƻ��6��������0���}�����s��Q"�tS�;����R��(�þ>Iᾣ���O��      ���R��8�
������Yؾ���ޥ����f���0�Z[�N8��ϐ���>�����JȤ��6H�a�ܻrF�����}:���:c";-�5;��?;Y�D;��F;�G;��G;2#H;cRH;�uH;H�H;£H;v�H;ĺH;�H;��H;�H;ĺH;v�H;��H;F�H;�uH;iRH;0#H;��G;�G;��F;T�D;��?;(�5;_";��:$�}:̖�rF�b�ܻ�6H�JȤ������>�ϐ��N8��Z[���0���f�ޥ������Yؾ����8�
�R��      �� ����R��N��/������0��4�s�ր:�g9��ʽ1Z����G��8�
.���5S���� 0X�t�D�nBd:�B�: ;��4;ʈ?;�~D;�F;yG;��G;P H;-PH;tH;�H;΢H;ǰH;.�H;q�H;6�H;n�H;.�H;ǰH;̢H;�H;tH;3PH;P H;��G;yG;�F;�~D;Ȉ?;��4; ;�B�:~Bd:|�D��/X���껭5S�
.���8���G�1Z���ʽg9�ր:�4�s��0�����/��N��R�����      GF�Wh����VVھ7�������~���S��#��o��8S��p₽2�6�o���hy��VFB��Eֻ�A?�̾	�mY�:���:g�";h46;\@;b�D;��F;�nG;��G;�H;@H;�fH;B�H;/�H;��H;гH;йH;��H;ʹH;ϳH;��H;,�H;?�H;�fH;@H;�H;��G;�nG;��F;_�D;[@;_46;d�";���:qY�:о	��A?��EֻVFB�hy��o���2�6�p₽8S���o���#��S��~������7��VVھ��Wh��      Vh���b���쾧*־�v��(���*��'�O�U� �s��r���؀�G�3���?ݜ�<�>�S�ѻޡ9�����!o�:>% ;tM#;C�6;LA@;��D;��F;qG;L�G;H;�@H;jgH;��H;��H;ީH;�H;��H;޻H;��H;�H;ީH;��H;��H;cgH;�@H;H;L�G;qG;��F;��D;JA@;<�6;nM#;:% ;#o�:����ޡ9�S�ѻ<�>�>ݜ���G�3��؀��r��s�U� �'�O�*��(����v���*־���b��      ���쾳�޾/5ʾL;���:��(�v��E�_'����q����u���+��W��A����4���Ļ9)�pj��{W�:b�;	%;�k7;$�@;��D;��F;�wG;T�G;5H;@CH;(iH;�H;��H;��H;��H;��H;u�H;��H;��H;��H;��H;�H;$iH;DCH;4H;U�G;�wG;��F;��D; �@;�k7;%;`�;�W�:�j��9)���Ļ��4��A���W缃�+���u�q�����_'��E�(�v��:��L;��/5ʾ��޾��      VVھ�*־/5ʾr��������M���9b��5�����ս����Xc���ʖռ�I��U�$�lT���Z�`\���:��;k�';�8;RA;�9E;��F;ƂG;��G;CH;
GH;lH;C�H;=�H;�H;ĵH;��H;Q�H;��H;ĵH;�H;8�H;B�H;lH;GH;CH;��G;łG;��F;�9E;RA;�8;h�';��;�:�\���Z�lT��V�$��I��ʖռ���Xc������ս���5��9b��M������r���/5ʾ�*־      7���v��M;������RP��E�r�z�H�U� ���5@��ѓ����K�a��վ���s�r���񕻞ܺ�4u9&�:"�;-�+;~�:;�"B;o�E;��F;אG;��G;/H;8LH;�oH;>�H;v�H;��H;7�H;ۼH;��H;ԼH;7�H;��H;r�H;9�H;�oH;<LH;.H;��G;ՐG;��F;n�E;�"B;x�:;,�+; �;&�:�4u9�ܺ��s����s��վ�a���K�ѓ��5@����U� �z�H�E�r�RP������M;���v��      ����(����:���M��E�r�&�O�#,�X�
��gٽpĥ���u�x1�h���)Ϥ���P�	[�.o�pp��@:c��:�P;>�/;9�<;C;�E;n!G;5�G;�G;�%H;�RH;�tH;��H;H�H;ٯH;�H;]�H;�H;V�H;�H;ԯH;D�H;��H;�tH;�RH;�%H;�G;4�G;r!G;�E;C;4�<;;�/;�P;e��:<:pp���.o�
[򻪎P�)Ϥ�h���x1���u�pĥ��gٽX�
�#,�&�O�E�r��M���:��(���      �~��*��(�v��9b�z�H�#,�MZ����7S��x^����N������μ�I���%+����۝.�x����j~:I��:-m;��3;�>;>�C;=PF;�FG;Q�G;��G;y/H;ZH;wzH;H�H;��H;_�H;!�H;,�H;��H;)�H;�H;]�H;��H;D�H;rzH;ZH;y/H;��G;P�G;�FG;;PF;8�C;�>;��3;)m;Q��:�j~:����ڝ.�����%+��I����μ�����N�x^��7S�����MZ�#,�z�H��9b�(�v�*��      �S�'�O��E��5�U� �X�
���罤9��'l���Xc���(��������[�����ݎ�Cܺp;9%��:/�	;Ed';e 8;<�@;�D;�F;jG;��G;NH;p:H;AbH;��H;�H;4�H;D�H;�H;9�H;��H;7�H;��H;D�H;/�H;�H;��H;HbH;q:H;OH;��G;jG;�F;x�D;<�@;e 8;Cd';3�	;!��:`;9Dܺ�ݎ������[��������(��Xc�'l���9�����X�
�U� ��5��E�'�O�      �#�U� �_'������gٽ7S��'l��N�j�C�3��i��վ�y���(���Ļ`A?���B��@:�[�:
Q;�.;��;;{tB;�E;�F;%�G;��G;�H;TFH;%kH;��H; �H;�H;i�H;�H;v�H;��H;r�H;�H;h�H;�H;�H;��H;*kH;VFH;�H;��G;%�G;��F;�E;{tB;��;;�.;Q;�[�:��@:��B�aA?���Ļ(�y����վ��i�C�3�N�j�'l��7S���gٽ����_'�U� �      �o��s��罫�ս4@��pĥ�x^���Xc�D�3���	�Ɍ˼�]��RFB��Z򻭜��kӺ ��8��:ܛ;�M#;u=5;?;K�C;|@F;:G;�G; �G;0'H;�RH;ztH;��H;~�H;.�H;��H;��H;��H;B�H;��H;��H;��H;(�H;x�H;��H;�tH;�RH;2'H;�G;�G;	:G;x@F;L�C;?;t=5;�M#;ܛ;��:`��8mӺ�����Z�RFB��]��Ɍ˼��	�C�3��Xc�x^��pĥ�5@����ս���s�      8S���r��q�����Г����u���N���(��i�ʌ˼�A����P�gs��:|�H����\:1�:r�;xn-;�:;�A;z,E;j�F;)oG;��G;�H;�7H;:_H;~H;�H;�H;w�H;�H;{�H;=�H;��H;=�H;{�H;�H;s�H;��H;�H;~H;@_H;�7H;�H;��G;,oG;h�F;|,E;��A;�:;�n-;r�;/�:�\:H���7|��gs���P��A��ʌ˼�i���(���N���u�ѓ�����r���r��      o₽�؀���u��Xc���K�x1�������վ��]����P����@T����9��o��3�9x&�:a�	;\%;F�5;��>;��C;�F;�!G;��G;��G;DH;`HH;�kH;��H;J�H;��H;��H;w�H;M�H;��H;��H;��H;L�H;z�H;��H;��H;M�H;��H;�kH;bHH;EH;��G;��G;�!G;�F;��C;��>;Q�5;^%;]�	;�&�:�3�9 �o���9�@T�������P��]���վ�����w1���K��Xc���u��؀�      2�6�F�3���+���`�i�����μ���y���QFB�fs�@T��(�D��{���:u9�q�:{��:�Y;�t0;��;;�B;�9E;�F;hG;ٿG;�G;z0H;�XH;'xH; �H;v�H;�H;��H;��H;�H;0�H;4�H;0�H;�H;��H;��H;��H;y�H;*�H;-xH;�XH;|0H;��G;ۿG;�gG;�F;�9E;�B;��;;�t0;zY;���:�q�:�:u9�{��'�D�?T��fs�QFB�y��������μh���b�����+�F�3�      l�����W�˖ռ�վ�+Ϥ��I����[�(��Z����9��{���;9QX�:ZX�::Q;B,;��8;�A@;BD;�@F;�,G;��G;��G;gH;�DH;hH;-�H;T�H;e�H;`�H;%�H;�H;��H;��H;f�H;��H;��H;�H; �H;[�H;j�H;\�H;7�H; hH;�DH;bH;��G;��G;�,G;�@F;BD;�A@;��8;<,;@Q;XX�:WX�:�;9�{����9���Z�(���[��I��)Ϥ��վ�̖ռ�W���      gy��?ݜ��A���I����s���P��%+������Ļ����6|��o�`:u9WX�:�+�:V;�);Ԅ6;u�>;�PC;d�E;��F;�xG;+�G;zH;e1H;XH;wH;��H;�H;�H;~�H;�H;B�H;��H;��H;��H;��H;��H;B�H;�H;z�H;�H;�H;��H;wH;XH;a1H;}H;,�G;�xG;��F;e�E;�PC;z�>;΄6;�);V;�+�:[X�:�:u9�o�2|�������Ļ����%+���P���s��I���A��?ݜ�      PFB�;�>���4�T�$�r��[�����ݎ�dA?�hӺ@����3�9�q�:ZX�:V;��';�=5;�=;�B;GE;K�F;�UG; �G;��G;UH;�HH;jH;��H;u�H;H�H;1�H;J�H;��H;A�H;�H;!�H;��H; �H;�H;@�H;��H;F�H;5�H;N�H;|�H;��H;jH;�HH;WH;��G;!�G;�UG;L�F;GE;�B;y�=;�=5;��';Z;ZX�:�q�:�3�9(���gӺ^A?��ݎ����[�u��U�$���4�8�>�      �EֻP�ѻ��ĻoT���񕻸.o�ԝ.�;ܺ��B� ��8�\:v&�:���:>Q;�);�=5;�:=;,#B;��D;�uF;�6G;ÚG;]�G;tH;�:H;^H;�zH;��H;a�H;ŲH;�H;��H;\�H;�H;m�H;2�H;��H;-�H;j�H;�H;X�H;��H;�H;ȲH;e�H;��H;�zH;^H;�:H;vH;Y�G;ĚG;�6G;�uF;��D;%#B;�:=;�=5;�);@Q;���:~&�:�\: ��8��B�9ܺٝ.��.o���rT����ĻL�ѻ      rA?�ء9�!9)��Z��ܺjp��@����;9�@:��:9�:Y�	;vY;<,;̈́6;v�=;!#B;��D;`XF;�!G;|�G;�G;�H;�.H;ySH;cqH;߉H;��H;c�H;��H;o�H;��H;��H;��H;��H;�H;��H;�H;�H;��H;��H;��H;r�H;ĹH;h�H;��H;މH;^qH;|SH;�.H;�H;�G;}�G;�!G;cXF;��D;"#B;t�=;Є6;<,;xY;Z�	;C�:��:�@:�;9p���fp��ܺ�Z�9)�ԡ9�      p�	�8����j���[���4u9h:�j~:-��:�[�:ߛ;y�;X%;�t0;��8;z�>;�B;��D;hXF;7G;_�G;��G;��G;�%H;KH;�iH;�H;��H;8�H;v�H;
�H;]�H;��H;��H;3�H;��H;��H;S�H;��H;}�H;2�H;��H;��H;`�H;�H;v�H;8�H;��H;�H;�iH;KH;�%H;��G;��G;b�G;8G;cXF;��D;�B;{�>;��8;�t0;\%;z�;ޛ;�[�:1��:�j~:P:�4u9�]���j��8���      aY�:o�:�W�:+�:&�:i��:e��:-�	;
Q;�M#;n-;N�5;��;;�A@;�PC;GE;�uF;�!G;b�G;��G;�G;H H;EH;�cH;8}H;u�H;��H;��H;��H;��H;��H;+�H;T�H;S�H;N�H;|�H;��H;u�H;K�H;S�H;R�H;(�H;��H;��H;��H;��H;��H;q�H;<}H;�cH;	EH;H H;�G;��G;c�G;�!G;�uF;GE;�PC;�A@;��;;O�5;�n-;�M#;Q;6�	;a��:u��:&�:��:oW�:�n�:      ���:,% ;F�;��;�;�P;+m;@d';�.;u=5;�:;��>;�B;BD;d�E;M�F;�6G;��G;��G;�G;tH;�AH;
`H;LyH;~�H;"�H;Q�H;�H;K�H;��H;��H;2�H;��H;B�H;��H;��H;F�H;��H;��H;A�H;��H;-�H;��H;��H;K�H;�H;M�H;�H;�H;IyH;`H;�AH;wH;�G;��G;��G;�6G;M�F;f�E;BD;�B;��>;�:;t=5; �.;=d';0m;�P;!�;��;P�;(% ;      \�";tM#;%;u�';*�+;>�/;��3;a 8;��;;?;�A;��C;�9E;�@F;��F;�UG;ĚG;$�G;��G;I H;�AH;�^H;GwH;�H;��H;�H;��H;.�H;��H;%�H;�H;��H;��H;��H;m�H;L�H;|�H;D�H;j�H;��H;��H;��H;�H;(�H;��H;-�H;��H;ݫH;��H;�H;@wH;�^H;�AH;I H;��G; �G;ǚG;�UG;��F;�@F;�9E;��C;��A;?;��;;k 8;��3;6�/;>�+;j�';%;jM#;      }46;B�6;�k7;*�8;v�:;@�<;+�>;H�@;�tB;U�C;�,E;�F;�F;�,G;�xG;%�G;_�G;�H;�%H;EH;`H;DwH;2�H;5�H;G�H;�H;��H;n�H;��H;��H;(�H;@�H;��H;]�H;��H;p�H;��H;k�H;��H;_�H;��H;<�H;*�H;��H;��H;n�H;��H;�H;K�H;3�H;*�H;EwH;`H;EH;�%H;�H;_�G;%�G;�xG;�,G;�F;�F;�,E;P�C;�tB;F�@;(�>;;�<;��:;(�8;�k7;#�6;      ^@;UA@;�@;RA;�"B;C;?�C;�D;�E;�@F;o�F;�!G;hG;��G;,�G;��G;vH;�.H;KH;�cH;IyH;�H;3�H;éH;�H;|�H;w�H;��H;�H;N�H;��H;J�H;9�H;��H;��H;_�H;��H;Z�H;��H;��H;9�H;I�H;��H;M�H;�H;��H;r�H;�H;	�H;��H;.�H;�H;GyH;�cH;KH;�.H;uH;��G;-�G;��G;hG;�!G;t�F;�@F;�E;��D;?�C;�
C;�"B;RA;�@;NA@;      ��D;��D;��D;�9E;h�E;)�E;FPF;�F;��F;:G;7oG;��G;ݿG;��G;H;]H;�:H;�SH;�iH;B}H;��H;��H;J�H;�H;=�H;��H;.�H;m�H;��H;(�H;��H;	�H;��H;��H;��H;%�H;c�H; �H;��H;��H;��H;�H;��H;+�H;��H;m�H;'�H;��H;?�H;	�H;J�H;��H;��H;<}H;�iH;�SH;�:H;]H;H;��G;޿G;��G;9oG;:G;��F;�F;HPF;!�E;r�E;�9E;��D;��D;      ��F;��F;��F;��F;��F;x!G;�FG;#jG;)�G;��G;��G;��G;�G;oH;e1H;�HH;^H;eqH;�H;p�H; �H;ګH;�H;|�H;��H;�H;�H;[�H;��H;��H;��H;��H;��H;��H;x�H;��H;	�H;��H;w�H;��H;��H;}�H;��H;��H;��H;Z�H;�H;�H;��H;z�H;�H;۫H; �H;n�H;��H;^qH;^H;�HH;e1H;iH;�G;��G;��G;�G;)�G;&jG;�FG;m!G;��F;��F;��F;��F;      �nG;qG;�wG;ǂG;̐G;1�G;_�G;��G;��G;"�G;�H;BH;y0H;�DH;XH;jH;�zH;�H;��H;��H;U�H;��H;��H;x�H;,�H;�H;=�H;��H;\�H;{�H;I�H;��H;��H;��H;6�H;��H;��H;��H;2�H;��H;��H;��H;K�H;z�H;\�H;��H;6�H;�H;-�H;t�H;��H;��H;T�H;��H;��H;܉H;�zH;jH;XH;�DH;y0H;EH;�H;�G;��G;��G;Z�G;0�G;�G;��G;�wG;qG;      ��G;I�G;N�G;��G;��G;��G;��G;LH;�H;7'H;�7H;gHH;�XH;"hH;wH;��H;��H;��H;8�H;��H;�H;*�H;j�H;��H;j�H;X�H;��H;9�H;v�H;@�H;��H;��H;��H;a�H;��H;�H;�H;��H;��H;c�H;��H;��H;��H;@�H;w�H;9�H;��H;[�H;o�H;��H;m�H;+�H;�H;��H;8�H;��H;��H;��H;wH;"hH;�XH;hHH;�7H;7'H;�H;NH;��G;��G;��G;��G;P�G;?�G;      �H;H;1H;OH;H;�%H;}/H;m:H;MFH;�RH;A_H;�kH;-xH;3�H;��H;z�H;g�H;j�H;z�H;¼H;N�H;��H;��H;�H;��H;��H;W�H;v�H;!�H;��H;��H;��H;S�H;��H;C�H;v�H;��H;r�H;C�H;��H;W�H;��H;��H;��H;"�H;v�H;S�H;��H;��H;	�H;��H;��H;K�H;��H;x�H;h�H;g�H;{�H;��H;1�H;*xH;�kH;D_H;�RH;OFH;m:H;}/H;�%H;+H;MH;1H;	H;      @H;�@H;HCH;GH;>LH;�RH;ZH;@bH;)kH;�tH;~H;��H;(�H;]�H;�H;H�H;ʲH;��H;�H;��H;��H;!�H;��H;H�H;*�H;��H;w�H;>�H;��H;��H;��H;g�H;��H;M�H;��H;��H;��H;��H;��H;M�H;��H;c�H;��H;��H;��H;>�H;t�H;��H;+�H;G�H;��H;"�H;��H;��H;�H;��H;ʲH;I�H;�H;[�H;'�H;��H;~H;�tH;(kH;FbH;ZH;�RH;>LH;GH;ICH;�@H;      �fH;{gH;.iH;lH;�oH;�tH;|zH;��H;��H;��H;��H;T�H;~�H;q�H;�H;:�H;�H;v�H;b�H;��H;��H;�H;&�H;��H;��H;��H;K�H;��H;��H;��H;g�H;�H;]�H;��H;��H;�H;'�H;�H;��H;��H;`�H; �H;g�H;��H;��H;��H;H�H;��H;��H;��H;,�H;�H;��H;��H;a�H;u�H;�H;8�H;�H;o�H;��H;U�H;�H;��H;��H;��H;�zH;�tH; pH;lH;/iH;}gH;      A�H;��H;�H;;�H;:�H;�H;L�H;�H;$�H;~�H;�H;��H;
�H;i�H;��H;M�H;��H;��H;��H;/�H;6�H;��H;=�H;H�H;	�H;}�H;��H;��H;��H;h�H;��H;s�H;��H;��H;&�H;@�H;@�H;@�H;$�H;��H;��H;o�H;��H;g�H;��H;��H;��H;�H;�H;B�H;A�H;��H;2�H;+�H;��H;��H;��H;O�H;��H;g�H;	�H;��H;�H;�H;#�H;�H;U�H;�H;E�H;<�H;�H;��H;      2�H;��H;��H;;�H;|�H;D�H;��H;.�H;�H;1�H;{�H;��H;�H;+�H;�H;��H;a�H;��H;��H;X�H;��H;��H;��H;6�H;��H;��H;��H;��H;Y�H;��H;[�H;��H;�H;5�H;T�H;v�H;}�H;v�H;Q�H;6�H;�H;��H;Z�H;��H;W�H;��H;��H;��H;��H;6�H;��H;��H;��H;U�H;��H;��H;b�H;��H;�H;+�H;�H;��H;}�H;2�H;�H;/�H;��H;=�H;��H;5�H;��H;��H;      ��H;ةH;��H;٫H;��H;ͯH;g�H;F�H;n�H;��H;�H;��H;��H;(�H;I�H;H�H;"�H;��H;7�H;W�H;G�H;��H;Y�H;��H;��H;��H;��H;d�H;��H;P�H;��H;��H;2�H;p�H;�H;��H;��H;��H;~�H;q�H;5�H;��H;��H;L�H;��H;`�H;��H;��H;��H;��H;`�H;��H;A�H;Q�H;6�H;��H;'�H;H�H;I�H;'�H;��H;��H;�H;��H;p�H;L�H;j�H;˯H;��H;ګH;��H;�H;      ̳H;#�H;ôH;ƵH;E�H;��H;*�H;~�H;�H;��H;��H;V�H;!�H;��H;��H;�H;q�H;��H;�H;O�H;��H;k�H;��H;��H;��H;p�H;-�H;��H;C�H;��H;��H;'�H;S�H;��H;��H;��H;��H;��H;��H;��H;W�H;'�H;��H;��H;?�H;��H;-�H;q�H;��H;��H;��H;j�H;��H;I�H;~�H;��H;v�H;�H;��H;��H;!�H;X�H;��H;��H;�H;��H;-�H;��H;E�H;ǵH;ŴH;'�H;      ͹H;��H;��H;��H;׼H;O�H;8�H;:�H;v�H;��H;F�H;��H;5�H;��H;��H;!�H;2�H;�H;��H;y�H;��H;G�H;h�H;P�H; �H;��H;��H;�H;y�H;��H;�H;D�H;{�H;��H;��H;��H;��H;��H;��H;��H;~�H;D�H;�H;��H;v�H;��H;��H;��H;!�H;Q�H;o�H;G�H;��H;u�H;��H; �H;6�H;#�H;��H;��H;5�H;��H;I�H;��H;y�H;?�H;<�H;R�H;ؼH;��H;��H;�H;      ȻH;ۻH;��H;N�H;�H;�H;��H;��H;��H;H�H;��H;��H;B�H;s�H;��H;��H;��H;��H;V�H;��H;O�H;��H;��H;��H;d�H;�H;��H;�H;��H;��H;$�H;D�H;~�H;��H;��H;��H;��H;��H;��H;��H;��H;C�H;$�H;��H;��H;�H;��H;�H;d�H;��H;��H;��H;J�H;��H;W�H;��H;��H;��H;��H;s�H;A�H;��H;��H;J�H;�H;��H;��H;�H;��H;M�H;��H;�H;      ιH;��H;��H;��H;׼H;U�H;7�H;:�H;v�H;��H;D�H;��H;6�H;��H;��H;!�H;0�H;�H;��H;y�H;��H;H�H;h�H;P�H;!�H;��H;��H;�H;z�H;��H;�H;F�H;}�H;��H;��H;��H;��H;��H;��H;��H;~�H;D�H;�H;��H;v�H;��H;��H;��H;!�H;Q�H;o�H;E�H;��H;u�H;��H;!�H;4�H;$�H;��H;��H;5�H;��H;I�H;��H;y�H;@�H;:�H;R�H;ۼH;��H;��H;�H;      ĳH;&�H;��H;��H;E�H;��H;,�H;��H;�H;��H;��H;V�H;"�H;��H;��H;�H;q�H;��H;�H;O�H;��H;k�H;��H;��H;��H;n�H;/�H;��H;E�H;��H;��H;'�H;T�H;��H;��H;��H;��H;��H;��H;��H;W�H;&�H;��H;��H;?�H;��H;-�H;q�H;��H;��H;��H;k�H;��H;I�H;~�H;��H;v�H;�H;��H;��H;!�H;Z�H;��H;��H;�H;��H;2�H;��H;I�H;��H;´H;)�H;      ��H;٩H;��H;ݫH;��H;ЯH;d�H;J�H;o�H;��H;�H;�H;��H;(�H;J�H;G�H;"�H;��H;6�H;U�H;E�H;��H;X�H;��H;��H;��H;��H;d�H;��H;Q�H;��H;��H;2�H;p�H;�H;��H;��H;��H;~�H;p�H;5�H;��H;��H;L�H;��H;`�H;��H;��H;��H;��H;`�H;��H;@�H;S�H;6�H;��H;%�H;I�H;J�H;'�H;��H;��H;�H;��H;p�H;N�H;k�H;ϯH;��H;ګH;��H;۩H;      2�H;��H;��H;6�H;v�H;F�H;��H;1�H;�H;1�H;{�H;��H;�H;+�H;�H;��H;_�H;��H;��H;X�H;��H;��H;��H;6�H;��H;��H;��H;��H;\�H;��H;[�H;��H;�H;5�H;S�H;x�H;}�H;v�H;S�H;5�H;�H;��H;Z�H;��H;S�H;��H;��H;��H;��H;3�H;��H;��H;��H;V�H;��H;��H;b�H;��H;�H;+�H;�H;��H;{�H;1�H;�H;4�H;��H;C�H;|�H;=�H;��H;��H;      3�H;��H;��H;:�H;6�H;��H;P�H;�H;#�H;~�H;�H;��H;�H;g�H;��H;M�H;��H;��H;��H;.�H;8�H;��H;=�H;E�H;�H;�H;��H;��H;��H;g�H;��H;p�H;��H;��H;'�H;?�H;@�H;?�H;#�H;��H;��H;o�H;��H;e�H;��H;��H;��H;��H;	�H;?�H;D�H;��H;/�H;,�H;��H;��H;��H;N�H;��H;g�H;
�H;��H;�H;�H;'�H;
�H;S�H;�H;7�H;:�H;�H;��H;      �fH;ygH;1iH;lH;�oH;�tH;|zH;��H;��H;��H;��H;U�H;~�H;o�H;	�H;8�H;�H;u�H;a�H;��H;��H; �H;&�H;��H;��H;��H;G�H;��H;��H;��H;g�H;�H;^�H;��H;��H;�H;&�H;�H;��H;��H;`�H;�H;e�H;��H;��H;��H;E�H;��H;��H;��H;-�H; �H;��H;��H;b�H;t�H;�H;8�H;�H;q�H;��H;W�H;��H;��H;��H;��H;�zH;�tH;pH;lH;6iH;{gH;      @H;�@H;BCH;GH;5LH;�RH;ZH;HbH;*kH;�tH;~H;��H;(�H;Y�H;�H;H�H;ȲH;��H;�H;��H;��H;#�H;��H;G�H;-�H;��H;w�H;@�H;��H;��H;��H;g�H;��H;O�H;��H;��H;��H;��H;��H;M�H;��H;e�H;��H;��H;��H;;�H;t�H;��H;(�H;C�H;��H;"�H;��H;��H;�H;��H;ʲH;K�H;�H;\�H;*�H;��H;~H;�tH;)kH;HbH;	ZH;�RH;>LH;GH;OCH;�@H;       H;H;BH;KH;H;�%H;{/H;m:H;UFH;�RH;A_H;�kH;-xH;4�H;��H;{�H;d�H;j�H;v�H;��H;N�H;��H;��H;�H;��H;��H;U�H;w�H;#�H;��H;��H;��H;U�H;��H;C�H;s�H;��H;s�H;C�H;��H;V�H;��H;��H;��H;�H;q�H;U�H;��H;��H;�H;��H;��H;K�H;��H;z�H;f�H;d�H;|�H;��H;3�H;,xH;�kH;B_H;�RH;TFH;q:H;/H;�%H;'H;HH;BH;H;      ��G;<�G;B�G;��G;��G;
�G;��G;RH;�H;7'H;�7H;gHH;�XH; hH;wH;��H;��H;��H;5�H;��H;�H;-�H;g�H;��H;o�H;T�H;��H;9�H;z�H;>�H;��H;��H;��H;a�H;��H;��H;�H;��H;��H;c�H;��H;��H;��H;=�H;t�H;4�H;��H;[�H;j�H;��H;o�H;+�H;�H;��H;8�H;��H;��H;��H;wH;"hH;�XH;gHH;�7H;6'H;�H;NH;��G;��G;��G;��G;P�G;<�G;      �nG;$qG;�wG;΂G;ېG;9�G;\�G;��G;��G;�G;�H;EH;v0H;�DH;XH;jH;�zH;�H;��H;��H;U�H;��H;��H;{�H;,�H;�H;9�H;��H;^�H;x�H;H�H;��H;��H;��H;4�H;��H;��H;��H;2�H;��H;��H;��H;K�H;x�H;Y�H;��H;9�H; �H;-�H;u�H;��H;��H;T�H;��H;��H;��H;�zH;jH;XH;�DH;w0H;GH;�H; �G;��G;��G;^�G;5�G;ߐG;ʂG;�wG;qG;      �F;��F;��F;��F;��F;|!G;~FG;$jG;*�G;�G;��G;��G;�G;iH;f1H;�HH;^H;eqH;��H;n�H;"�H;ګH;�H;|�H;��H;�H;�H;Z�H;��H;��H;��H;��H;��H;��H;x�H;��H;
�H;��H;u�H;��H;��H;��H;��H;��H;��H;X�H;�H;�H;��H;{�H;�H;۫H; �H;q�H;�H;bqH;^H;�HH;j1H;kH;�G;��G;��G;��G;%�G;"jG;�FG;m!G;��F;��F;��F;��F;      ��D;��D;��D;�9E;g�E;)�E;HPF;�F;��F;:G;6oG;��G;ۿG;��G;�H;]H;�:H;�SH;�iH;?}H;��H;��H;G�H;�H;?�H;��H;)�H;m�H;��H;'�H;��H;�H;��H;��H;��H;"�H;c�H;!�H;��H;��H;��H;�H;��H;*�H;��H;j�H;,�H;��H;=�H;�H;M�H;��H;��H;C}H;�iH;�SH;�:H;^H;�H;��G;�G;��G;6oG;:G;��F;�F;FPF;!�E;o�E;�9E;��D;��D;      <@;@A@;�@;RA;�"B;C;?�C;�D; �E;|@F;q�F;�!G;�gG;��G;-�G;��G;vH;�.H;KH;�cH;JyH;�H;.�H;éH;�H;x�H;u�H;��H;�H;K�H;��H;M�H;:�H;��H;��H;[�H;��H;\�H;��H;��H;<�H;J�H;��H;N�H;�H;��H;u�H;�H;�H;éH;3�H;�H;JyH;�cH;KH;�.H;vH;��G;-�G;��G;�gG;�!G;q�F;~@F;�E;{�D;?�C; C;�"B;4RA;�@;(A@;      o46;>�6;�k7;1�8;r�:;:�<;#�>;F�@;�tB;P�C;�,E;�F;�F;�,G;�xG;(�G;`�G;�H;�%H;EH;
`H;GwH;-�H;4�H;J�H;�H;��H;m�H;��H;��H;)�H;A�H;��H;]�H;��H;p�H;��H;n�H;��H;\�H;��H;A�H;,�H;��H;��H;k�H;��H;�H;H�H;5�H;/�H;EwH;`H;EH;�%H;�H;b�G;'�G;�xG;�,G;�F;�F;�,E;R�C;�tB;J�@;$�>;;�<;r�:;-�8;�k7;'�6;      `�";xM#;%;m�';*�+;A�/;��3;e 8;��;;?;��A;��C;�9E;�@F;��F;�UG;ĚG;$�G;��G;J H;�AH;�^H;BwH;�H;��H;֫H;��H;-�H;��H;#�H;�H;��H;��H;��H;j�H;G�H;|�H;H�H;i�H;��H;��H;��H;#�H;(�H;��H;+�H;��H;ޫH;��H;�H;EwH;�^H;�AH;L H;��G; �G;ŚG;�UG;��F;�@F;�9E;��C;��A;?;��;;h 8;��3;-�/;A�+;_�';%;jM#;      ���:E% ;X�;��;�;Q;-m;@d';�.;r=5;�:;��>;�B;BD;i�E;P�F;�6G;��G;��G;�G;wH;�AH;`H;JyH;�H;�H;M�H;�H;K�H;��H;��H;2�H;��H;E�H;��H;��H;G�H;��H;��H;@�H;��H;/�H;��H;��H;I�H;�H;Q�H; �H;�H;MyH;`H;�AH;wH;�G;��G;��G;�6G;P�F;k�E;BD;�B;��>;�:;u=5;�.;Dd';2m;�P;"�;��;f�;1% ;      �Y�:%o�:{W�:+�:&�:u��:g��:7�	;Q;�M#;�n-;N�5;��;;�A@;�PC;!GE;�uF;�!G;c�G;��G;�G;I H;EH;�cH;<}H;p�H;��H;��H;üH;��H;��H;,�H;U�H;U�H;N�H;w�H;��H;w�H;K�H;P�H;R�H;)�H;��H;��H;¼H;��H;��H;u�H;9}H;�cH;EH;I H;�G;��G;c�G;�!G;�uF;!GE;�PC;�A@;��;;N�5;�n-;�M#;Q;0�	;a��:c��:&�:�:W�:o�:      p�	�(����j���[���4u9d:�j~:+��:�[�:ޛ;y�;[%;�t0;��8;}�>;�B;��D;eXF;7G;a�G;��G;��G;�%H;KH;�iH;��H;��H;7�H;w�H;�H;^�H;��H;��H;3�H;�H;��H;S�H;��H;~�H;2�H;��H;��H;`�H;�H;v�H;7�H;��H;�H;�iH;	KH;�%H;��G;��G;c�G;8G;dXF;��D;�B;}�>;��8;�t0;Y%;y�;ޛ;�[�:3��:�j~:`:�4u9 \���j�� ���      �A?�С9�&9)��Z��ܺ\p��P��� <9�@:��:;�:Z�	;xY;<,;ф6;y�=;"#B;��D;aXF;�!G;�G; �G;�H;�.H;|SH;_qH;܉H;��H;h�H;��H;r�H;��H;��H;��H;��H;�H;��H;�H;�H;��H;��H;��H;t�H;��H;f�H;��H;߉H;_qH;xSH;�.H;�H;�G;|�G;�!G;cXF;��D;!#B;u�=;ф6;<,;uY;Y�	;A�:��:�@:�;9P���fp���ܺ�Z�.9)�Ρ9�      �EֻP�ѻ��ĻlT���񕻶.o�؝.�;ܺ��B����8�\:~&�:���:>Q;�);�=5;�:=;(#B;��D;�uF;�6G;ĚG;_�G;tH;�:H;^H;�zH;��H;g�H;ĲH;	�H;��H;\�H;�H;m�H;0�H;��H;0�H;j�H;�H;X�H;��H;�H;ǲH;d�H;��H;�zH;^H;�:H;vH;`�G;ÚG;�6G;�uF;��D;%#B;�:=;�=5;�);>Q;���:z&�:�\:���8��B�9ܺڝ.��.o���pT����ĻL�ѻ      PFB�;�>���4�S�$�s��[�����ݎ�cA?�jӺ(����3�9�q�:ZX�:\;��';�=5;|�=;�B;GE;P�F;�UG;$�G;��G;ZH;�HH;jH;��H;|�H;H�H;4�H;H�H;��H;D�H;�H;�H;��H; �H;�H;>�H;��H;F�H;4�H;K�H;z�H;��H;jH;�HH;UH;��G;%�G;�UG;H�F;GE;�B;x�=;�=5;��';X;ZX�:�q�:�3�9(���jӺcA?��ݎ����[�u��T�$���4�:�>�      gy��?ݜ��A���I����s���P��%+������Ļ����4|��o��:u9[X�:�+�:\;�);Є6;x�>;�PC;h�E;��F;�xG;+�G;~H;f1H;XH;wH;��H;�H;�H;~�H;�H;C�H;��H;��H;��H;��H;��H;C�H;�H;z�H;�H;�H;��H; wH;XH;b1H;zH;-�G;�xG;��F;a�E;�PC;u�>;̈́6;�);T;�+�:WX�:`:u9�o�6|�������Ļ����%+���P���s��I���A��?ݜ�      l�����W�˖ռ�վ�)Ϥ��I����[�(��Z����9��{���;9]X�:dX�:>Q;<,;��8;�A@;BD;�@F;�,G;��G;��G;hH;�DH;hH;4�H;V�H;j�H;`�H;"�H;�H;��H;��H;f�H;��H;��H;�H;!�H;[�H;g�H;Y�H;3�H;hH;�DH;dH;��G;��G;�,G;�@F;BD;�A@;��8;<,;>Q;VX�:WX�:�;9�{����9���Z�(���[��I��)Ϥ��վ�˖ռ�W���      2�6�F�3���+���`�i�����μ���y���QFB�fs�?T��&�D��{���:u9�q�:��:zY;�t0;��;;�B;�9E;�F;hG;ݿG;�G;y0H;�XH;.xH;$�H;y�H;�H;��H;��H;�H;0�H;4�H;0�H;�H;��H;��H;��H;w�H;'�H;-xH;�XH;y0H;��G;׿G;hG;�F;�9E;�B;��;;�t0;xY;}��:�q�:�:u9�{��*�D�@T��fs�RFB�y��������μh���b�����+�F�3�      o₽�؀���u��Xc���K�w1�������վ��]����P����?T����9���o��3�9z&�:Z�	;\%;K�5;��>;��C;�F;�!G;��G;��G;DH;`HH;�kH;��H;N�H;��H;��H;z�H;M�H;��H;��H;��H;J�H;x�H;��H;��H;L�H;��H;�kH;^HH;BH;��G;��G;�!G;�F;��C;��>;N�5;[%;Z�	;z&�:�3�9 �o���9�@T�������P��]���վ�����w1���K��Xc���u��؀�      8S���r��r�����Г����u���N���(��i�ʌ˼�A����P�fs��6|�8����\:+�:p�;~n-;�:;��A;�,E;k�F;-oG;��G;�H;�7H;>_H;~H;�H;�H;v�H;�H;{�H;=�H;��H;?�H;z�H;�H;t�H;�H;�H;~H;@_H;�7H;�H;��G;)oG;m�F;�,E;��A;ޞ:;~n-;o�;+�:�\:H���8|��gs���P��A��ʌ˼�i���(���N���u�ѓ�����r���r��      �o��s��罫�ս4@��pĥ�x^���Xc�C�3���	�Ɍ˼�]��RFB��Z򻬜��gӺ���8��:ܛ;�M#;x=5;?;O�C;~@F;	:G;�G;�G;0'H;�RH;|tH;��H;{�H;-�H;��H;��H;��H;B�H;��H;��H;��H;+�H;z�H;��H;}tH;�RH;0'H;�G;�G;:G;~@F;R�C;?;p=5;�M#;ٛ;��:`��8mӺ�����Z�RFB��]��Ɍ˼��	�C�3��Xc�x^��pĥ�5@����ս���s�      �#�U� �_'������gٽ7S��'l��N�j�C�3��i��վ�y���(���Ļ\A?���B���@:�[�:Q;
�.;��;;tB;�E;��F;&�G;��G;�H;VFH;&kH;��H;�H;�H;k�H;�H;s�H;��H;r�H;�H;i�H;�H;�H;��H;(kH;UFH;�H;��G;(�G;��F;�E;tB;��;;�.;Q;�[�:��@:��B�aA?���Ļ(�z����վ��i�C�3�N�j�'l��7S���gٽ����_'�U� �      �S�&�O��E��5�U� �X�
���罤9��'l���Xc���(��������[�����ݎ�Bܺ ;9)��:0�	;Hd';h 8;@�@;��D;�F;jG;��G;LH;q:H;AbH;��H;�H;4�H;F�H;~�H;9�H;��H;7�H;�H;F�H;1�H;�H;��H;HbH;q:H;NH;��G;jG;�F;�D;@�@;e 8;Cd';4�	;��:`;9@ܺ�ݎ������[��������(��Xc�'l���9�����X�
�U� ��5��E�&�O�      �~��*��(�v��9b�z�H�#,�LZ����7S��x^����N������μ�I���%+����ٝ.������j~:M��:/m;��3;�>;>�C;=PF;�FG;P�G;��G;y/H;ZH;wzH;G�H;��H;`�H;�H;,�H;��H;)�H;!�H;`�H;��H;E�H;tzH;ZH;{/H;��G;S�G;�FG;=PF;?�C;�>;��3;)m;W��:�j~:����؝.�����%+��I����μ�����N�x^��7S�����MZ�#,�z�H��9b�(�v�*��      ����(����:���M��E�r�&�O�#,�X�
��gٽpĥ���u�x1�h���)Ϥ���P�	[�.o�vp��D:g��:�P;=�/;:�<;C;�E;n!G;4�G;�G;�%H;�RH;�tH;��H;F�H;ׯH;�H;[�H;�H;[�H;�H;ׯH;D�H;��H;�tH;�RH;�%H;�G;5�G;u!G;�E;C;9�<;:�/;�P;i��:8:tp���.o�
[򻪎P�)Ϥ�h���x1���u�pĥ��gٽX�
�#,�&�O�E�r��M���:��(���      8���v��M;������RP��E�r�z�H�T� ���5@��Г����K�a��վ���s�r���񕻥ܺ�4u9&�:$�;/�+;|�:;�"B;o�E;��F;ԐG;��G;/H;5LH;�oH;:�H;r�H;��H;2�H;ڼH;��H;ּH;4�H;��H;r�H;9�H;�oH;<LH;/H;��G;ڐG;��F;n�E;�"B;|�:;-�+;�;&�:�4u9�ܺ��r����s��վ�a���K�ѓ��5@����U� �z�H�E�r�RP������M;���v��      VVھ�*־/5ʾr��������M���9b��5�����ս����Xc���˖ռ�I��U�$�lT���Z�`\���:�;j�';�8;RA;�9E;��F;ÂG;��G;AH;GH;lH;C�H;9�H;�H;ĵH;��H;Q�H;��H;õH;�H;9�H;C�H;lH;GH;CH;��G;ƂG;��F;�9E;RA;�8;h�';��;�:�\���Z�lT��U�$��I��ʖռ���Xc������ս���5��9b��M������r���/5ʾ�*־      ���쾳�޾/5ʾL;���:��(�v��E�_'����q����u���+��W��A����4���Ļ9)�pj��W�:d�;%;�k7;$�@;��D;��F;�wG;T�G;4H;>CH;*iH;�H;��H;��H;��H;��H;u�H;��H;��H;��H;��H;�H;&iH;DCH;5H;U�G;�wG;��F;��D;$�@;�k7;%;`�;�W�:xj��9)���Ļ��4��A���W缃�+���u�q�����_'��E�(�v��:��L;��/5ʾ��޾��      Vh���b���쾧*־�v��(���*��'�O�U� �s��r���؀�G�3���?ݜ�<�>�S�ѻߡ9�����%o�:?% ;tM#;C�6;LA@;��D;��F;qG;L�G;H;�@H;hgH;��H;��H;ީH;�H;��H;�H;��H;�H;ߩH;��H;��H;cgH;�@H;H;L�G;qG;��F;��D;LA@;<�6;nM#;;% ;'o�:����ޡ9�T�ѻ<�>�>ݜ���G�3��؀��r��s�U� �'�O�*��(����v���*־���b��      ���^�T_ݾ��ɾj*��쫖�{x�&G�P,�����b��]@{���/�����䙼�J;�M�ͻ��4�W���:6;��#;�6;[@;3�D;��F;�lG;��G;7H;�:H;�bH;߀H;,�H;/�H;ٱH;��H;ܹH;�H;رH;/�H;*�H;ۀH;�bH;�:H;6H;��G;�lG;��F;3�D;[@;�6;��#;2;��:W���4�M�ͻ�J;��䙼����/�]@{��b�����P,�&G�{x�쫖�i*����ɾT_ݾ^�      ^�3���:پ{�žg�����9t�p�C�������㪫�W`w�F-����*`����7�5Sɻ�K/��xƹ���:�/;�f$;�7;�~@;K�D;\�F;�nG;��G;"H;�;H;jcH;p�H;��H;q�H;�H;.�H;"�H;*�H;	�H;o�H;��H;m�H;dcH;�;H;#H;��G;�nG;f�F;K�D;�~@;�7;�f$;�/;���:�xƹ�K/�5Sɻ��7�)`�����F-�W`w�㪫�������p�C�9t���g���{�ž�:پ3��      U_ݾ�:پ�V;+���Ƥ�La����g��$:��Z�oݽ�ƣ�zl�e.%��߼g���9.�ʴ��LV�`1p��@�:x;N(&;4�7;:�@;�
E;��F;kuG;$�G;OH;�=H;MeH;ĂH;u�H;M�H;��H;��H;��H;��H;��H;M�H;r�H;ÂH;GeH;�=H;OH;&�G;kuG;��F;�
E;6�@;.�7;L(&;x;�@�:�1p�MV�ʴ���9.�g���߼e.%�zl��ƣ�oݽ�Z��$:���g�La���Ƥ�+���V;�:پ      ��ɾ{�ž+��qת�쫖�!�����T��J+�:��2̽�s���yZ����Mμfy����\Ϩ�N,� �6��:��
;_�(;WN9;�A;NE;3�F;�G;��G;|H;�AH;1hH;�H;A�H;թH;ͳH;��H;x�H;��H;ϳH;ԩH;=�H;�H;-hH;�AH;|H;��G;�G;9�F;~NE;��A;ON9;\�(;��
;��: �6N,�\Ϩ���fy��Mμ����yZ��s���2̽:��J+���T�!���쫖�qת�+��|�ž      j*��g����Ƥ�쫖��/��>�c��G=�����zｐж��ɇ�Q�C�
��""��q;k��&��-��l�˺8Y�9v��:9;�h,;�	;;�PB;e�E;� G;ߌG;��G;hH;GH;OlH; �H;��H;��H;;�H;�H;ּH;�H;<�H;��H;��H;��H;JlH;GH;hH;��G;ߌG;� G;d�E;�PB;�	;;�h,;9;~��: Y�9o�˺�-���&�p;k�""��
��Q�C��ɇ��ж��z�����G=�>�c��/��쫖��Ƥ�g���      쫖���La��!���>�c�p�C�z#���RvϽ����zl�dg*����
���I���軽\c�퀺�t,:���:��;�_0;h�<;�1C;��E;w#G;V�G;�G; H;�MH;6qH;��H;}�H;ޭH;-�H;��H;_�H;��H;,�H;ۭH;{�H;��H;5qH;�MH; H;�G;S�G;|#G;��E;�1C;c�<;�_0;�;���:�t,:	퀺�\c�����I��
�����dg*�zl�����RvϽ��z#�p�C�>�c�!���La����      {x�9t���g���T��G=�z#�6�oݽ�b������AG����ލǼgy��I�$�d����$��uƹQ��:�&�:�� ;O4;w�>;PD;�[F;�FG;��G;�G;�)H;_UH;�vH;��H;�H;��H;m�H;��H;,�H;��H;l�H;��H;�H;��H;�vH;fUH;�)H;�G;~�G;�FG;�[F;ND;q�>;M4;�� ;�&�:O��:�uƹ�$�e���I�$�gy��ލǼ���AG������b��nݽ6�z#��G=���T���g�9t�      %G�p�C��$:��J+������oݽ]���.I���yZ��"����ҫ��bT��� �M����˺�m9=ٶ:g�;`(;�8;g�@;��D;�F;AhG;��G;�H;/5H;�]H;e}H;�H;��H;V�H;ɻH;��H;7�H;��H;̻H;V�H;��H;�H;c}H;�]H;15H;�H;��G;DhG;�F;��D;d�@;�8;	`(;l�;;ٶ:�m9��˺M���� �bT�ҫ������"��yZ�-I��]���oݽ������J+��$:�p�C�      P,�����Z�:��z�RvϽ�b��-I��f]a�F-�g� � "��v�{�D�!�������4��P(�oQ:�L�:��;֊/;�'<;ݟB;��E;��F;��G;��G;4H;<AH;gH;M�H;6�H;ҪH;��H;��H;��H;T�H;��H;��H;��H;̪H;3�H;O�H;gH;@AH;6H;��G;��G;��F;��E;ݟB;�'<;֊/;�;�L�:�nQ:�P(���4�����D�!�v�{� "��h� �F-�f]a�-I���b��RvϽ�z�:��Z����      ������oݽ�2̽�ж����������yZ�F-�շ�-aļXO���J;����x�|���º�N@9ǂ�:>�;�f$;��5;�N?;:D;�LF;�:G;��G;��G;�!H;�MH;�pH;��H;ӟH;2�H;�H;B�H;v�H;��H;t�H;B�H;�H;-�H;͟H;��H;�pH;�MH;�!H;��G;��G;�:G;�LF;;D;�N?;��5;�f$;?�;ł�:�N@9��ºv�|���軾J;�XO��-aļշ�F-��yZ����������ж��2̽oݽ���      �b��㪫��ƣ��s���ɇ�zl�BG��"�h� �-aļa���I��C��ۙ�@�uƹV�k:���:�;>>.;
;;��A;�AE;^�F;mG;��G;��G;U2H;�ZH;�zH;֒H;��H;��H;[�H;-�H; �H;�H;�H;.�H;[�H;��H;��H;ؒH;�zH;�ZH;X2H;��G;��G;mG;\�F;�AE;��A;
;;J>.;�;���:f�k:uƹ>��ۙ��C��I�a��-aļh� ��"�BG�zl��ɇ��s���ƣ�㪫�      \@{�W`w�zl��yZ�Q�C�dg*�������!"��XO���I�=|�7Ϩ�jK/�p$T�<Q:X��:��;�(&;�#6;�%?;��C;r#F;�#G;�G;��G;�H;)CH;�gH;}�H;X�H;n�H;�H;��H;�H;��H;��H;��H;�H;��H;�H;g�H;[�H;��H;�gH;*CH;�H;��G;"�G;�#G;w#F;��C;�%?;�#6;�(&;��;d��:@Q:l$T�gK/�7Ϩ�<|��I�XO�� "����鼮��cg*�R�C��yZ�zl�V`w�      ��/�E-�e.%����	�����ލǼҫ��v�{��J;��C�8Ϩ�FO:�����X[�9���:r;��;;.1;�'<;�5B;�NE;�F;1fG;�G;.�G;�*H;�SH;�tH; �H;��H; �H;O�H;z�H;��H;�H;�H;�H;��H;y�H;J�H;�H;��H;(�H;�tH;�SH;�*H;*�G;�G;1fG;�F;�NE;�5B;(<;A.1;�;v;���:h[�9����DO:�6Ϩ��C��J;�t�{�ѫ��ލǼ��������e.%�E-�      ������߼Nμ "���
��gy��aT�D�!���軺ۙ�mK/������m9�A�:���:0�;D�,;�N9;@@;�^D;�LF;T.G;�G;��G;�H;�?H;dH;�H;n�H;�H;��H;��H;��H;��H;��H;y�H;��H;��H;��H;��H;��H;	�H;v�H;�H;dH;�?H;�H;��G;�G;Z.G;�LF;�^D;F@;�N9;@�,;6�;���:�A�: m9����hK/��ۙ����C�!�`T�gy���
��""��Oμ�߼���      �䙼*`��h��fy��n;k��I�I�$��� �����u�|�<��$T�H[�9�A�:j��:"�;�);+7;��>;�tC;�E;��F;�uG;�G;��G;�+H;�SH;�sH;��H;a�H;�H;̻H;��H;7�H;q�H;��H;��H;��H;n�H;7�H;��H;ȻH;�H;g�H;��H;�sH;�SH;�+H;��G;�G;�uG;��F;�E;�tC;��>;$7;�);"�;h��:�A�:X[�9t$T�:�u�|������� �I�$��I�r;k�fy��h��*`��      �J;���7��9.����&����^���M����4���ºuƹ0Q:���:���:"�;��(;��5;��=;��B;�[E;C�F;�TG;��G;��G;�H;�CH;fH;ɁH;u�H;��H;��H;��H;��H;U�H;��H;>�H;�H;<�H;��H;T�H;��H;��H;��H;��H;y�H;ˁH;fH;�CH;�H;��G;��G;�TG;G�F;�[E;��B;��=;��5;��(;$�;���:���:@Q:�tƹ��º��4�M��`�����軪&����9.���7�      G�ͻ2Sɻδ��^Ϩ��-���\c��$���˺�P(� O@9n�k:X��:t;5�;�);��5;L�=;*QB;kE;�F;%8G;C�G;C�G;�	H;U5H;�YH;AwH;؎H;��H;ӰH;��H;��H;T�H;!�H;��H;u�H;�H;q�H;~�H;#�H;P�H;��H;��H;ְH;��H;َH;BwH;�YH;[5H;�	H;C�G;E�G;'8G;�F;lE;!QB;L�=;��5;�);5�;t;^��:v�k:�N@9�P(���˺�$��\c��-��bϨ�Դ��-Sɻ      ��4��K/�PV�B,�P�˺퀺xuƹ�m9oQ:т�:���:��;|�;A�,;$7;��=;QB;��D;�cF;$G;̇G;��G;��G;x)H;�NH;�mH;܆H;ŚH;%�H;�H;�H;��H;��H;��H;��H;w�H;�H;u�H;��H;��H;��H;��H;�H;�H;(�H;ŚH;܆H;�mH;�NH;v)H;��G;��G;͇G;$G;�cF;��D; QB;��=;$7;>�,;|�;��;���:͂�:oQ:m9�uƹ�쀺N�˺J,�HV��K/�      HV�0yƹ�1p� (�6(Y�9�t,:e��:Eٶ:�L�:A�;�;�(&;?.1;�N9;��>;��B;lE;�cF;�G;*�G;��G;��G;V H;�EH;�eH;�H;��H;ҥH;��H;��H;�H;��H;��H;R�H;��H;J�H;��H;G�H;��H;Q�H;��H;��H;�H;��H;��H;ԥH;��H;�H;�eH;�EH;P H;��G;��G;-�G;�G;�cF;nE;��B;��>;�N9;>.1;�(&;�;C�;�L�:Iٶ:a��:�t,:8Y�9 �6�1p�(yƹ      ���:���:�@�:3��:r��:���:�&�:g�;��;�f$;H>.;�#6;(<;G@;�tC;�[E;�F;&$G;-�G;��G;�G;�H;�?H;�_H;�yH;^�H;�H;��H;0�H;v�H;��H;N�H;q�H;��H;��H;�H;g�H;��H;��H;��H;p�H;J�H;��H;v�H;0�H;��H;�H;Z�H;�yH;�_H;�?H;�H;�G;��G;.�G;!$G;�F;�[E;�tC;C@;(<;�#6;J>.;�f$;��;n�;�&�:��:z��:��:�@�:���:      X;�/;�w;�
;9;��;�� ;`(;Պ/;��5;
;;�%?;�5B;�^D;�E;G�F;%8G;؇G;��G;�G;�H;�<H;�[H;�uH;��H;U�H;:�H;>�H;��H;��H;��H;i�H;�H;��H;|�H;�H;��H;x�H;|�H;��H;�H;d�H;��H;��H;��H;>�H;7�H;T�H;��H;�uH;�[H;�<H;�H;�G;��G;ӇG;'8G;F�F;�E;�^D;�5B;�%?;
;;��5;ъ/;`(;�� ;�;9;�
;x;�/;      ��#;�f$;Z(&;i�(;�h,;�_0;J4;�8;�'<;�N?;��A;��C;�NE;�LF;��F;�TG;D�G;��G;��G;�H;�<H;nZH;�sH;��H;��H;��H;ԵH;ɿH;��H;�H;:�H;3�H;T�H;v�H;��H;��H;�H;��H;��H;v�H;Q�H;/�H;>�H;�H;��H;˿H;еH;��H;��H;��H;�sH;mZH;�<H;�H;��G;��G;G�G;�TG;��F;�LF;�NE;��C;��A;�N?;�'<;�8;M4;�_0;�h,;^�(;N(&;�f$;      /�6;�7;.�7;dN9;�	;;m�<;��>;p�@;�B;BD;�AE;y#F;�F;b.G;�uG;��G;G�G;��G;V H;�?H;�[H;�sH;7�H;X�H;�H;*�H;��H;%�H;��H;$�H;N�H;��H;B�H;.�H;=�H;��H;0�H;��H;:�H;/�H;?�H;��H;R�H;$�H;��H;(�H;��H;*�H;�H;T�H;1�H;�sH;�[H;�?H;V H;��G;H�G;��G;�uG;^.G;�F;}#F;�AE;=D;�B;q�@;��>;j�<;�	;;`N9;+�7;�7;      [@;�~@;,�@;��A;�PB;�1C;RD;��D;��E;�LF;b�F;�#G;1fG;�G;�G;��G;�	H;)H;�EH;�_H;�uH;�H;U�H;d�H;;�H;�H;(�H;��H;Q�H;��H;�H;��H;��H;j�H;i�H; �H;B�H;��H;g�H;j�H;��H;��H;�H;��H;Q�H;��H;$�H;�H;>�H;`�H;P�H;�H;�uH;�_H;�EH;x)H;�	H;��G;�G;�G;1fG; $G;e�F;�LF;��E;��D;SD;�1C;�PB;��A;/�@;�~@;      V�D;I�D;�
E;uNE;`�E;��E;�[F;ޱF;��F;�:G;mG;%�G;�G;��G;��G;�H;_5H;�NH;�eH;�yH;��H;��H;�H;B�H;��H;��H;)�H;��H;��H;y�H;P�H;��H;R�H;z�H;z�H;��H;�H;��H;x�H;|�H;O�H;��H;U�H;z�H;��H;��H;#�H;��H;��H;@�H;�H;��H;��H;�yH;�eH;�NH;a5H;�H;��G;��G;�G;+�G;mG;;G;��F;�F;�[F;��E;h�E;pNE;�
E;I�D;      ��F;a�F;��F;/�F;� G;#G;�FG;NhG;��G;��G;��G;��G;1�G;�H;�+H;�CH;�YH;�mH;�H;Y�H;T�H;��H;%�H;�H;��H;��H;4�H;��H;�H;�H;[�H;�H;��H;~�H;]�H;��H;��H;��H;[�H;~�H;��H;�H;[�H;�H;�H;��H;.�H;��H;��H;�H;%�H;��H;T�H;V�H;�H;�mH;�YH;�CH;�+H;�H;1�G;��G;��G;��G;��G;PhG;�FG;t#G;� G;:�F;��F;d�F;      �lG;�nG;juG;�G;ՌG;P�G;��G;~�G;��G;��G;��G;�H;�*H;�?H;�SH;fH;EwH;�H;��H;�H;>�H;ѵH;�H;+�H;(�H;4�H;T�H;��H;��H;(�H;�H;h�H;��H;m�H;��H;\�H;x�H;U�H;��H;n�H;��H;d�H;�H;(�H;��H;��H;M�H;7�H;*�H;&�H;�H;ҵH;>�H;�H;��H;چH;EwH;fH;�SH;�?H;�*H;�H;��G;��G;��G;��G;��G;L�G;�G;�G;kuG;�nG;      ��G;��G;�G;��G;��G;�G;�G;�H;8H;�!H;[2H;0CH;�SH;dH;�sH;ʁH;؎H;ŚH;ԥH;��H;A�H;ȿH;!�H;��H;��H;��H;��H;��H;�H;��H;d�H;��H;t�H;6�H;|�H;��H;�H;��H;|�H;9�H;t�H;��H;d�H;��H;�H;��H;��H;��H;��H;��H;"�H;ȿH;>�H;��H;ѥH;��H;؎H;ˁH;�sH;dH;�SH;0CH;_2H;�!H;8H;�H;�G;��G;��G;��G; �G;��G;      3H;H;LH;�H;ZH; H;*H;+5H;6AH;�MH;�ZH;�gH;�tH;�H;��H;x�H;��H;,�H;��H;0�H;��H;��H;��H;P�H;��H;�H;��H;�H;��H;L�H;q�H;��H;3�H;��H;�H;L�H;V�H;F�H;�H;��H;6�H;��H;s�H;J�H;��H;�H;��H;�H;��H;L�H;��H;��H;��H;-�H;��H;(�H;��H;y�H;��H;�H;�tH;�gH;�ZH;�MH;9AH;+5H;*H; H;dH;�H;LH;H;      �:H;|;H;�=H;�AH;GH;�MH;cUH;�]H;gH;�pH;�zH;��H;'�H;x�H;d�H;��H;װH;�H;��H;s�H;��H;�H;�H;��H;y�H;�H;&�H;��H;J�H;��H;j�H;)�H;��H;1�H;��H;��H;��H;��H;��H;1�H;��H;%�H;j�H;��H;J�H;��H;!�H;�H;z�H;��H;"�H;�H;��H;p�H;��H;�H;װH;��H;d�H;u�H;'�H;��H;�zH;�pH;gH;�]H;cUH;�MH;GH;�AH;�=H;{;H;      �bH;{cH;QeH;3hH;MlH;9qH; wH;f}H;P�H;��H;��H;b�H;ǡH;�H;�H;��H;��H;�H;�H;��H;��H;>�H;O�H;�H;S�H;[�H;�H;h�H;t�H;p�H;;�H;��H;'�H;��H;��H;��H;�H;��H;��H;��H;*�H;��H;;�H;m�H;s�H;d�H;�H;^�H;V�H;�H;T�H;>�H;��H;��H;�H;�H;��H;��H;�H;�H;ɡH;d�H;��H;��H;S�H;i}H;	wH;/qH;WlH;1hH;SeH;}cH;      ހH;t�H;ĂH;߄H;��H;��H;�H;�H;9�H;ӟH;��H;r�H;&�H;��H;ϻH;��H;��H;��H;��H;S�H;o�H;4�H;��H;��H;��H;�H;d�H;��H;��H;*�H;��H;<�H;��H;��H;�H;9�H;-�H;9�H;�H;��H;��H;:�H;��H;)�H;��H;��H;b�H;�H;��H;��H;��H;6�H;i�H;N�H;��H;��H;��H;��H;һH;��H;&�H;r�H;��H;ӟH;9�H;�H;�H;��H;�H;�H;̂H;{�H;      ,�H;��H;��H;A�H;��H;{�H;�H;��H;˪H;2�H;��H;�H;V�H;��H;��H;��H;X�H;��H;��H;w�H;�H;U�H;?�H;��H;S�H;��H;��H;z�H;9�H;��H;&�H;��H;��H;�H;Q�H;b�H;/�H;b�H;N�H;�H;��H;��H;%�H;��H;7�H;w�H;��H;��H;V�H;��H;C�H;T�H;�H;s�H;��H;��H;Z�H;��H;��H;��H;V�H;�H;��H;3�H;ΪH;��H;�H;u�H;��H;:�H;��H;��H;      -�H;k�H;O�H;ͩH;��H;ҭH;��H;W�H;��H;��H;h�H;��H;��H;��H;>�H;\�H;(�H;��H;V�H;��H;��H;y�H;+�H;a�H;w�H;z�H;i�H;9�H;��H;4�H;��H;��H;�H;I�H;h�H;o�H;��H;m�H;e�H;I�H;�H;��H;��H;0�H;��H;4�H;g�H;{�H;z�H;`�H;0�H;w�H;��H;��H;U�H;��H;-�H;\�H;>�H;��H;��H;��H;i�H;��H;��H;\�H;��H;ҭH;��H;ͩH;X�H;x�H;      ձH;�H;��H;гH;L�H;%�H;w�H;˻H;��H;M�H;7�H;)�H;��H;��H;x�H;��H;��H;��H;��H;��H;��H;��H;6�H;[�H;t�H;T�H;��H;{�H;�H;��H;��H;�H;Q�H;i�H;p�H;��H;��H;��H;m�H;i�H;S�H;�H;��H;��H;�H;v�H;��H;U�H;v�H;[�H;;�H;��H;z�H;��H;��H;��H;��H;�H;v�H;��H;��H;*�H;;�H;M�H;��H;ϻH;z�H;(�H;J�H;ӳH;��H;�H;      ��H;,�H;��H;��H;�H;��H;��H;��H;��H;�H;
�H;��H;�H;��H;��H;>�H;w�H;v�H;K�H; �H;��H;��H;��H;��H;��H;��H;W�H;��H;O�H;��H;��H;?�H;h�H;s�H;��H;��H;��H;��H;��H;w�H;j�H;=�H;��H;��H;L�H;��H;Y�H;��H;��H;��H;��H;��H;}�H;��H;J�H;y�H;{�H;A�H;��H;��H;�H;��H;�H;��H;�H;��H;��H;��H;�H;��H;��H;:�H;      �H;�H;κH;u�H;мH;`�H;3�H;9�H;Z�H;��H; �H;��H;,�H;��H;��H;&�H;)�H;�H;��H;l�H;��H;�H;.�H;8�H;�H;��H;u�H;�H;Z�H;��H;�H;1�H;1�H;��H;��H;��H;��H;��H;��H;��H;5�H;/�H;�H;��H;V�H;�H;u�H;��H;�H;8�H;3�H;�H;��H;h�H;��H;�H;)�H;'�H;��H;��H;,�H;��H;!�H;��H;^�H;=�H;5�H;_�H;ѼH;r�H;ϺH;(�H;      ��H;-�H;��H;��H;�H;��H;��H;��H;��H;�H;�H;��H;	�H;��H;��H;>�H;w�H;v�H;K�H; �H;��H;��H;��H;��H;��H;��H;W�H;��H;P�H;��H;��H;?�H;i�H;t�H;��H;��H;��H;��H;��H;v�H;j�H;=�H;��H;��H;L�H;��H;W�H;��H;��H;��H;��H;��H;}�H;��H;J�H;y�H;z�H;A�H;��H;��H;�H;��H;�H;�H;�H;��H;��H;��H;	�H;��H;��H;5�H;      ͱH;�H;��H;ȳH;L�H;#�H;x�H;ͻH;��H;M�H;8�H;)�H;��H;��H;y�H;��H;��H;��H;��H;��H;��H;��H;6�H;[�H;v�H;T�H;��H;{�H;�H;��H;��H;�H;P�H;i�H;p�H;��H;��H;��H;o�H;i�H;U�H;�H;��H;��H;�H;u�H;��H;X�H;s�H;Z�H;;�H;��H;y�H;��H;��H;��H;��H;�H;v�H;��H;��H;,�H;8�H;M�H;��H;ԻH;~�H;"�H;M�H;ȳH;��H;�H;      ,�H;j�H;O�H;ѩH;��H;׭H;��H;Z�H;��H;��H;i�H;��H;��H;��H;@�H;[�H;+�H;��H;V�H;��H;��H;|�H;+�H;c�H;|�H;z�H;j�H;9�H;��H;4�H;��H;��H;�H;I�H;f�H;m�H;��H;o�H;e�H;G�H;�H;��H;��H;0�H;��H;4�H;g�H;}�H;w�H;]�H;0�H;y�H;��H;��H;V�H;��H;+�H;]�H;@�H;��H;��H;��H;h�H;��H;��H;^�H;��H;ԭH;��H;˩H;W�H;k�H;      -�H;��H;~�H;=�H;��H;|�H;�H;��H;˪H;3�H;��H;�H;V�H;��H;��H;��H;W�H;��H;��H;w�H;�H;U�H;<�H;��H;W�H;��H;��H;z�H;;�H;��H;%�H;��H;��H;�H;P�H;c�H;/�H;b�H;P�H;�H;��H;��H;%�H;��H;3�H;u�H;��H;��H;R�H;��H;F�H;T�H;
�H;t�H;��H;��H;Z�H;��H;��H;��H;W�H;�H;��H;3�H;ϪH;��H;�H;y�H;��H;D�H;��H;��H;      ΀H;z�H;��H;݄H;��H;��H;�H;�H;6�H;ҟH;��H;q�H;$�H;��H;һH;��H;��H;��H;��H;P�H;p�H;6�H;��H;��H;��H;�H;b�H;��H;��H;)�H;��H;;�H;��H;��H;�H;6�H;-�H;8�H;�H;��H;��H;;�H;��H;(�H;��H;��H;`�H;�H;��H;��H;��H;6�H;h�H;N�H;��H;��H;��H;��H;лH;��H;&�H;r�H;��H;ԟH;<�H;�H;
�H;��H;��H;ބH;��H;q�H;      �bH;{cH;TeH;.hH;SlH;9qH;�vH;e}H;Q�H;��H;ߒH;d�H;ǡH;�H;�H;��H;��H;�H;�H;��H;��H;@�H;O�H;�H;V�H;X�H;�H;e�H;w�H;n�H;;�H;��H;'�H;��H;��H;��H;�H;��H;��H;��H;*�H;��H;:�H;k�H;p�H;b�H;�H;\�H;R�H;�H;U�H;@�H;��H;��H;�H;�H;��H;��H;�H;�H;ǡH;f�H;ߒH;��H;Q�H;l}H;wH;6qH;]lH;;hH;[eH;|cH;      �:H;�;H;�=H;�AH;
GH;�MH;bUH;�]H;gH;�pH;�zH;��H;'�H;v�H;g�H;��H;ְH;�H;��H;r�H;��H;�H;�H;��H;|�H;�H;$�H;��H;M�H;��H;j�H;)�H;��H;1�H;��H;��H;��H;��H;��H;1�H;��H;(�H;j�H;��H;H�H;��H;!�H;�H;w�H;��H;%�H;�H;��H;p�H;��H;�H;װH;��H;g�H;v�H;'�H;��H;�zH;�pH;gH;^H;fUH;�MH;GH;�AH;�=H;{;H;      >H;H;]H;�H;PH; H;*H;+5H;?AH;�MH;�ZH;�gH;�tH;�H;��H;y�H;��H;-�H;��H;-�H;��H;��H;��H;P�H;��H;�H;��H;�H;��H;I�H;q�H;��H;4�H;��H;�H;J�H;V�H;I�H;�H;��H;6�H;��H;s�H;J�H;��H;	�H;��H;�H;��H;I�H;��H;��H;��H;/�H;��H;(�H;��H;y�H;��H;�H;�tH;�gH;�ZH;�MH;=AH;15H;*H; H;cH;�H;]H;H;      ��G;��G;�G;��G;��G;�G;�G;�H;6H;�!H;[2H;-CH;�SH;dH;�sH;ˁH;؎H;ŚH;ХH;��H;A�H;ɿH;�H;��H;��H;��H;��H;��H;�H;��H;e�H;��H;r�H;7�H;{�H;��H;�H;��H;{�H;7�H;u�H;��H;g�H;��H;�H;��H;��H;��H;��H;��H;'�H;ȿH;<�H;��H;ҥH;��H;َH;ˁH;�sH;dH;�SH;/CH;\2H;�!H;8H;�H;�G;�G;��G;��G; �G;��G;      �lG;�nG;euG;�G;�G;Y�G;��G;��G;��G;��G;��G;�H;�*H;�?H;�SH;fH;DwH;��H;��H;�H;>�H;ҵH;��H;+�H;(�H;1�H;Q�H;��H;��H;'�H;�H;i�H;��H;m�H;��H;W�H;x�H;W�H;��H;n�H;��H;g�H;�H;'�H;��H;��H;P�H;8�H;)�H;'�H;�H;ԵH;<�H; �H;��H;܆H;EwH;fH;�SH;�?H;�*H;�H;��G;��G;��G;��G;��G;S�G;�G;�G;kuG;�nG;      ��F;c�F;��F;/�F;� G;�#G;�FG;PhG;��G;��G;��G;��G;1�G;�H; ,H;�CH;�YH;�mH;�H;U�H;U�H;��H;"�H;�H;��H;��H;1�H;��H;�H;�H;Z�H;�H;��H;~�H;\�H;��H;��H;��H;[�H;~�H;��H;�H;^�H;�H;�H;��H;1�H;��H;��H;�H;'�H;��H;T�H;Y�H;�H;�mH;�YH;�CH;,H;�H;3�G;��G;��G;��G;��G;LhG;�FG;u#G;� G;-�F;��F;R�F;      U�D;F�D;�
E;wNE;^�E;��E;�[F;߱F;��F;;G;mG;)�G;�G;��G;��G;�H;_5H;�NH;�eH;�yH;��H;��H;�H;A�H;��H;��H;%�H;��H;��H;v�H;S�H;��H;O�H;z�H;z�H;��H;�H;��H;x�H;|�H;R�H;��H;V�H;y�H;��H;��H;&�H;��H;��H;@�H;��H;��H;��H;�yH;�eH;�NH;a5H;�H;��G;��G;�G;(�G;mG;�:G;��F;߱F;�[F;��E;g�E;qNE;�
E;F�D;      �Z@;�~@;)�@;�A;�PB;�1C;RD;��D; �E;�LF;c�F; $G;/fG;�G;�G;��G;�	H;})H;�EH;�_H;�uH;�H;P�H;c�H;>�H;�H;&�H;��H;S�H;��H;	�H;��H;��H;j�H;h�H;��H;B�H;��H;g�H;h�H;��H;��H;�H;��H;S�H;��H;'�H;�H;=�H;e�H;U�H;��H;�uH;�_H;�EH;z)H;�	H;��G;�G;�G;0fG;�#G;c�F;�LF;��E;��D;RD;�1C;QB;�A;(�@;�~@;      $�6;�7;�7;jN9;�	;;h�<;~�>;m�@;�B;>D;�AE;z#F;�F;_.G;�uG;��G;G�G;��G;V H;�?H;�[H;�sH;3�H;W�H;�H;"�H;��H;%�H;��H; �H;Q�H;��H;A�H;.�H;=�H;��H;3�H;��H;:�H;,�H;A�H;��H;T�H;%�H;��H;$�H;�H;*�H;�H;W�H;5�H;�sH;�[H;�?H;X H;��G;H�G;��G;�uG;].G;�F;y#F;�AE;?D;�B;q�@;�>;h�<;�	;;gN9;�7;�7;      ��#;�f$;P(&;_�(;�h,;�_0;O4;�8;�'<;�N?;��A;��C;�NE;�LF;��F;�TG;D�G;��G;��G;�H;�<H;nZH;�sH;��H;��H;��H;ѵH;˿H;��H;�H;>�H;4�H;R�H;w�H;��H;��H;�H;��H;��H;u�H;T�H;2�H;@�H;�H;��H;ɿH;ҵH;��H;��H;��H;�sH;pZH;�<H;�H;��G;��G;C�G;�TG;��F;�LF;�NE;��C;��A;�N?;�'<;�8;I4;�_0;�h,;T�(;P(&;�f$;      N;�/;
x;��
;9;��;�� ;`(;֊/;��5;
;;�%?;�5B;�^D;�E;I�F;'8G;ՇG;��G;�G;�H;�<H;�[H;�uH;��H;Q�H;5�H;<�H;��H;��H;��H;i�H;
�H;��H;|�H;{�H;��H;}�H;z�H;��H;�H;h�H;��H;��H;��H;<�H;:�H;U�H;��H;�uH;�[H;�<H;�H;�G;��G;чG;%8G;G�F;�E;�^D;�5B;�%?;
;;��5;֊/;`(;�� ;��;9;��
;x;�/;      +��:���:�@�:/��:t��: ��:�&�:o�;�;�f$;J>.;�#6;(<;E@;�tC;�[E;�F;%$G;-�G;��G;�G;�H;�?H;�_H;�yH;W�H;�H;��H;2�H;r�H;��H;N�H;t�H;��H;��H;��H;h�H;��H;��H;��H;q�H;M�H;��H;u�H;0�H;��H; �H;\�H;�yH;�_H;�?H;�H;�G;��G;.�G;!$G;�F;�[E;�tC;E@;(<;�#6;J>.;�f$;�;i�;�&�:���:���:��:�@�:���:      PV�0yƹ�1p� &�6Y�9�t,:_��:Eٶ:�L�:A�;�;�(&;>.1;�N9;��>;��B;kE;�cF;�G;,�G;��G;��G;V H;�EH;�eH;�H;��H;ѥH;��H;��H;�H;��H;��H;T�H;��H;H�H;��H;H�H;��H;Q�H;��H;��H;�H;��H;��H;ѥH;��H;�H;�eH;�EH;V H;��G;��G;.�G;�G;�cF;lE;��B;��>;�N9;>.1;�(&;�;@�;�L�:Kٶ:c��:�t,: Y�9 $�6�1p�yƹ      ��4��K/�UV�E,�L�˺�쀺�uƹ@m9oQ:˂�:���:��;}�;@�,;'7;��=;QB;��D;�cF;$G;͇G;��G;��G;w)H;�NH;�mH;؆H;ĚH;)�H;�H;�H;��H;��H;��H;��H;v�H;�H;w�H;��H;��H;��H;��H;�H;�H;(�H;ĚH;܆H;�mH;�NH;x)H;��G;��G;̇G;$G;�cF;��D;QB;��=;)7;>�,;|�;��;���:͂�:oQ:@m9�uƹ�쀺S�˺J,�]V��K/�      G�ͻ2Sɻϴ��\Ϩ��-���\c��$���˺�P(��N@9n�k:`��:v;3�;�);��5;M�=;$QB;jE;�F;)8G;D�G;D�G;�	H;\5H;�YH;AwH;ՎH;��H;ѰH;��H;��H;T�H;$�H;��H;u�H;!�H;u�H;~�H;!�H;Q�H;��H;��H;԰H;��H;ՎH;BwH;�YH;W5H;�	H;G�G;D�G;"8G;�F;kE;#QB;L�=;��5; �);5�;t;Z��:r�k:�N@9�P(���˺�$��\c��-��`Ϩ�Ӵ��/Sɻ      �J;���7��9.����&����_���M����4���º�tƹHQ:���:���:&�;��(;��5;��=;��B;�[E;I�F;�TG;��G;��G;�H;�CH;fH;ɁH;y�H;��H;��H;��H;��H;V�H;��H;<�H;�H;<�H;��H;U�H;��H;��H;��H;��H;x�H;ɁH;fH;�CH;�H;��G;��G;�TG;@�F;�[E;��B;��=;��5;��(;$�;���:���:0Q: uƹ��º��4�M��c�����軫&����9.���7�      �䙼)`��i��fy��o;k��I�I�$��� �����t�|�<�x$T�X[�9�A�:p��:$�;�);'7;��>;�tC;�E;��F;�uG;�G;��G;�+H;�SH;�sH;��H;b�H;�H;̻H;��H;9�H;o�H;��H;��H;��H;n�H;9�H;��H;ȻH;�H;b�H;��H;�sH;�SH;�+H;��G;�G;�uG;��F;�E;�tC;��>;$7;�);"�;h��:�A�:H[�9�$T�<�x�|������� �I�$��I�r;k�gy��i��*`��      ������߼Nμ "���
��gy��`T�C�!���軺ۙ�iK/�����0m9�A�:���:3�;>�,;�N9;C@;�^D;�LF;Z.G;�G;��G;�H;�?H;dH;�H;q�H;	�H;��H;��H;��H;��H;��H;z�H;��H;��H;��H;��H;��H;�H;u�H;�H;dH;�?H;�H;��G;�G;^.G;�LF;�^D;F@;�N9;@�,;3�;���:�A�: m9����jK/��ۙ����D�!�`T�hy���
��#"��Nμ�߼���      ��/�E-�e.%����	�����ލǼѫ��v�{��J;��C�7Ϩ�DO:������[�9���:t;��;>.1;(<;�5B;�NE;�F;4fG;�G;.�G;�*H;�SH;�tH;"�H;��H; �H;M�H;~�H;��H;�H;�H;�H;��H;z�H;L�H;�H;��H;%�H;�tH;�SH;�*H;,�G;�G;1fG;�F;�NE;�5B;(<;;.1;}�;t;���:p[�9����GO:�8Ϩ��C��J;�u�{�ѫ��ލǼ��������f.%�E-�      \@{�W`w�zl��yZ�Q�C�dg*������� "��XO���I�<|�7Ϩ�hK/�d$T�DQ:\��:��;�(&;�#6;�%?;��C;y#F;�#G;$�G;��G;�H;)CH;�gH;~�H;\�H;j�H;�H;��H;�H;��H;��H;��H;�H;��H;�H;h�H;Y�H;��H;�gH;(CH;�H;��G;�G;�#G;y#F;��C;�%?;�#6;�(&;��;\��:4Q:l$T�jK/�8Ϩ�=|��I�XO�� "����鼮��cg*�R�C��yZ�zl�V`w�      �b��㪫��ƣ��s���ɇ�zl�BG��"�h� �-aļa���I��C��ۙ�<�uƹZ�k:���:�;D>.;
;;��A;�AE;_�F;mG;��G;��G;Y2H;�ZH;�zH;ْH;��H;��H;^�H;-�H;�H;�H;�H;-�H;\�H;��H;��H;֒H;�zH;�ZH;X2H;��G;��G;mG;_�F;�AE;��A;
;;F>.;�;���:b�k: uƹ?��ۙ��C��I�a��-aļh� ��"�BG�zl��ɇ��s���ƣ�㪫�      ������oݽ�2̽�ж����������yZ�F-�շ�,aļXO���J;����v�|���º�N@9Â�:>�;�f$;��5;�N?;;D;�LF;�:G;��G;��G;�!H;�MH;�pH;��H;ϟH;0�H;�H;B�H;v�H;��H;v�H;B�H;�H;/�H;͟H;��H;�pH;�MH;�!H;��G;��G;�:G;�LF;?D;�N?;��5;�f$;=�;���:�N@9��ºv�|���軿J;�XO��-aļշ�F-��yZ����������ж��2̽oݽ���      P,�����Z�:��z�RvϽ�b��-I��f]a�F-�h� � "��u�{�D�!�������4��P(��nQ:�L�:�;ڊ/;�'<;ߟB;��E;��F;��G;��G;5H;?AH;gH;P�H;5�H;ѪH;��H;��H;��H;V�H;��H;��H;��H;̪H;3�H;O�H;gH;@AH;5H;��G;��G;��F; �E;��B;�'<;ӊ/;�;�L�:�nQ:�P(���4�����D�!�v�{� "��h� �F-�f]a�-I���b��RvϽ�z�:��Z����      %G�p�C��$:��J+������oݽ]���-I���yZ��"����ҫ��bT��� �M����˺`m9?ٶ:i�;`(;�8;i�@;��D;�F;AhG;�G;�H;/5H;�]H;f}H;�H;��H;V�H;ɻH;��H;7�H;��H;̻H;U�H;��H;�H;e}H;�]H;15H;�H;�G;BhG;߱F;��D;g�@;�8;`(;l�;;ٶ:�m9��˺M���� �bT�ҫ������"��yZ�-I��]���oݽ������J+��$:�p�C�      {x�9t���g���T��G=�z#�6�oݽ�b������AG����ލǼgy��I�$�d����$��uƹQ��:�&�:�� ;O4;v�>;OD;�[F;�FG;~�G;�G;�)H;_UH;�vH;��H;�H;��H;l�H;��H;-�H;��H;l�H;��H;�H;��H;�vH;eUH;*H;�G;��G;�FG;�[F;RD;w�>;L4;�� ;�&�:M��:�uƹ�$�d���I�$�gy��ލǼ���AG������b��nݽ6�z#��G=���T���g�9t�      뫖���La��!���>�c�p�C�z#���RvϽ����zl�dg*����
���I���軼\c�퀺�t,:���:��;�_0;h�<;�1C;��E;t#G;S�G;�G; H;�MH;;qH;��H;|�H;ޭH;,�H;��H;_�H;��H;,�H;ܭH;{�H;��H;6qH;�MH; H;�G;S�G;|#G;��E;�1C;f�<;�_0;�;���:�t,:퀺�\c�����I��
�����dg*�zl�����RvϽ��z#�p�C�>�c�!���La����      j*��g����Ƥ�쫖��/��>�c��G=�����zｐж��ɇ�Q�C�
��""��p;k��&��-��s�˺0Y�9|��:9;�h,;�	;;�PB;g�E;� G;܌G;��G;hH;GH;OlH;��H;��H;��H;8�H;�H;ּH;�H;;�H;��H;��H;��H;LlH;GH;jH;��G;�G;� G;e�E;�PB;�	;;�h,;9;���: Y�9k�˺�-���&�p;k�#"��
��Q�C��ɇ��ж��z�����G=�>�c��/��쫖��Ƥ�g���      ��ɾ{�ž+��qת�쫖�!�����T��J+�:��2̽�s���yZ����Mμfy����\Ϩ�N,�  �6��: �
;^�(;VN9;�A;NE;/�F;�G;��G;|H;�AH;3hH;�H;?�H;ԩH;ͳH;��H;y�H;��H;ͳH;ҩH;?�H;�H;0hH;�AH;|H;��G;�G;9�F;~NE;�A;RN9;\�(;��
;��: �6K,�[Ϩ���fy��Nμ����yZ��s���2̽:��J+���T�!���쫖�qת�+��|�ž      U_ݾ�:پ�V;+���Ƥ�La����g��$:��Z�oݽ�ƣ�zl�e.%��߼g���9.�ʴ��LV�p1p��@�:x;L(&;4�7;:�@;�
E;��F;juG;$�G;OH;�=H;NeH;ĂH;s�H;L�H;��H;��H;��H;��H;��H;L�H;r�H;ÂH;IeH;�=H;OH;'�G;luG;��F;�
E;9�@;.�7;L(&;x;�@�:�1p�LV�ʴ���9.�g���߼e.%�zl��ƣ�oݽ�Z��$:���g�La���Ƥ�+���V;�:پ      ^�3���:پ{�žg�����9t�p�C�������㪫�W`w�F-����*`����7�5Sɻ�K/��xƹ���:�/;�f$;�7;�~@;K�D;Z�F;�nG;��G;"H;�;H;jcH;o�H;��H;q�H;	�H;-�H;$�H;*�H;	�H;q�H;��H;o�H;dcH;�;H;#H;��G;�nG;g�F;J�D;�~@;�7;�f$;�/;���:�xƹ�K/�6Sɻ��7�)`�����F-�W`w�㪫�������p�C�9t���g���{�ž�:پ4��      GF�Wh����UVھ7�������~���S��#��o��7S��p₽1�6�n���hy��VFB��Eֻ�A?�̾	�pY�:���:h�";i46;_@;`�D;��F;�nG;��G;�H;@H;�fH;A�H;.�H;��H;гH;йH;��H;˹H;гH;��H;.�H;A�H;�fH;@H;�H;��G;�nG;��F;_�D;Y@;a46;h�";���:rY�:Ծ	��A?��EֻVFB�hy��n���1�6�p₽7S���o���#��S��~������7��UVھ��Wh��      Vh���b���쾧*־�v��(���*��'�O�U� �s��r���؀�F�3���>ݜ�<�>�Q�ѻޡ9�����%o�:>% ;tM#;C�6;OA@;��D;��F;qG;M�G;H;�@H;hgH;��H;��H;ީH;�H;��H;޻H;��H;�H;ܩH;��H;��H;cgH;�@H;H;L�G;qG;��F;��D;JA@;<�6;pM#;<% ;)o�:����ޡ9�P�ѻ<�>�>ݜ���F�3��؀��r��s�U� �'�O�*��)����v���*־���b��      ���쾳�޾/5ʾL;���:��(�v��E�_'����q����u���+��W��A����4���Ļ9)�`j��}W�:b�;%;�k7;$�@;��D;��F;�wG;W�G;4H;=CH;*iH;�H;��H;��H;��H;��H;r�H;��H;��H;��H;��H;�H;#iH;DCH;4H;U�G;�wG;��F;��D; �@;�k7;%;`�;�W�:�j��9)���Ļ��4��A���W缃�+���u�p�����_'��E�(�v��:��L;��/5ʾ��޾��      UVھ�*־/5ʾr��������M���9b��5�����ս����Xc���ʖռ�I��U�$�kT���Z�`\���:�;n�';�8;RA;�9E;��F;ƂG;��G;CH;
GH;lH;C�H;;�H;�H;��H;��H;P�H;��H;ĵH;�H;8�H;A�H;lH;GH;CH;��G;ÂG;��F;�9E;RA;�8;h�';��;�:�\���Z�kT��U�$��I��ʖռ���Xc������ս���5��9b��M������r���/5ʾ�*־      7���v��L;������RP��D�r�z�H�U� ���5@��ѓ����K�a��վ���s�q���񕻛ܺ�4u9&�:"�;0�+;��:;�"B;n�E;��F;ՐG;��G;/H;5LH;�oH;;�H;u�H;��H;4�H;ؼH;��H;ԼH;7�H;��H;q�H;9�H;�oH;<LH;.H;��G;ԐG;��F;n�E;�"B;z�:;,�+;!�;&�:�4u9�ܺ��r����s��վ�`���K�ѓ��5@����U� �z�H�D�r�SP������L;���v��      ����)����:���M��D�r�&�O�#,�X�
��gٽpĥ���u�v1�h���)Ϥ���P�[�.o�np��@:e��:�P;>�/;=�<;C;�E;n!G;7�G;�G;�%H;�RH;�tH;��H;G�H;ׯH;�H;[�H;�H;V�H;�H;ԯH;C�H;�H;�tH;�RH;�%H;�G;4�G;t!G;�E;C;6�<;;�/;�P;k��:<:np���.o�	[򻨎P�)Ϥ�g���v1���u�pĥ��gٽX�
�#,�&�O�D�r��M���:��)���      �~��*��(�v��9b�z�H�#,�MZ����6S��x^����N������μ�I���%+����ڝ.�p����j~:K��:/m;��3;�>;>�C;=PF;�FG;S�G;��G;x/H;ZH;uzH;E�H;��H;]�H;�H;*�H;��H;'�H;�H;]�H;��H;B�H;rzH;ZH;y/H;��G;N�G;�FG;=PF;;�C;�>;��3;+m;S��:�j~:����ڝ.�����%+��I����μ�����N�x^��6S�����MZ�#,�z�H��9b�(�v�*��      �S�&�O��E��5�U� �X�
���罤9��'l���Xc���(��������[�����ݎ�@ܺp;9&��:0�	;Gd';f 8;>�@;��D;�F;jG;��G;OH;q:H;AbH;��H;�H;2�H;B�H;}�H;7�H;��H;6�H;�H;C�H;/�H; �H;��H;HbH;r:H;OH;��G;jG;�F;z�D;>�@;e 8;Cd';6�	;&��:p;9?ܺ�ݎ������[��������(��Xc�'l���9�����X�
�U� ��5��E�'�O�      �#�U� �_'������gٽ6S��'l��N�j�B�3��i��վ�y���(���Ļ\A?���B��@:�[�:Q;�.;��;;tB;�E;��F;&�G;��G;�H;TFH;%kH;��H;�H;�H;g�H;
�H;s�H;��H;p�H;�H;h�H;�H;�H;��H;*kH;VFH;�H;��G;&�G;��F;�E;tB;��;;�.;Q;�[�:��@:��B�\A?���Ļ(�y����վ��i�B�3�N�j�'l��6S���gٽ����_'�U� �      �o��s��罪�ս4@��pĥ�x^���Xc�B�3���	�Ɍ˼�]��RFB��Z򻬜��fӺ ��8��:ޛ;�M#;w=5;?;M�C;~@F;:G;�G; �G;0'H;�RH;ytH;��H;|�H;-�H;��H;��H;��H;A�H;��H;��H;��H;(�H;x�H;��H;�tH;�RH;0'H;�G;�G;	:G;y@F;O�C;?;t=5;�M#;ޛ;��:���8gӺ�����Z�QFB��]��Ɍ˼��	�B�3��Xc�x^��pĥ�5@����ս���s�      7S���r��q�����Г����u���N���(��i�Ɍ˼�A����P�fs��7|�0����\:8�:p�;xn-;�:;��A;},E;k�F;-oG;��G;�H;�7H;:_H;	~H;�H;�H;t�H;�H;x�H;;�H;��H;<�H;z�H;�H;s�H; �H;�H;~H;@_H;�7H;�H;��G;/oG;h�F;~,E;��A;�:;�n-;u�;4�:�\:0���6|��fs���P��A��Ɍ˼�i���(���N���u�ѓ�����q���r��      o₽�؀���u��Xc���K�v1�������վ��]����P����?T����9���o��3�9z&�:a�	;\%;G�5;��>;��C;�F;�!G;��G;��G;EH;`HH;�kH;��H;J�H;��H;��H;u�H;J�H;��H;��H;��H;J�H;x�H;��H;��H;M�H;��H;�kH;bHH;DH;��G;��G;�!G;�F;��C;��>;Q�5;^%;^�	;�&�:�3�9��o���9�>T�������P��]���վ�ߤ���v1���K��Xc���u��؀�      1�6�E�3���+���`�h�����μ���y���PFB�es�?T��)�D��{���:u9�q�:��:�Y;�t0;��;;�B;�9E;�F;hG;ٿG;�G;z0H;�XH;'xH; �H;v�H;�H;��H;��H;�H;/�H;3�H;/�H;�H;��H;��H;��H;z�H;(�H;-xH;�XH;z0H;��G;޿G;hG;�F;�9E;�B;��;;�t0;|Y;���:�q�:�:u9�{��(�D�=T��es�QFB�x��������μh���a�����+�D�3�      k�����W�˖ռ�վ�*Ϥ��I����[�(��Z����9��{���;9UX�:\X�:;Q;B,;��8;�A@;BD;�@F;�,G;��G;��G;gH;�DH;hH;-�H;R�H;e�H;^�H;$�H;�H;��H;��H;e�H;��H;��H;�H; �H;[�H;j�H;\�H;5�H; hH;�DH;aH;��G;��G;�,G;�@F;BD;�A@;��8;<,;DQ;ZX�:YX�:�;9�{����9���Z�(���[��I��)Ϥ��վ�˖ռ�W���      fy��>ݜ��A���I����s���P��%+������Ļ����4|��o��:u9WX�:�+�:Z;�);Մ6;w�>;�PC;e�E;��F;�xG;+�G;zH;e1H;XH; wH;��H;�H;��H;~�H;�H;A�H;��H;��H;��H;��H;��H;B�H;�H;z�H;�H;�H;��H;wH;XH;a1H;~H;,�G;�xG;��F;h�E;�PC;z�>;΄6;�);X;�+�:[X�:�:u9��o�2|�������Ļ����%+���P���s��I���A��>ݜ�      PFB�:�>���4�S�$�q��
[�����ݎ�aA?�aӺ ����3�9�q�:^X�:Z;��';�=5;��=;�B;GE;L�F;�UG;!�G;��G;SH;�HH;jH;��H;u�H;H�H;0�H;H�H;��H;@�H;�H; �H;��H;�H;�H;>�H;��H;D�H;5�H;L�H;{�H;��H;jH;�HH;YH;��G;"�G;�UG;M�F;!GE;�B;{�=;�=5;��';\;ZX�:�q�:�3�9 ���^ӺZA?��ݎ����[�t��T�$���4�7�>�      �EֻM�ѻ��ĻlT���񕻶.o�ԝ.�9ܺ��B�@��8�\:z&�:���:AQ;�);�=5;�:=;,#B;��D;�uF;�6G;ĚG;\�G;uH;�:H;^H;�zH;��H;`�H;ŲH;�H;��H;\�H;�H;m�H;2�H;��H;-�H;j�H;�H;X�H;��H;�H;ǲH;e�H;��H;�zH;^H;�:H;uH;\�G;ŚG;�6G;�uF;��D;$#B;�:=;�=5;�);BQ;���:~&�:�\: ��8x�B�3ܺ؝.��.o���pT����ĻH�ѻ      pA?�ء9� 9)��Z��ܺhp��0����;9�@:��::�:Y�	;yY;<,;΄6;x�=;!#B;��D;cXF;�!G;|�G;�G;�H;�.H;ySH;cqH;߉H;��H;c�H;��H;o�H;��H;��H;��H;��H;�H;��H;�H;�H;��H;��H;��H;t�H;ùH;f�H;��H;߉H;\qH;|SH;�.H;�H; �G;�G;�!G;dXF;��D;"#B;u�=;ф6;<,;yY;\�	;D�:��:�@: <9X���dp��}ܺ�Z�9)�ԡ9�      l�	� ���xj���[���4u9t:�j~:.��:�[�:ߛ;z�;\%;�t0;��8;{�>;	�B;��D;kXF;7G;a�G;��G;��G;�%H;KH;�iH;�H;��H;8�H;v�H;�H;[�H;��H;��H;3�H;�H;��H;S�H;��H;~�H;2�H;��H;��H;^�H;�H;v�H;7�H;��H;�H;�iH;KH;�%H;��G;��G;c�G;:G;cXF;��D;�B;~�>;��8;�t0;^%;|�;ߛ;�[�:0��:�j~:X:5u9 ]���j�����      bY�:!o�:�W�:/�:&�:m��:i��:/�	;Q;�M#;�n-;O�5;��;;�A@;�PC;"GE;�uF;�!G;c�G;��G;�G;H H;EH;�cH;8}H;u�H;��H;��H;��H;��H;��H;,�H;T�H;S�H;N�H;z�H;��H;u�H;K�H;Q�H;R�H;)�H;��H;��H;��H;��H;��H;q�H;<}H;�cH;	EH;I H;�G;��G;f�G;�!G;�uF;GE;�PC;�A@;��;;Q�5;�n-;�M#;Q;7�	;a��:w��:&�:�:uW�:o�:      ���:.% ;F�;��;�;�P;,m;@d';�.;w=5;�:;��>;�B;BD;f�E;O�F;�6G;��G;��G;�G;uH;�AH;`H;LyH;|�H;"�H;Q�H;�H;K�H;��H;��H;1�H;��H;@�H;��H;��H;C�H;��H;��H;A�H;��H;+�H;��H;��H;K�H;�H;M�H;�H;�H;IyH;`H;�AH;xH;�G;��G;��G;�6G;L�F;h�E;
BD;�B;��>;�:;u=5; �.;>d';2m;�P;!�;��;R�;,% ;      _�";xM#;%;v�';,�+;=�/;��3;a 8;��;;?;��A;��C;�9E;�@F;��F;�UG;ŚG;$�G;��G;J H;�AH;�^H;GwH;�H;��H;�H;��H;.�H;��H;%�H;�H;��H;��H;��H;m�H;K�H;y�H;E�H;m�H;��H;��H;��H;�H;&�H;��H;-�H;��H;ݫH;��H;�H;@wH;�^H;�AH;J H;��G;!�G;ǚG;�UG;��F;�@F;�9E;��C;�A;?;��;;i 8;��3;7�/;?�+;k�';	%;lM#;      }46;B�6;�k7;*�8;x�:;@�<;,�>;H�@;�tB;S�C;�,E;�F;�F;�,G;�xG;'�G;`�G;�H;�%H;EH;
`H;EwH;2�H;5�H;G�H;�H;��H;n�H;��H;��H;(�H;@�H;��H;]�H;��H;o�H;��H;i�H;��H;`�H;��H;=�H;*�H;��H;��H;n�H;��H;�H;J�H;1�H;,�H;EwH;`H;EH;�%H;�H;b�G;$�G;�xG;�,G;�F;�F;�,E;O�C;�tB;J�@;(�>;>�<;��:;)�8;�k7;&�6;      _@;VA@;�@;RA;�"B;C;?�C;~�D;�E;�@F;n�F;�!G;hG;��G;-�G;��G;vH;�.H;KH;�cH;JyH;�H;3�H;ĩH;�H;~�H;x�H;��H;�H;N�H;��H;J�H;:�H;��H;��H;^�H;��H;X�H;��H;��H;9�H;I�H;��H;M�H;�H;��H;q�H;~�H;�H;��H;-�H;�H;IyH;�cH;KH;�.H;vH;��G;/�G;��G;�gG;�!G;q�F;@F;�E;��D;?�C;�
C;�"B;RA;�@;OA@;      ��D;��D;��D;�9E;h�E;(�E;HPF;�F;��F;:G;6oG;��G;޿G;��G;~H;]H;�:H;�SH;�iH;B}H;��H;��H;K�H;�H;=�H;��H;-�H;m�H;��H;+�H;��H;	�H;��H;��H;��H;%�H;c�H; �H;��H;��H;��H;�H;��H;+�H;��H;m�H;%�H;��H;?�H;	�H;H�H;��H;��H;?}H;�iH;�SH;�:H;\H;H;��G;�G;��G;9oG;:G;��F;�F;HPF;!�E;r�E;�9E;��D;��D;      ��F;��F;��F;��F;��F;t!G;�FG;#jG;)�G;�G;��G;��G;�G;oH;e1H;�HH;^H;fqH;�H;q�H; �H;ګH;�H;~�H;��H;
�H;�H;[�H;��H;��H;��H;��H;��H;��H;x�H;��H;�H;��H;w�H;��H;��H;�H;��H;��H;��H;Z�H;�H;�H;��H;z�H;�H;۫H;�H;p�H;�H;aqH;^H;�HH;e1H;iH;�G;��G;��G;�G;,�G;'jG;�FG;j!G;��F;��F;��F;��F;      �nG;qG;�wG;ƂG;̐G;1�G;^�G;��G;��G;"�G;�H;BH;y0H;�DH;XH;jH;�zH;�H;��H;��H;V�H;��H;��H;z�H;,�H;�H;=�H;��H;]�H;{�H;K�H;��H;��H;��H;4�H;��H;��H;��H;3�H;��H;��H;��H;K�H;{�H;Z�H;��H;6�H;�H;-�H;t�H;��H;��H;U�H;��H;��H;މH;�zH;jH;XH;�DH;w0H;EH;�H;�G;��G;��G;X�G;-�G;�G;��G;�wG;qG;      ��G;H�G;P�G;��G;��G;��G;��G;LH;�H;7'H;�7H;hHH;�XH;#hH; wH;��H;��H;��H;:�H;��H;�H;*�H;j�H;��H;j�H;X�H;��H;;�H;w�H;@�H;��H;��H;��H;a�H;��H; �H;�H;��H;��H;d�H;��H;��H;��H;A�H;v�H;9�H;��H;Z�H;m�H;��H;k�H;+�H;�H;��H;8�H;��H;��H;��H;wH; hH;�XH;gHH;�7H;6'H;�H;NH;��G;��G;��G;��G;N�G;?�G;      �H;H;1H;OH;H;�%H;|/H;j:H;MFH;�RH;A_H;�kH;-xH;3�H;��H;z�H;e�H;l�H;{�H;¼H;N�H;��H;��H;�H;��H;��H;Y�H;w�H;"�H;��H;��H;��H;V�H;��H;E�H;v�H;��H;r�H;E�H;��H;W�H;��H;��H;��H;"�H;v�H;R�H;��H;��H;�H;��H;��H;K�H;��H;x�H;h�H;g�H;{�H;��H;1�H;*xH;�kH;B_H;�RH;OFH;m:H;|/H;�%H;+H;KH;/H;H;      @H;�@H;HCH;GH;>LH;�RH;ZH;?bH;(kH;~tH;~H;��H;'�H;]�H;�H;I�H;ʲH;��H;�H;��H;��H;"�H;��H;H�H;*�H;��H;z�H;A�H;��H;��H;��H;h�H;��H;O�H;��H;��H;��H;��H;��H;O�H;��H;e�H;��H;��H;��H;>�H;t�H;��H;+�H;F�H;��H;#�H;��H;��H;�H;��H;ȲH;K�H;�H;[�H;(�H;��H;~H;�tH;(kH;FbH;ZH;�RH;>LH;	GH;ICH;�@H;      �fH;xgH;.iH;lH;�oH;�tH;~zH;��H;��H;��H;��H;T�H;~�H;o�H;�H;8�H;�H;x�H;b�H;��H;��H;�H;(�H;��H;��H;��H;K�H;��H;��H;��H;h�H;�H;`�H;��H;��H;	�H;(�H;�H;��H;��H;a�H;�H;h�H;��H;��H;��H;H�H;��H;��H;��H;*�H;�H;��H;��H;a�H;u�H;�H;8�H;�H;o�H;��H;U�H;��H;��H;��H;��H;�zH;�tH;pH;lH;/iH;{gH;      C�H;��H;�H;>�H;:�H;�H;N�H;�H;$�H;~�H;�H;��H;	�H;h�H;�H;M�H;��H;��H;��H;/�H;8�H;��H;?�H;F�H;�H;�H;��H;��H;��H;j�H;��H;v�H;��H;��H;'�H;B�H;B�H;B�H;$�H;��H;��H;p�H;��H;j�H;��H;��H;��H;��H;�H;A�H;A�H;��H;2�H;,�H;��H;��H;��H;O�H;��H;g�H;	�H;��H;�H;~�H;$�H;�H;S�H;�H;E�H;>�H;�H;��H;      0�H;��H;��H;;�H;}�H;C�H;��H;.�H;�H;/�H;z�H;��H;�H;+�H;�H;��H;a�H;��H;��H;Y�H;��H;��H;��H;5�H;��H;��H;��H;��H;\�H; �H;]�H;��H;�H;6�H;U�H;x�H;~�H;x�H;S�H;8�H;�H;��H;[�H;��H;W�H;��H;��H;��H;��H;5�H;��H;��H;��H;U�H;��H;��H;b�H;��H;�H;+�H;�H;��H;}�H;1�H;�H;/�H;��H;=�H;��H;5�H;��H;��H;      ��H;ةH;��H;٫H;��H;˯H;f�H;F�H;n�H;��H;�H;��H;��H;'�H;H�H;G�H;!�H;��H;7�H;W�H;E�H;��H;Y�H;��H;��H;��H;��H;d�H;��H;Q�H;��H;��H;4�H;q�H;��H;��H;��H;��H;�H;s�H;6�H;��H;��H;O�H;��H;`�H;��H;��H;��H;��H;`�H;��H;@�H;Q�H;6�H;��H;'�H;H�H;I�H;(�H;��H;�H;�H;��H;r�H;L�H;k�H;̯H;��H;׫H;��H;�H;      ̳H;%�H;ôH;ƵH;E�H;��H;)�H;~�H;�H;��H;��H;V�H;�H;��H;��H;�H;q�H;��H;�H;O�H;��H;j�H;��H;��H;��H;n�H;-�H;��H;F�H;��H;��H;(�H;U�H;��H;��H;��H;��H;��H;��H;��H;W�H;(�H;��H;��H;A�H;��H;/�H;r�H;��H;��H;��H;i�H;��H;I�H;~�H;��H;v�H;�H;��H;��H;�H;X�H;��H;��H;�H;��H;,�H;��H;E�H;ɵH;ƴH;&�H;      ˹H;��H;��H;��H;ּH;O�H;7�H;9�H;u�H;��H;F�H;��H;5�H;��H;��H;!�H;2�H;�H;��H;y�H;��H;G�H;g�H;P�H; �H;��H;��H;�H;z�H;��H;�H;F�H;~�H;��H;��H;��H;��H;��H;��H;��H;��H;F�H;�H;��H;v�H; �H;��H;��H; �H;Q�H;n�H;G�H;��H;u�H;��H; �H;6�H;$�H;��H;��H;5�H;��H;I�H;��H;y�H;?�H;<�H;R�H;ڼH;��H;��H;�H;      ȻH;ۻH;��H;P�H;~�H;�H;��H;��H;��H;F�H;��H;��H;A�H;q�H;��H;��H;��H;��H;W�H;��H;N�H;��H;��H;��H;c�H;�H;��H;�H;��H;��H;&�H;F�H;��H;��H;��H;��H;��H;��H;��H;��H;��H;F�H;&�H;��H;��H;�H;��H;�H;c�H;��H;��H;�H;H�H;��H;W�H;��H;��H;��H;��H;t�H;A�H;��H;��H;I�H;�H;��H;��H;�H;��H;N�H;��H;�H;      ˹H;��H;��H;��H;׼H;T�H;4�H;7�H;s�H;��H;D�H;��H;6�H;��H;��H;!�H;2�H;�H;��H;y�H;��H;H�H;g�H;P�H; �H;��H;��H;�H;|�H;��H;�H;G�H;�H;��H;��H;��H;��H;��H;��H;��H;��H;F�H;�H;��H;v�H;��H;��H;��H; �H;P�H;n�H;E�H;��H;u�H;��H;!�H;4�H;$�H;��H;��H;5�H;��H;I�H;��H;y�H;?�H;:�H;R�H;ݼH;��H;��H;�H;      ³H;'�H;��H;��H;E�H;��H;*�H;��H;�H;��H;��H;V�H;!�H;��H;��H;�H;q�H;��H;~�H;N�H;��H;k�H;��H;��H;��H;m�H;/�H;��H;E�H;��H;��H;*�H;U�H;��H;��H;��H;��H;��H;��H;��H;X�H;(�H;��H;��H;A�H;��H;-�H;t�H;��H;��H;��H;j�H;��H;I�H;~�H;��H;v�H;�H;��H;��H;�H;Z�H;��H;��H;�H;��H;2�H;��H;H�H;��H;´H;'�H;      ��H;שH;��H;۫H;��H;ϯH;c�H;J�H;n�H;��H;�H;�H;��H;'�H;J�H;G�H;$�H;��H;7�H;U�H;G�H;��H;Y�H;��H;��H;��H;��H;d�H;��H;Q�H;��H;��H;5�H;q�H;��H;��H;��H;��H;�H;p�H;5�H;��H;��H;M�H;��H;`�H;��H;��H;��H;��H;`�H;��H;>�H;S�H;7�H;��H;%�H;H�H;J�H;'�H;��H;�H;�H;��H;r�H;M�H;k�H;ͯH;��H;׫H;��H;٩H;      0�H;��H;��H;6�H;v�H;D�H;��H;1�H;�H;1�H;z�H;��H;�H;+�H;�H;��H;a�H;��H;��H;X�H;��H;��H;��H;5�H;��H;��H;��H;��H;]�H; �H;]�H;��H;�H;6�H;U�H;z�H;~�H;w�H;T�H;5�H;�H;��H;[�H;��H;U�H;��H;��H;��H;��H;3�H;��H;��H;��H;V�H;��H;��H;a�H;��H;�H;+�H;�H;��H;{�H;/�H;�H;4�H;��H;@�H;|�H;=�H;��H;��H;      1�H;��H;��H;8�H;4�H;��H;P�H;�H;!�H;|�H;�H;��H;�H;g�H;��H;N�H;��H;��H;��H;.�H;8�H;��H;<�H;E�H;�H;}�H;��H;��H;��H;h�H;��H;s�H;��H;��H;(�H;@�H;B�H;B�H;&�H;��H;��H;r�H;��H;g�H;��H;��H;��H;��H;	�H;?�H;D�H;��H;/�H;,�H;��H;��H;��H;N�H;��H;g�H;
�H;��H;�H;�H;'�H;
�H;S�H;�H;:�H;;�H;�H;��H;      �fH;xgH;/iH;lH;�oH;�tH;|zH;��H;��H;��H;��H;U�H;~�H;o�H;�H;8�H;�H;x�H;b�H;��H;��H; �H;&�H;��H;��H;��H;G�H;��H;��H;��H;h�H;�H;`�H;��H;��H;�H;'�H;�H;��H;��H;a�H;�H;g�H;��H;��H;��H;G�H;��H;��H;��H;-�H;�H;��H;��H;b�H;u�H;�H;8�H;	�H;o�H;~�H;W�H;��H;��H;��H;��H;�zH;�tH;pH;lH;6iH;ygH;      @H;�@H;BCH;GH;3LH;�RH;ZH;GbH;*kH;�tH;~H;��H;(�H;\�H;�H;I�H;ʲH;��H;�H;��H;��H;#�H;��H;G�H;*�H;��H;v�H;@�H;��H;��H;��H;h�H;��H;O�H;��H;��H;��H;��H;��H;O�H;��H;g�H;��H;��H;��H;=�H;t�H;��H;*�H;D�H;��H;#�H;��H;��H;�H;��H;ʲH;I�H;�H;\�H;(�H;��H;~H;�tH;)kH;HbH;ZH;�RH;>LH;GH;SCH;�@H;      H;H;BH;HH;H;�%H;y/H;m:H;UFH;�RH;A_H;�kH;-xH;3�H;��H;{�H;d�H;m�H;x�H;��H;N�H;��H;��H;�H;��H;��H;S�H;v�H;#�H;��H;��H;��H;W�H;��H;C�H;s�H;��H;s�H;C�H;��H;Y�H;��H;��H;��H;�H;s�H;S�H;��H;��H;�H;��H;��H;K�H;��H;z�H;f�H;d�H;|�H;��H;3�H;-xH;�kH;D_H;�RH;UFH;q:H;/H;�%H;'H;FH;BH;�H;      ��G;>�G;B�G;��G;��G;�G;��G;PH;�H;7'H;�7H;gHH;�XH;#hH;wH;��H;��H;��H;7�H;��H;�H;+�H;g�H;��H;m�H;S�H;��H;7�H;x�H;>�H;��H;��H;��H;a�H;��H;��H;�H;��H;��H;d�H;��H;��H;��H;@�H;v�H;6�H;��H;X�H;l�H;��H;o�H;+�H;߹H;��H;:�H;��H;��H;��H;wH;"hH;�XH;eHH;�7H;6'H;�H;NH;��G;��G;��G;��G;P�G;>�G;      �nG;"qG;�wG;ЂG;ؐG;9�G;\�G;��G;��G;�G;�H;EH;w0H;�DH;XH;jH;�zH;�H;��H;��H;V�H;��H;��H;{�H;,�H;�H;8�H;��H;]�H;z�H;I�H;��H;��H;��H;4�H;��H;��H;��H;2�H;��H;��H;��H;L�H;{�H;Z�H;��H;9�H;�H;-�H;w�H;��H;��H;T�H;��H;��H;߉H;�zH;jH;XH;�DH;w0H;EH;�H; �G;��G;��G;a�G;5�G;ߐG;͂G;�wG;qG;      ��F;��F;��F;��F;��F;|!G;�FG;'jG;-�G;�G;��G;��G;�G;lH;f1H;�HH;^H;eqH;�H;p�H;"�H;ګH;�H;{�H;��H;�H;�H;X�H;��H;��H;��H;��H;��H;��H;x�H;��H;
�H;��H;u�H;��H;��H;��H;��H;��H;��H;X�H;�H;�H;��H;{�H;�H;ګH; �H;q�H;�H;aqH;^H;�HH;j1H;kH;�G;��G;��G;��G;&�G;"jG;�FG;n!G;��F;��F;��F;�F;      �D;��D;��D;�9E;g�E;+�E;FPF;�F;��F;:G;6oG;��G;ݿG;��G;�H;^H;�:H;�SH;�iH;?}H;��H;��H;G�H;�H;?�H;��H;'�H;l�H;��H;'�H;��H;�H;��H;��H;��H;"�H;c�H;"�H;��H;��H;��H;	�H;��H;*�H;��H;i�H;*�H;��H;=�H;�H;N�H;��H;��H;C}H;�iH;�SH;�:H;]H;�H;��G;�G;��G;6oG;:G;��F;�F;IPF;!�E;q�E;�9E;��D;��D;      @@;>A@;�@; RA;�"B;C;?�C;�D; �E;|@F;o�F;�!G;�gG;��G;/�G;��G;uH;�.H;KH;�cH;LyH;�H;.�H;éH;�H;w�H;t�H;��H;�H;J�H;��H;M�H;:�H;��H;��H;\�H;��H;^�H;��H;��H;=�H;L�H;��H;M�H;�H;��H;w�H;~�H;�H;ƩH;3�H;�H;JyH;�cH;KH;�.H;vH;��G;0�G;��G;�gG;�!G;r�F;~@F;�E;{�D;?�C;C;�"B;3RA;�@;(A@;      p46;>�6;�k7;4�8;v�:;;�<;%�>;F�@;�tB;P�C;�,E;�F;�F;�,G;�xG;(�G;`�G;�H;�%H;EH;`H;EwH;-�H;5�H;J�H;�H;��H;m�H;��H;��H;*�H;C�H;��H;_�H;��H;p�H;��H;n�H;��H;\�H;��H;A�H;/�H;��H;��H;m�H;��H;�H;H�H;5�H;0�H;GwH;
`H;EH;�%H;�H;c�G;(�G;�xG;�,G;�F;�F;�,E;S�C;�tB;J�@;%�>;;�<;t�:;/�8;�k7;)�6;      c�";xM#;%;m�';,�+;D�/;��3;e 8;��;;?;��A;��C;�9E;�@F;��F;�UG;ŚG;$�G;��G;J H;�AH;�^H;AwH;�H;��H;٫H;��H;-�H;��H;#�H;�H;��H;��H;��H;j�H;G�H;|�H;I�H;k�H;��H;��H;��H;"�H;(�H;��H;+�H;��H;ޫH;��H;�H;GwH;�^H;�AH;L H;��G;#�G;ĚG;�UG;��F;�@F;�9E;��C;��A;?;��;;i 8;��3;/�/;B�+;a�';%;jM#;      ���:D% ;X�;��;�;Q;/m;@d';�.;t=5;�:;��>;�B;BD;i�E;P�F;�6G;��G;��G;�G;uH;�AH;`H;LyH;�H;�H;K�H;߹H;K�H;��H;��H;2�H;��H;D�H;��H;��H;D�H;��H;��H;A�H;��H;/�H;��H;��H;I�H;߹H;Q�H; �H;~�H;NyH;
`H;�AH;uH;�G;��G;��G;�6G;O�F;k�E;BD;�B;��>;�:;u=5;�.;Ed';3m;�P;$�;��;f�;0% ;      �Y�:)o�:�W�:+�:&�:u��:i��:9�	;Q;�M#;�n-;O�5;��;;�A@;�PC;"GE;�uF;�!G;c�G;��G;�G;J H;EH;�cH;<}H;p�H;��H;��H;üH;��H;��H;+�H;U�H;U�H;N�H;v�H;��H;w�H;K�H;P�H;T�H;+�H;��H;��H;¼H;��H;��H;t�H;9}H;�cH;EH;I H;�G;��G;e�G;�!G;�uF;!GE;�PC;�A@;��;;O�5;�n-;�M#;Q;2�	;c��:c��:&�:�:�W�:o�:      p�	�(���pj���[���4u9l:�j~:0��:�[�:ߛ;y�;^%;�t0;��8;�>;�B;��D;gXF;7G;c�G;��G;��G;�%H;KH;�iH;��H;��H;4�H;w�H;�H;^�H;��H;��H;3�H;��H;��H;S�H;��H;~�H;2�H;��H;��H;`�H;
�H;v�H;5�H;��H;�H;�iH;
KH;�%H;��G;��G;e�G;8G;dXF;��D;�B;~�>;��8;�t0;\%;z�;ޛ;�[�:4��:�j~:h:�4u9�[���j�� ���      ~A?�С9�$9)��Z�xܺVp��@��� <9 �@:��:>�:]�	;yY;<,;ӄ6;{�=;"#B;��D;aXF;�!G;��G;!�G;�H;�.H;|SH;^qH;ىH;��H;h�H;��H;r�H;��H;��H;��H;��H;�H;��H;�H;}�H;��H;��H;��H;t�H;��H;f�H;��H;߉H;_qH;ySH;�.H;�H;!�G;}�G;�!G;cXF;��D;!#B;v�=;ӄ6;<,;xY;Z�	;D�:��:�@:<9@���`p���ܺ�Z�-9)�С9�      �EֻO�ѻ��ĻlT���񕻶.o�ם.�6ܺ��B� ��8�\:�&�:���:AQ;�);�=5;�:=;'#B;��D;�uF;�6G;ŚG;_�G;vH;�:H;^H;�zH;��H;e�H;ĲH;	�H;��H;\�H;�H;m�H;0�H;��H;0�H;j�H;�H;X�H;��H;�H;ǲH;d�H;��H;�zH;^H;�:H;vH;b�G;ŚG;�6G;�uF;��D;%#B;�:=;�=5;�);AQ;���:~&�:�\: ��8x�B�5ܺڝ.��.o���oT����ĻJ�ѻ      PFB�:�>���4�S�$�r��[�����ݎ�_A?�cӺ����3�9�q�:^X�:^;��';�=5;}�=;�B;GE;P�F;�UG;'�G;��G;YH;�HH;jH;��H;{�H;I�H;4�H;J�H;��H;B�H;�H; �H;��H; �H;�H;>�H;��H;F�H;3�H;I�H;z�H;��H;jH;�HH;SH;��G;(�G;�UG;I�F;GE;�B;{�=;�=5;��';\;\X�:�q�:�3�9���cӺ_A?��ݎ����[�t��S�$���4�:�>�      fy��>ݜ��A���I����s���P��%+������Ļ����2|� �o��:u9]X�:�+�:\;�);ӄ6;z�>;�PC;k�E;��F;�xG;-�G;~H;f1H;XH;wH;��H;�H;�H;}�H;�H;C�H;��H;��H;��H;��H;��H;B�H;�H;{�H;�H;�H;��H; wH;XH;b1H;zH;0�G;�xG;��F;d�E;�PC;w�>;΄6;�);X;�+�:WX�:�:u9�o�4|�������Ļ����%+���P���s��I���A��>ݜ�      l�����W�˖ռ�վ�)Ϥ��I����[�(��Z����9��{�� <9_X�:dX�:@Q;<,;��8;�A@;BD;�@F;�,G;��G;��G;hH;�DH;hH;3�H;V�H;j�H;`�H;"�H;�H;��H;��H;e�H;��H;��H;�H; �H;[�H;g�H;[�H;4�H;hH;�DH;dH;��G;��G;�,G;�@F;BD;�A@;��8;<,;@Q;\X�:WX�:�;9�{����9���Z�(���[��I��)Ϥ��վ�˖ռ�W���      1�6�E�3���+���`�h�����μ���y���PFB�es�>T��'�D��{�� ;u9�q�:���:}Y;�t0;��;;�B;�9E;�F;hG;ݿG;�G;y0H;�XH;-xH;$�H;y�H;�H;��H;��H;�H;/�H;3�H;/�H;�H;��H;��H;��H;w�H;'�H;-xH;�XH;w0H;�G;ٿG;hG;�F;�9E;�B;��;;�t0;yY;���:�q�:�:u9�{��)�D�?T��es�QFB�y��������μh���a�����+�E�3�      o₽�؀���u��Xc���K�v1����ߤ��վ��]����P����>T����9���o��3�9~&�:Z�	;^%;M�5;��>;��C;�F;�!G;��G;��G;BH;`HH;�kH;��H;M�H;��H;��H;x�H;J�H;��H;��H;��H;J�H;w�H;��H;��H;L�H;��H;�kH;`HH;AH;��G;��G;�!G;�F;��C;��>;N�5;[%;^�	;~&�:�3�9��o���9�?T�������P��]���վ�ߤ���v1���K��Xc���u��؀�      7S���r��r�����Г����u���N���(��i�Ɍ˼�A����P�es��4|�(����\:0�:r�;~n-;�:;��A;�,E;m�F;/oG;��G;�H;�7H;>_H;~H;�H;�H;t�H;�H;x�H;?�H;��H;=�H;z�H;�H;q�H; �H;�H;~H;A_H;�7H;�H;��G;)oG;n�F;�,E;��A;ޞ:;n-;p�;0�:�\:0���7|��fs���P��A��Ɍ˼�i���(���N���u�ѓ�����q���r��      �o��s��罪�ս4@��pĥ�x^���Xc�B�3���	�Ȍ˼�]��QFB��Z򻪜��cӺ���8��:ܛ;�M#;y=5;?;P�C;~@F;
:G;�G;�G;0'H;�RH;}tH;��H;z�H;-�H;��H;��H;��H;A�H;��H;��H;��H;*�H;x�H;��H;~tH;�RH;/'H;�G;�G;:G;@F;R�C;?;q=5;�M#;ۛ;��:���8gӺ�����Z�QFB��]��Ɍ˼��	�B�3��Xc�x^��pĥ�5@����ս���s�      �#�U� �_'������gٽ6S��'l��N�j�B�3��i��վ�y���(���ĻZA?���B���@:�[�:Q;
�.;��;;�tB;�E;��F;(�G;��G;�H;VFH;&kH;��H;�H;�H;i�H;�H;u�H;��H;s�H;�H;h�H;�H;�H;��H;(kH;VFH;�H;��G;)�G;��F; �E;�tB;��;;�.;Q;�[�:��@:��B�\A?���Ļ(�y����վ��i�B�3�N�j�'l��6S���gٽ����_'�U� �      �S�&�O��E��5�T� �X�
���罤9��(l���Xc���(��������[�����ݎ�=ܺ@;9(��:2�	;Hd';f 8;@�@;��D;�F;jG;��G;LH;p:H;@bH;��H;�H;2�H;D�H;~�H;7�H;��H;7�H;~�H;D�H;.�H;�H;��H;FbH;r:H;NH;��G;jG;�F;��D;@�@;e 8;Cd';6�	;$��:�;9;ܺ�ݎ������[��������(��Xc�'l���9�����X�
�U� ��5��E�&�O�      �~��*��(�v��9b�z�H�#,�MZ����6S��x^����N������μ�I���%+����؝.������j~:O��:0m;��3;�>;>�C;>PF;�FG;N�G;��G;y/H;ZH;wzH;E�H;��H;_�H;�H;*�H;��H;'�H;�H;]�H;��H;D�H;tzH;ZH;{/H;��G;P�G;�FG;=PF;>�C;�>;��3;+m;W��:�j~:����؝.�����%+��I����μ�����N�x^��6S�����MZ�#,�z�H��9b�(�v�*��      ����(����:���M��D�r�&�O�#,�X�
��gٽpĥ���u�v1�g���)Ϥ���P�[�.o�rp��D:i��:�P;>�/;;�<;C;�E;m!G;4�G;�G;�%H;�RH;�tH;��H;F�H;ׯH;�H;[�H;�H;[�H;�H;֯H;C�H;��H;�tH;�RH;�%H;�G;4�G;u!G;�E;C;:�<;;�/;�P;m��:<:pp���.o�[򻨎P�)Ϥ�g���v1���u�pĥ��gٽX�
�#,�&�O�D�r��M���:��)���      7���v��L;������RP��D�r�z�H�T� ���5@��Г����K�`��վ���s�q���񕻡ܺ�4u9&�:$�;-�+;��:;�"B;o�E;��F;ԐG;��G;.H;4LH;�oH;:�H;t�H;��H;3�H;ڼH;��H;ԼH;6�H;��H;q�H;:�H;�oH;<LH;/H;��G;אG;��F;n�E;�"B;|�:;-�+;!�;&�:�4u9�ܺ��q����s��վ�a���K�ѓ��5@����U� �z�H�D�r�RP������L;���v��      UVھ�*־/5ʾr��������M���9b��5�����ս����Xc���ʖռ�I��U�$�kT���Z� \���:�;k�';�8;RA;�9E;��F;G;��G;AH;	GH;lH;C�H;8�H;�H;��H;��H;S�H;��H;õH;ޫH;9�H;B�H;lH;GH;CH;��G;łG;��F;�9E;RA;�8;j�';��;�:`\���Z�jT��T�$��I��ʖռ���Xc������ս���5��9b��M������r���/5ʾ�*־      ���쾳�޾/5ʾL;���:��(�v��E�_'����q����u���+��W��A����4���Ļ9)�`j��W�:d�;%;�k7;&�@;��D;��F;�wG;W�G;4H;=CH;(iH;�H;��H;��H;��H;��H;s�H;��H;��H;��H;��H;�H;$iH;DCH;4H;W�G;�wG;��F;��D;$�@;�k7;%;`�;�W�:pj��9)���Ļ��4��A���W缃�+���u�q�����`'��E�(�v��:��L;��/5ʾ��޾��      Vh���b���쾦*־�v��(���*��'�O�U� �s��r���؀�F�3���>ݜ�<�>�Q�ѻޡ9�����'o�:@% ;tM#;C�6;OA@;��D;��F;qG;M�G;H;�@H;ggH;��H;��H;ީH;�H;��H;�H;��H;�H;ީH;��H;��H;cgH;�@H;H;L�G;qG;��F;��D;KA@;>�6;pM#;<% ;+o�:����ܡ9�R�ѻ<�>�>ݜ���F�3��؀��r��s�U� �'�O�*��(����v���*־���b��      1�$��� ����#��@��'�þ�*��0Dx���=�����Pν���"'K��c���o�V����E^���S��w[:���:e;,�4;H`?;�mD;T�F;LvG;�G;>H;aOH;�sH;��H;{�H;��H;�H;S�H;&�H;O�H;�H;��H;x�H;��H;�sH;kOH;=H;�G;OvG;^�F;�mD;B`?;#�4;e;���:�w[:��S�E^����n�V����c�!'K�����Pν�����=�0Dx��*��'�þ@��#������� �      �� ����R��O��/������0��4�s�ր:�g9��ʽ1Z����G��8�
.���5S�����/X�x�D�vBd:�B�:
 ;��4;ˈ?;�~D;�F;yG;��G;P H;*PH;tH;�H;̢H;ưH;+�H;q�H;5�H;m�H;,�H;ưH;ˢH;�H;tH;3PH;Q H;��G;yG;�F;�~D;ǈ?;��4; ;�B�:~Bd:x�D��/X���껭5S�	.���8���G�1Z���ʽg9�ր:�4�s��0�����/��O��R�����      ���R��8�
������Yؾ���ޥ����f���0�Z[�N8��ΐ���>�����IȤ��6H�`�ܻrF�����}:��:f";2�5;��?;T�D;��F;
�G;��G;2#H;bRH;�uH;F�H;£H;w�H;ĺH;�H;��H;�H;ĺH;v�H;��H;E�H;�uH;gRH;2#H;��G;	�G;��F;T�D;��?;+�5;b";��:$�}:̖�rF�`�ܻ�6H�HȤ������>�ΐ��N8��Z[���0���f�ޥ������Yؾ����8�
�R��      #��N������<I�(�þ�R��;���tS��Q"��s������}��0��켈�����6�F�ƻ6}*� �����:~x;\%;�l7;ݳ@;��D;��F;��G;��G;�'H;�UH;^xH;M�H;F�H;��H;��H;��H;x�H;��H;��H;��H;C�H;K�H;ZxH;�UH;�'H;��G;��G;��F;��D;س@;�l7;X%;{x;��:���4}*�F�ƻ��6��������0���}�����s��Q"�sS�;����R��(�þ<Iᾣ���O��      @��/�待Yؾ(�þ
Ī�|쏾�k�ր:�~�z�ؽ�����c�\y���Ҽ����C� �h�(�� #(7I�:��
;��(;�_9;��A;h\E;o�F;��G;��G;�.H;�ZH;�{H;�H;I�H;Q�H;�H;��H;v�H;��H;�H;P�H;G�H;�H;�{H;�ZH;�.H;��G;��G;s�F;g\E;��A;}_9;��(;��
;O�: !(7(��h�C� �������Ҽ\y��c�����z�ؽ~�ր:��k�|쏾
Ī�(�þ�Yؾ/��      '�þ�������R��|쏾4�s��H�����������ΐ����D��c�����;�f�R,�����P��P�9ϳ�:�;$j-;R�;;u�B;��E;]G;��G;��G;�6H;�`H;X�H;L�H;ԩH;N�H;��H;S�H;��H;O�H;��H;K�H;ѩH;J�H;V�H;�`H;�6H;��G;��G;bG;��E;p�B;K�;;"j-;�;ӳ�:@�9�P�����S,�;�f������c���D�ΐ�������������H�4�s�|쏾�R��������      �*���0��ޥ��;����k��H��#%�Z[��Pνt��`�f�1/%���伅���s�=��?ػ�FL���D�l�R:��:6�;82;��=;��C;h0F;GGG;��G;&H;�?H;�gH;��H;*�H;��H;��H;��H;��H;r�H;��H;��H;��H;��H;'�H;��H;�gH;�?H;#H;��G;LGG;h0F;��C;��=;42;2�;��:d�R:��D��FL��?ػs�=��������1/%�`�f�t���PνZ[��#%��H��k�;���ޥ���0��      0Dx�4�s���f�sS�ր:����Z[��7ս�榽��}���;��8�T�����r����9G�����̬�%��:�;�}$;ń6;�?;��D;ȔF;�pG;��G;�H;"JH;@oH;:�H;v�H;��H;7�H;��H;��H;&�H;��H;��H;9�H;��H;s�H;:�H;GoH;$JH;�H;��G;�pG;ȔF;�D;�?;Ƅ6;�}$;�;%��:�̬���9G�������r�T����8���;���}��榽�7սZ[����ր:�sS���f�4�s�      ��=�ր:���0��Q"�~������Pν�榽?����G�0����Ҽ ��GE:�;�ܻ�D^�����hi:A��:�;8|,;��:;N�A;BiE;��F;�G;��G;�(H;4UH;{wH;p�H;#�H;��H;�H;��H;��H;�H;��H;��H;�H;��H;!�H;o�H;�wH;5UH;�(H;~�G;�G;��F;>iE;O�A;��:;8|,;�;C��:`i:�����D^�9�ܻFE:� ����Ҽ1����G�?���榽�Pν����~��Q"���0�ր:�      ���g9�Z[��s�z�ؽ���t����}���G���~��/c��U�V�D,��*����������:��:T ;e�3;�0>;ƚC;�F;�8G;-�G;lH;�7H;�`H;�H;�H;��H;K�H;��H;G�H;��H;�H;��H;I�H;��H;H�H;��H;�H;�H;�`H;�7H;iH;*�G;�8G;�F;ǚC;�0>;b�3;X ;��:��:�������*��D,�U�V�/c��������G���}�t�����z�ؽ�s�Z[�g9�      �Pν�ʽN8���������ΐ��`�f���;�1����AȤ�2�f�(��Kߵ�Qo5���D�4�-:H��:�>;�+;�_9;�A;h�D;#�F;�vG;��G;H;tGH;XlH;��H;��H;��H;-�H;��H;��H;�H;$�H;�H;��H;��H;*�H;�H;��H;ǈH;alH;vGH;H;��G;�vG;�F;i�D;�A;�_9;�+;�>;F��:L�-:��D�Oo5�Iߵ�'��2�f�AȤ���0����;�`�f�͐���������N8���ʽ      ���1Z��ΐ����}��c���D�1/%��8���Ҽ/c��1�f�����ƻz/X�P������9�:>�;�";��3;>>;BYC;u�E;�G;�G;c�G;�,H; WH;xH;��H;/�H;�H;�H;��H;0�H;E�H;.�H;E�H;1�H;��H;�H;�H;2�H;��H;xH;WH;�,H;b�G;�G;�G;y�E;HYC;>>;��3;�";=�;�:���9N���x/X��ƻ���1�f�/c����Ҽ�8�1/%���D��c���}�ΐ��1Z��      !'K���G��>��0�[y��c����S��� ��T�V�'���ƻ�od�z�º �(7�4�:���:��;�P.;ҡ:;zA;-�D;ɨF;NnG;8�G;�H;�@H;"fH;]�H;,�H;��H;ԸH;��H;��H;��H;{�H;7�H;{�H;��H;��H;��H;ѸH;��H;3�H;d�H;$fH;�@H;�H;>�G;MnG;ʨF;0�D;zA;ݡ:;�P.;��;���:�4�: �(7t�º�od��ƻ'��T�V� ��R�����伔c�\y��0��>���G�      �c��8���������Ҽ����������r�GE:�C,�Iߵ�|/X���º�Ƭ�p�}:	�:�;K�);$m7;�?;��C;F;V)G;�G;E�G;�)H;�SH;�tH;\�H;{�H;�H;��H;��H;��H;�H;��H;L�H;��H;�H;��H;��H;��H;�H;��H;f�H;�tH;�SH;�)H;J�G;�G;\)G;
F;��C;�?;(m7;H�);�;�:t�}:@Ƭ�~�ºy/X�Gߵ�C,�EE:���r�����������Ҽ�켵����8�      ��
.��IȤ���������:�f�r�=����:�ܻ�*��Mo5�\��� ~(7x�}:�n�:-�;�>&;��4;��=;��B;�E;�F;��G;��G;*H;�AH;�eH;<�H;јH;X�H;ڷH;g�H; �H;��H;k�H;��H;Q�H;��H;j�H;��H;�H;d�H;ݷH;]�H;ؘH;@�H;�eH;}AH;1H;��G;��G;�F;�E;��B;��=;��4;�>&;,�;�n�:��}: �(7T���Ko5��*��6�ܻ���r�=�8�f���������JȤ�	.��      h�V��5S��6H���6�B� �S,��?ػ4G���D^������D����9�4�:	�:-�;�%;��3;�<;VB;�E;�F;�XG;��G;E H;h0H;LWH;YvH;�H;z�H;��H;��H;��H;p�H;N�H;��H;��H;8�H;��H;��H;N�H;m�H;��H;��H;��H;�H;�H;\vH;GWH;l0H;E H; �G;�XG;�F;�E;XB;�<;��3;�%;0�;	�:�4�:���9��D�����D^�4G���?ػP,�E� ���6��6H��5S�      ��ﻩ��d�ܻF�ƻc󩻶���FL� ������@��P�-:�:���:�;�>&;��3;R9<;�A;۰D;BZF;5G;��G;��G;i!H;+JH;/kH;��H;��H;c�H;��H;��H;��H;��H;��H;��H;c�H;��H;_�H;��H;��H;��H;��H;��H;��H;g�H;��H;��H;*kH;2JH;j!H;��G;��G;5G;HZF;ݰD;�A;U9<;��3;�>&;�;���:�:`�-:`������ ���FL����g�I�ƻi�ܻ���      �D^��/X�rF�(}*����P��|�D� ̬�li:��:L��:9�;��;H�);��4;�<;�A;'�D;v9F;�G;o�G;C�G;=H;?H;ZaH;}H;|�H;v�H;��H;�H;��H;b�H;�H;�H;��H;&�H;��H;%�H;��H;�H;{�H;_�H;��H;�H;��H;v�H;|�H;}H;^aH;?H;:H;F�G;o�G;�G;w9F;#�D;�A;�<;��4;F�);��;9�;X��:��:xi:�ˬ���D��P����/}*��qF��/X�      8�S���D�Ė����� "(7��9��R:3��:G��: ��:�>;�";�P.;(m7;��=;YB;ݰD;�9F; G;�G;R�G;�H;�6H;iYH;�uH;�H;�H;��H;��H;��H;�H;��H;�H;6�H;`�H;��H;��H;��H;^�H;5�H;�H;��H; �H;��H;��H;��H;�H;�H;�uH;lYH;�6H;�H;U�G;�G; G;v9F;߰D;UB;��=;(m7;�P.;�";�>;��:M��:3��:��R:��9 $(7(���Ė���D�      jw[:nBd:8�}:��:E�:׳�:�:�;�;X ;�+;��3;١:;�?;��B;�E;HZF;�G;�G;p�G;>H;T1H;�SH;`pH;ׇH;H�H;�H;y�H;��H;��H;��H;��H;p�H;"�H;��H;�H;Y�H;�H;��H;!�H;p�H;��H;��H;��H;��H;|�H;�H;D�H;ڇH;`pH;�SH;T1H;BH;p�G;�G;�G;HZF;�E;��B;�?;١:;��3;�+;W ;�;�;�:��:K�:��:�}:BBd:      &��:�B�:���:rx;��
;�;2�;�}$;6|,;e�3;�_9;:>;zA;��C;�E;�F;!5G;v�G;U�G;>H;�/H;�PH;mH;H�H;��H;��H;n�H;��H;��H;�H;\�H;��H;��H;��H;i�H;K�H;��H;D�H;k�H;��H;��H;��H;]�H;�H;��H;��H;i�H;��H;��H;E�H;�lH;�PH;�/H;>H;W�G;r�G;!5G;�F;�E;��C;zA;;>;�_9;c�3;4|,;�}$;7�;�;��
;px;؆�:�B�:      e; ;r";h%;��(;"j-;42;��6;��:;�0>;�A;BYC;0�D;F;�F;�XG;��G;I�G;�H;U1H;�PH;�kH;u�H;{�H;1�H;.�H;ּH;��H;��H;�H;k�H;��H;v�H;p�H;��H;`�H;��H;Z�H;��H;n�H;u�H;��H;n�H;�H;��H;��H;мH;+�H;4�H;x�H;m�H;�kH;�PH;U1H;�H;F�G;��G;�XG;�F;F;.�D;DYC;�A;�0>;��:;Ʉ6;82;j-;��(;Z%;f"; ;      ?�4;��4;)�5;�l7;}_9;V�;;��=;�?;V�A;˚C;q�D;|�E;ͨF;`)G;��G;�G;��G;EH;�6H;�SH; mH;r�H;��H;
�H;��H;P�H;"�H;2�H;��H;��H;�H;��H;3�H;��H;��H;a�H;��H;\�H;��H;��H;/�H;��H;�H;�H;��H;3�H;�H;O�H;��H;�H;��H;r�H;mH;�SH;�6H;=H;��G;�G;��G;])G;̨F;~�E;p�D;ƚC;V�A;�?;��=;S�;;�_9;�l7;&�5;��4;      H`?;Ԉ?;��?;ٳ@;��A;v�B;��C;�D;7iE;�F;#�F;�G;NnG;�G;��G;I H;j!H;?H;lYH;^pH;H�H;v�H;�H;E�H;��H;&�H;A�H;�H;��H;s�H;S�H;��H;��H;��H;��H;=�H;N�H;7�H;��H;��H;��H;��H;U�H;r�H;��H;�H;<�H;&�H;��H;A�H;�H;x�H;E�H;[pH;iYH;?H;m!H;I H;��G;�G;MnG;�G;&�F;�F;>iE;��D;��C;d�B;��A;ӳ@;��?;ˈ?;      �mD;�~D;P�D;��D;c\E;��E;u0F;ƔF;��F;�8G;�vG;�G;>�G;P�G;1H;s0H;6JH;haH;�uH;�H;��H;6�H;��H;��H;��H;��H;j�H;�H;��H;��H;^�H;A�H;��H;��H;��H;��H;*�H;��H;��H;��H;��H;;�H;_�H;��H;��H;�H;d�H;��H;��H;��H;��H;6�H;��H;އH;�uH;caH;6JH;r0H;2H;M�G;?�G;��G;�vG;�8G;��F;ȔF;s0F;��E;m\E;��D;P�D;�~D;      J�F;�F;��F;��F;h�F;`G;PGG;�pG;�G;1�G;��G;g�G;�H;*H;AH;OWH;0kH;}H;�H;E�H;��H;(�H;L�H;&�H;��H;0�H;��H;��H;��H;�H;�H;��H;��H;��H;;�H;��H;��H;��H;9�H;��H;��H;��H;�H;�H;��H;�H;��H;2�H;��H;#�H;K�H;)�H;��H;B�H;�H;}H;2kH;NWH;AH;*H;�H;i�G;��G;2�G;�G;�pG;NGG;XG;}�F;��F;��F;�F;      avG;yG;�G;��G;��G;��G;��G;��G;}�G;kH;H;�,H;�@H;�SH;�eH;\vH;��H;��H;�H;�H;p�H;ӼH;#�H;F�H;g�H;��H;c�H;]�H;��H;��H;`�H;��H;��H;A�H;��H;&�H;%�H; �H;��H;B�H;��H;��H;`�H;��H;��H;[�H;]�H;��H;j�H;@�H;"�H;ּH;p�H;�H;�H;{�H;��H;[vH;�eH;�SH;�@H;�,H;!H;kH;~�G;��G;��G;��G;ǝG;��G;�G;�xG;      �G;��G;��G;��G;��G;��G;1H;�H;�(H;�7H;xGH;	WH;$fH;�tH;<�H;�H;��H;v�H;��H;x�H;��H;�H;/�H;�H;�H;}�H;]�H;��H;��H;g�H;��H;��H;W�H;��H;P�H;��H;��H;��H;O�H;��H;W�H;��H;��H;e�H;��H;��H;V�H;�H;�H;�H;/�H;��H;��H;v�H;��H;s�H;��H;�H;:�H;�tH;%fH;WH;}GH;�7H;�(H;�H;0H;��G;��G;��G;��G;��G;      9H;E H;/#H;(H;u.H;�6H;�?H;JH;+UH;�`H;`lH;xH;a�H;b�H;ԘH;�H;j�H;��H;�H;��H;��H;��H;��H;��H;��H;��H;��H;��H;4�H;��H;��H;P�H;��H;s�H;��H;��H;��H;��H;��H;u�H;��H;K�H;��H;��H;1�H;��H;��H;��H;��H;��H;��H;��H;��H;��H;�H;��H;h�H;��H;֘H;`�H;^�H;xH;blH;�`H;.UH;JH;�?H;6H;�.H; (H;-#H;H H;      `OH; PH;mRH;�UH;�ZH;�`H;�gH;=oH;}wH;�H;ƈH;��H;3�H;��H;Y�H;��H;��H;�H;��H;��H;�H;�H;{�H;o�H;��H;�H;��H;g�H;��H;��H;I�H;��H;h�H;��H;��H;�H;5�H;�H;��H;��H;h�H;��H;I�H;��H;��H;d�H;��H;�H;��H;k�H;}�H;	�H;�H;��H;��H;�H;��H;��H;Y�H;��H;3�H;��H;ǈH;�H;wH;DoH;�gH;�`H;�ZH;�UH;kRH;"PH;      �sH;)tH;�uH;`xH;�{H;X�H;��H;=�H;s�H;�H;��H;8�H;��H;��H;�H;��H;��H;��H;#�H;�H;d�H;p�H;�H;S�H;_�H;�H;`�H;��H;��H;P�H;��H;l�H;��H;�H;Z�H;e�H;\�H;b�H;X�H;�H;��H;i�H;��H;O�H;��H;��H;]�H;�H;b�H;R�H;�H;n�H;`�H;��H;#�H;��H;��H;��H;�H;��H;��H;;�H;��H;�H;t�H;A�H;��H;O�H;�{H;^xH;�uH;,tH;      ��H;
�H;F�H;J�H;�H;B�H;3�H;v�H;(�H;��H;��H;�H;۸H;��H;g�H;��H;��H;f�H;��H;��H;��H;��H;��H;��H;@�H;��H;��H;��H;O�H;��H;e�H;��H;�H;[�H;��H;��H;��H;��H;��H;\�H;�H;��H;d�H;��H;L�H;��H;��H;��H;A�H;��H;��H;��H;��H;��H;��H;g�H;��H;��H;i�H;��H;ڸH;�H;��H;��H;(�H;y�H;8�H;C�H;��H;J�H;P�H;�H;      ��H;٢H;ϣH;F�H;P�H;ѩH;��H;��H;��H;N�H;2�H;�H;��H;��H;"�H;s�H;��H;��H;�H;v�H;��H;w�H;/�H;��H;��H;��H;��H;]�H;��H;n�H;��H;�H;S�H;��H;��H;��H;��H;��H;��H;��H;T�H;�H;��H;i�H;��H;W�H;��H;��H;��H;��H;3�H;w�H;��H;u�H;�H;��H;��H;v�H;$�H;��H;��H;�H;4�H;O�H;��H;��H;��H;˩H;V�H;@�H;٣H;٢H;      |�H;��H;v�H;��H;S�H;D�H;��H;;�H;��H;��H; �H;��H;��H;��H;��H;U�H;��H;!�H;<�H;%�H;��H;p�H;��H;��H;��H;��H;=�H;��H;s�H;��H;	�H;\�H;��H;��H;��H;��H;��H;��H;��H;��H;��H;[�H;	�H;��H;o�H;��H;;�H;��H;��H;��H;��H;p�H;��H;�H;;�H;"�H;��H;V�H;��H;��H;��H;��H;�H;��H;��H;>�H;��H;C�H;[�H;��H;��H;̰H;      �H;@�H;ѺH;��H;�H;��H;��H;��H;��H;R�H;��H;<�H;��H;�H;r�H;��H;��H;��H;a�H;��H;n�H;��H;��H;��H;��H;2�H;��H;P�H;��H;�H;T�H;��H;��H;��H;��H;��H;��H;��H;��H;��H;��H;��H;Q�H;��H;��H;L�H;��H;3�H;��H;��H;��H;��H;i�H;��H;^�H;��H;��H;��H;r�H;�H;��H;>�H;��H;S�H;��H;��H;��H;��H;�H;��H;ҺH;?�H;      N�H;k�H;�H;��H;��H;E�H;��H;��H;��H;��H;�H;L�H;��H;��H;��H;��H;e�H;#�H;��H;�H;N�H;]�H;Z�H;,�H;��H;��H;"�H;��H;��H;&�H;b�H;��H;��H;��H;��H;��H;��H;��H;��H;��H;��H;��H;a�H; �H;��H;��H;"�H;��H;��H;/�H;_�H;[�H;H�H;�H;��H;)�H;f�H;��H;��H;��H;��H;L�H;�H;��H;��H;��H;�H;I�H;��H;��H;�H;{�H;      +�H;2�H;��H;w�H;r�H;��H;{�H;)�H;�H;�H;3�H;<�H;D�H;Z�H;[�H;?�H;��H;��H;��H;b�H;��H;��H;��H;D�H;)�H;��H; �H;��H;��H;?�H;Z�H;��H;��H;��H;��H;��H;��H;��H;��H;��H;��H;��H;X�H;9�H;��H;��H;"�H;��H;(�H;F�H;��H;��H;��H;]�H;��H;��H;��H;A�H;[�H;[�H;D�H;>�H;5�H;�H;�H;-�H;�H;��H;u�H;x�H;��H;;�H;      O�H;o�H;�H;��H;��H;K�H;��H;��H;��H;��H;�H;K�H;��H;��H;��H;��H;e�H;&�H;��H;�H;O�H;^�H;Z�H;,�H;��H;��H;"�H;��H;��H;$�H;b�H;��H;��H;��H;��H;��H;��H;��H;��H;��H;��H;��H;a�H;�H;��H;��H; �H;��H;��H;.�H;_�H;Z�H;H�H;�H;��H;)�H;f�H;��H;��H;��H;��H;L�H;�H;��H;��H;��H;�H;H�H;��H;��H;�H;x�H;      ߹H;C�H;˺H;��H;�H;��H;��H;��H;��H;R�H;��H;<�H;��H;�H;t�H;��H;��H;��H;^�H;��H;p�H;��H;��H;��H;��H;0�H;��H;P�H;��H;�H;T�H;��H;��H;��H;��H;��H;��H;��H;��H;��H;��H;��H;S�H;��H;��H;J�H;��H;6�H;��H;��H;��H;��H;g�H;��H;`�H;��H;��H;��H;q�H;�H;��H;?�H;��H;R�H;��H;��H;��H;��H;�H;��H;ѺH;A�H;      |�H;��H;v�H;��H;S�H;G�H;��H;>�H;��H;��H;�H;��H;��H;��H;��H;U�H;��H;"�H;;�H;#�H;��H;q�H;��H;��H;��H;��H;>�H;��H;u�H;��H;�H;\�H;��H;��H;��H;��H;��H;��H;��H;��H;��H;[�H;�H;��H;n�H;��H;;�H;��H;��H;��H;��H;p�H;��H;!�H;;�H;!�H;��H;X�H;��H;��H;��H;��H; �H;��H;��H;@�H;��H;F�H;]�H;��H;�H;��H;      �H;ߢH;̣H;C�H;L�H;ԩH;��H;��H;��H;N�H;3�H;�H;��H;��H;%�H;t�H;��H;��H;�H;w�H;��H;w�H;.�H;��H;��H;��H;��H;\�H;��H;o�H;��H;�H;Q�H;��H;��H;��H;��H;��H;��H;��H;S�H;�H;��H;i�H;��H;V�H;��H;��H;��H;��H;6�H;v�H;��H;u�H;�H;��H;��H;v�H;$�H;��H;��H;�H;3�H;N�H;��H;��H;��H;ΩH;R�H;J�H;ڣH;آH;      ��H;�H;5�H;F�H;�H;S�H;4�H;y�H;&�H;��H;��H;�H;ظH;��H;j�H;��H;��H;g�H;��H;��H;��H;��H;��H;��H;A�H;��H;��H;��H;R�H;��H;e�H;��H;�H;Z�H;��H;��H;��H;��H;��H;[�H;�H;��H;b�H;��H;K�H;��H;��H;��H;@�H;��H;��H;��H;��H;��H;��H;g�H;��H;��H;i�H;��H;ڸH;�H;��H;��H;*�H;|�H;:�H;F�H;�H;G�H;<�H;�H;      �sH;)tH;�uH;ZxH;�{H;X�H;��H;;�H;s�H;�H;��H;;�H;��H;��H;�H;��H;��H;��H;"�H;��H;d�H;p�H;�H;S�H;_�H;	�H;[�H;��H;��H;O�H;��H;n�H;��H;�H;[�H;c�H;\�H;e�H;X�H;�H;��H;k�H;��H;L�H;��H;��H;]�H;�H;_�H;P�H;�H;p�H;^�H;��H;%�H;��H;��H;��H;�H;��H;��H;;�H;��H;�H;t�H;D�H;��H;V�H;�{H;exH;�uH;*tH;      nOH;)PH;dRH;�UH;�ZH;�`H;�gH;GoH;�wH;�H;ǈH;��H;3�H;��H;\�H;��H;��H;�H;��H;��H;�H;�H;w�H;l�H;��H;�H;��H;d�H;��H;��H;K�H;��H;g�H;��H;��H;�H;5�H;�H;��H;��H;i�H;��H;K�H;�H;��H;a�H;��H;�H;��H;i�H;��H;	�H;�H;��H;��H;߾H;��H;��H;[�H;��H;3�H;��H;ǈH;�H;wH;GoH;�gH;�`H;�ZH;�UH;wRH; PH;      GH;E H;@#H;�'H;m.H;�6H;�?H;JH;4UH;�`H;`lH;xH;`�H;b�H;טH;��H;h�H;��H; �H;��H;��H;��H;��H;��H;��H;��H;��H;��H;4�H;��H;��H;R�H;��H;u�H;��H;��H;��H;��H;��H;s�H;��H;O�H;��H;��H;0�H;��H;��H;��H;��H;��H;��H;��H;��H;��H;�H;��H;h�H;��H;טH;b�H;a�H;xH;blH;�`H;5UH;"JH;�?H;�6H;~.H;�'H;>#H;? H;      !�G;��G;��G;��G;��G;��G;0H;�H;�(H;�7H;yGH;WH;$fH;�tH;?�H;�H;��H;w�H;��H;x�H;��H;��H;,�H;�H;�H;v�H;X�H;��H;��H;b�H;��H;��H;V�H;��H;Q�H;��H;��H;��H;P�H;��H;Y�H;��H;��H;d�H;��H;��H;Y�H;}�H;�H;�H;6�H;��H;��H;x�H;��H;q�H;��H;�H;@�H;�tH;%fH;WH;{GH;�7H;�(H;�H;/H;��G;��G;��G;��G;��G;      OvG;yG;�G;��G;��G;��G;��G;��G;~�G;iH;H;�,H;�@H;�SH;�eH;]vH;��H;��H;�H;�H;r�H;ּH;�H;F�H;h�H;��H;^�H;\�H;��H;��H;^�H;��H;��H;B�H;��H;"�H;%�H;"�H;��H;D�H;��H;��H;a�H;��H;��H;[�H;^�H;��H;k�H;A�H;)�H;ּH;p�H;�H;�H;|�H;��H;]vH;�eH;�SH;�@H;�,H;!H;kH;�G;��G;��G;��G;ŝG;��G;
�G;	yG;      B�F;�F;��F;��F;n�F;iG;IGG;�pG;�G;0�G;��G;j�G;�H;*H;�AH;OWH;/kH;}H;�H;D�H;��H;(�H;H�H;&�H;��H;,�H;��H;��H;��H;�H;�H;��H;��H;��H;;�H;��H;��H;��H;9�H;��H;��H;��H;�H;�H;��H;|�H;��H;2�H;��H;%�H;P�H;(�H;��H;E�H;�H;}H;3kH;OWH;�AH;*H;�H;i�G;��G;4�G;�G;�pG;LGG;\G;v�F;��F;��F;�F;      �mD;�~D;M�D;��D;a\E;��E;r0F;ǔF;��F;�8G;�vG;�G;<�G;M�G;4H;s0H;6JH;haH;�uH;��H;��H;8�H;��H;��H;��H;��H;d�H;�H;��H;��H;^�H;B�H;��H;��H;��H;��H;(�H;��H;��H;��H;��H;B�H;c�H;��H;��H;�H;g�H;��H;��H;��H;��H;8�H;��H;�H;�uH;caH;7JH;r0H;6H;O�G;?�G;�G;�vG;�8G;��F;ȔF;s0F;��E;k\E;��D;O�D;�~D;      )`?;��?;��?;�@;��A;~�B;��C;��D;EiE;�F;'�F;�G;KnG;�G;��G;I H;j!H;?H;hYH;]pH;H�H;w�H;�H;C�H;��H;�H;=�H;�H;��H;p�H;U�H;��H;��H;��H;��H;9�H;O�H;:�H;��H;��H;��H;��H;Y�H;s�H;��H;�H;A�H;&�H;��H;E�H;�H;w�H;H�H;`pH;jYH;?H;m!H;K H;��G;�G;MnG;�G;'�F;�F;?iE;�D;��C;r�B;��A;�@;��?;��?;      1�4;��4;�5;�l7;z_9;P�;;��=;
�?;[�A;ɚC;m�D;~�E;̨F;`)G;��G;�G;��G;DH;�6H;�SH;mH;r�H;��H;�H;��H;I�H;�H;2�H;��H;z�H;�H;��H;2�H;��H;��H;a�H;��H;a�H;��H;��H;2�H;��H;�H;��H;��H;2�H;#�H;O�H;��H;
�H;��H;t�H;mH;�SH;�6H;?H;��G;�G;��G;])G;ͨF;{�E;l�D;ɚC;V�A;�?;��=;R�;;y_9;�l7;�5;��4;      e; ;f";\%;��(;(j-;82;Ƅ6;��:;�0>;�A;FYC;.�D;	F;�F;�XG;��G;I�G;�H;U1H;�PH;�kH;p�H;x�H;5�H;%�H;ѼH;��H;��H;�H;n�H;��H;u�H;p�H;��H;[�H;��H;]�H;��H;m�H;v�H;��H;r�H;�H;��H;��H;ּH;.�H;2�H;~�H;u�H;�kH;�PH;X1H;�H;G�G;��G;�XG;�F;
F;0�D;BYC;�A;�0>;��:;Ʉ6;22;j-;�(;N%;f";  ;      ��:�B�:��:yx;��
;�;4�;�}$;:|,;b�3;�_9;=>;zA;��C;�E;�F;5G;v�G;U�G;>H;�/H;�PH;�lH;F�H;��H;��H;g�H;��H;��H;�H;]�H;��H;��H;��H;j�H;G�H;��H;H�H;j�H;��H;��H;��H;`�H;�H;��H;��H;l�H;��H;��H;I�H;mH;�PH;�/H;AH;X�G;u�G;!5G;�F;�E;��C;zA;:>;�_9;e�3;8|,;�}$;9�;�;��
;wx;���:�B�:      �w[:�Bd: �}:��:E�:��:�:�;�;X ;�+;��3;ܡ:;�?;��B;�E;FZF;�G;�G;p�G;BH;W1H;�SH;^pH;ۇH;D�H;ݪH;v�H;��H;��H;��H;��H;s�H;"�H;��H;�H;\�H;�H;��H;�H;r�H;��H;��H;��H;��H;x�H;�H;H�H;هH;dpH;�SH;U1H;AH;r�G;�G;�G;FZF;�E;��B;�?;ڡ:;��3;�+;W ;�;�;�:ϳ�:O�:��:(�}:bBd:      4�S���D����І�� (7��9��R:/��:O��:��:�>;�";�P.;(m7;��=;YB;ݰD;z9F;G;�G;W�G;�H;�6H;iYH;�uH;�H;�H;��H;��H;��H;�H;��H;�H;8�H;a�H;��H;��H;��H;^�H;6�H;�H;��H;"�H;��H;��H;��H;�H;�H;�uH;mYH;�6H;�H;W�G;�G;G;w9F;ݰD;UB;��=;'m7;�P.;�";�>;��:M��:3��:��R:��9 (7І��ؖ���D�      �D^��/X�rF�.}*����P��|�D�@ˬ��i:��:R��::�;��;H�);��4;�<;�A;$�D;v9F;�G;q�G;E�G;?H;?H;^aH;}H;x�H;t�H;��H;�H;��H;`�H;�H;�H;��H;&�H;��H;(�H;��H;�H;�H;_�H;��H;�H;��H;t�H;|�H;}H;ZaH;?H;?H;E�G;n�G;�G;v9F;$�D;�A;�<;��4;E�);��;9�;X��:��:|i:�ˬ���D��P����2}*�rF��/X�      ��ﻫ��d�ܻE�ƻc󩻶���FL��������P��X�-:�:���:�;�>&;��3;U9<;�A;ڰD;EZF;!5G;��G;��G;l!H;2JH;-kH;��H;��H;h�H;��H;��H;��H;��H;��H;��H;c�H;��H;c�H;��H;��H;��H;��H;��H;��H;h�H;��H;��H;,kH;/JH;o!H;��G;��G;5G;HZF;۰D;�A;T9<;��3;�>&;�;���:�:T�-:`������ ���FL����h�I�ƻi�ܻ���      i�V��5S��6H���6�C� �P,��?ػ3G���D^������D����9�4�:�:1�;�%;��3;�<;SB;�E;�F;�XG;�G;F H;l0H;LWH;XvH;�H;~�H;��H;��H;��H;p�H;T�H;��H;��H;8�H;��H;��H;M�H;m�H;��H;��H;��H;~�H;�H;XvH;KWH;h0H;F H;�G;�XG;��F;�E;SB;�<;��3;�%;0�;	�:�4�:���9��D�����D^�4G���?ػQ,�E� ���6��6H��5S�      ��	.��JȤ���������9�f�r�=����9�ܻ�*��Ko5�X��� �(7|�}:�n�:.�;�>&;��4;��=;��B;�E;�F;��G;��G;/H;�AH;�eH;=�H;טH;Y�H;޷H;g�H; �H;��H;j�H;��H;Q�H;��H;j�H;��H;�H;c�H;ݷH;Y�H;ؘH;<�H;�eH;~AH;-H;��G;��G;�F;�E;��B;��=;��4;�>&;,�;�n�:x�}: ~(7X���Mo5��*��8�ܻ���s�=�8�f���������JȤ�
.��      �c��8���������Ҽ����������r�FE:�C,�Hߵ�z/X�~�º@Ƭ���}:�:�;F�);%m7;�?;��C;	F;[)G;�G;L�G;*H;�SH;�tH;b�H;�H;�H;��H;��H;��H;�H;��H;M�H;��H;�H;��H;��H;��H;�H;��H;c�H;�tH;�SH;�)H;E�G;�G;])G;	F;��C;�?;#m7;H�);�;	�:t�}:�Ƭ���ºz/X�Hߵ�C,�FE:���r�����������Ҽ�켴����8�      !'K���G��>��0�[y��c����R��� ��T�V�&���ƻ�od�v�º �(7�4�:���:��;�P.;֡:;zA;-�D;̨F;QnG;>�G;�H;�@H;"fH;c�H;/�H;��H;ָH;��H;��H;��H;}�H;7�H;}�H;��H;��H;��H;ѸH;��H;0�H;c�H;"fH;�@H;�H;8�G;OnG;ͨF;.�D;zA;ڡ:;�P.;��;���:�4�: �(7x�º�od��ƻ'��U�V� ��R�����伔c�\y��0��>���G�      ���1Z��ΐ����}��c���D�1/%��8���Ҽ/c��1�f�����ƻy/X�N������9�:9�;�";��3;B>;BYC;{�E;�G;�G;e�G;�,H;WH;xH;��H;4�H;�H;�H;��H;0�H;D�H;0�H;E�H;0�H;��H;�H;�H;1�H;��H;xH; WH;�,H;c�G;�G;�G;|�E;DYC;:>;��3;�";<�;�:���9N���{/X��ƻ���1�f�/c����Ҽ�8�1/%���D��c���}�ΐ��1Z��      �Pν�ʽN8���������ΐ��`�f���;�1����AȤ�2�f�'��Jߵ�No5���D�<�-:D��:�>;�+;�_9;�A;j�D;#�F;�vG;��G;H;vGH;^lH;ÈH;��H;��H;-�H;��H;��H;�H;%�H;�H;��H;��H;*�H;�H;��H;ňH;`lH;uGH;H;��G;�vG;$�F;l�D;�A;�_9;�+;�>;D��:D�-:��D�Oo5�Kߵ�(��2�f�AȤ���1����;�`�f�ΐ���������N8���ʽ      ���g9�Z[��s�z�ؽ���t����}���G���~��/c��U�V�D,��*����������:��:V ;i�3;�0>;ɚC;�F;�8G;+�G;iH;�7H;�`H;
�H;�H;��H;K�H;��H;G�H;��H;�H;��H;G�H;��H;H�H;��H;�H;�H;�`H;�7H;fH;+�G;�8G;�F;ʚC;�0>;_�3;X ;��:��:�������*��D,�U�V�/c��������G���}�t�����{�ؽ�s�Z[�g9�      ��=�ր:���0��Q"�~������Pν�榽?����G�0����Ҽ ��GE:�9�ܻ�D^�����\i:E��:�;<|,;��:;Q�A;BiE;��F;�G;�G;�(H;4UH;|wH;q�H;!�H;��H;�H;��H;��H;�H;��H;��H;�H;��H;!�H;o�H;}wH;5UH;�(H;~�G;�G;��F;EiE;O�A;��:;4|,;�;A��:`i:�����D^�:�ܻGE:� ����Ҽ1����G�?���榽�Pν����~��Q"���0�ր:�      0Dx�4�s���f�sS�ր:����Z[��7ս�榽��}���;��8�T�����r����8G����@ͬ�)��:�;�}$;Ƅ6;�?;��D;˔F;�pG;��G;�H;!JH;@oH;;�H;v�H;��H;9�H;��H;��H;&�H;��H;��H;7�H;��H;s�H;:�H;EoH;$JH;�H;��G;�pG;ǔF;��D;�?;ń6;�}$;�;#��:�̬���9G�������r�T����8���;���}��榽�7սZ[����ր:�sS���f�4�s�      �*���0��ޥ��;����k��H��#%�Z[��Pνt��`�f�1/%���伅���s�=��?ػ�FL���D�l�R:��:4�;62;��=;��C;h0F;GGG;��G;#H;�?H;�gH;��H;*�H;��H;��H;~�H;��H;t�H;��H;��H;��H;��H;*�H;��H;�gH;�?H;%H;��G;MGG;f0F;��C;��=;42;0�;�:d�R:��D��FL��?ػs�=��������1/%�`�f�t���PνZ[��#%��H��k�;���ޥ���0��      '�þ�������R��{쏾5�s��H�����������ΐ����D��c�����;�f�R,�����P��P�9ӳ�:�;!j-;R�;;v�B;��E;[G;��G;��G;�6H;�`H;[�H;M�H;ԩH;O�H;��H;R�H;��H;R�H;��H;N�H;ҩH;L�H;W�H;�`H;�6H;��G;��G;cG;��E;w�B;O�;;!j-;�;׳�:H�9�P�����R,�;�f������c���D�ΐ�������������H�5�s�|쏾�R��������      @��/�待Yؾ(�þ
Ī�|쏾�k�ր:�~�z�ؽ�����c�\y���Ҽ����B� �g�*�� "(7M�:��
;��(;�_9;��A;j\E;l�F;��G;��G;�.H;�ZH;�{H;�H;H�H;S�H;�H;��H;v�H;��H;�H;O�H;G�H;�H;�{H;�ZH;�.H;��G;��G;u�F;g\E;��A;~_9;��(;��
;Q�: !(7&��h�B� �������Ҽ\y��c�����z�ؽ~�ր:��k�|쏾
Ī�(�þ�Yؾ/��      #��O������<I�(�þ�R��;���tS��Q"��s������}��0��켇�����6�E�ƻ6}*�������:~x;Z%;�l7;ܳ@;��D;��F;��G;��G;�'H;�UH;`xH;M�H;D�H;��H;��H;��H;z�H;��H;��H;��H;D�H;M�H;]xH;�UH;�'H;��G;��G;��F;��D;ܳ@;�l7;X%;{x;��:���2}*�D�ƻ��6��������0���}�����s��Q"�sS�;����R��(�þ<Iᾣ���O��      ���R��8�
������Yؾ���ޥ����f���0�Z[�N8��ΐ���>�����IȤ��6H�`�ܻrF�����}:���:c";0�5;��?;V�D;��F;	�G;��G;0#H;`RH;�uH;F�H;��H;v�H;úH;�H;��H;�H;ĺH;v�H;��H;E�H;�uH;gRH;2#H;��G;
�G;��F;T�D;��?;+�5;b";��:,�}:Ȗ�rF�`�ܻ�6H�HȤ������>�ΐ��N8��Z[���0���f�ޥ������Yؾ����8�
�R��      �� ����R��N��/������0��4�s�ր:�g9��ʽ1Z����G��8�
.���5S�����/X�p�D�zBd:�B�: ;��4;ˈ?;�~D;�F;yG;��G;O H;*PH;tH;�H;̢H;ưH;,�H;o�H;6�H;n�H;,�H;ǰH;ˢH;�H;tH;3PH;P H;��G;yG;�F;�~D;ǈ?;��4; ;�B�:�Bd:��D��/X���껭5S�	.���8���G�1Z���ʽg9�ր:�4�s��0�����/��N��R�����      EEb�`]��N��7����s� ���˾��(�j��!,�o���K��Bm�*��6,˼��x�Z���1�����`�:t�:�;�1;:,>;e�C;VwF;�G;n H;�>H;�hH;,�H;A�H;�H;��H;��H;�H;l�H;�H;��H;��H;�H;@�H;)�H;�hH;�>H;p H;��G;_wF;e�C;6,>;�1;�;t�:l�:
����1��Z����x�6,˼*��Bm�K��o����!,�(�j�����˾s� �����7��N�`]�      `]�d�W��TI�v3��D�������Ǿv����f�7)�$��r;���Fi��k���Ǽ�[t�L�	�(Ȅ�X��ܠ:��:��;.J2;VZ>;'	D;>F;8�G;�H;�?H;viH;ÈH;��H;Q�H;�H;��H;5�H;��H;1�H;��H;�H;P�H;��H;��H;{iH;�?H;�H;8�G;FF;'	D;PZ>;(J2;��;��:�:X��'Ȅ�L�	��[t���Ǽ�k��Fi�r;��$��7)��f�v�����Ǿ�����D�v3��TI�d�W�      �N��TI���;�/�'�l��쾀���x󐾴Z��K ��s�@����&^���"����g����̨u�� ���2<:��:�
;>g3;��>;WBD;x�F;ޔG;kH;BH;\kH;.�H;��H;	�H;��H;A�H;��H;"�H;��H;A�H;��H;�H;��H;)�H;ckH;BH;lH;ߔG;��F;WBD;��>;7g3;�
;��:�2<:� ��ʨu������g��"����&^�@����s潥K ��Z�x󐾀�����l�/�'���;��TI�      �7�v3�/�'����s� ��{Ծ���G���y�F�����ӽ���^�L�Iv��뮼OT����PV���=�f)i:z��:�z ;�$5;��?;�D;��F;�G;sH;dFH;rnH;b�H;K�H;J�H;��H;	�H;1�H;��H;-�H;�H;��H;H�H;J�H;^�H;xnH;fFH;rH;�G;��F;�D;��?;{$5;�z ;v��:v)i:��=��PV���OT��뮼Iv�^�L�����ӽ���y�F�G�������{Ծs� ����/�'�v3�      ����D�l�s� �U�ݾj���U͓��f��>/�����'���섽N�6�}t�w��\�:�$Tʻw.� ۷�Ft�:�;��$;�Y7;T�@;�	E;��F;+�G;�H;LH;�rH;��H;��H;��H;��H;�H;$�H;��H;!�H;�H;��H;��H;��H;��H;�rH;	LH;�H;)�G;��F;�	E;M�@;�Y7;��$;�;Nt�:(۷�x.�$Tʻ]�:�w��}t�N�6��섽�'������>/��f�U͓�j���V�ݾs� �l��D�      s� ��������{Ծj���v���Y�x��SC��^��޽?���w�e�'��B�Ѽ#G������R����� ޤ8ɇ�:�Y;H�);��9;��A;��E;�G;�G;@!H;
SH;�wH;I�H;Y�H;�H;��H;I�H;V�H;��H;R�H;K�H;��H;�H;Y�H;G�H;�wH;
SH;A!H;
�G;�G;��E;��A;��9;E�);�Y;χ�:�ݤ8����R�����#G��B�Ѽ'��w�e�?����޽�^��SC�Y�x�v���j����{Ծ�쾟���      ��˾��Ǿ�������U͓�Y�x���J��K �l���������?����뮼(�[����3|��W����:C�:�';d/;Cg<;�C;GF;�NG;��G;-H;:[H;�}H;��H;��H;��H;�H;��H;��H;��H;��H;��H;�H;��H;��H;��H;�}H;=[H;-H;��G;�NG;FF;�C;@g<;b/;�';I�:��:�W��3|����'�[��뮼���?������l����K ���J�Y�x�U͓����������Ǿ      ��v���x�G����f��SC��K �mn����Ž���
�Z��k�}ռ,X��_y-�)���l.�`��P�:�+�:�;4;�>;�D;�wF;�G;��G;�9H;'dH;T�H;��H;2�H;H�H;��H;~�H;+�H;E�H;)�H;��H;��H;E�H;/�H;~�H;Z�H;*dH;�9H;��G;�G;�wF;�D;�>;4;{�;�+�:�P�:X��k.�)���^y-�,X��}ռ�k�
�Z������Žmn���K ��SC��f�G���x�v���      (�j��f��Z�y�F��>/��^�l�����ŽF ���Fi��Q+�zt�lT��l�W�����1��$Ⱥ8X�9yP�:�Y;��(;��8;�A;�E;��F;<�G;sH;�FH;�mH;j�H;��H;�H;H�H;��H;`�H;��H;��H;��H;a�H;��H;D�H;�H;��H;o�H;�mH;�FH;pH;8�G;��F;�E;�A;��8;��(;�Y;yP�:(X�9 Ⱥ�1�����l�W�lT��yt�Q+��Fi�F ����Žl����^��>/�x�F��Z��f�      �!,�7)��K ��������޽������Fi��0����鷼��x�����.��M�(����
+i:z��:(�;��0;8�<;tC;��E;�<G;��G;�$H;:TH;�wH;ǒH;�H;!�H;X�H;�H;c�H;s�H;O�H;q�H;f�H;�H;U�H;�H;�H;ΒH;�wH;;TH;�$H;��G;�<G;��E;uC;:�<;��0;.�;~��:+i:���N�(��.�������x�鷼����0��Fi�������޽�������K �7)�      n���$��s��ӽ�'��?������	�Z��Q+�����"��G����0���׻ƕb�4W���X�9ء�:`;�*';�Y7;�#@;�D;�F;�G;��G;8H;�aH;́H;5�H;z�H;H�H;l�H;x�H;W�H;%�H;�H;&�H;Z�H;y�H;i�H;F�H;|�H;<�H;ҁH;�aH;8H;��G;�G;ߖF;	�D;�#@;�Y7;�*';"`;ԡ�:Y�92W��ŕb���׻��0�G���"������Q+�	�Z����>����'���ӽ�s�$��      J��r;��@�������섽v�e��?��k�zt�鷼G���e7�����Ǆ�j0� �t� u�:,�:n;m1;D�<;L�B;�E;�G;��G;3H;QJH;3oH;ҋH;��H;�H;m�H;��H;��H;j�H;��H;��H;��H;j�H;��H;��H;k�H;�H;��H;ۋH;4oH;QJH;0H;��G;�G;�E;O�B;E�<;x1;p;�+�:*u�:��t�h0��Ǆ���껂e7�G��鷼yt��k��?�v�e��섽���@���r;��      Bm��Fi��&^�^�L�N�6�'����}ռlT����x���0����������ط��n`:��:�;�*;�8;��@;�D;E�F;�}G;z�G;l1H;�[H;C|H;��H;��H;Y�H;��H;��H;^�H;h�H;��H;E�H;��H;g�H;^�H;��H;��H;]�H;��H;��H;F|H;�[H;h1H;�G;�}G;H�F;"�D;��@;(�8;�*;�;��:o`:hط��������껽�0���x�lT��}ռ��&��O�6�_�L��&^��Fi�      )���k��Iv�{t�C�Ѽ�뮼+X��l�W������׻�Ǆ��� ��5<:\��:�Y;�t%;�$5;�Z>;�`C;��E;*G;B�G;�H;�GH;ElH;ǈH;ӞH;��H;��H;n�H;��H;��H;K�H;F�H;�H;F�H;J�H;��H;��H;m�H;��H;��H;ܞH;ʈH;ElH;�GH;�H;A�G;*G;��E;�`C;�Z>;�$5;�t%;�Y;\��:5<:������Ǆ���׻���j�W�+X���뮼B�Ѽ}t�Jv���k�      4,˼��Ǽ�"���뮼w��#G��&�[�\y-�����.��ĕb�p0㺈ط�5<:�L�:�\;r�!;�J2;�g<;/0B;CE;�F;'�G;��G;^4H;v\H;�{H;~�H;v�H;/�H;��H;�H;i�H;$�H;&�H;��H;��H;��H;%�H;$�H;h�H;�H;��H;5�H;|�H;��H;�{H;r\H;b4H;��G;(�G;�F;CE;80B;�g<;�J2;x�!;�\;�L�:5<:�ط�l0���b��.�����\y-�&�[�!G��w���뮼�"����Ǽ      ��x��[t���g�LT�\�:�������$����1��J�(�.W��@�t��n`:\��:�\;{ ;��0;T;;�<A;��D;�wF;�cG;-�G;�!H;�MH;YoH;J�H;Z�H;��H;e�H;9�H;��H;/�H;D�H;��H;m�H;��H;k�H;��H;D�H;,�H;��H;=�H;i�H;��H;]�H;M�H;RoH;�MH;�!H;0�G;�cG;�wF;��D;�<A;N;;��0;{ ;�\;\��:�n`:��t�*W��I�(��1��$���������^�:�NT���g��[t�      V��I�	������Tʻ�R��3|�d.�Ⱥ���0Y�9$u�:��:�Y;v�!;��0;Օ:;��@;�BD;f2F;Z8G;��G;�H;@@H;�cH;��H;I�H;�H;�H;!�H;d�H;��H;��H;@�H;��H;��H;W�H;��H;�H;B�H;��H;��H;i�H;$�H;�H;�H;K�H;��H;�cH;B@H;�H;��G;[8G;j2F;�BD;��@;ؕ:;��0;x�!;�Y;��:(u�:8Y�9���Ⱥd.�3|��R��#Tʻ�����G�	�      �1��"Ȅ�̨u��PV�i.����zW��0��@X�9+i:ܡ�:�+�:�;�t%;�J2;K;;��@;]D;�F;G;X�G;hH;Z5H;VZH;xH;�H;��H;�H;�H;-�H;?�H;��H;�H;��H;�H;2�H;��H;/�H;�H;��H;��H;��H;C�H;3�H;�H;�H;��H;�H;
xH;UZH;U5H;jH;Z�G;	G;�F;ZD;��@;H;;�J2;�t%;�;�+�:衼:+i:hX�9��W�����f.��PV�¨u�#Ȅ�      إ��*X��� ��l�=� ۷��ߤ8��:�P�:�P�:���:'`;n;�*;�$5;�g<;�<A;�BD;�F;�G;X�G;A�G;w-H;�RH;-qH;��H;��H;Q�H;�H;�H;��H;��H;��H;'�H;��H;r�H;j�H;��H;g�H;p�H;��H;$�H;��H;��H;��H;�H;�H;Q�H;��H;��H;/qH;�RH;z-H;C�G;Z�G;�G;�F;�BD;�<A;�g<;�$5;�*;p;*`;���:�P�:�P�:��: ߤ8۷���=�� ��,X��      L�:ؠ:�2<:�)i:Ft�:χ�:]�:�+�:�Y;.�;�*';v1;$�8;�Z>;80B;��D;j2F;G;Z�G;��G;W)H;\NH;JlH; �H;8�H;X�H;q�H;�H;Z�H;��H;�H; �H;�H;/�H;��H;��H;��H;��H;��H;.�H;�H;��H;�H;��H;Z�H;�H;p�H;U�H;<�H; �H;HlH;]NH;Y)H;��G;\�G;
G;j2F;��D;:0B;�Z>;$�8;w1;�*';.�;�Y;�+�:W�:݇�:Jt�:^)i:�2<:��:      ��:���:���:f��:�;�Y;�';x�;��(;��0;�Y7;@�<;��@;�`C;CE;�wF;Z8G;b�G;C�G;U)H;�LH;�iH;�H;/�H;z�H;��H;��H;9�H;��H;��H;��H;-�H;��H;o�H;��H;}�H;��H;v�H;��H;n�H;��H;)�H;��H;��H;��H;9�H;��H;��H;|�H;.�H;�H;�iH;�LH;W)H;C�G;^�G;[8G;�wF;CE;�`C;��@;A�<;�Y7;��0;~�(;w�;�';�Y;�;f��:��:���:      �;��;;�z ;��$;G�);`/;4;��8;<�<;$@;K�B;!�D;��E;�F;�cG;��G;nH;{-H;^NH;�iH;�H;��H;��H;��H;��H;z�H;w�H;�H;��H;H�H;�H;�H;��H;��H;F�H;��H;@�H;��H;��H;�H;�H;K�H;��H;�H;w�H;v�H;��H;��H;��H;��H;�H;�iH;^NH;{-H;kH;��G;�cG;�F;��E;!�D;L�B;$@;:�<;��8;4;d/;C�);��$;�z ; ;��;      ,�1;,J2;5g3;�$5;�Y7;��9;Sg<;�>;�A;yC;�D;	�E;I�F;*G;*�G;3�G;�H;_5H;�RH;HlH;	�H;��H; �H;��H;^�H;?�H;3�H;	�H;��H;��H;a�H;��H;^�H;��H;��H;�H;I�H;��H;��H;��H;[�H;��H;d�H;��H;��H;�H;/�H;>�H;`�H;��H;��H;��H;�H;HlH;�RH;Z5H;�H;1�G;*�G;*G;H�F;
�E;�D;tC;�A; �>;Mg<;��9;�Y7;�$5;2g3;J2;      9,>;^Z>;��>;��?;I�@;��A;�C;�D;�E;��E;�F;�G;�}G;E�G;��G;�!H;C@H;]ZH;/qH;�H;.�H;��H;��H;��H;��H;��H;�H;��H;��H;��H;<�H;�H;��H;z�H;@�H;��H;��H;��H;=�H;z�H;�H;�H;=�H;��H;��H;��H;�H;��H;��H;�H;��H;��H;.�H;�H;-qH;XZH;E@H;�!H;��G;A�G;�}G;�G;�F;��E;�E;�D;�C;��A;S�@;��?;��>;VZ>;      ��C;%	D;QBD;�D;�	E;��E;QF;�wF;��F;�<G;��G;��G;�G;�H;e4H;�MH;dH;xH;��H;C�H;��H;��H;d�H;��H;"�H;��H;��H;P�H;W�H;��H;��H;Z�H;z�H;2�H;��H;>�H;?�H;8�H;��H;3�H;u�H;T�H;��H;��H;R�H;M�H;��H;��H;$�H;��H;`�H;��H;��H;?�H;��H;xH;dH;�MH;f4H;�H;��G;��G;��G;�<G;��F;�wF;QF;��E;�	E;�D;QBD;%	D;      KwF;BF;}�F;��F;��F;�G;�NG;
�G;9�G;��G;��G;6H;n1H;�GH;u\H;\oH;��H;�H;��H;U�H;��H;��H;<�H;��H;��H;A�H;�H;�H;��H;{�H;	�H;H�H;)�H;��H;g�H;��H;��H;��H;d�H;��H;(�H;D�H;	�H;y�H;��H;�H;
�H;C�H;��H;��H;:�H;��H;��H;S�H;��H;�H;��H;YoH;v\H;�GH;n1H;7H;��G;��G;<�G;�G;�NG;}G;��F;��F;z�F;EF;      �G;?�G;ڔG;�G; �G;
�G;��G;��G;mH;�$H;8H;PJH;�[H;HlH;�{H;M�H;O�H;�H;U�H;q�H;��H;w�H;4�H;#�H;��H;�H;��H;Z�H;A�H;��H;(�H;�H;��H;~�H;��H;��H;�H;��H;��H;~�H;��H;�H;(�H;��H;;�H;U�H;��H;�H;��H;�H;3�H;x�H;��H;p�H;S�H;��H;N�H;M�H;�{H;ClH;�[H;QJH;8H;�$H;oH;��G;��G;�G;5�G;�G;۔G;*�G;      p H;�H;eH;yH;�H;@!H;-H;�9H;�FH;BTH;�aH;:oH;E|H;͈H;}�H;]�H;�H;�H;�H;�H;:�H;u�H;�H;��H;J�H;
�H;W�H;O�H;��H;��H;��H;��H;p�H;��H;�H;X�H;\�H;T�H;�H;��H;n�H;��H;��H;��H;��H;L�H;S�H;�H;O�H;��H;�H;u�H;9�H;�H;�H;�H;�H;]�H;~�H;͈H;F|H;:oH;�aH;ATH;�FH;�9H;-H;5!H;�H;wH;eH;�H;      �>H;|?H;BH;tFH;�KH;
SH;A[H;#dH;�mH;�wH;ҁH;ًH;��H;ٞH;y�H;��H;!�H;�H;�H;[�H;��H;�H;��H;��H;R�H;�H;9�H;��H;�H;��H;��H;e�H;��H;/�H;i�H;��H;��H;��H;h�H;1�H;��H;`�H;��H;��H;�H;��H;4�H;��H;U�H;��H;��H;�H;��H;X�H;�H;�H;!�H;��H;y�H;؞H;��H;ًH;ׁH;�wH;�mH;&dH;>[H;SH;LH;rFH;BH;}?H;      �hH;jiH;gkH;nnH;�rH;�wH;�}H;S�H;m�H;̒H;:�H;��H;��H;��H;0�H;g�H;%�H;/�H;��H;��H;��H;��H;}�H;��H;��H;q�H;��H;��H;��H;��H;i�H;��H;�H;v�H;��H;��H;��H;��H;��H;v�H;�H;��H;i�H;��H;��H;��H;��H;v�H;��H;��H;~�H;��H;��H;��H;��H;/�H;%�H;h�H;2�H;��H;��H;��H;=�H;ђH;m�H;W�H;�}H;�wH;�rH;qnH;gkH;miH;      1�H;ԈH;3�H;d�H;��H;K�H;��H;��H;��H;�H;��H;�H;c�H;��H;��H;@�H;n�H;G�H;��H;�H;��H;K�H;a�H;=�H;��H;	�H;)�H;��H;��H;p�H;��H;*�H;��H;��H;��H;��H;��H;��H;��H;��H;��H;'�H;��H;o�H;��H;��H;$�H;�H;��H;:�H;d�H;K�H;��H;�H;��H;F�H;p�H;A�H;��H;��H;d�H;�H;��H;�H;��H;��H;��H;A�H;��H;d�H;5�H;ֈH;      H�H;��H;��H;J�H;��H;P�H;��H;2�H;�H;!�H;M�H;r�H;��H;w�H;�H;��H;��H;��H;��H;�H;3�H;�H;��H;�H;W�H;C�H;�H;��H;b�H;��H;#�H;w�H;��H;��H;��H;��H;�H;��H;��H;��H;��H;v�H;!�H;��H;^�H;��H; �H;F�H;Z�H;�H;��H;�H;/�H;�H;��H;��H;��H;��H;�H;u�H;��H;t�H;Q�H;"�H;�H;5�H;��H;P�H;��H;J�H;��H;��H;      �H;]�H;�H;M�H;�H;�H;��H;D�H;A�H;Z�H;o�H;��H;��H;��H;k�H;3�H;��H;�H;,�H;�H;��H;"�H;]�H;~�H;z�H;&�H;��H;u�H;��H;!�H;~�H;��H;��H;��H;�H;�H;��H;�H;�H;��H;��H;��H;}�H;�H;��H;o�H;��H;)�H;{�H;~�H;`�H;!�H;��H;�H;,�H;�H;��H;6�H;n�H;��H;��H;��H;s�H;[�H;F�H;E�H;��H;�H;
�H;F�H;�H;^�H;      �H;�H;��H;��H;��H;��H;��H;��H;��H;�H;��H;��H;h�H;��H;*�H;I�H;G�H;�H;��H;6�H;v�H;��H;��H;r�H;2�H;��H;z�H;��H;/�H;x�H;��H;��H;��H;��H;(�H;0�H;�H;0�H;'�H;��H;��H;��H;��H;v�H;+�H;��H;y�H;��H;4�H;q�H;��H;��H;q�H;/�H;��H;�H;L�H;K�H;+�H;��H;g�H;��H;��H;�H;��H;��H;��H;��H; �H;��H;��H;�H;      ��H;��H;L�H;�H;�H;D�H;��H;��H;d�H;m�H;b�H;t�H;u�H;T�H;-�H;��H;��H;�H;t�H;��H;��H;��H;~�H;2�H;��H;^�H;��H;�H;j�H;��H;��H;��H;�H;)�H;�H;'�H;F�H;(�H;�H;+�H;�H;��H;��H;��H;e�H;�H;��H;a�H;��H;3�H;��H;��H;��H;��H;r�H;�H;��H;��H;-�H;T�H;u�H;u�H;e�H;p�H;i�H;��H;��H;D�H;�H;�H;O�H;��H;      �H;0�H;��H;.�H;�H;L�H;��H;.�H;��H;z�H;-�H;��H;��H;J�H;��H;m�H;��H;0�H;k�H;��H;��H;D�H;��H;��H;7�H;��H;��H;X�H;��H;��H;��H;��H;�H;3�H;)�H;�H;2�H;�H;(�H;7�H;�H;��H;��H;��H;��H;T�H;��H;��H;7�H;��H;�H;C�H;{�H;��H;j�H;5�H;��H;o�H;��H;M�H;��H;��H;0�H;{�H;��H;/�H;��H;N�H;"�H;-�H;��H;?�H;      q�H;��H;9�H;��H;��H;��H;��H;H�H;��H;R�H;�H;��H;P�H;�H;��H;��H;b�H;��H;��H;��H;��H;��H;I�H;��H;A�H;��H;�H;b�H;��H;��H;��H;�H;�H;�H;G�H;/�H; �H;2�H;F�H;�H;�H;�H;��H;��H;��H;^�H;�H;��H;?�H;��H;O�H;��H;��H;��H;��H;��H;b�H; �H;��H;�H;P�H;��H;�H;T�H;��H;K�H;��H;��H;��H;��H;:�H;��H;      �H;5�H;��H;.�H; �H;P�H;��H;,�H;��H;z�H;,�H;��H;��H;M�H;��H;m�H;��H;0�H;k�H;��H;��H;D�H;��H;��H;7�H;��H;��H;W�H;��H;��H;��H;��H;�H;5�H;,�H;�H;2�H;�H;(�H;6�H;�H;��H;��H;��H;��H;S�H;��H;��H;7�H;��H;�H;@�H;{�H;��H;j�H;5�H;��H;o�H;��H;L�H;��H;��H;0�H;x�H;��H;0�H;��H;N�H;%�H;1�H;��H;<�H;      ��H;��H;E�H;�H;�H;@�H;��H;��H;e�H;n�H;b�H;t�H;s�H;T�H;.�H;��H;��H;�H;t�H;��H;��H;��H;~�H;2�H;��H;[�H;��H;�H;j�H;��H;��H;��H;�H;)�H;�H;(�H;F�H;)�H;�H;+�H;�H;��H;��H;��H;e�H;	�H;��H;a�H;��H;2�H;��H;��H;��H;��H;r�H;�H;��H;��H;,�H;T�H;u�H;w�H;b�H;n�H;g�H;��H;��H;=�H;�H;�H;M�H;��H;      �H;�H;��H;��H;��H;��H;��H;��H;��H;�H;��H;��H;g�H;��H;-�H;I�H;J�H;�H;��H;3�H;v�H;��H;��H;r�H;3�H;��H;z�H;��H;1�H;x�H;��H;��H;��H;��H;)�H;/�H;�H;0�H;'�H;��H;��H;��H;��H;t�H;(�H;��H;y�H;��H;0�H;n�H;��H;��H;m�H;0�H;��H;�H;J�H;L�H;-�H;��H;g�H;��H;��H;�H;��H;��H;��H;��H;�H;��H;��H;�H;      �H;b�H;�H;G�H; �H;�H;��H;H�H;C�H;Z�H;p�H;��H;��H;��H;o�H;4�H;��H;�H;+�H;
�H;��H;!�H;Z�H;~�H;{�H;!�H;��H;s�H;��H;!�H;}�H;��H;��H;��H;�H;	�H;��H;�H;�H;��H;��H;��H;}�H;�H;��H;n�H;��H;(�H;z�H;}�H;b�H;�H;��H;�H;+�H;�H;��H;6�H;n�H;��H;��H;��H;s�H;X�H;D�H;H�H;��H;�H;�H;N�H; �H;[�H;      7�H;��H;��H;C�H;��H;`�H;��H;6�H;�H; �H;M�H;r�H;��H;u�H;�H;��H;��H;��H;��H;�H;4�H;	�H;��H;�H;Z�H;@�H; �H;��H;e�H;��H;!�H;w�H;��H;��H;��H;��H;�H;��H;��H;��H;��H;v�H; �H;��H;^�H;��H;��H;F�H;X�H;�H;��H;	�H;-�H; �H;��H;��H;��H;��H;�H;u�H;��H;t�H;O�H;"�H;�H;6�H;��H;S�H;��H;F�H;��H;��H;      %�H;ԈH;3�H;^�H;��H;I�H;��H;��H;��H;�H;��H;�H;c�H;��H;��H;A�H;p�H;G�H;��H;�H;��H;M�H;`�H;<�H;��H;�H;$�H;��H;��H;o�H;��H;*�H;��H;��H;��H;��H;��H;��H;��H;��H;��H;(�H;��H;l�H;��H;��H;$�H;�H;��H;9�H;g�H;M�H;��H;�H;��H;F�H;q�H;A�H;��H;��H;d�H;�H;��H;�H;��H;��H;��H;G�H;��H;k�H;:�H;ԈH;      �hH;siH;akH;znH;�rH;�wH;�}H;[�H;q�H;ϒH;:�H;��H;��H;��H;5�H;h�H;%�H;0�H;��H;��H;��H;��H;z�H;��H;��H;o�H;��H;��H;��H;��H;k�H;��H;�H;v�H;��H;��H;��H;��H;��H;v�H;�H;��H;i�H;��H;��H;��H;��H;u�H;��H;��H;��H;��H;��H;��H;��H;-�H;%�H;i�H;3�H;��H;��H;��H;=�H;ђH;n�H;[�H;�}H;�wH;�rH;|nH;rkH;liH;      �>H;z?H;#BH;oFH;�KH;SH;=[H;&dH;�mH;�wH;ҁH;ًH;��H;ٞH;|�H;��H;�H;�H;�H;X�H;��H;�H;��H;��H;S�H;z�H;6�H;��H;�H;��H;��H;e�H;��H;/�H;i�H;��H;��H;��H;h�H;/�H;��H;b�H;��H;��H;�H;��H;6�H;��H;S�H;��H;��H;�H;��H;[�H;�H;�H;�H;��H;|�H;ڞH;��H;ًH;ՁH;�wH;�mH;)dH;B[H;
SH;LH;mFH;!BH;s?H;      y H;�H;[H;zH;�H;L!H;-H;�9H;�FH;ATH;�aH;9oH;E|H;ΈH;��H;]�H;�H;�H;�H; �H;:�H;v�H;�H;��H;M�H;�H;S�H;L�H;��H;��H;��H;��H;n�H;��H;�H;U�H;^�H;W�H;�H;��H;p�H;��H;��H;��H;��H;I�H;T�H;�H;L�H;��H;�H;v�H;7�H;�H;�H;�H;�H;]�H;��H;ΈH;F|H;:oH;�aH;ATH;�FH;�9H;-H;:!H;�H;wH;gH;�H;      �G;E�G;ܔG;��G;.�G;�G;��G;��G;oH;�$H;8H;TJH;�[H;FlH;�{H;N�H;N�H;�H;S�H;p�H;��H;x�H;/�H;#�H;��H;
�H;��H;W�H;@�H;��H;%�H;�H;��H;~�H;��H;��H;�H;��H;��H;��H;��H;�H;)�H;��H;;�H;U�H;��H;�H;��H; �H;9�H;z�H;��H;r�H;T�H;��H;N�H;N�H;�{H;FlH;�[H;QJH;8H;�$H;oH;��G;��G;
�G;5�G;��G;�G;6�G;      AwF;AF;��F;��F;��F;�G;�NG;�G;@�G;��G;��G;9H;p1H;�GH;w\H;\oH;��H;�H;��H;T�H;��H;��H;8�H;��H;��H;<�H;
�H;�H;��H;u�H;�H;H�H;(�H;��H;g�H;��H;��H;��H;d�H;��H;)�H;H�H;�H;x�H;��H;�H;�H;C�H;��H;��H;?�H;��H;��H;U�H;��H;�H;��H;\oH;z\H;�GH;o1H;7H;��G;��G;8�G;
�G;�NG;�G;��F;��F;m�F;1F;      ��C;!	D;PBD;�D;�	E;��E;RF;�wF;��F;�<G;��G;��G;��G;�H;i4H;�MH;dH;xH;��H;@�H;��H;��H;^�H;��H;$�H;��H;��H;M�H;V�H;��H;��H;X�H;w�H;3�H;��H;;�H;A�H;;�H;��H;4�H;z�H;Z�H;��H;��H;S�H;J�H;��H;��H;$�H;��H;e�H;��H;��H;@�H;ÉH;xH;dH;�MH;j4H;�H;��G;��G;��G;�<G;��F;�wF;RF;��E;�	E;�D;QBD;#	D;      ,>;CZ>;��>;��?;D�@; �A;�C;�D;�E;��E;�F;�G;�}G;E�G;��G;�!H;C@H;]ZH;-qH;�H;/�H;��H;��H;�H;��H;��H;�H;��H;��H;��H;<�H;�H;�H;{�H;=�H;��H;��H;��H;=�H;z�H;��H;�H;A�H;��H;��H;��H;�H;��H;��H;��H;��H;��H;/�H; �H;/qH;[ZH;E@H;�!H;��G;E�G;�}G;�G;�F;��E;�E;�D;�C;��A;\�@;ů?;��>;.Z>;      �1;$J2;)g3;�$5;~Y7;��9;Jg<;�>;�A;vC;�D;
�E;H�F;*G;.�G;5�G;�H;^5H;�RH;HlH;�H;��H;��H;��H;`�H;7�H;-�H;	�H;��H;{�H;a�H;��H;[�H;��H;��H;�H;L�H;�H;��H;��H;`�H;��H;g�H;��H;��H;�H;4�H;>�H;^�H;��H;��H;��H;�H;IlH;�RH;Z5H;�H;3�G;.�G;*G;I�F;�E;�D;vC;�A; �>;Kg<;��9;~Y7;�$5;)g3;J2;      �;��; ;�z ;��$;L�);e/;4;��8;:�<;$@;Q�B;!�D;��E;�F;�cG;��G;lH;z-H;^NH;�iH;�H;��H;��H;��H;��H;t�H;v�H;�H;��H;H�H;�H;�H;��H;��H;A�H;��H;D�H;��H;��H;�H;�H;N�H;��H;�H;v�H;z�H;��H;��H;��H;��H;�H;�iH;`NH;{-H;kH;��G;�cG;�F;��E;!�D;L�B; $@;:�<;��8;4;^/;6�);��$;�z ;;��;      ��:��:��:t��:�;�Y;�';{�;��(;��0;�Y7;B�<;��@;�`C;CE;�wF;[8G;a�G;A�G;W)H;�LH;�iH;�H;/�H;{�H;��H;��H;7�H;��H;��H;��H;-�H;��H;o�H;��H;x�H;��H;z�H;��H;k�H;��H;-�H;��H;��H;��H;7�H;��H;��H;z�H;0�H;�H;�iH;�LH;Y)H;D�G;^�G;Z8G;�wF;CE;�`C;��@;>�<;�Y7;��0;��(;�;�';�Y;�;t��:%��:���:      ��:�:�2<:�)i:Ft�:݇�:a�:�+�:�Y;,�;�*';w1;'�8;�Z>;;0B;�D;j2F;G;Y�G;��G;Y)H;^NH;IlH; �H;<�H;S�H;j�H;�H;Z�H;��H;�H;��H;�H;0�H;��H;��H;��H;��H;��H;,�H;�H; �H;�H;��H;[�H;�H;q�H;W�H;9�H;$�H;JlH;]NH;[)H;��G;Z�G;
G;j2F;��D;;0B;�Z>;&�8;v1;�*';,�;�Y;�+�:W�:ˇ�:Nt�:v)i:�2<:Р:      ֥��.X��� ��t�=�@۷��ߤ8��:�P�:�P�:���:'`;p;�*;�$5;�g<;�<A;�BD;�F;�G;Y�G;C�G;z-H;�RH;+qH;��H;��H;M�H;�H;
�H;��H;��H;��H;%�H;��H;r�H;h�H;��H;h�H;p�H;��H;'�H;��H;��H;��H;�H;�H;Q�H;��H;��H;1qH;�RH;z-H;D�G;\�G;�G;�F;�BD;�<A;�g<;�$5;�*;n;'`;���:�P�:�P�:��:`ߤ8@۷�x�=�� ��$X��      �1��Ȅ�Ϩu��PV�d.����~W�����xX�9+i:⡼:�+�:�;�t%;�J2;N;;��@;\D;�F;G;Z�G;hH;Z5H;XZH;xH;�H;��H;�H;�H;*�H;A�H;��H; �H;��H;�H;2�H;��H;3�H;�H;��H; �H;��H;C�H;2�H;�H;�H;��H;�H;xH;XZH;[5H;jH;X�G;
G;�F;ZD;��@;K;;�J2;�t%;�;�+�:桼:+i:hX�9 ��W�����e.��PV�بu� Ȅ�      V��J�	������Tʻ�R��	3|�c.�Ⱥ���8Y�9*u�:��:�Y;|�!;��0;ؕ:;��@;�BD;h2F;[8G;��G;�H;C@H;�cH;��H;H�H;�H;�H;�H;g�H;��H;��H;C�H;��H;��H;Z�H;��H;��H;@�H;��H;��H;i�H;"�H;�H;�H;I�H;��H;�cH;C@H;�H;��G;X8G;l2F;�BD;��@;ؕ:;��0;z�!;�Y;��:$u�:8Y�9���Ⱥc.�3|��R��$Tʻ�����I�	�      ��x��[t���g�MT�\�:�������#����1��K�(�*W����t��n`:\��:�\;{ ;��0;O;;�<A;��D;�wF;�cG;1�G;�!H;�MH;WoH;H�H;Y�H;��H;e�H;:�H;��H;-�H;E�H;��H;k�H;��H;k�H;��H;B�H;,�H;��H;<�H;g�H;��H;Z�H;H�H;VoH;�MH;�!H;3�G;�cG;�wF;��D;�<A;N;;��0;{ ;�\;Z��:�n`:��t�,W��K�(��1��$���������_�:�MT���g��[t�      5,˼��Ǽ�"���뮼w��"G��&�[�\y-�����.����b�p0㺀ط�5<:�L�:�\;v�!;�J2;�g<;40B;CE;�F;,�G;��G;b4H;v\H;�{H;��H;y�H;0�H;��H;�H;h�H;&�H;&�H;��H;��H;��H;%�H;&�H;h�H;�H;��H;2�H;|�H;~�H;�{H;u\H;a4H;��G;+�G;�F;CE;70B;�g<;�J2;v�!;�\;�L�:5<:�ط�p0�Õb��.�����\y-�'�[�"G��w���뮼�"����Ǽ      )���k��Iv�{t�B�Ѽ�뮼+X��k�W������׻�Ǆ������ 5<:d��:�Y;�t%;�$5;�Z>;�`C;��E;*G;E�G;�H;�GH;BlH;ɈH;؞H;��H;��H;n�H;��H;��H;J�H;E�H;�H;H�H;H�H;��H;��H;k�H;��H;��H;ٞH;ɈH;BlH;�GH;�H;G�G;*G;��E;�`C;�Z>;�$5;�t%;�Y;Z��:5<:������Ǆ���׻���k�W�*X���뮼A�Ѽ}t�Iv���k�      Bm��Fi��&^�^�L�N�6�'����}ռlT����x���0���������Xط�o`:��:�;�*;!�8;�@;�D;I�F;�}G;�G;l1H;�[H;C|H;��H;��H;\�H;��H;��H;a�H;h�H;��H;E�H;��H;g�H;^�H;��H;��H;Z�H;��H;��H;C|H;�[H;k1H;z�G;�}G;I�F;�D;��@;&�8;�*;�;��:�n`:`ط��������껽�0���x�lT��}ռ��&��O�6�_�L��&^��Fi�      J��r;��@�������섽v�e��?��k�yt�鷼G���e7�����Ǆ�d0㺀�t�$u�:�+�:n;t1;I�<;N�B;�E;�G;��G;3H;NJH;3oH;֋H;��H;�H;k�H;��H;��H;i�H;��H;��H;��H;i�H;��H;��H;j�H;�H;��H;ڋH;3oH;MJH;3H;��G;�G;
�E;L�B;A�<;v1;l;�+�:$u�:��t�f0��Ǆ���껂e7�G��鷼zt��k��?�v�e��섽���@���r;��      n���$��s��ӽ�'��?������	�Z��Q+�����"��G����0���׻ĕb�2W���X�9ҡ�:`;�*';�Y7;�#@;�D;�F;��G;��G;8H;�aH;ЁH;6�H;}�H;H�H;l�H;{�H;W�H;&�H;�H;&�H;X�H;y�H;i�H;F�H;z�H;9�H;ҁH;�aH;8H;��G;�G;�F;
�D;�#@;�Y7;�*';`;ԡ�:Y�94W��ƕb���׻��0�G���"������Q+�
�Z����>����'���ӽ�s�$��      �!,�7)��K ��������޽������Fi��0����鷼��x�����.��M�(�����*i:z��:)�;��0;:�<;vC;��E;�<G;��G;�$H;:TH;�wH;ʒH;�H; �H;X�H;�H;c�H;q�H;O�H;q�H;d�H;�H;U�H;�H;�H;˒H;�wH;;TH;�$H;��G;�<G;��E;vC;8�<;��0;.�;x��:+i:���N�(��.�������x�鷼����0��Fi�������޽�������K �7)�      (�j��f��Z�x�F��>/��^�l�����ŽF ���Fi��Q+�yt�lT��l�W�����1��$ȺX�9yP�:�Y;��(;��8;�A;�E;��F;8�G;pH;�FH;�mH;m�H;��H;�H;H�H;��H;^�H;��H;��H;��H;`�H;��H;D�H;�H;��H;m�H;�mH;�FH;oH;;�G;��F;�E;�A;��8;��(;�Y;wP�:8X�9"Ⱥ�1�����l�W�lT��zt�Q+��Fi�F ����Žl����^��>/�x�F��Z��f�      ��v���x�G����f��SC��K �mn����Ž���
�Z��k�}ռ,X��_y-�(���k.�x��P�:�+�:��;4;�>;�D;�wF; �G;��G;�9H;&dH;T�H;��H;2�H;H�H;��H;~�H;+�H;E�H;)�H;�H;��H;E�H;/�H;��H;X�H;*dH;�9H;��G;�G;�wF;�D;�>;4;{�;�+�:�P�:P��i.�)���^y-�,X��}ռ�k�
�Z������Žmn���K ��SC��f�G���x�v���      ��˾��Ǿ�������U͓�Y�x���J��K �l���������?����뮼'�[����3|��W����:E�:�';b/;Cg<;�C;GF;�NG;��G;-H;;[H;�}H;��H;��H;��H;��H;��H;��H;��H;��H;��H;�H;��H;��H;��H;�}H;>[H;-H;��G;�NG;DF;�C;Cg<;a/;�';O�:��:�W��3|����'�[��뮼���?������l����K ���J�Z�x�U͓����������Ǿ      s� ��������{Ծj���v���Y�x��SC��^��޽?���w�e�'��B�Ѽ#G������R����� ޤ8χ�:�Y;E�);��9;��A;��E;G;
�G;@!H;	SH;�wH;N�H;Z�H;�H;��H;I�H;V�H;��H;V�H;K�H;��H;�H;Z�H;H�H;�wH;SH;C!H;
�G;�G;��E;��A;��9;E�);�Y;Ӈ�:�ݤ8����R�����#G��B�Ѽ'��w�e�?����޽�^��SC�Y�x�v���j����{Ծ�쾟���      ����D�l�s� �U�ݾj���U͓��f��>/�����'���섽N�6�}t�w��\�:�$Tʻy.� ۷�Jt�:�;��$;�Y7;T�@;�	E;��F;'�G;�H;LH;�rH;��H;��H;��H;��H;�H;%�H;��H;!�H;�H;�H;��H;��H;��H;�rH;
LH;�H;+�G;��F;�	E;S�@;�Y7;��$;�;Nt�:(۷�t.�$Tʻ\�:�w��}t�N�6��섽�'������>/��f�U͓�j���V�ݾs� �l��D�      �7�v3�/�'����s� ��{Ծ���H���y�F�����ӽ���^�L�Iv��뮼OT����PV���=�n)i:|��:�z ;�$5;��?;�D;��F;�G;rH;dFH;qnH;d�H;K�H;H�H;��H;	�H;1�H;��H;.�H;	�H;��H;J�H;M�H;`�H;znH;fFH;sH;�G;��F;�D;��?;}$5;�z ;z��:�)i:��=��PV���OT��뮼Iv�^�L�����ӽ���y�F�G�������{Ծs� ����/�'�v3�      �N��TI���;�/�'�l��쾀���x󐾴Z��K ��s�@����&^���"����g����̨u�� ���2<:#��:�
;<g3;��>;XBD;w�F;ܔG;kH;BH;\kH;/�H;��H;�H;��H;?�H;��H;"�H;��H;B�H;��H;�H;��H;)�H;ckH;BH;nH;�G;��F;WBD;��>;5g3;�
;��:�2<:� ��ʨu������g��"����&^�@����s潥K ��Z�x󐾀�����l�/�'���;��TI�      `]�d�W��TI�v3��D�������Ǿv����f�7)�$��r;���Fi��k���Ǽ�[t�L�	�(Ȅ�X���:��:��;.J2;VZ>;'	D;=F;8�G;�H;�?H;viH;ÈH;��H;Q�H;�H;��H;4�H;��H;1�H;��H;�H;P�H;��H;��H;{iH;�?H;�H;:�G;HF;%	D;QZ>;(J2;��;��:�:X��'Ȅ�L�	��[t���Ǽ�k��Fi�r;��$��7)��f�v�����Ǿ�����D�v3��TI�d�W�      �?��|h��=v��� ��6�X��O/�0y�@�;ఖ��+X��� �ѽ����^n;�Y�������B(�ך��N����e9!�:�;�Y.;W�<;eWC;�ZF;��G;�/H;1jH;8�H;F�H;�H;'�H;��H;W�H;��H;��H;��H;V�H;��H;%�H;�H;C�H;?�H;4jH;0H;��G;�ZF;fWC;S�<;�Y.;�;#�:�e9P��՚���B(�����Y��^n;����� �ѽ���+X�ఖ�@�;0y��O/�6�X�� ��=v��|h��      |h��/���a�����y�VvS�pM+��v�9ɾ�����T�]�\ν����w\8�����x��%�J���l�뺐�9x-�:k�;��.; �<;�nC;�dF;�G;�1H;�jH;��H;��H;ɵH;g�H;��H;b�H;��H;��H;��H;d�H;��H;f�H;ɵH;��H;��H;�jH;�1H;�G;�dF;�nC;�<;��.;j�;v-�:��9l��I���%��x�����w\8�����\ν]��T�����9ɾ�v�pM+�VvS���y�a���/���      =v��a���V ��`�h�6E�W��i���{㼾|���nH�҈�x�ý�Ȅ��s/��o��#����� J�� кx	�9[g�:�l;(0;!]=;ڲC;ـF;q�G;6H;mH;'�H;��H;|�H;��H;@�H;��H;�H;��H; �H;��H;=�H;��H;|�H;��H;,�H; mH;6H;p�G;�F;ڲC;]=; 0;�l;]g�:�	�9(к J������#���o��s/��Ȅ�x�ý҈��nH�|��{㼾i���W��6E�`�h�V ��a���      � ����y�`�h���N��O/����B�߾B���*|��6�p}�䳽hSt�;�!�nrμ?F{��_��X����X:0��:�Z;�2;�O>;oD;,�F;{�G;=H;�pH;��H;H�H;ɷH;��H;��H;[�H;z�H;\�H;v�H;[�H;��H;��H;ɷH;D�H;��H;�pH;=H;y�G;1�F;mD;�O>;�2;�Z;.��:t:ȓ���X���_�?F{�mrμ;�!�hSt�䳽p}��6��*|�B��B�߾����O/���N�`�h���y�      6�X�VvS�6E��O/��S�HW����������KS\��� ���9����Y�y��΃����]������b���Y�P�Y:��:f`;=�4;�?;;�D;��F;�G;FH;FuH;H;��H;��H;�H;��H;�H;�H;��H;�H;�H;��H;�H;�H;��H;ƓH;FuH;FH;�G;��F;;�D;�?;6�4;f`;��:`�Y:��Y��b�������]�΃��y���Y�9����彑� �LS\���������HW���S��O/�6E�VvS�      �O/�pM+�W�����HW��9ɾ@���Mw�� :�i��v�ý�L��[n;�\���qv���E<��˻��-���py�:�^;�%;��7;x�@;5E;�"G;�G;8PH;�zH;��H;X�H;x�H;��H;��H;	�H;��H;��H;��H;
�H;��H;��H;x�H;T�H;H;�zH;8PH;�G;�"G;5E;r�@;��7;�%;�^;vy�:����-��˻�E<�qv��[���Zn;��L��v�ýi��� :��Mw�@��9ɾHW�����W��pM+�      0y��v�i���B�߾����@��>����nH���B὜u����d�/O�grμH"�����	����뺐r89c;�:b�;�+;Y|:;{7B;��E;�aG;rH;�ZH;e�H;*�H;��H;�H;F�H;B�H;�H;��H;t�H;��H;�H;B�H;E�H;�H;��H;0�H;f�H;�ZH;kH;bG;��E;v7B;T|:;�+;`�;k;�:�r89���	�����H"��grμ.O���d��u��B����nH�?���@������B�߾i����v�      @�;9ɾ{㼾B�������Mw��nH�����Z�
䳽ʕ��p\8�l#������^N�I���b��Hx�P5:��:3�;��0;!]=;A�C;�[F;؞G;�)H;�eH;s�H;!�H;;�H;��H;�H;��H;'�H;��H;l�H;��H;+�H;��H;�H;��H;:�H;(�H;s�H;�eH;�)H;؞G;�[F;:�C;]=;��0;.�;��:H5:�Hx� �b�I��
^N�����l#��p\8�ʕ��
䳽�Z񽯯��nH��Mw�����B��{㼾9ɾ      ఖ�����|���*|�KS\�� :����Z�k$������ �K�u���Oļ����������:&����M/�:�^;��#;�G6;<�?;��D;I�F;��G;@H;�pH;��H;t�H;�H;I�H;.�H;j�H;n�H;��H;x�H;��H;q�H;k�H;,�H;K�H;�H;w�H;ޏH;�pH;@H;��G;H�F;��D;>�?;�G6;��#;�^;M/�:���8&������������Oļu�� �K�����k$���Z���� :�KS\��*|�|������      �+X��T��nH��6��� �i��B�
䳽�����mR����ټ�����E<��?ݻ.d\������ :�d�:��;*�,;|�:;\7B;��E;qLG;0H;\SH;�{H;|�H;�H;�H;<�H;R�H;�H;��H;��H;��H;��H;��H;�H;Q�H;:�H;�H;�H;��H;�{H;WSH;,H;qLG;��E;\7B;|�:;'�,;��;�d�: !:����.d\��?ݻ�E<�����
ټ����mR�����
䳽B�i���� ��6��nH��T�      ��]�ӈ�p}���v�ý�u��ɕ�� �K�����o�hv���&R���R^��p�� �>����:aB;<";i�4;��>;BD;��F;�G;�)H;gdH;r�H;�H;_�H;&�H;*�H;~�H;��H;�H;
�H;��H;�H;�H;��H;~�H;*�H;(�H;c�H;�H;r�H;fdH;�)H;�G;��F;DD;��>;i�4;D";dB;��: t>�r��Q^�����&R�gv���o���� �K�ɕ���u��v�ý��p}�ӈ�]�      ��ѽ\νx�ý䳽8����L����d�p\8�u��
ټgv����Y��_�����6���[���Y:]��:Lm;�r-;�:;p�A;-oE;�"G;K�G;XGH;�sH;�H;��H;�H;"�H;�H;��H;u�H;|�H;'�H;��H;'�H;~�H;{�H;��H;�H;&�H;�H;��H;�H;�sH;XGH;M�G;�"G;3oE;q�A;�:;�r-;Pm;c��:��Y:�[�4�������_���Y�gv��
ټt��p\8���d��L��9���䳽x�ý\ν      ���������Ȅ�iSt��Y�Zn;�.O�k#���Oļ�����&R��_������N3�ąY� 4:�:د;�?&;�G6;�X?;�D;'xF;��G;-!H;�^H;��H;�H;íH;;�H;��H;��H;��H;�H;��H;P�H;�H;P�H;��H;	�H;��H;��H;�H;E�H;ɭH;�H;��H;�^H;1!H;��G;)xF;�D;�X?;�G6;�?&;֯;�:4:��Y��N3������_��&R������Oļk#��.O�Zn;��Y�iSt��Ȅ�����      \n;�w\8��s/�;�!�x��]���frμ��������E<��������N3�4Hx���9��:�^;U ;*2;d�<;�B;��E;'5G;�G;*FH;|qH;��H;>�H;��H;F�H;��H;��H;��H;��H;�H;n�H;�H;n�H;�H;��H;��H;��H;��H;P�H;��H;A�H;��H;vqH;-FH;�G;+5G;��E;��B;l�<;.2;U ;�^;��:��9(Hx��N3��������E<��������grμ[���y��<�!��s/�v\8�      V������o�mrμ̓��qv��G"��^N�����?ݻP^��:��̅Y���9��:��:��;R�.;||:;�>A;��D;&�F;��G;�)H;aH;�H;u�H;۬H;,�H;�H;/�H;W�H;��H;�H;O�H;��H;��H;��H;N�H;�H;��H;V�H;2�H;�H;2�H;߬H;u�H;�H;aH;�)H;��G;)�F;��D;�>A;�|:;N�.;��;ަ�:��:��9��Y�6��O^���?ݻ���^N�G"��pv��΃��nrμ�o����      �����x���#��<F{���]��E<����D�뻤���)d\�l�뺤[��3:��:��:}[;d�,;��8;!@;�0D;r[F;{G;�
H;>PH;vH;ݐH;6�H;�H;�H;]�H;q�H;��H;��H;t�H;o�H;��H;��H;��H;m�H;s�H;��H;��H;t�H;c�H;#�H;��H;8�H;ԐH;vH;=PH;�
H;{G;v[F;�0D;!@;��8;i�,;{[;��:��:�3:�[�h��)d\�����D�뻟���E<���]�<F{��#���x��      �B(��%�����_�|����˻�����b�2&����� l>���Y:�:�^;��;i�,;
`8;c�?;��C;pF;�FG;B�G;�?H;kH;�H;��H;�H;L�H;��H;b�H;k�H;�H;u�H;��H;��H;}�H;��H;x�H;~�H;��H;p�H;�H;o�H;c�H;��H;O�H;�H;��H;��H; kH;�?H;C�G;�FG;wF;��C;\�?;`8;h�,;��;�^;�:��Y: `>�����/&���b� 	���˻����_�����%�      ǚ��C��� J���X���b���-�����Hx����!:��:W��:ү;T ;M�.;��8;X�?;��C;��E;.#G;��G;�1H;�aH;C�H;m�H;o�H;��H;��H;S�H;�H;(�H;0�H;��H;�H;��H;3�H;��H;0�H;~�H;�H;��H;-�H;,�H;�H;U�H;��H;��H;i�H;q�H;@�H;�aH;�1H;��G;1#G;��E;��C;\�?;��8;N�.;Q ;ѯ;Y��:��:!:@���Hx������-�
�b��X��J��D���      ����� к������Y����@s89d5:U/�:�d�:hB;Lm;�?&;02;�|:;!@;��C;��E;sG;��G;N(H;�ZH;czH;2�H;ʤH;��H;\�H;��H;��H;U�H;��H;��H;B�H;$�H;C�H;��H;u�H;��H;@�H;!�H;@�H;��H;��H;Z�H;��H;��H;Z�H;��H;ΤH;2�H;^zH;�ZH;R(H;��G;sG;��E;³C;!@;�|:;.2;�?&;Lm;iB;�d�:W/�:d5: s89�����Y�ʓ��"к���      ��e9��9�	�9�:L�Y:vy�:};�:��:�^;��;E";�r-;�G6;i�<;�>A;�0D;uF;7#G;��G;�$H;UWH;�vH;k�H;6�H;7�H;o�H;�H;��H;q�H;0�H;��H;x�H;��H;!�H;�H;��H;��H;��H;�H; �H;��H;u�H;��H;0�H;o�H;��H;�H;n�H;<�H;6�H;g�H;�vH;WWH;�$H;��G;3#G;tF;�0D;�>A;e�<;�G6;�r-;G";��;�^;��:w;�:�y�:\�Y:`:�	�90�9      Y�:Z-�:%g�:��:��:�^;a�;-�;��#;)�,;g�4;�:;X?;�B;��D;w[F;�FG;��G;Q(H;SWH;_uH;��H;�H;�H;�H;��H;��H;��H;��H;��H;��H;��H;��H;��H;��H;Q�H;L�H;J�H;��H;��H;��H;��H;��H;��H;��H;��H;��H;��H;�H;�H;	�H;��H;buH;UWH;R(H;��G;�FG;u[F;��D;�B;�X?;�:;l�4;'�,;��#;*�;e�;�^;��: ��:Ag�:X-�:      �;u�;�l;[;f`;�%;�+;��0;�G6;�:;��>;p�A;�D;��E;)�F;{G;G�G;�1H;�ZH;�vH;��H;@�H;��H;ŸH;~�H;M�H;��H;��H;��H;��H;3�H;4�H;��H;��H;d�H;��H;��H;��H;a�H;��H;��H;.�H;4�H;��H;��H;��H;��H;K�H;��H;øH;��H;A�H;��H;�vH;�ZH;�1H;I�G;{G;)�F;��E;�D;p�A;��>;|�:;�G6;��0;�+;�%;x`;�Z;�l;m�;      �Y.;��.;0;�2;2�4;��7;e|:;(]=;B�?;`7B;HD;2oE;*xF;55G;��G;�
H;�?H;�aH;czH;i�H;�H;��H;C�H;��H;\�H;��H;��H;��H;�H;��H;��H;X�H;R�H;?�H;��H;�H;?�H;�H;��H;A�H;N�H;U�H;��H;��H;�H;��H;��H;��H;a�H;��H;>�H;��H;�H;j�H;ezH;�aH;�?H;�
H;��G;/5G;*xF;4oE;ID;Z7B;F�?;+]=;`|:;��7;A�4;�2;0;��.;      V�<;)�<;]=;�O>;�?;{�@;}7B;@�C;�D;��E;��F;�"G;��G;�G;�)H;BPH;!kH;H�H;2�H;5�H;�H;��H;��H;2�H;*�H;-�H;?�H;��H;�H;5�H;��H;
�H;�H;��H;?�H;{�H;��H;t�H;<�H;��H;�H;�H;��H;3�H;�H;��H;;�H;0�H;-�H;.�H;��H;¸H;�H;2�H;0�H;C�H;"kH;APH;�)H; �G;��G;�"G;��F;��E;��D;F�C;y7B;h�@;�?;�O>;]=; �<;      �WC;�nC;ӲC;fD;7�D;$5E;��E;�[F;K�F;uLG;��G;R�G;1!H;4FH;aH;vH;��H;y�H;ؤH;C�H;�H;��H;c�H;6�H;��H; �H;;�H;��H;��H;��H;��H;��H;��H;1�H;��H;��H;��H;��H;��H;/�H;��H;��H;��H;��H;��H;��H;6�H;��H;��H;2�H;a�H;��H;�H;>�H;פH;v�H; �H;vH;aH;1FH;3!H;U�G;��G;tLG;N�F;�[F;��E;5E;B�D;lD;ӲC;�nC;      �ZF;�dF;��F;'�F;��F;�"G;bG;��G;��G;5H;�)H;\GH;�^H;�qH;	�H;ސH;��H;p�H;��H;n�H;��H;G�H;��H;3�H;��H;�H;��H;��H;h�H;��H;��H;��H; �H;t�H;��H;�H;�H;�H;��H;t�H; �H;��H;��H;��H;c�H;��H;��H;!�H;��H;-�H;��H;J�H;��H;l�H;��H;l�H;��H;ߐH;	�H;}qH;�^H;^GH;�)H;3H;��G;�G;bG;�"G;��F;3�F;݀F;�dF;      �G;�G;j�G;}�G;�G;	�G;zH;�)H;�?H;ZSH;gdH;�sH;��H;��H;t�H;9�H;�H;��H;`�H;�H;��H;��H;��H;E�H;9�H;��H;��H;=�H;~�H;��H;^�H;��H;p�H;��H;�H;6�H;Q�H;/�H;��H;��H;o�H;��H;[�H;��H;x�H;8�H;�H;��H;;�H;>�H;��H;��H;��H;�H;]�H;��H;�H;9�H;t�H;��H;��H;�sH;hdH;YSH;@H;�)H;tH;�G;�G;t�G;k�G;ܪG;      0H;�1H;6H;=H;�EH;7PH;�ZH;�eH;�pH;�{H;t�H;�H;�H;E�H;ڬH;��H;M�H;��H;��H;��H;��H;��H;��H;��H;��H;��H;9�H;u�H;\�H;J�H;��H;b�H;��H;	�H;A�H;V�H;A�H;R�H;@�H;�H;��H;^�H;��H;I�H;W�H;q�H;5�H;��H;��H;��H;��H;��H;��H;��H;��H;��H;L�H;��H;۬H;C�H;�H;�H;x�H;�{H;�pH;�eH;�ZH;-PH;
FH;=H;6H;�1H;      *jH;�jH;mH;�pH;5uH;�zH;j�H;o�H;֏H;}�H;
�H;��H;ɭH;��H;-�H;$�H;��H;Y�H;��H;r�H;��H;��H;�H;�H;��H;e�H;x�H;]�H;S�H;��H;M�H;��H;��H;0�H;`�H;g�H;X�H;c�H;]�H;2�H;��H;��H;N�H;��H;M�H;Y�H;q�H;c�H;��H;�H;�H;��H;��H;o�H;��H;W�H;��H;&�H;-�H;��H;ʭH;��H;�H;��H;ڏH;s�H;h�H;�zH;DuH;�pH;mH;�jH;      7�H;��H;0�H;��H;ēH;��H;-�H;#�H;u�H;�H;b�H;�H;B�H;P�H;�H;`�H;i�H;�H;S�H;.�H;��H;��H;��H;3�H;��H;��H;��H;I�H;��H;C�H;��H;��H;0�H;Y�H;d�H;z�H;��H;x�H;b�H;X�H;,�H;��H;��H;@�H;��H;I�H;}�H;��H;��H;.�H;��H;��H;��H;-�H;T�H;�H;f�H;c�H;�H;N�H;C�H;�H;f�H;�H;w�H;'�H;1�H;��H;ƓH;��H;0�H;��H;      J�H;��H;��H;I�H;��H;W�H;��H;>�H;�H;�H;/�H;-�H;�H;��H;5�H;x�H;v�H;2�H;��H;��H;��H;6�H;��H;��H;��H;��H;^�H;��H;S�H;��H;��H;$�H;[�H;i�H;��H;��H;{�H;~�H;�H;j�H;Y�H;"�H;��H;��H;M�H;��H;Z�H;��H;��H;��H;��H;6�H;��H;��H;��H;0�H;v�H;z�H;6�H;��H;
�H;0�H;0�H;�H;�H;D�H;��H;M�H;��H;I�H;��H;��H;      ��H;ѵH;~�H;ȷH;}�H;o�H;��H;��H;P�H;<�H;.�H;�H;��H;��H;X�H;��H;�H;6�H;��H;~�H;��H;5�H;V�H;�H;��H;��H;��H;c�H;��H;��H;�H;<�H;d�H;��H;��H;��H;��H;��H;��H;��H;d�H;:�H;�H;��H;��H;a�H;��H;��H;��H;�H;Y�H;6�H;��H;{�H;��H;7�H;�H;��H;X�H;��H;��H;�H;4�H;?�H;P�H;��H;��H;q�H;��H;ɷH;��H;εH;      ,�H;p�H;	�H;��H;�H;��H;H�H;�H;)�H;T�H;��H;��H;��H;��H;��H;��H;z�H;��H;K�H;��H;��H;��H;R�H;�H;��H;�H;q�H;��H;��H;3�H;V�H;f�H;z�H;��H;��H;��H;��H;��H;��H;��H;w�H;f�H;U�H;/�H;��H;��H;m�H; �H;��H;�H;U�H;��H;��H;��H;K�H;��H;}�H;��H;��H;��H;��H;��H;��H;U�H;-�H;�H;H�H;~�H; �H;��H;�H;r�H;      ��H;��H;>�H;��H;��H;��H;I�H;��H;n�H;�H;��H;�H;�H;��H;�H;x�H;��H;�H;*�H;)�H;��H;��H;?�H;��H;-�H;q�H;��H;�H;0�H;[�H;c�H;��H;��H;��H;��H;��H;��H;��H;��H;��H;��H;��H;c�H;X�H;,�H;�H;��H;s�H;/�H;��H;E�H;��H;��H;"�H;(�H;�H;��H;z�H;�H;��H;�H;�H;��H;�H;q�H;��H;N�H;��H;��H;��H;H�H;��H;      P�H;u�H;��H;b�H;+�H;�H;�H;-�H;u�H;��H;$�H;��H;��H;�H;V�H;r�H;��H;��H;D�H;
�H;��H;d�H;��H;5�H;��H;��H;��H;@�H;b�H;g�H;{�H;��H;��H;��H;��H;��H;��H;��H;��H;��H;��H;��H;z�H;b�H;[�H;<�H;��H;��H;��H;5�H;��H;b�H;��H;�H;D�H;��H;��H;v�H;X�H;�H;��H;��H;'�H;��H;z�H;/�H;�H;�H;,�H;c�H;��H;v�H;      ��H;��H;�H;w�H;�H;��H;��H;��H;��H;��H;�H;,�H;Q�H;r�H;��H;��H;~�H;2�H;��H;��H;V�H;��H;�H;l�H;��H;�H;0�H;U�H;k�H;�H;~�H;��H;��H;��H;��H;��H;��H;��H;��H;��H;��H;��H;|�H;z�H;f�H;Q�H;/�H;�H;��H;o�H;�H;��H;P�H;��H;��H;7�H;��H;��H;��H;t�H;S�H;*�H;�H;��H;��H;��H;��H;��H;�H;v�H;�H;��H;      ��H;��H;��H;^�H;��H;��H;y�H;l�H;}�H;��H;��H;��H;�H;�H;��H;��H;��H;��H;{�H;��H;W�H;��H;B�H;��H;��H;�H;M�H;H�H;_�H;��H;w�H;��H;��H;��H;��H;��H;��H;��H;��H;��H;��H;��H;w�H;��H;X�H;C�H;M�H;	�H;��H;��H;F�H;��H;P�H;��H;{�H;��H;��H;��H;��H;�H;�H;��H;��H;��H;�H;r�H;��H;��H;��H;_�H;��H;��H;      ��H;��H;��H;y�H;�H;��H;��H;��H;��H;��H;�H;,�H;T�H;u�H;��H;��H;�H;3�H;��H;��H;W�H;��H;�H;l�H;��H;�H;0�H;U�H;m�H;~�H;~�H;��H;��H;��H;��H;��H;��H;��H;��H;��H;��H;��H;|�H;x�H;f�H;O�H;.�H;�H;��H;m�H;�H;��H;P�H;��H;��H;7�H;��H;��H;��H;r�H;T�H;*�H;�H;��H;��H;��H;��H;��H;�H;z�H;�H;��H;      F�H;w�H;��H;[�H;)�H;��H;�H;/�H;u�H;��H;$�H;��H;��H;�H;X�H;t�H;��H;��H;D�H;
�H;��H;d�H;��H;4�H;��H;��H;��H;@�H;`�H;f�H;z�H;��H;��H;��H;��H;��H;��H;��H;��H;��H;��H;��H;z�H;`�H;[�H;9�H;��H;��H;��H;4�H;��H;d�H;��H;�H;D�H;��H;��H;v�H;V�H;�H;��H;��H;$�H;��H;w�H;4�H;�H;��H;0�H;\�H;��H;y�H;      ��H;��H;;�H;��H;��H;��H;G�H;��H;p�H;�H;��H;�H;�H;��H;�H;z�H;��H;�H;*�H;(�H;��H;��H;>�H;��H;.�H;o�H;��H;�H;0�H;[�H;c�H;��H;��H;��H;��H;��H;��H;��H;��H;��H;��H;��H;b�H;X�H;)�H;�H;��H;s�H;.�H;��H;E�H;��H;��H;$�H;*�H;�H;��H;}�H;�H;��H;�H;�H;��H;�H;r�H;��H;O�H;��H;��H;��H;D�H;��H;      ,�H;x�H;�H;��H;�H;��H;E�H;�H;*�H;T�H;��H;��H;��H;��H;��H;��H;}�H;��H;I�H;��H;��H;��H;N�H;�H;��H;�H;m�H;��H;��H;3�H;U�H;c�H;x�H;��H;��H;��H;��H;��H;��H;��H;w�H;f�H;U�H;.�H;��H;��H;m�H;�H;��H;��H;V�H;��H;��H;��H;H�H;��H;|�H;��H;��H;��H;��H;��H;��H;R�H;,�H;�H;M�H;�H;�H;��H;�H;p�H;      v�H;ԵH;q�H;·H;{�H;�H;��H;��H;O�H;<�H;/�H;�H;��H;��H;[�H;��H;�H;7�H;��H;|�H;��H;6�H;U�H;�H;��H;��H;��H;c�H;��H;��H;�H;:�H;f�H;�H;��H;��H;��H;��H;��H;��H;d�H;:�H;�H;��H;��H;^�H;��H;��H;��H;�H;\�H;6�H;��H;z�H;��H;4�H;�H;��H;Z�H;��H;��H;�H;/�H;?�H;R�H;��H;��H;r�H;�H;ŷH;w�H;εH;      ?�H;��H;��H;D�H;��H;W�H;��H;@�H;�H;�H;-�H;0�H;�H;��H;6�H;z�H;w�H;0�H;��H;��H;��H;7�H;��H;��H;��H;��H;X�H;��H;S�H;��H;��H;$�H;[�H;i�H;��H;�H;{�H;��H;�H;j�H;\�H;$�H;��H;��H;L�H;��H;X�H;��H;��H;��H;��H;9�H;��H;��H;��H;0�H;w�H;z�H;7�H;��H;�H;/�H;-�H;�H;�H;D�H;��H;T�H;��H;P�H;��H;��H;      H�H;��H;,�H;��H;��H;ƗH;,�H;+�H;x�H;�H;b�H;�H;C�H;N�H;�H;b�H;g�H;�H;S�H;.�H;��H;��H;��H;0�H;��H;��H;��H;I�H;��H;B�H;��H;��H;+�H;Y�H;d�H;x�H;��H;z�H;b�H;Y�H;/�H;��H;��H;@�H;��H;F�H;�H;��H;��H;-�H;��H;��H;��H;-�H;U�H;�H;f�H;b�H;�H;N�H;B�H;�H;e�H;�H;u�H;*�H;0�H;��H;ɓH;��H;=�H;��H;      ;jH;�jH;,mH;�pH;.uH; {H;f�H;r�H;ޏH;}�H;�H;��H;ʭH;��H;2�H;&�H;��H;\�H;��H;o�H;��H;��H;�H;�H;��H;^�H;r�H;Z�H;Q�H;��H;L�H;��H;��H;0�H;_�H;f�H;X�H;f�H;]�H;0�H;��H;��H;N�H;��H;M�H;V�H;t�H;e�H;��H;�H;�H;��H;��H;q�H;��H;W�H;��H;'�H;2�H;��H;ɭH;��H;�H;|�H;��H;u�H;j�H;�zH;>uH;�pH;,mH;�jH;      0H;�1H;6H;=H;�EH;FPH;�ZH;�eH;�pH;�{H;w�H;�H;�H;E�H;ݬH;��H;M�H;��H;��H;��H;��H;��H;��H;��H;��H;��H;5�H;r�H;\�H;E�H;��H;a�H;��H;�H;?�H;T�H;C�H;U�H;?�H;�H;��H;a�H;��H;H�H;W�H;p�H;5�H;��H;��H;��H;��H;��H;��H;��H;��H;��H;O�H;��H;ݬH;B�H;�H;�H;x�H;�{H;�pH;�eH;�ZH;1PH;FH;=H;6H;�1H;      �G;��G;m�G;��G;�G;�G;{H;�)H;@H;ZSH;jdH;�sH;��H;��H;u�H;;�H;�H;��H;]�H;�H;��H;��H;��H;C�H;9�H;��H;�H;9�H;|�H;��H;Z�H;��H;m�H;��H;�H;2�H;O�H;2�H;��H;��H;q�H;��H;^�H;��H;z�H;8�H;�H;��H;:�H;A�H;��H;��H;��H;�H;^�H;��H;�H;<�H;w�H;��H;��H;�sH;hdH;YSH;@H;�)H;H;�G;�G;��G;q�G;�G;      �ZF;�dF;�F;%�F;��F;�"G;�aG;�G;��G;6H;�)H;bGH;�^H;qH;�H;ߐH;��H;q�H;��H;n�H;��H;G�H;��H;0�H;��H;�H;��H;��H;h�H;��H;��H;��H;�H;s�H;��H;�H;�H;�H;��H;t�H;�H;��H;��H;��H;c�H;��H;��H;!�H;��H;0�H;��H;H�H;��H;l�H;��H;l�H;��H;ߐH;�H;}qH;�^H;\GH;�)H;5H;��G;ߞG;�aG;�"G;��F;'�F;ЀF;�dF;      �WC;�nC;ӲC;jD;5�D;*5E;��E;�[F;P�F;uLG;��G;U�G;3!H;2FH;aH;vH;��H;y�H;פH;?�H;�H;��H;_�H;3�H;��H;��H;6�H;��H;��H;��H;��H;��H;��H;/�H;��H;��H;��H;��H;��H;2�H;��H;��H;��H;��H;��H;��H;:�H; �H;��H;3�H;e�H;��H;�H;A�H;ؤH;u�H;��H;vH;aH;2FH;4!H;R�G;��G;tLG;L�F;�[F;��E;5E;@�D;hD;ҲC;�nC;      8�<;�<;]=;�O>;߁?;��@;7B;D�C;��D;��E;��F;�"G;��G;�G;�)H;DPH;"kH;J�H;0�H;2�H;�H;��H;��H;/�H;-�H;'�H;:�H;��H;�H;1�H;��H;
�H;�H;��H;=�H;x�H;��H;z�H;<�H;��H;�H;�H;��H;5�H;�H;��H;?�H;.�H;,�H;2�H;��H;��H;�H;5�H;3�H;D�H;$kH;BPH;�)H;�G;��G;�"G;��F;��E;��D;<�C;{7B;x�@;��?;�O>;]=;��<;      �Y.;��.;0;�2;1�4;��7;_|:;+]=;G�?;_7B;ED;4oE;*xF;25G;��G;�
H;�?H;�aH;dzH;g�H;�H;��H;>�H;��H;a�H;��H;��H;��H;�H;��H;��H;V�H;N�H;?�H;��H;�H;B�H;�H;��H;>�H;R�H;Y�H;��H;��H;�H;��H;��H;��H;^�H;��H;B�H;��H;�H;k�H;ezH;�aH;�?H;�
H;��G;/5G;*xF;2oE;ED;]7B;E�?;+]=;^|:;��7;1�4;�2;0;��.;      �;u�;�l;�Z;d`;�%;�+;��0;�G6;}�:;��>;t�A;�D;��E;,�F;{G;G�G;�1H;�ZH;�vH;��H;A�H;��H;øH;��H;G�H;��H;��H;��H;��H;3�H;2�H;��H;��H;a�H;��H;��H;��H;a�H;��H;��H;4�H;9�H;��H;��H;��H;��H;K�H;�H;ƸH;��H;A�H;��H;�vH;�ZH;�1H;G�G;{G;*�F;��E;�D;n�A;��>;|�:;�G6;��0;�+;�%;|`;�Z;�l;h�;      M�:�-�:Mg�:.��:��:�^;b�;0�;��#;'�,;l�4;�:;�X?;�B;��D;w[F;�FG;��G;Q(H;SWH;_uH;��H;
�H;�H;�H;��H;��H;��H;��H;��H;��H;��H;��H;��H;��H;M�H;M�H;O�H;��H;��H;��H;��H;��H;��H;��H;��H;��H;��H;�H;�H;�H;��H;buH;VWH;R(H;��G;�FG;u[F;��D;�B;�X?;�:;l�4;)�,;��#;3�;g�;�^;��:4��:_g�:\-�:       �e9��9�	�9�:P�Y:�y�:�;�:��:�^;��;J";�r-;�G6;i�<;�>A;�0D;tF;5#G;��G;�$H;WWH;�vH;i�H;5�H;<�H;l�H;��H;��H;n�H;*�H;��H;w�H;��H;"�H;�H;��H;��H;��H;�H;�H;��H;x�H;��H;-�H;q�H;��H;�H;o�H;8�H;;�H;m�H;�vH;WWH;�$H;��G;4#G;tF;�0D;�>A;e�<;�G6;�r-;H";��;�^;��:y;�:ry�:h�Y:t:�	�9x�9      �����"к������Y���� s89l5:]/�:�d�:iB;Mm;�?&;02;�|:; !@;��C;��E;rG;��G;Q(H;�ZH;czH;0�H;ΤH;��H;W�H;��H;��H;S�H;��H;��H;A�H;$�H;D�H;��H;u�H;��H;C�H;#�H;A�H;��H;��H;X�H;��H;��H;\�H;��H;ʤH;5�H;dzH;�ZH;Q(H;��G;sG;��E;��C;!@;�|:;-2;�?&;Lm;hB;�d�:[/�:l5: s89�����Y�����,кz��      Ϛ��?���"J���X��	�b���-���뺴Hx� ��!:��:Y��:ӯ;R ;R�.;��8;[�?;��C;��E;0#G;��G;�1H;�aH;A�H;q�H;j�H;��H;��H;U�H;�H;*�H;-�H;��H;�H;�H;2�H;��H;3�H;}�H;�H;��H;/�H;,�H;�H;U�H;��H;��H;l�H;m�H;C�H;�aH;�1H;��G;3#G;��E;��C;Z�?;��8;R�.;P ;ү;Y��:��:!:0���Hx������-��b��X��%J��@���      �B(� %�����_�|����˻�����b�1&����� `>���Y:�:�^;��;l�,;`8;_�?;��C;sF;�FG;C�G;�?H; kH;��H;��H;�H;J�H;��H;]�H;l�H;�H;s�H;��H;��H;{�H;��H;{�H;~�H;��H;r�H;�H;o�H;c�H;��H;J�H;�H;��H;��H;!kH;�?H;C�G;�FG;wF;��C;^�?;`8;k�,;��;�^;�:��Y: h>�����.&���b� 	���˻�����_�����%�      �����x���#��<F{���]��E<����C�뻣���)d\�h�뺐[� 4:��:��:�[;e�,;��8;!@;�0D;w[F;{G;�
H;?PH;vH;ېH;4�H;�H; �H;]�H;q�H;��H;��H;t�H;o�H;��H;��H;��H;m�H;s�H;��H;��H;s�H;`�H;!�H;��H;4�H;ڐH;vH;>PH;�
H;{G;r[F;�0D;!@;��8;f�,;}[;��:��:�3:�[�j��+d\�����D�뻠���E<���]�<F{��#���x��      W������o�mrμ̓��pv��G"��^N�����?ݻP^��9����Y���9��:��:��;O�.;|:;�>A;��D;&�F;��G;�)H;aH;�H;p�H;۬H;/�H;�H;2�H;V�H;��H;�H;O�H;��H;��H;��H;O�H;�H;��H;T�H;0�H;�H;2�H;ݬH;q�H;	�H;aH;�)H;��G;)�F;��D;�>A;~|:;N�.;��;ަ�:��:��9ȅY�9��P^���?ݻ���^N�G"��pv��΃��nrμ�o����      \n;�v\8��s/�;�!�x��\���grμ��������E<��������N3�(Hx��9�:�^;T ;-2;e�<;��B;��E;)5G;�G;.FH;|qH;��H;>�H;��H;I�H;��H;��H;��H;��H;�H;m�H;�H;p�H;�H;��H;��H;��H;��H;M�H;��H;A�H;��H;xqH;)FH;�G;/5G;��E;�B;k�<;)2;T ;�^;��:��90Hx��N3��������E<��������grμ[���y��;�!��s/�v\8�      ���������Ȅ�hSt��Y�Zn;�.O�k#���Oļ�����&R��_������N3���Y�4:�:կ;�?&;�G6;�X?;�D;*xF;��G;1!H;�^H;��H;�H;ǭH;?�H;�H;��H;��H;�H;��H;P�H;�H;P�H;��H;	�H;��H;��H; �H;A�H;ɭH;�H;��H;�^H;,!H;��G;+xF;�D;~X?;�G6;�?&;ӯ;�: 4:��Y��N3������_��&R������Oļk#��.O�Zn;��Y�iSt��Ȅ�����       �ѽ\νx�ý䳽8����L����d�o\8�t��
ټgv����Y��_�����4���[���Y:U��:Mm;�r-;�:;p�A;2oE;�"G;N�G;YGH;�sH;�H;��H;�H;(�H;�H;��H;y�H;~�H;&�H;��H;'�H;|�H;v�H;��H;�H;#�H;�H;��H;�H;�sH;XGH;J�G;�"G;3oE;p�A;
�:;�r-;Im;Y��:��Y:�[�4�������_���Y�gv��
ټt��p\8���d��L��9���䳽x�ý\ν      ��]�ӈ�p}���v�ý�u��ɕ�� �K�����o�hv���&R���P^��p�� �>����:_B;A";m�4;��>;HD;��F;�G;�)H;cdH;q�H;	�H;a�H;)�H;-�H;��H;��H;�H;�H;��H;�H;�H;��H;}�H;(�H;%�H;a�H;�H;q�H;adH;�)H;�G;��F;GD;��>;e�4;@";^B;��: |>�r��R^�����&R�hv���o���� �K�ɕ���u��v�ý��p}�ӈ�]�      �+X��T��nH��6��� �i��B�
䳽�����mR����
ټ�����E<��?ݻ-d\������ :�d�:��;-�,;z�:;`7B;��E;qLG;/H;WSH;�{H;�H;�H;�H;:�H;R�H;�H;��H;��H;��H;��H;��H;
�H;O�H;9�H;�H;�H;��H;�{H;VSH;/H;nLG;��E;_7B;z�:;$�,;��;�d�: !:����.d\��?ݻ�E<�����ټ����mR�����
䳽B�i���� ��6��nH��T�      ఖ�����|���*|�KS\�� :����Z�k$������ �K�u���Oļ����������8&����I/�:�^;��#;�G6;>�?;��D;K�F;��G; @H;�pH;��H;u�H;�H;I�H;0�H;m�H;p�H;��H;z�H;��H;p�H;j�H;,�H;I�H;�H;u�H;�H;�pH;�?H;��G;I�F;��D;?�?;�G6;��#;�^;G/�:���8&������������Oļu�� �K�����k$���Z���� :�LS\��*|�|������      @�;9ɾ{㼾B�������Mw��nH�����Z�
䳽ʕ��p\8�l#������^N�H���b��Hx�P5:��:3�;��0;$]=;C�C;�[F;՞G;�)H;�eH;r�H;#�H;=�H;��H;�H;��H;(�H;��H;l�H;��H;*�H;��H;�H;~�H;;�H;'�H;u�H;�eH;�)H;ٞG;�[F;A�C;!]=;��0;.�;��:H5:�Hx���b�I��
^N�����l#��p\8�ʕ��
䳽�Z񽰯��nH��Mw�����B��{㼾9ɾ      0y��v�i���B�߾����@��>����nH���B὜u����d�/O�grμH"�����	����뺐r89i;�:d�;�+;W|:;|7B;��E;�aG;mH;�ZH;e�H;,�H;��H;�H;H�H;E�H;�H;��H;t�H;��H;�H;D�H;E�H;�H;��H;.�H;f�H;�ZH;nH;bG;��E;{7B;X|:;�+;`�;o;�:pr89��� 	�����H"��grμ/O���d��u��B����nH�?���@������B�߾i����v�      �O/�pM+�W�����HW��9ɾ@���Mw�� :�i��v�ý�L��Zn;�\���qv���E<��˻��-� ��ry�:�^;�%;��7;y�@;5E;�"G;�G;7PH;�zH;��H;Z�H;y�H;��H;��H;	�H;��H;��H;��H;
�H;��H;��H;y�H;V�H;��H;�zH;:PH;�G;�"G;5E;y�@;��7;�%;�^;xy�:����-��˻�E<�qv��[���Zn;��L��v�ýi��� :��Mw�@��9ɾHW�����W��pM+�      6�X�VvS�6E��O/��S�HW����������KS\��� ���9����Y�y��΃����]������b���Y�\�Y:��:f`;<�4;�?;<�D;��F;�G;FH;CuH;��H;��H;�H;�H;��H;�H;�H;��H;�H;�H;��H;�H;�H;��H;ƓH;GuH;FH;�G;��F;9�D;�?;8�4;f`;��:`�Y:��Y��b�������]�΃��z���Y�9����彑� �LS\���������HW���S��O/�6E�VvS�      � ����y�`�h���N��O/����B�߾B���*|��6�p}�䳽hSt�;�!�mrμ?F{��_��X����`:4��:�Z;�2;�O>;oD;'�F;v�G;=H;�pH;��H;I�H;ɷH;��H;��H;[�H;z�H;^�H;w�H;[�H;��H;��H;˷H;G�H;��H;�pH;=H;z�G;1�F;mD;�O>;�2;�Z;0��:x:ȓ���X���_�>F{�mrμ;�!�hSt�䳽p}��6��*|�B��B�߾����O/���N�`�h���y�      =v��b���V ��`�h�6E�W��j���{㼾|���nH�҈�x�ý�Ȅ��s/��o��#�����!J��"к�	�9]g�:�l;'0;!]=;ܲC;׀F;m�G;6H;mH;'�H;��H;~�H;��H;>�H;��H;�H;��H;�H;��H;>�H;��H;|�H;��H;,�H; mH;6H;q�G;�F;ܲC;]=; 0;�l;]g�:�	�9"к J������#���o��s/��Ȅ�x�ý҈��nH�|��{㼾j���W��6E�`�h�W ��b���      |h��/���b�����y�VvS�pM+��v�9ɾ�����T�]�\ν����w\8�����x��%�J���h�뺘�9v-�:k�;��.; �<;�nC;�dF;�G;�1H;�jH;��H;��H;ʵH;g�H;��H;d�H;��H;��H;��H;e�H;��H;f�H;ʵH;��H;��H;�jH;�1H;�G;�dF;�nC;�<;��.;j�;v-�:��9n��I���%��x�����w\8�����\ν]��T�����9ɾ�v�pM+�VvS���y�a���/���      dܿ2�ֿ�aǿ=^��/���Xo���7����iþ�(���-=��` �
A���_�0]�-p����I�N�ѻ~�)� �R���:2�
;�*;$�:;��B;�HF;'�G;�lH;�H;t�H;=�H;��H;}�H;M�H;|�H;�H;��H;�H;|�H;L�H;{�H;��H;<�H;|�H;��H;�lH;*�G;IF;��B; �:;�*;0�
;��:��R�~�)�L�ѻ��I�-p��0]��_�
A���` ��-=��(���iþ����7�Xo�/���=^���aǿ2�ֿ      2�ֿCpѿ�¿������_Xi�ϕ3��
�UD��Fl��A�9�.���R��\� �cx��.�E��ͻ�$�� �㍨:@�;P�*;6�:;�B;�TF;��G;(nH;��H;��H;k�H;��H;��H;[�H;�H; �H;��H;�H;��H;Z�H;��H;��H;g�H;ŷH;��H;)nH;��G;�TF;�B;4�:;H�*;>�;卨:� ��$��ͻ.�E�cx�� �\��R��.��A�9�El��UD���
�ϕ3�_Xi��������¿Cpѿ      �aǿ�¿����������"Y��f'�����6o���.}��k/����#ڟ� <Q�,#�ע��(;�*���4�� a7��:��;v,;��;;�C;�vF;�G;�rH;�H;��H;�H;��H;��H;��H;��H;M�H;��H;F�H;��H;��H;��H;��H;�H;��H; �H;�rH;�G;wF;�C;��;;o,;�;�: ]7�6��(����(;�ע�,#� <Q�#ڟ�����k/��.}�6o�������f'��"Y�����������¿      =^������k���Xo���@�(�#�޾����9ce�/����ڽ󻒽�f@������R���O*�FG��
����C^94��:;`d.;�<;��C;��F;��G;�yH;��H;�H;�H;��H;i�H;��H;��H;��H;�H;{�H;��H;��H;h�H;��H;�H;�H;��H;�yH;��G;��F;��C;��<;Yd.;;2��:0D^9���DG���O*��R�������f@�󻒽��ڽ/��9ce�����#�޾(���@�Xo�k�������      /����������Xo��!J�K�#��\��UD������zPH�����b��C��� +���ټ'����运����t�:,��:G�;�Y1;>;�0D;�F;aH;F�H;ĨH;�H;[�H;��H;�H;b�H;H�H;��H;_�H;��H;I�H;a�H;	�H;��H;W�H;�H;ŨH;E�H;aH;��F;�0D;>;�Y1;G�;(��:��:���运���'����ټ� +�C���b�����zPH�����UD���\��K�#��!J�Xo��������      Xo�_Xi��"Y���@�K�#��
��о�A���i���(�}��tr��
�_��5��ɺ�n�`��<��^�d�P�\�d�X:�P�:�`;α4;��?;��D;x8G;m0H;��H;m�H;r�H;�H;��H;��H;��H;��H;�H;��H;�H;��H;��H;��H;��H;�H;w�H;m�H;��H;j0H;|8G;��D;��?;ȱ4;�`;�P�:d�X:T�\�]�d��<��n�`��ɺ��5�
�_�tr��}����(��i��A���о�
�K�#���@��"Y�_Xi�      ��7�ϕ3��f'�(��\���о�����.}��-=�{
���Ľ[��*:�����������7� GĻ��$��N��ǿ�:�{;�D&;�+8;JA;�E;��G;}LH;�H;u�H;2�H;��H;��H;��H;��H;�H;��H;�H;~�H;�H;��H;��H;��H;��H;6�H;x�H;�H;wLH;��G;�E;JA;�+8;�D&;�{;Ϳ�: O����$�GĻ��7���������*:�[����Ľ{
��-=��.}������о�\��(��f'�ϕ3�      ���
�����#�޾VD���A���.}�(�D�ht���ڽ�!��\����Y�ļ�
v�;��ſ���Iɺ(S�9���:(;�-;��;;��B;iIF;��G;fH;��H;�H;,�H;��H;c�H;��H;Z�H;��H;��H;g�H;��H;��H;\�H;��H;c�H;��H;1�H;�H;��H;fH;��G;iIF;��B;��;;�-;(;���:S�9�IɺĿ��:���
v�Y�ļ���\��!����ڽht�(�D��.}��A��VD��#�޾�����
�      �iþUD��6o�����������i��-=�ht�����R��gys�y +����v񗼑(;�&�ѻ�s@�ą!�4j:�P�:��;�D3;5�>;FD;��F;�	H;;|H;��H;q�H;4�H;��H;��H;��H;�H;.�H;n�H;��H;m�H;/�H;�H;��H;��H;��H;7�H;t�H;��H;:|H;�	H;��F;FD;5�>;�D3;��;�P�:4j:ȅ!��s@�%�ѻ�(;�v����y +�gys��R�����ht��-=��i���������6o��UD��      �(��Fl���.}�9ce�yPH���(�{
���ڽ�R����{�B�6�� �+p��[�`�ʨ��,��8IҺ�L^9���:ޣ;�~(;2�8;�IA;|E;jG;�=H;B�H;լH;�H;]�H;%�H;h�H;��H;��H;��H;��H;J�H;��H;��H;��H;��H;i�H;&�H;b�H; �H;֬H;B�H;�=H;jG;|E;�IA;2�8;�~(;�;���:�L^9.IҺ�,��ʨ�[�`�+p��� �A�6���{��R����ڽ{
���(�zPH�9ce��.}�El��      �-=�A�9��k/�/�����}��Ľ�!��gys�B�6�##��ɺ��vz����<^��`�$��~�T�r:��:��;�Y1;�H=;+xC;)wF;�G;�eH;H�H;��H;��H;��H;P�H;��H;��H;��H;c�H;w�H;��H;y�H;e�H;��H;��H;��H;Q�H;��H;��H;��H;H�H;�eH;�G;%wF;+xC;I=;�Y1;��;	��:X�r:x~�`�$�:^������vz��ɺ�##�B�6�gys��!����Ľ}���/���k/�A�9�      �` �~.�����ڽ�b��tr��Z��\�y +�� ��ɺ�>��O*�?ͻ�5R�ǅ���:6��:��;�);�t8;f�@;Z*E;n8G;?$H;@�H;A�H;�H;�H;��H;k�H;`�H; �H;M�H;��H;��H; �H;��H;��H;Q�H;�H;^�H;n�H;��H;&�H;�H;>�H;>�H;A$H;k8G;_*E;g�@;�t8;�);��;6��:�:�ƅ��5R�>ͻ�O*�=��ɺ�� �x +�\�Z��tr���b����ڽ���~.��      
A���R��#ڟ�����C��
�_�*:�������*p���vz��O*��4ֻk������094�:1;T� ;�D3;K�=;��C;�kF;��G;�\H;��H;N�H; �H;7�H;��H;v�H;��H;��H;�H;��H;W�H;��H;W�H;��H;
�H;��H;��H;z�H;��H;>�H; �H;L�H;��H;�\H;��G;�kF;��C;K�=;�D3;V� ;1;D�:��09���k��4ֻ�O*��vz�*p����輢��*:�	�_�C������#ڟ��R��      �_�\�<Q��f@�~ +��5�����X�ļv�Z�`����@ͻ
k��Hɺ �6�E�:�P�:,�;�d.;I�:;%�A;)|E;zNG;E'H;��H;ǥH;[�H;��H;#�H;H�H;W�H;3�H;��H;��H;�H;��H;��H;��H;�H;��H;��H;3�H;\�H;O�H;*�H;��H;[�H;��H;�H;C'H;NG;+|E;%�A;Q�:;�d.;-�;�P�:I�: ~6��Hɺk�>ͻ���Z�`�u�X�ļ�����5� +��f@� <Q�\�      /]� �,#������ټ�ɺ������
v��(;�ʨ�:^���5R�"��� �6����:���:��;-�*;�+8;�!@;Y�D;c�F;��G;�eH;~�H;��H;��H;��H;��H;��H;�H;r�H;��H;e�H;}�H;.�H;Y�H;+�H;z�H;e�H;��H;p�H;!�H;��H;��H;��H;��H;��H;��H;�eH;��G;d�F;[�D;�!@;�+8;'�*;��;���:���: 6�����5R�8^��ʨ��(;��
v������ɺ���ټ����,#� �      *p��bx��	ע��R��&��n�`���7�8��&�ѻ�,��]�$� ǅ���09K�:���:�;�~(;�Z6;��>;ϨC;�HF;ܠG;�DH;I�H;��H;��H;�H;)�H;�H;��H;��H;��H;��H;�H;��H;��H;��H;��H;��H;�H;��H;��H;��H;��H;�H;,�H;�H;��H;��H;F�H;�DH;ޠG;�HF;ըC;��>;�Z6;�~(;�;���:K�:��09 ǅ�Z�$��,��"�ѻ8����7�k�`�'���R��	ע�`x��      �I�+�E��(;��O*����<��GĻ�����s@� IҺP~��:D�:�P�:��;�~(;�5;�>;:C;4�E;zcG;;$H;�{H;;�H;�H;��H;��H;:�H;��H;�H;W�H;��H;O�H;��H;A�H;��H;��H;��H;=�H;��H;J�H;��H;Z�H; �H;��H;=�H;��H;��H;�H;:�H;�{H;;$H;}cG;9�E;;C;�>;�5;�~(;�;�P�:D�:��:@~�$IҺ�s@�����GĻ�<�����O*��(;�*�E�      ?�ѻ�ͻ'���;G��⿐�V�d���$��Iɺ��!� M^9`�r:,��:
1;,�;)�*;�Z6;�>;?�B;��E;�8G;�	H; nH;�H;L�H;��H;d�H;��H;��H;H�H;��H;��H;v�H;��H;��H;��H;�H;!�H;�H;��H;��H;��H;t�H;��H;�H;I�H;��H;��H;a�H;��H;F�H;�H;nH;�	H;�8G;��E;;�B;�>;�Z6;)�*;+�;
1;2��:|�r:�L^9��!��Iɺ��$�V�d�޿��>G��"����ͻ      e�)�!�$�3����������\��N��hS�904j:���:��:��;X� ;�d.;�+8;��>;:C;��E;�)G;��G;dH;��H;��H;_�H;��H;7�H;��H;��H;��H;��H;��H;J�H;{�H;`�H; �H;7�H;I�H;4�H;��H;]�H;x�H;F�H;��H;��H;��H;��H;��H;2�H;��H;_�H;��H;��H;dH;��G;�)G;��E;=C;��>;�+8;�d.;Y� ;��;��:���:<4j:`S�9�N��(�\�������2��#�$�      0�R� � V7�0E^9��:p�X:㿙:���:�P�:�;��;�);�D3;P�:;�!@;֨C;8�E;�8G;��G;�`H;r�H;�H;�H;{�H;<�H;3�H;M�H;^�H;��H;��H;��H;�H;��H;��H;0�H;n�H;c�H;h�H;,�H;��H;��H;	�H;��H;��H;��H;`�H;J�H;0�H;?�H;{�H;�H;�H;u�H;�`H;��G;�8G;7�E;ӨC;�!@;M�:;�D3;�);��;�;�P�:���:ݿ�:��X:��:D^9 `7�� �      ��:���:��:&��:��:�P�:�{;(;��;�~(;�Y1;�t8;I�=;$�A;Y�D;�HF;zcG;�	H;dH;o�H;I�H;ֶH;3�H;��H;��H;=�H;I�H;��H;#�H;��H;~�H;��H;U�H;��H;H�H;��H;��H;��H;H�H;��H;R�H;��H;~�H;��H;!�H;��H;E�H;:�H;��H;��H;/�H;ضH;L�H;q�H;dH;�	H;}cG;�HF;\�D;!�A;I�=;�t8;�Y1;�~(;��;(;�{;�P�:.��:&��:��:Í�:      0�
;L�;�;;D�;�`;�D&;�-;�D3;4�8;I=;d�@;��C;.|E;e�F;�G;?$H;nH;��H;�H;ڶH;��H;9�H;�H;g�H;��H;��H;u�H;k�H;�H; �H;��H;��H;�H;e�H;��H;��H;��H;c�H;�H;��H;��H; �H;�H;i�H;u�H;��H;��H;k�H;�H;5�H;��H;ܶH;�H;��H;nH;A$H;�G;g�F;*|E;��C;g�@;
I=;4�8;�D3;�-;�D&;�`;\�;;��;C�;      �*;L�*;n,;kd.;�Y1;ֱ4;,8;��;;<�>;�IA;3xC;_*E;�kF;�NG;��G;�DH;�{H; �H;��H;�H;0�H;7�H;��H;��H;��H;_�H;�H;��H;��H;��H;��H;p�H;��H;;�H;��H;��H;��H;��H;��H;;�H;��H;k�H;��H;��H;��H;��H;�H;a�H;��H;��H;��H;9�H;3�H;�H;��H;�H;�{H;�DH;��G;�NG;�kF;a*E;5xC;�IA;A�>;��;;�+8;ϱ4;�Y1;ld.;k,;6�*;      "�:;@�:;��;;�<;�>;��?;JA;��B;FD;|E;(wF;n8G;��G;I'H;�eH;M�H;;�H;P�H;`�H;x�H;��H;�H;��H;��H;�H;��H;��H;6�H;y�H;q�H;�H;��H;�H;]�H;�H;��H;��H;��H;|�H;]�H;�H;��H;�H;o�H;s�H;6�H;��H;��H;�H;��H;��H;�H;��H;v�H;_�H;J�H;<�H;M�H;�eH;C'H;��G;m8G;+wF;|E;FD;��B;JA;��?;>;��<;��;;5�:;      ңB;�B;�C;��C;�0D;��D;��E;iIF;��F;jG;$�G;H$H;�\H;�H;��H;��H;%�H;��H;��H;H�H;��H;m�H;��H;#�H;��H;s�H;��H;F�H;-�H;��H;��H;��H;/�H;t�H;��H;��H;��H;��H;��H;t�H;)�H;��H;��H;��H;&�H;E�H;��H;t�H;��H;�H;��H;p�H;��H;B�H;��H;��H;'�H;¨H;��H;�H;�\H;I$H;'�G;jG;��F;mIF;��E;��D;�0D;��C;�C;�B;      �HF;�TF;wF;��F;s�F;~8G;��G;��G;�	H;�=H; fH;B�H;��H;ΥH;��H;��H;��H;h�H;6�H;0�H;>�H;��H;a�H;��H;p�H;��H;%�H;�H;��H;G�H;��H;#�H;7�H;r�H;��H;��H;��H;��H;��H;q�H;3�H;�H;��H;C�H;��H;�H; �H;��H;t�H;��H;\�H;��H;>�H;/�H;5�H;d�H;��H;��H;��H;˥H;��H;C�H;fH;�=H;�	H;��G;��G;t8G;��F;��F;�vF;�TF;      ;�G;��G;�G;��G;VH;j0H;�LH;fH;7|H;C�H;J�H;@�H;I�H;]�H;��H;�H;��H;��H;��H;M�H;N�H;��H;�H;��H;��H;#�H;��H;��H;R�H;��H;��H;3�H;R�H;u�H;��H;��H;��H;��H;��H;v�H;N�H;-�H;��H;��H;J�H;��H;��H;'�H;��H;��H;�H;��H;N�H;L�H;��H;��H;��H;�H;��H;X�H;K�H;B�H;M�H;C�H;;|H;fH;}LH;d0H;nH;��G;�G;��G;      �lH;(nH;�rH;�yH;<�H;��H;�H;��H;��H;ݬH;��H;��H;��H;��H;��H;-�H;=�H;��H;��H;]�H;��H;r�H;��H;7�H;?�H;�H;��H;6�H;��H;��H;�H;=�H;a�H;e�H;�H;��H;��H;��H;}�H;e�H;^�H;7�H;�H;��H;��H;3�H;��H;�H;B�H;3�H;��H;s�H;��H;]�H;��H;��H;=�H;-�H;��H;��H;�H;��H;��H;ܬH;��H;��H;�H;��H;I�H;�yH;�rH;nH;      �H;��H;�H;��H;��H;i�H;{�H;�H;i�H;�H;��H;&�H;>�H;)�H;��H;�H;��H;N�H;��H;��H;*�H;g�H;��H;w�H;&�H;��H;K�H;��H;��H;�H;)�H;L�H;a�H;e�H;d�H;o�H;m�H;k�H;c�H;g�H;a�H;H�H;,�H;�H;��H;��H;D�H;��H;'�H;r�H;��H;f�H;&�H;��H;��H;L�H;��H;�H;��H;)�H;>�H;&�H;��H;!�H;p�H;�H;{�H;g�H;ŨH;��H;�H;��H;      t�H;��H;��H;�H;�H;q�H;4�H;-�H;4�H;b�H;��H;��H;��H;T�H;��H;��H;$�H;�H;��H;��H;��H;�H;��H;p�H;��H;<�H;��H;��H;�H;%�H;A�H;D�H;R�H;d�H;N�H;\�H;q�H;Z�H;I�H;d�H;N�H;A�H;@�H;"�H;�H;��H;��H;A�H;��H;l�H;��H;�H;��H;��H;��H;�H;$�H;��H;��H;Q�H;��H;��H;��H;f�H;7�H;0�H;8�H;p�H;�H;�H;��H;��H;      A�H;�H;�H;%�H;Z�H;�H;��H;��H;��H;*�H;U�H;u�H;�H;a�H;&�H;��H;a�H;��H;��H;��H;��H;#�H;��H;�H;��H;��H;��H;�H;0�H;G�H;V�H;O�H;A�H;@�H;a�H;O�H;/�H;L�H;]�H;B�H;@�H;O�H;V�H;E�H;*�H;	�H;��H;��H;��H;�H;��H;!�H;��H;��H;��H;��H;b�H;��H;&�H;a�H;��H;x�H;W�H;-�H;��H;��H;��H;��H;h�H;#�H;�H;�H;      ��H;��H;��H;��H;��H;��H;�H;d�H;��H;i�H;��H;g�H;��H;:�H;u�H;��H;��H;|�H;P�H;�H;��H;��H;n�H;��H;��H;�H;/�H;=�H;L�H;E�H;I�H;V�H;>�H;7�H;K�H;,�H;%�H;/�H;H�H;9�H;@�H;V�H;H�H;D�H;G�H;9�H;,�H;!�H;��H;��H;r�H;��H;��H;�H;O�H;}�H;��H;��H;u�H;:�H;��H;h�H;��H;l�H;��H;f�H;	�H;��H;��H;��H;��H;��H;      ��H;��H;�H;l�H;�H;��H;��H;��H;��H;��H;��H;�H; �H;��H;��H;��H;V�H;�H;��H;��H;_�H;��H;��H;�H;/�H;3�H;R�H;g�H;h�H;U�H;;�H;@�H;G�H;>�H;!�H;�H;K�H;�H;�H;A�H;D�H;B�H;:�H;P�H;a�H;a�H;O�H;4�H;0�H;�H;��H;��H;Y�H;��H;��H;�H;W�H;��H;��H;��H;�H;�H;��H;��H;��H;��H;��H;��H;�H;g�H;�H;��H;      F�H;X�H;��H;��H;c�H;��H;��H;\�H;�H;��H;��H;V�H;�H;��H;k�H;�H;��H;��H;d�H;��H;��H;#�H;:�H;W�H;r�H;n�H;q�H;g�H;g�H;g�H;:�H;:�H;@�H;(�H;�H;�H;%�H;�H;�H;)�H;@�H;:�H;:�H;d�H;a�H;c�H;o�H;o�H;t�H;V�H;>�H;"�H;��H;��H;d�H;�H;��H;�H;k�H;��H;�H;V�H;��H;��H;�H;]�H;��H;��H;m�H;��H;��H;b�H;      u�H;��H;��H;��H;V�H;��H;!�H;��H;3�H;��H;n�H;��H;��H;�H;��H;��H;H�H;��H;�H;4�H;N�H;d�H;��H;u�H;��H;��H;��H;�H;g�H;P�H;Y�H;L�H;!�H;�H;#�H;�H;��H;�H;"�H;�H;"�H;O�H;W�H;K�H;`�H;y�H;��H;��H;��H;u�H;��H;a�H;H�H;-�H; �H;��H;J�H;��H;��H;�H;��H;��H;q�H;��H;7�H;��H;&�H;��H;W�H;��H;��H;��H;      �H;�H;J�H;~�H;��H;�H;��H;��H;k�H;��H;~�H;��H;X�H;��H;/�H;��H;��H;�H;9�H;n�H;��H;��H;��H;��H;��H;��H;��H;��H;q�H;`�H;K�H;0�H;#�H;�H;�H;�H;�H;�H;�H;"�H;#�H;3�H;I�H;\�H;m�H;��H;��H;��H;��H;��H;��H;��H;��H;j�H;9�H;
�H;��H;��H;.�H;��H;X�H;��H;��H;��H;q�H;��H;��H;�H;��H;~�H;I�H;+�H;      ��H;��H;��H;�H;\�H;��H;�H;h�H;��H;L�H;��H;*�H;��H;�H;b�H;��H;��H;(�H;N�H;k�H;��H;��H;��H;��H;��H;��H;��H;��H;r�H;x�H;,�H;)�H;P�H;%�H;��H;�H;��H;�H;��H;&�H;S�H;,�H;,�H;t�H;k�H;��H;��H;��H;��H;��H;��H;��H;��H;h�H;O�H;,�H;��H;��H;`�H;	�H;��H;*�H;��H;M�H;��H;m�H;!�H;��H;_�H;�H;��H;��H;      �H;!�H;D�H;�H;��H;�H;��H;��H;k�H;��H;}�H;��H;Z�H;��H;/�H;��H;��H;�H;9�H;n�H;��H;��H;��H;��H;��H;��H;��H;��H;r�H;^�H;K�H;2�H;%�H;�H;�H;�H;�H;�H;�H;!�H;#�H;3�H;I�H;Z�H;m�H;��H;��H;��H;��H;��H;��H;��H;��H;j�H;9�H;
�H;��H;��H;.�H;��H;Z�H;��H;��H;��H;q�H;��H;��H;�H;��H;��H;L�H;'�H;      m�H;��H;��H;��H;V�H;��H;!�H;��H;3�H;��H;n�H;��H;��H;�H;��H;��H;G�H;��H; �H;2�H;N�H;d�H;��H;r�H;��H;��H;��H;}�H;g�H;N�H;W�H;L�H;!�H;�H;#�H;�H;��H;�H;#�H;�H;#�H;L�H;W�H;I�H;`�H;x�H;��H;��H;��H;t�H;��H;c�H;G�H;/�H; �H;��H;J�H;��H;��H;�H;��H;��H;n�H;��H;6�H;��H;*�H;��H;Z�H;��H;��H;��H;      F�H;W�H;��H;��H;e�H;��H;��H;^�H;�H;��H;��H;U�H;�H;��H;l�H;�H;��H;�H;c�H;��H;��H;#�H;:�H;Y�H;t�H;k�H;r�H;g�H;h�H;g�H;:�H;:�H;@�H;(�H;�H;�H;%�H;�H;�H;(�H;A�H;:�H;9�H;c�H;^�H;c�H;o�H;q�H;q�H;S�H;>�H;#�H;��H;��H;f�H;�H;��H;�H;l�H;��H;�H;U�H;��H;��H;�H;`�H;��H;��H;l�H;��H;��H;W�H;      ��H;��H;�H;g�H;�H;��H;��H;��H;��H;��H;��H;�H;�H;��H;��H;��H;V�H;�H;�H;��H;_�H;��H;��H;�H;0�H;-�H;O�H;g�H;h�H;U�H;:�H;=�H;E�H;=�H;�H;�H;K�H;�H;�H;@�H;B�H;A�H;:�H;O�H;^�H;`�H;N�H;4�H;-�H;�H;��H;��H;V�H;��H;��H;�H;V�H;��H;��H;��H;�H;�H;��H;��H;��H;��H;��H;��H;�H;o�H;�H;��H;      z�H;��H;��H;��H;��H;��H;�H;g�H;��H;i�H;��H;g�H;��H;;�H;w�H;��H;��H;|�H;M�H;�H;��H;��H;n�H;��H;��H;�H;*�H;=�H;O�H;D�H;H�H;U�H;>�H;6�H;K�H;*�H;%�H;/�H;H�H;9�H;>�H;V�H;G�H;B�H;G�H;7�H;*�H;�H;��H;��H;t�H;��H;��H;�H;O�H;|�H;��H;��H;u�H;:�H;��H;h�H;��H;j�H;��H;g�H;�H;��H;��H;��H;��H;��H;      5�H;�H;�H;�H;a�H;�H;��H;��H;��H;*�H;U�H;x�H;~�H;c�H;(�H;��H;b�H;��H;��H;��H;��H;#�H;��H;�H;��H;��H;��H;
�H;/�H;E�H;U�H;O�H;@�H;@�H;a�H;N�H;/�H;N�H;]�H;B�H;@�H;O�H;U�H;B�H;)�H;�H;��H;��H;��H;�H;��H;#�H;��H;��H;��H;��H;d�H;��H;'�H;a�H;�H;x�H;W�H;,�H;��H;��H;��H; �H;m�H;)�H;�H;~�H;      ��H;��H;��H;�H;�H;|�H;5�H;4�H;9�H;c�H;��H;��H;��H;R�H;��H;��H;$�H;�H;��H;��H;��H;�H;��H;m�H;��H;:�H;��H;��H;�H;!�H;@�H;B�H;N�H;d�H;L�H;Z�H;q�H;Z�H;K�H;d�H;O�H;B�H;@�H;"�H;
�H;��H;��H;C�H;��H;i�H;��H;�H;��H;��H;��H;�H;$�H;��H;��H;Q�H;��H;��H;��H;f�H;6�H;3�H;6�H;m�H;�H;"�H;��H;��H;      ��H;��H;*�H;��H;��H;p�H;{�H;�H;v�H;�H;��H;(�H;>�H;*�H;��H;�H;��H;P�H;��H;��H;+�H;i�H;��H;w�H;(�H;��H;F�H;��H;��H;
�H;(�H;L�H;`�H;e�H;c�H;m�H;m�H;m�H;c�H;e�H;a�H;L�H;,�H;�H;��H;��H;F�H;��H;'�H;r�H;��H;i�H;&�H;��H;��H;L�H;��H;�H;��H;)�H;@�H;%�H;��H;�H;s�H;�H;}�H;j�H;��H;��H;*�H;~�H;      �lH;nH;�rH;�yH;8�H;��H;��H;��H;��H;߬H;��H;��H; �H;��H;��H;-�H;=�H;��H;��H;]�H;��H;s�H;��H;6�H;B�H;�H;��H;3�H;��H;��H;�H;:�H;]�H;d�H;}�H;��H;��H;��H;}�H;g�H;c�H;:�H;	�H;��H;��H;2�H;��H;�H;?�H;4�H;��H;s�H;��H;]�H;��H;��H;=�H;-�H;��H;��H; �H;��H;��H;ܬH;��H;��H;�H;��H;I�H;�yH;�rH;nH;      -�G;��G;�G;��G;gH;t0H;�LH;fH;;|H;C�H;L�H;E�H;K�H;[�H;��H;�H;��H;��H;��H;L�H;O�H;��H;�H;��H;��H;�H;��H;��H;O�H;��H;��H;0�H;N�H;t�H;��H;��H;��H;��H;��H;x�H;R�H;3�H;��H;��H;K�H;��H;��H;'�H;��H;��H;�H;��H;L�H;O�H;��H;��H;��H;�H;��H;Z�H;I�H;A�H;L�H;B�H;:|H;fH;�LH;k0H;lH;��G;�G;��G;      �HF;�TF;	wF;�F;z�F;�8G;��G;��G;�	H;�=H;fH;G�H;��H;˥H;��H;��H;��H;i�H;6�H;0�H;@�H;��H;Z�H;��H;q�H;��H; �H;�H;��H;A�H;��H;!�H;3�H;q�H;��H;��H;��H;��H;��H;r�H;6�H;#�H;��H;D�H;��H;	�H;#�H;��H;q�H;��H;a�H;��H;>�H;0�H;6�H;b�H;��H;��H;��H;˥H;��H;B�H;fH;�=H;�	H;��G;��G;u8G;��F;��F;�vF;�TF;      ΣB;�B;�C;��C;�0D;��D; �E;jIF;��F;jG;'�G;I$H;�\H;�H;��H;¨H;%�H;��H;��H;C�H;��H;p�H;��H;!�H;��H;l�H;��H;C�H;*�H;��H;��H;��H;*�H;r�H;��H;��H;��H;��H;��H;v�H;/�H;��H;��H;��H;'�H;B�H;��H;t�H;��H; �H;��H;p�H;��H;C�H;��H;��H;'�H;��H;��H;�H;�\H;F$H;#�G;jG;��F;jIF;��E;��D;�0D;��C;�C;�B;       �:;$�:;�;;�<;�>;ʧ?;JA;��B;FD;|E;+wF;p8G;��G;F'H;�eH;P�H;;�H;P�H;_�H;v�H;��H;�H;��H;��H;�H;��H;��H;4�H;v�H;m�H;�H;��H;�H;]�H;|�H;��H;��H;��H;|�H;^�H;�H;��H;�H;q�H;u�H;3�H;��H;��H;�H;��H;��H;�H;��H;y�H;`�H;M�H;>�H;O�H;�eH;E'H;��G;k8G;)wF;|E;FD;��B;JA;��?;>;�<;}�;;�:;      �*;D�*;g,;ud.;�Y1;ϱ4;�+8;��;;D�>;�IA;.xC;a*E;�kF;�NG;��G;�DH;�{H; �H;��H;�H;2�H;9�H;��H;��H;��H;Z�H;�H;��H;��H;��H;��H;n�H;��H;;�H;��H;��H;��H;��H;��H;:�H;��H;q�H;��H;��H;��H;��H;�H;a�H;��H;��H;��H;9�H;5�H;�H;��H;�H;�{H;�DH;��G;�NG;�kF;\*E;.xC;�IA;?�>;��;;�+8;α4;�Y1;vd.;e,;/�*;      0�
;N�;��;;E�;�`;�D&;�-;�D3;4�8;
I=;j�@;��C;+|E;j�F;�G;?$H;nH;��H;�H;ڶH;��H;5�H;�H;m�H;��H;��H;u�H;i�H;�H;�H;��H;��H;�H;c�H;��H;��H;��H;a�H;�H;��H;��H;$�H;
�H;j�H;s�H;��H;��H;i�H;#�H;9�H;��H;ݶH;�H;��H;nH;?$H;�G;g�F;+|E;��C;f�@;I=;3�8;�D3;�-;�D&;�`;\�; ;��;B�;      ��:�:��:4��:��:�P�:�{;(;��;�~(;�Y1;�t8;K�=;$�A;]�D;�HF;{cG;�	H;dH;q�H;H�H;ٶH;/�H;��H;��H;7�H;D�H;��H; �H;��H;~�H;��H;R�H;��H;G�H;��H;��H;��H;G�H;��H;V�H;��H;��H;��H;!�H;��H;H�H;:�H;��H;��H;3�H;ٶH;L�H;r�H;dH;�	H;{cG;�HF;]�D;#�A;I�=;�t8;�Y1;�~(;��;(;�{;�P�:6��::��:�:ύ�:      ��R�� � Y7� E^9��:��X:鿙:���:�P�:�;��;�);�D3;N�:;�!@;רC;7�E;�8G;��G;�`H;r�H;�H;�H;{�H;?�H;/�H;H�H;]�H;��H;��H;��H;�H;��H;��H;/�H;j�H;d�H;k�H;,�H;��H;��H;�H;��H;��H;��H;^�H;M�H;3�H;>�H;�H;�H;�H;u�H;�`H;��G;�8G;7�E;ըC;�!@;L�:;�D3;�);��;�;�P�:���:ۿ�:h�X:��:�D^9 Y7�� �      c�)�!�$�1����������\��N��`S�9@4j:���:��:��;Y� ;�d.;�+8;��>;:C;��E;�)G;��G;dH;��H;��H;]�H;��H;3�H;��H;��H;��H;��H;��H;H�H;{�H;`�H;��H;6�H;I�H;6�H;��H;]�H;{�H;J�H;��H;��H;��H;��H;��H;5�H;��H;c�H;��H;��H;dH;��G;�)G;��E;:C;��>;�+8;�d.;V� ;��;��:���:44j:`S�9�N��$�\��������8���$�      F�ѻ�ͻ(���>G��ݿ��L�d���$��Iɺ��!� M^9t�r:2��:
1;+�;-�*;�Z6;�>;<�B;��E;�8G;�	H;nH;�H;J�H;��H;a�H;��H;��H;H�H;��H;��H;u�H;��H;��H;��H;�H;"�H;�H;��H;��H;��H;u�H;��H;�H;I�H;��H;��H;b�H;��H;J�H;�H;nH;�	H;�8G;��E;<�B;�>;�Z6;*�*;)�;1;,��:|�r:�L^9��!��Iɺ��$�R�d�޿��@G��,����ͻ      �I�,�E��(;��O*����<��GĻ�����s@� IҺH~���:D�:�P�:�;�~(;�5;�>;8C;5�E;{cG;;$H;�{H;;�H;�H;��H;��H;9�H;��H;�H;X�H;��H;O�H;��H;@�H;��H;��H;��H;?�H;��H;J�H;��H;]�H; �H;��H;:�H;��H;��H;�H;<�H;�{H;=$H;ycG;9�E;8C;�>;�5;�~(;�;�P�:D�:�:P~�(IҺ�s@�����GĻ�<�����O*��(;�+�E�      *p��bx��	ע��R��&��k�`���7�8��#�ѻ�,��Z�$��ƅ���09K�:���:�;�~(;�Z6;��>;ШC;�HF;ޠG;�DH;L�H;��H;��H;�H;(�H;�H;��H;��H;��H;��H;�H;��H;��H;��H;��H;��H;�H;��H;��H;��H;��H;�H;*�H;�H;��H;��H;K�H;�DH;ޠG;�HF;ըC;��>;�Z6;�~(;�;���:I�:��09ǅ�[�$��,��$�ѻ8����7�l�`�(���R��ע�bx��      /]� �,#������ټ�ɺ������
v��(;�ɨ�9^���5R���� 6����:���:��;)�*;�+8;�!@;[�D;d�F;��G;�eH;��H;��H;��H;��H;��H;��H; �H;r�H;��H;g�H;{�H;)�H;X�H;)�H;{�H;g�H;��H;p�H; �H;��H;��H;��H;��H;��H;�H;�eH;��G;e�F;X�D;�!@;�+8;'�*;��;���:���: �6� ����5R�:^��ʨ��(;��
v������ɺ���ټ����,#� �      �_�\� <Q��f@�~ +��5�����X�ļu�Z�`����>ͻk��Hɺ |6�Q�:�P�:+�;�d.;L�:;*�A;*|E;NG;G'H;�H;ȥH;X�H;��H;&�H;K�H;\�H;3�H;��H;��H;�H;��H;��H;��H;�H;��H;��H;3�H;Z�H;O�H;*�H;��H;X�H;ǥH;��H;I'H;�NG;*|E;#�A;P�:;�d.;,�;�P�:K�: 6��Hɺk�@ͻ���Z�`�v�X�ļ�����5� +��f@�<Q�\�      
A���R��#ڟ�󻒽C��
�_�*:�������*p���vz��O*��4ֻk������09>�:1;T� ;�D3;O�=;��C;�kF;��G;�\H;��H;H�H;��H;=�H;��H;x�H;��H;��H;
�H;��H;W�H;��H;W�H;��H;
�H;��H;��H;x�H;��H;@�H; �H;I�H;��H;�\H;��G;�kF;��C;F�=;�D3;R� ;1;>�:��09���k��4ֻ�O*��vz�+p����輣��*:�
�_�C������#ڟ��R��      �` �~.�����ڽ�b��tr��Z��\�x +�� ��ɺ�=��O*�>ͻ�5R��ƅ���:*��:��;�); u8;f�@;_*E;p8G;D$H;@�H;=�H;�H;"�H;��H;o�H;`�H;�H;Q�H;��H;��H;!�H;��H;��H;O�H; �H;^�H;n�H;��H;(�H;�H;=�H;?�H;>$H;n8G;a*E;g�@;�t8;�);��;2��:�:ǅ��5R�@ͻ�O*�>��ɺ�� �x +�\�Z��tr���b����ڽ���~.��      �-=�A�9��k/�/�����}��Ľ�!��gys�B�6�##��ɺ��vz����:^��`�$��~�L�r:��:��;�Y1;I=;.xC;(wF;�G;�eH;E�H;��H;��H;��H;S�H;��H;��H;��H;d�H;z�H;��H;y�H;d�H;��H;��H;��H;P�H;��H;��H;��H;E�H;�eH;�G;(wF;.xC;�H=;�Y1;��;��:X�r:�~�a�$�;^������vz��ɺ�##�B�6�gys��!����Ľ}���/���k/�A�9�      �(��El���.}�9ce�yPH���(�{
���ڽ�R����{�A�6�� �+p��\�`�ʨ��,��2IҺ�L^9���:�;�~(;2�8;�IA;|E;jG;�=H;A�H;լH;�H;`�H;(�H;h�H;��H;��H;��H;��H;L�H;��H;��H;��H;��H;f�H;%�H;_�H;!�H;֬H;?�H;�=H;jG;|E;�IA;0�8;�~(;�;���:�L^9.IҺ�,��ʨ�[�`�+p��� �B�6���{��R����ڽ{
���(�zPH�9ce��.}�El��      �iþUD��6o�����������i��-=�ht�����R��gys�y +����v񗼐(;�$�ѻ�s@�ԅ!�4j:�P�:��;�D3;7�>;FD;��F;�	H;:|H;��H;t�H;6�H;��H;��H;��H;�H;.�H;n�H;��H;m�H;/�H;�H;��H;��H;��H;6�H;v�H;��H;:|H;�	H;��F;FD;8�>;�D3;��;�P�:4j:ą!��s@�&�ѻ�(;�v����y +�gys��R�����ht��-=��i���������6o��UD��      ���
�����#�޾UD���A���.}�(�D�ht���ڽ�!��\����Y�ļ�
v�:��Ŀ���Iɺ(S�9���: (;�-;��;;��B;jIF;��G;fH;��H;�H;-�H;��H;d�H;��H;]�H;��H;��H;h�H;��H;��H;Y�H;��H;c�H;��H;1�H;�H;��H;fH;��G;hIF;��B;��;;�-;(;���:S�9�Iɺÿ��;���
v�Y�ļ���\��!����ڽht�(�D��.}��A��VD��#�޾�����
�      ��7�ϕ3��f'�(��\���о�����.}��-=�{
���Ľ[��*:�����������7�GĻ��$� O��Ϳ�:�{;�D&;�+8;JA;�E;��G;wLH;�H;v�H;4�H;��H; �H;��H;��H;�H;��H;�H;��H;�H;��H;��H; �H;��H;6�H;y�H;�H;{LH;��G;�E;JA;�+8;�D&;�{;ѿ�:�N����$�GĻ��7���������*:�[����Ľ{
��-=��.}������о�\��(��f'�ϕ3�      Xo�_Xi��"Y���@�K�#��
��о�A���i���(�}��ur��
�_��5��ɺ�n�`��<��_�d�P�\�h�X:�P�:�`;α4;��?;��D;u8G;j0H;��H;k�H;u�H;�H;��H;��H;��H;��H;�H;��H;�H;��H;��H;��H;��H;�H;w�H;m�H;��H;k0H;~8G;��D;��?;̱4;�`;�P�:p�X:\�\�]�d��<��n�`��ɺ��5�
�_�ur��}����(��i��A���о�
�K�#���@��"Y�_Xi�      /����������Xo��!J�K�#��\��VD������zPH�����b��C��� +���ټ'����꿐�
�����:.��:E�;�Y1;	>;�0D;y�F;^H;C�H;¨H;
�H;[�H;��H;	�H;e�H;E�H;��H;_�H;��H;H�H;_�H;�H;��H;X�H;�H;ŨH;H�H;dH;��F;�0D;	>;�Y1;H�;,��:��:���濐���'����ټ� +�C���b�����zPH�����UD���\��K�#��!J�Xo��������      =^������k���Xo���@�(�#�޾����9ce�/����ڽ󻒽�f@������R���O*�FG����� D^94��:;^d.; �<;��C;�F;��G;�yH;��H;�H; �H;��H;i�H;��H;��H;��H;�H;~�H;��H;��H;i�H;��H;�H; �H;��H;�yH;��G;��F;��C; �<;Zd.;;4��:PD^9���CG���O*��R�������f@�󻒽��ڽ/��9ce�����#�޾(���@�Xo�k�������      �aǿ�¿����������"Y��f'�����6o���.}��k/����#ڟ� <Q�,#�ע��(;�*���3�� `7��:�;u,;��;;�C;�vF;�G;�rH;�H;��H;�H;��H;��H;��H;��H;L�H;��H;G�H;��H;��H;��H;��H;�H;��H;�H;�rH;�G;wF;�C;��;;o,;�;�: \7�2��'����(;�ע�,#� <Q�#ڟ�����k/��.}�6o�������f'��"Y�����������¿      2�ֿCpѿ�¿������_Xi�ϕ3��
�UD��Fl��A�9�.���R��\� �cx��.�E��ͻ�$�� �卨:@�;P�*;8�:;�B;�TF;��G;&nH;��H;��H;k�H;��H;��H;[�H;��H;�H;��H;�H;��H;[�H;��H;��H;g�H;ŷH;��H;)nH;��G;�TF;�B;5�:;H�*;>�;卨:� ��$��ͻ.�E�cx�� �\��R��.��A�9�Fl��UD���
�ϕ3�_Xi��������¿Cpѿ      �� $������꿯�ſ�ޞ�%3s��2�>����� j���xHͽƸ����'�@<ͼp�n�b���:Q^��-.�x��:pW;dS%;io8;��A;DF;�H;{�H;��H;��H; �H;�H;#�H;��H;��H;��H;�H;��H;��H;��H;"�H;�H;�H;��H;��H;~�H;�H; DF;��A;eo8;]S%;nW;~��:�-.�;Q^�`���p�n�@<ͼ��'�Ƹ��xHͽ�� j���=����2�%3s��ޞ���ſ������ $�       $�������忇�����cm�U�-�����Ph��Vde�!-�֪ɽ�v��'�$�~�ɼxmj�4���X����ņ:jx;�%;6�8;HB;#RF;�H;�H;�H;��H;E�H;�H;�H;x�H;��H;��H;�H;��H;��H;u�H;�H;�H;A�H;��H;�H;�H;�H;-RF;FB;2�8;�%;jx;�ņ:���X�2���xmj�~�ɼ'�$��v��֪ɽ!-�Vde�Ph������U�-�cm��������忝����      ����������ԿLw�����:�\�"����k��Y0X�����;����w����������]����F�����ɒ:��;�';��9;�oB;�zF;�!H;u�H;��H;�H;p�H;�H;�H;��H;��H;��H;��H;��H;��H;}�H;�H;�H;k�H;	�H;��H;u�H;�!H;�zF;�oB;��9;�';��;�ɒ:����F��黩�]����������w��;�����Y0X�k�����"�:�\����Lw���Կ��𿝏�      ������Կp���ޞ�_F�g�C�-E�"�;�I��D���"��e�c�{��֯���J��ѻʢ)��K�'��:�
;�M*;p�:;�C;͸F;�8H;/�H;K�H;[�H;��H;�H;�H;��H;��H;��H;��H;��H;��H;�H;�H;�H;��H;_�H;M�H;-�H;�8H;ӸF;�C;l�:;�M*;�
;'��:K�ʢ)��ѻ��J��֯�{�e�c�"����D��I��"�;-E�g�C�_F��ޞ�p���Կ��      ��ſ���Lw���ޞ�����>�W�5�%�����hɰ��|x�e{+�ѱ����J��  �Ͷ��X�1�'���+�` 
9��:��;�-;��<;`�C;�G;�TH;'�H;��H;��H;��H;+�H;�H;e�H;��H;u�H;��H;q�H;��H;c�H;�H;+�H;��H;��H;��H;'�H;�TH;�G;]�C;��<;߷-;��;��:� 
9+�&���X�1�Ͷ���  ��J���ѱ�e{+��|x�hɰ�����5�%�>�W������ޞ�Lw�����      �ޞ�������_F�>�W�W�-���?Kɾ�G����O����ƽǸ��̈́-���ۼㄼ34�ǐ��ζ�,]:���:�;��1;�c>;F�D;{\G;.sH;x�H;7�H;D�H;��H;J�H;�H;I�H;j�H;]�H;��H;Z�H;h�H;D�H;
�H;K�H;��H;J�H;7�H;x�H;,sH;\G;E�D;�c>;z�1;�;��:4]:�ζ�ǐ�34�ㄼ��ۼ̈́-�Ǹ��ƽ�����O��G��?Kɾ��W�-�>�W�_F�������      %3s�cm�:�\�g�C�5�%����TҾj��	 j��C(����]P����[�{������Y�6��_X�T�<��k::��:�� ;؟5;4R@;8uE;ѲG;�H; �H;��H;��H;!�H;F�H;	�H;A�H;N�H;9�H;n�H;6�H;L�H;@�H;�H;D�H;�H;��H;��H; �H;�H;ղG;8uE;0R@;ԟ5;�� ;0��:�k:X�<�_X�5����Y����{���[�\P����콪C(�	 j�j���TҾ��5�%�g�C�:�\�cm�      �2�U�-�"�-E�����?Kɾj����s�8�5���t㻽�v��z0��;��+���*����06� AS�MM�:R�	;r�(;��9;�/B;JDF;"H;��H;]�H;��H;��H;M�H;c�H;��H;�H;�H;�H;:�H;�H;�H;�H;��H;`�H;J�H;��H;��H;]�H;��H;#H;KDF;�/B;��9;r�(;L�	;WM�:@AS�-6�����*��+���;�z0��v��t㻽��8�5���s�j��?Kɾ����-E�"�U�-�      =����������"�;hɰ��G��	 j�8�5��	�ΪɽX����J�r���沼��]�����	x�L	��$n:���:�v;��/;h-=;��C;�F;�HH;|�H;��H;��H;�H;}�H;f�H;��H;��H;��H;��H;�H;��H;��H;��H;��H;f�H;{�H;�H;��H;��H;z�H;�HH;�F;��C;j-=;��/;�v;���:(n:L	���	x������]��沼r���J�X���Ϊɽ�	�8�5�	 j��G��hɰ�"�;��徶���      ��Ph��k���I���|x���O��C(��Ϊɽ����QDX�F��%<ͼㄼ�X!��s���W��uK���:�y; �#;�H6;R@;�PE;h�G;]�H;��H;�H;��H;}�H;��H;T�H;��H;��H;��H;��H;��H;��H;��H;��H;��H;R�H;��H;��H;��H;�H;��H;Y�H;k�G;�PE;R@;�H6;��#;�y;!��:puK��W��s���X!�ㄼ%<ͼF��QDX�����Ϊɽ��C(���O��|x��I��k��Ph��       j�Vde�Y0X�D�e{+�������t㻽Y���QDX������ۼʾ����;�B>ۻX�P�y��>":���:��;·-;��;;��B;ozF;�H;a�H;X�H;��H;��H;��H;��H;N�H;��H;|�H;r�H;��H;\�H;��H;r�H;|�H;��H;K�H;��H;��H;��H;��H;W�H;]�H;�H;kzF;��B;��;;·-;��;���:�>":@�y�X�A>ۻ��;�ɾ����ۼ���QDX�X���t㻽��콂��e{+�D�Y0X�Vde�      ��!-������б�ƽ\P���v���J�F����ۼ��a�J������+��|rѺ`(
9�M�:��;v $;��5;��?;`�D;@\G;�eH;��H;��H;��H;��H;��H;��H;5�H;T�H;<�H;5�H;G�H;�H;G�H;3�H;=�H;R�H;2�H;��H;�H;��H;��H;��H;��H;�eH;@\G;d�D;��?;��5;� $;��;�M�:�(
9|rѺ�+������`�J�
����ۼF���J��v��\P��ƽѱ轂����!-�      xHͽ֪ɽ�;��"����Ǹ����[�z0�r��$<ͼɾ��`�J�����j��w*� ��:Bb�:9�;��/;�L<;�C;mF;o�G;ۡH;��H;��H;��H;�H;2�H;��H;�H;�H;��H;��H;��H;��H;��H;��H;��H;�H;�H;��H;8�H;�H;��H;��H;��H;�H;o�G;mF;�C;�L<;��/;=�;>b�:���:��t*��j�����`�J�ɾ��$<ͼq��z0���[�Ƹ����"���;��֪ɽ      Ÿ���v����w�e�c��J�̈́-�z��;缃沼ㄼ��;������j���5�0��?Q:<��:Si;�M*;h�8;g�@;�PE;�uG;iH;��H;��H;��H;��H;��H;T�H;��H;��H;��H;��H;��H;��H;��H;��H;��H;��H;��H;��H;��H;\�H;��H; �H;��H;��H;��H;iH;�uG;�PE;g�@;p�8;�M*;Si;J��:?Q:�깟5��j��������;�ㄼ�沼�;�{�̄-��J�e�c���w��v��      ��'�'�$����{��  ���ۼ����+����]��X!�@>ۻ�+��w*�0����>:���:��;%�%;ҟ5;|�>;�(D;��F;W!H;�H;*�H;��H;��H;��H;��H;L�H;��H;��H;j�H;p�H;J�H;6�H;Q�H;4�H;I�H;p�H;j�H;��H;��H;Q�H;��H;��H;��H;��H;+�H;�H;X!H;��F;�(D;��>;ԟ5;!�%;�;���:��>:(��u*��+��>>ۻ�X!���]��+�������ۼ�  �{����'�$�      =<ͼ|�ɼ�����֯�̶��ㄼ��Y��*�����s��X�xrѺ0�?Q:���:��
;8�#;S�3;wc=;�#C;DF;��G;�H;��H;��H;�H;��H;5�H;��H;F�H;o�H;G�H;�H;2�H;��H;��H;��H;��H;��H;2�H;�H;F�H;s�H;I�H;�H;8�H;��H;�H;��H;��H;��H;��G;DF;�#C;xc=;M�3;<�#;��
;���:?Q:P�|rѺX��s������*���Y�ㄼͶ���֯�����{�ɼ      k�n�tmj���]���J�V�1�14�0������	x��W�(�y��(
9���:J��:�;<�#;>�2;�<;QpB;�E;��G;�eH;��H;�H;��H;��H;��H;��H;�H;*�H;�H;��H;��H;��H;��H;��H;��H;��H;��H;��H;��H;��H;�H;+�H;�H;��H;��H;��H;��H;�H;��H;�eH;��G;�E;QpB;�<;A�2;<�#;�;J��:���:�(
9$�y��W��	x����2��04�V�1���J���]�smj�      R���,������ѻ ���ǐ�QX�$6�B	�� uK�?":�M�:8b�:Pi;$�%;M�3;�<;00B;��E;X\G;�HH;$�H;z�H;@�H;��H;�H;�H;��H;��H;��H;��H;��H;��H;C�H;8�H;8�H;�H;5�H;4�H;C�H;��H;��H;��H;��H;��H;��H;�H;�H;��H;<�H;v�H;%�H;�HH;]\G;��E;,0B;�<;L�3;$�%;Pi;8b�:�M�:$?":uK�8	��"6�VX�ǐ�����ѻ��.���      #Q^�X��F���)�+��ζ�(�<��>S�@n:)��:Ž�:��;=�;�M*;֟5;zc=;QpB;��E;�JG;08H;M�H;g�H;��H;�H;d�H;��H;u�H;��H;��H;��H;v�H;[�H;7�H;��H;��H;��H;��H;��H;��H;��H;5�H;Z�H;v�H;��H;��H;��H;p�H;��H;i�H;�H;��H;h�H;P�H;68H;�JG;��E;TpB;tc=;؟5;�M*;?�;��;ɽ�:)��:Ln:@?S�8�<��ζ�+�̢)��F�X�      �-.���X�� ~K�� 
9@]:H�k:UM�:���:�y;��;~ $;��/;n�8;��>;�#C;�E;`\G;48H;��H;��H; �H;p�H;�H;j�H;5�H;��H;��H;��H;e�H;�H;��H;��H;��H;�H;v�H;]�H;q�H;{�H;��H;��H;��H;�H;a�H;��H;��H;��H;0�H;m�H;�H;l�H; �H;��H;��H;68H;\\G;
�E;�#C;��>;l�8;��/;� $;��;�y;���:[M�:8�k:X]:� 
9K����<��      ���:�ņ:�ɒ:��:��: ��:2��:M�	;�v;�#;��-;��5;~L<;g�@;�(D;DF;��G;�HH;P�H;��H;��H;+�H;��H;@�H;��H;p�H;��H;��H;C�H;�H;��H;��H;U�H;H�H;�H;�H;�H;	�H;�H;G�H;R�H;��H;��H;�H;A�H;��H;��H;l�H;�H;;�H;��H;,�H;��H;��H;P�H;�HH;��G;DF;�(D;c�@;�L<;��5;Ʒ-; �#;�v;M�	;@��:���:��:��:�ɒ:�ņ:      pW;vx;��;"�
;��;�;�� ;r�(;��/;�H6;��;;��?;�C;�PE;��F;��G;�eH;+�H;l�H;�H;/�H;��H;�H;��H;C�H;h�H;l�H;L�H;��H;��H;��H;0�H;��H;��H;��H;��H;��H;��H;��H;��H;��H;*�H;��H;��H;��H;L�H;h�H;e�H;H�H;��H;�H;��H;/�H;�H;k�H;(�H;�eH;��G;��F;�PE;�C;��?;��;;�H6;��/;x�(;�� ;�;��;�
;��;nx;      {S%;�%;��';�M*;޷-;��1;�5;��9;q-=;R@;��B;f�D;mF;�uG;[!H;��H;��H;��H;��H;m�H;��H;�H;��H;J�H;a�H;Z�H;�H;��H;��H;|�H;
�H;��H;��H;�H;p�H;Y�H;:�H;U�H;k�H;��H;��H;��H;
�H;y�H;��H;��H;�H;]�H;e�H;H�H;��H;�H;��H;m�H;��H;y�H;��H;�H;Y!H;�uG;mF;f�D;��B;R@;t-=;�9;�5;��1;�-;�M*;��';��%;      fo8;<�8;��9;p�:;{�<;�c>;5R@;�/B;��C;�PE;lzF;A\G;o�G;iH;�H;��H;�H;E�H;�H;�H;>�H;��H;I�H;T�H;L�H;-�H;��H;��H;V�H;��H;��H;��H;G�H;�H;�H;�H;��H;	�H;�H;�H;C�H;��H;��H;��H;P�H;��H;��H;0�H;O�H;Q�H;C�H;��H;>�H;�H;
�H;?�H;�H;��H;�H;iH;m�G;A\G;pzF;�PE;��C;�/B;2R@;�c>;��<;m�:;��9;2�8;      ��A;CB;�oB;�C;W�C;V�D;CuE;KDF;�F;o�G;�H;�eH;�H;��H;1�H;��H;��H;��H;q�H;t�H;�H;H�H;i�H;V�H;�H;��H;��H;\�H;��H;��H;b�H;3�H;��H;��H;��H;��H;��H;��H;��H;��H;��H;,�H;b�H;��H;��H;Z�H;��H;��H;�H;S�H;e�H;I�H;�H;o�H;p�H;��H;��H;��H;1�H;��H;�H;�eH;�H;o�G;"�F;NDF;CuE;L�D;e�C;�C;�oB;EB;      DF;-RF;�zF;̸F;�G;�\G;ֲG;-H;�HH;c�H;c�H;��H;��H;��H;��H;�H;��H;�H;��H;1�H;r�H;d�H;[�H;3�H;��H;x�H;K�H;��H;��H;U�H;�H;��H;��H;��H;h�H;U�H;b�H;P�H;c�H;��H;��H;��H;�H;R�H;��H;��H;G�H;{�H;��H;0�H;X�H;e�H;p�H;0�H;��H;�H;��H;�H;��H;��H;��H;��H;g�H;c�H;�HH;.H;ղG;x\G;�G;ӸF;�zF;*RF;      �H; H;�!H;�8H;�TH;,sH;!�H;��H;|�H;��H;[�H;��H;��H;��H;��H;��H;��H; �H;w�H;��H;��H;i�H;�H;��H;��H;I�H;��H;{�H;@�H;	�H;��H;��H;X�H;9�H;$�H;�H;�H;��H;�H;;�H;T�H;��H;��H;�H;9�H;x�H;��H;N�H;��H;��H;�H;l�H;��H;��H;u�H;�H;��H;��H;��H;��H;��H;��H;[�H;��H;~�H;��H;�H;'sH;�TH;�8H;�!H;�H;      ��H;�H;n�H;6�H;�H;z�H;-�H;]�H;�H;�H;�H;��H;��H;�H;��H;:�H;��H;��H;��H;��H;��H;I�H;��H;��H;V�H;��H;x�H;M�H;��H;��H;i�H;?�H;�H;��H;��H;��H;��H;��H;��H;��H;�H;<�H;i�H;��H;��H;J�H;r�H;��H;W�H;��H;��H;I�H;��H;��H;��H;��H;��H;:�H;��H; �H;��H;��H;�H;�H;�H;`�H;-�H;o�H;*�H;6�H;q�H;��H;      ��H;�H;��H;[�H;��H;3�H;��H;��H;��H;��H;��H;��H;�H;��H;��H;�H; �H;��H;��H;��H;H�H;��H;��H;U�H;��H;��H;7�H;��H;��H;c�H;-�H;��H;��H;��H;��H;��H;w�H;��H;��H;��H;��H;��H;-�H;b�H;��H;��H;2�H;��H;��H;O�H;��H;��H;E�H;��H;��H;��H; �H;�H;��H;��H;�H;��H;��H;��H;��H;��H;��H;1�H;��H;\�H;��H;�H;      ��H;��H;�H;S�H;��H;D�H;��H;��H;�H;��H;��H;�H;6�H;_�H;N�H;I�H;/�H;��H;��H;e�H;
�H;��H;v�H;��H;��H;M�H;�H;��H;e�H;&�H;��H;��H;��H;��H;a�H;F�H;:�H;E�H;]�H;��H;��H;��H;��H;#�H;_�H;��H;��H;O�H;��H;��H;y�H;��H;�H;b�H;��H;��H;/�H;L�H;M�H;\�H;8�H;�H;��H;��H;�H;��H;��H;C�H;��H;X�H;�H;��H;      &�H;[�H;w�H;��H;��H;��H;'�H;T�H;��H;��H;��H;��H;��H;��H;��H;x�H;#�H;��H;z�H;%�H;��H;��H;	�H;��H;_�H;	�H;��H;o�H;2�H;��H;��H;~�H;s�H;:�H;�H;"�H; �H;�H;�H;<�H;r�H;}�H;��H;��H;-�H;j�H;��H;�H;c�H;��H;�H;��H;��H;�H;z�H;��H;#�H;x�H;��H;��H;��H;��H;��H;��H;��H;W�H;/�H;��H;��H;��H;y�H;[�H;      �H;�H;�H;�H;$�H;A�H;J�H;d�H;k�H;T�H;O�H;9�H;�H;��H;��H;J�H;��H;��H;`�H;��H;��H;0�H;��H;��H;0�H;��H;��H;@�H;��H;��H;y�H;]�H;<�H;�H;��H;��H;��H;��H;��H;�H;>�H;[�H;w�H;��H;��H;=�H;��H;��H;2�H;��H;��H;0�H;��H;��H;^�H;��H;��H;M�H;��H;��H;�H;7�H;T�H;V�H;j�H;c�H;O�H;D�H;3�H;�H; �H;�H;      /�H;#�H;)�H;�H;�H;�H;�H;��H;��H;��H;��H;X�H;�H;��H;m�H;�H;��H;��H;;�H;��H;`�H;�H;��H;D�H;��H;��H;X�H;�H;��H;��H;n�H;<�H;��H;��H;��H;��H;��H;��H;��H;��H;��H;?�H;l�H;��H;��H;�H;U�H;��H;��H;F�H;��H;�H;Z�H;��H;<�H;��H;��H;!�H;o�H;��H;�H;X�H;��H;��H;��H;��H;	�H;��H;"�H;�H;2�H;#�H;      |�H;v�H;�H;{�H;d�H;>�H;E�H;�H;��H;��H;��H;C�H;�H;��H;w�H;9�H;��H;H�H;��H;��H;O�H;��H;�H;�H;��H;��H;5�H;��H;��H;��H;4�H;�H;��H;��H;��H;��H;��H;��H;��H;��H;��H;
�H;5�H;��H;��H;��H;4�H;��H;��H;�H;��H;��H;K�H;��H;��H;M�H;��H;;�H;v�H;��H;�H;A�H;��H;��H;��H;�H;K�H;>�H;k�H;{�H;��H;��H;      ��H;��H;��H;��H;��H;c�H;U�H;!�H;��H;��H;|�H;@�H;�H;��H;S�H;��H;��H;8�H;��H;��H;�H;��H;m�H;�H;��H;_�H;�H;��H;��H;b�H;�H;��H;��H;��H;��H;��H;��H;��H;��H;��H;��H;��H;�H;^�H;��H;��H;�H;b�H;��H;�H;p�H;��H;�H;|�H;��H;>�H;��H;��H;S�H;��H;�H;A�H;�H;��H;��H;#�H;Y�H;c�H;��H;��H;��H;��H;      ��H;��H;��H;��H;j�H;V�H;@�H;�H;��H;��H;��H;K�H;��H;��H;8�H;��H;��H;5�H;��H;u�H;�H;��H;R�H;�H;��H;J�H;��H;��H;��H;I�H;�H;��H;��H;��H;��H;��H;��H;��H;��H;��H;��H;��H;�H;E�H;��H;��H;��H;M�H;��H;�H;X�H;��H;�H;t�H;��H;<�H;��H;��H;9�H;��H;��H;J�H;��H;��H;��H;�H;G�H;W�H;m�H;��H;��H;��H;      �H;�H;
�H;��H;��H;��H;r�H;;�H;�H;��H;f�H;$�H;��H;��H;Z�H;��H;��H;�H;��H;d�H;�H;��H;<�H;��H;��H;^�H;�H;��H;}�H;?�H;�H;��H;��H;��H;��H;��H;y�H;��H;��H;��H;��H;��H;�H;;�H;w�H;��H;�H;a�H;��H;��H;?�H;��H;	�H;`�H;��H;�H;��H;��H;\�H;��H;��H;"�H;j�H;��H;�H;@�H;y�H;��H;��H;��H;
�H;�H;      ��H;��H;��H;��H;k�H;Z�H;@�H;�H;��H;��H;��H;K�H;��H;��H;6�H;��H;��H;5�H;��H;u�H;�H;��H;R�H;�H;��H;J�H;��H;��H;��H;H�H;�H;��H;��H;��H;��H;��H;��H;��H;��H;��H;��H;��H;�H;C�H;��H;��H;��H;N�H;��H;�H;X�H;��H;�H;t�H;��H;<�H;��H;��H;9�H;��H;��H;K�H;��H;��H;��H;"�H;G�H;V�H;q�H;��H;��H;��H;      ��H;��H;��H;��H;��H;^�H;S�H;#�H;��H;��H;|�H;@�H;�H;��H;U�H;��H;��H;:�H;��H;��H;!�H;��H;m�H;�H;��H;^�H;�H;��H;��H;a�H;�H;��H;��H;��H;��H;��H;��H;��H;��H;��H;��H;��H;�H;[�H;��H;��H;�H;b�H;��H;�H;p�H;��H;�H;}�H;��H;>�H;��H;��H;Q�H;��H;�H;C�H;|�H;��H;��H;)�H;]�H;]�H;��H;��H;��H;��H;      |�H;u�H;}�H;|�H;e�H;B�H;D�H;�H;��H;��H;��H;C�H;�H;��H;x�H;8�H;��H;J�H;��H;��H;O�H;��H;�H;�H;��H;��H;6�H;��H;��H;��H;4�H;�H;��H;��H;��H;��H;��H;��H;��H;��H;��H;
�H;4�H;��H;��H;��H;4�H;��H;��H;�H;��H;��H;I�H;��H;��H;L�H;��H;<�H;x�H;��H;�H;D�H;��H;��H;��H;�H;L�H;@�H;n�H;}�H;��H;u�H;      -�H;)�H;*�H;�H;�H;�H;�H;��H;��H;��H;��H;[�H;�H;��H;q�H;�H;��H;��H;>�H;��H;^�H;�H;��H;F�H;��H;��H;U�H;�H;��H;��H;l�H;;�H;��H;��H;��H;��H;��H;��H;��H;��H;��H;?�H;n�H;��H;��H;�H;U�H;��H;��H;C�H;��H;�H;W�H;��H;?�H;��H;��H;!�H;o�H;��H;�H;Y�H;��H;��H;��H;��H;�H;�H;�H;"�H;3�H;#�H;      �H;�H;�H;�H;$�H;Q�H;M�H;f�H;j�H;T�H;R�H;9�H;�H;��H;��H;M�H;��H;��H;`�H;��H;��H;3�H;��H;��H;2�H;��H;�H;@�H;��H;��H;v�H;Z�H;<�H;�H;��H;��H;��H;��H;��H;�H;<�H;[�H;v�H;��H;��H;<�H;�H;��H;0�H;��H;��H;2�H;��H;��H;a�H;��H;��H;M�H;��H;��H;�H;<�H;T�H;X�H;n�H;f�H;O�H;D�H;)�H;�H;�H;�H;      �H;[�H;w�H;��H;��H;��H;&�H;T�H;��H;��H;��H;��H;��H;��H;��H;z�H;#�H;��H;z�H;"�H;��H;��H;
�H;��H;c�H;�H;��H;j�H;2�H;��H;��H;}�H;r�H;:�H;�H; �H; �H;"�H;�H;<�H;r�H;~�H;��H;��H;+�H;i�H;��H;�H;_�H;��H;�H;��H;��H;"�H;}�H;��H;$�H;z�H;��H;��H;��H;��H;��H;��H;��H;W�H;+�H;��H;��H;��H;~�H;Z�H;      ��H;��H;
�H;_�H;��H;O�H;��H;��H;�H;��H;��H;�H;8�H;^�H;Q�H;L�H;/�H;��H;��H;g�H;�H;��H;v�H;��H;��H;H�H;�H;��H;e�H;$�H;��H;��H;��H;��H;`�H;C�H;8�H;F�H;]�H;��H;��H;��H;��H;#�H;^�H;��H;�H;Q�H;��H;��H;|�H;��H;�H;b�H;��H;��H;/�H;L�H;N�H;a�H;9�H;�H;��H;��H;�H;��H;��H;A�H;��H;e�H;�H;��H;      ��H;�H;	�H;Y�H;��H;:�H;��H;��H;��H;��H;��H;��H;�H;��H;��H;�H;�H;��H;��H;��H;I�H;��H;��H;U�H;��H;��H;3�H;��H;��H;a�H;+�H;��H;��H;��H;��H;��H;v�H;��H;��H;��H;��H;��H;.�H;b�H;��H;��H;3�H;��H;��H;N�H;��H;��H;E�H;��H;��H;��H;�H;�H;��H;��H;�H;��H;��H;��H;��H;��H;��H;4�H;��H;Y�H;	�H;�H;      ��H;��H;f�H;8�H;�H;��H;.�H;g�H;�H;�H;�H;��H;��H;�H;��H;;�H;��H;��H;��H;��H;��H;J�H;��H;��H;W�H;��H;t�H;J�H;��H;��H;h�H;=�H;�H;��H;��H;��H;��H;��H;��H;��H;�H;=�H;j�H;��H;��H;G�H;t�H;��H;U�H;��H;��H;I�H;��H;��H;��H;��H;��H;;�H;��H;�H;��H;��H;�H;�H;�H;`�H;-�H;s�H;*�H;6�H;s�H;��H;      �H;H;�!H;�8H;�TH;5sH;"�H;��H;�H;��H;[�H;��H;��H;��H;��H;��H;��H;"�H;v�H;��H;��H;l�H;�H;��H;��H;E�H;��H;z�H;=�H;�H;��H;��H;T�H;6�H;!�H;��H;�H;��H;!�H;;�H;W�H;��H;��H;�H;9�H;w�H;��H;N�H;��H;��H; �H;n�H;��H;��H;v�H;�H;��H;��H;��H;��H;��H;��H;[�H;��H;~�H;��H;%�H;.sH;�TH;�8H;�!H;�H;      DF;,RF;�zF;ŸF;�G;�\G;ϲG;0H;�HH;c�H;g�H;��H;��H;��H;��H;�H;��H;�H;��H;0�H;u�H;d�H;W�H;1�H;��H;r�H;G�H;��H;��H;Q�H;�H;��H;��H;��H;f�H;S�H;e�H;U�H;e�H;��H;��H;��H;�H;T�H;��H;��H;I�H;{�H;��H;1�H;[�H;e�H;r�H;1�H;��H;�H;��H;�H;��H;��H;��H;��H;g�H;c�H;�HH;)H;ѲG;y\G;�G;ʸF;~zF;RF;      ��A;BB;�oB;�C;Y�C;Y�D;DuE;MDF;#�F;p�G;�H;�eH;�H;��H;5�H;��H;��H;��H;q�H;q�H;�H;I�H;e�H;V�H;�H;��H;��H;Y�H;��H;��H;`�H;0�H;��H;��H;��H;��H;��H;��H;��H;��H;��H;3�H;g�H;��H;��H;W�H;��H;��H;�H;T�H;i�H;J�H;�H;r�H;r�H;��H;��H;��H;7�H;��H;�H;�eH;�H;o�G;�F;MDF;BuE;L�D;b�C;�C;�oB;BB;      Fo8;$�8;��9;w�:;{�<;�c>;5R@;�/B;��C;�PE;ozF;D\G;o�G;iH;�H;��H;�H;E�H;�H;�H;@�H;��H;C�H;T�H;O�H;'�H;��H;��H;S�H;��H;��H;��H;F�H;�H;�H;�H;��H;�H;�H;�H;J�H;��H;��H;��H;S�H;��H;��H;.�H;L�H;V�H;H�H;��H;@�H;�H;�H;C�H;�H;��H;�H;iH;o�G;A\G;pzF;�PE;��C;�/B;4R@;�c>;��<;��:;��9;�8;      eS%;�%;��';�M*;ڷ-;��1;��5;�9;x-=;R@;��B;f�D;mF;�uG;^!H;��H;��H;~�H;��H;m�H;��H;�H;��H;J�H;e�H;T�H;�H;��H;��H;v�H;
�H;��H;��H;�H;n�H;Y�H;=�H;X�H;m�H;��H;��H;��H;�H;}�H;��H;��H;�H;[�H;b�H;I�H;��H;�H;��H;q�H;��H;{�H;��H;��H;^!H;�uG;
mF;f�D;��B;R@;r-=;��9;ޟ5;��1;ڷ-;�M*;��';��%;      nW;xx;��;�
;��;�;�� ;x�(;��/;�H6;��;;��?;�C;�PE;��F;��G;�eH;+�H;k�H;�H;/�H;��H;�H;��H;I�H;a�H;k�H;M�H;��H;��H;��H;-�H;��H;��H;��H;��H;��H;��H;��H;��H;��H;0�H;��H;��H;��H;L�H;l�H;h�H;E�H;��H;�H;��H;2�H;�H;k�H;*�H;�eH;��G;��F;�PE;�C;��?;��;;�H6;��/;x�(;�� ;r;��;�
;��;nx;      ���:Ɔ:�ɒ:'��:��:��::��:P�	;�v;��#;ķ-;��5;�L<;e�@;�(D;DF;��G;�HH;P�H;��H;��H;,�H;��H;@�H;�H;k�H;��H;��H;A�H;�H;��H;��H;S�H;I�H;�H;�H;�H;�H;�H;E�H;U�H;��H;��H;�H;A�H;��H;��H;n�H; �H;A�H;��H;,�H;��H;��H;P�H;�HH;��G;DF;�(D;e�@;�L<;��5;ķ-;�#;�v;S�	;:��:���:�:-��:�ɒ:�ņ:      t-.����p��0~K�� 
9\]:P�k:kM�:���:�y;��;� $;��/;n�8;��>;�#C;
�E;_\G;48H;��H;��H;�H;o�H;�H;n�H;.�H;��H;��H;��H;`�H;�H;��H;��H;��H;}�H;r�H;^�H;t�H;|�H;��H;��H;��H;"�H;d�H;��H;��H;��H;3�H;k�H;�H;q�H;�H;��H;��H;48H;_\G;�E;�#C;��>;j�8;��/;~ $;��;�y;���:[M�:8�k:<]:� 
9�~K�p����      "Q^�X��F�¢)�+��ζ�8�<��>S�Pn:)��:Ž�:��;?�;�M*;ڟ5;zc=;QpB;��E;�JG;38H;P�H;j�H;��H;�H;j�H;��H;o�H;��H;��H;��H;v�H;[�H;7�H;��H;��H;��H;��H;��H;��H;��H;7�H;]�H;z�H;��H;��H;��H;s�H;��H;d�H;�H;��H;h�H;P�H;48H;�JG;��E;QpB;uc=;؟5;�M*;=�;��;Ž�:'��:Dn:�>S�D�<��ζ�+���)��F�	X�      X���(������ѻ���ǐ�QX�6�4	�� uK�?":�M�:8b�:Pi;'�%;P�3;�<;-0B;��E;[\G;�HH;'�H;{�H;B�H;��H;�H;�H;��H;��H;��H;��H;��H;��H;E�H;5�H;5�H;�H;7�H;4�H;C�H;��H;��H;��H;��H;��H;��H;�H;�H;��H;@�H;}�H;%�H;�HH;]\G;��E;-0B;�<;M�3;'�%;Oi;8b�:�M�: ?": uK�4	��6�VX�ǐ�����ѻ ��*���      l�n�umj���]���J�U�1�04�0������	x��W�$�y��(
9���:F��:�;>�#;A�2;�<;OpB;�E;��G;�eH;��H;�H;��H;��H;��H;��H;�H;'�H;�H;��H;��H;��H;��H;��H;��H;��H;��H;��H;��H;��H;�H;+�H;�H;��H;��H;��H;��H;�H;��H;�eH;��G;�E;OpB;�<;?�2;<�#;�;F��:���:�(
9(�y��W��	x����2��04�W�1���J���]�tmj�      =<ͼ}�ɼ�����֯�̶��ㄼ��Y��*�����s��X�xrѺ0�?Q:���:��
;8�#;O�3;uc=;�#C;DF;��G;��H;��H;��H;�H;��H;4�H; �H;D�H;q�H;G�H;�H;6�H;��H;��H;��H;��H;��H;1�H;�H;D�H;s�H;I�H;�H;8�H;��H;�H;��H;��H;��H;��G;DF;�#C;tc=;M�3;:�#;��
;���:?Q:P�|rѺX��s������*���Y�ㄼͶ���֯�����}�ɼ      ��'�'�$����{��  ���ۼ����+����]��X!�>>ۻ�+��u*�(����>:���:��;"�%;ҟ5;��>;�(D;��F;_!H;�H;-�H;��H;��H;��H;��H;M�H;��H;��H;j�H;q�H;J�H;2�H;Q�H;4�H;I�H;p�H;j�H;��H;��H;N�H;��H;��H;��H;��H;*�H;�H;\!H;��F;�(D;��>;П5;!�%;��;���:��>:@��w*��+��@>ۻ�X!���]��+�������ۼ�  �{����'�$�      Ÿ���v����w�e�c��J�̈́-�{��;缃沼ㄼ��;������j���5���?Q:D��:Pi;�M*;j�8;l�@;�PE;�uG;iH;��H;��H;��H;��H;��H;W�H;��H;��H;��H;��H;��H;��H;��H;��H;��H;��H;��H;��H;��H;\�H;��H; �H;��H;��H;��H;iH;�uG;�PE;c�@;n�8;�M*;Ri;F��:?Q:(�깟5��j��������;�ㄼ�沼�;�{�̄-��J�e�c���w��v��      xHͽ֪ɽ�;��"����Ǹ����[�z0�r��$<ͼɾ��`�J�����j��s*� ����::b�:;�;��/;�L<;�C;
mF;p�G;ߡH;��H;��H;��H;�H;4�H;��H;�H;�H;��H;��H;��H;��H;��H;��H;��H;�H;�H;��H;6�H; �H;��H;��H;��H;ݡH;o�G;mF;�C;|L<;��/;9�;:b�:���:0�s*��j�����`�J�ɾ��$<ͼr��z0���[�Ǹ����"���;��ժɽ      ��!-������б�ƽ\P���v���J�F����ۼ
��`�J������+��vrѺ�(
9�M�:��;| $;��5;��?;f�D;C\G;�eH;��H;��H;��H;��H;��H;��H;2�H;U�H;=�H;3�H;D�H;�H;G�H;3�H;=�H;T�H;2�H;��H;�H;��H;��H;��H;��H;�eH;A\G;h�D;��?;��5;~ $;��;�M�:�(
9|rѺ�+������a�J�����ۼF���J��v��\P��ƽѱ轂����!-�       j�Vde�Y0X�D�e{+�������t㻽Y���QDX������ۼɾ����;�@>ۻX�P�y��>":���:��;Ʒ-;��;;��B;ozF;�H;a�H;T�H;��H;��H;��H;��H;M�H;��H;~�H;q�H;��H;]�H;��H;r�H;~�H;��H;M�H;��H;��H;��H;�H;T�H;`�H;�H;ozF;��B;��;;��-;��;���:�>":D�y�X�B>ۻ��;�ʾ����ۼ���QDX�Y���t㻽��콂��e{+�D�Y0X�Vde�      ��Ph��k���I���|x���O��C(��Ϊɽ����QDX�F��%<ͼㄼ�X!��s���W��uK�!��:�y;�#;�H6;R@;�PE;l�G;]�H;��H;�H;��H;��H;��H;R�H;��H;��H;��H;��H;��H;��H;��H;��H;��H;R�H;��H;��H;��H;
�H;��H;]�H;h�G;�PE;R@;�H6;��#;�y;��:puK��W��s���X!�ㄼ%<ͼF��QDX�����Ϊɽ��C(���O��|x��I��k��Ph��      =����������"�;hɰ��G��	 j�8�5��	�ΪɽX����J�r���沼��]�����	x�P	��(n:���:�v;��/;j-=;��C;�F;�HH;z�H;��H;��H;�H;~�H;f�H;��H;��H;��H;��H;�H;��H;��H;��H;��H;g�H;}�H;�H;��H;��H;|�H;�HH;�F;��C;k-=;��/;�v;���:$n:H	���	x������]��沼r���J�X���Ϊɽ�	�8�5�	 j��G��hɰ�"�;��徶���      �2�U�-�"�-E�����?Kɾj����s�8�5���t㻽�v��z0��;��+���*����16� AS�QM�:S�	;r�(;��9;�/B;KDF; H;��H;\�H;��H;��H;N�H;c�H;��H;�H;�H;�H;:�H;�H;�H;�H;��H;b�H;M�H;��H;��H;]�H;��H;#H;JDF;�/B;��9;t�(;M�	;[M�:@AS�+6�����*��+���;�z0��v��t㻽��8�5���s�j��?Kɾ����-E�"�U�-�      %3s�cm�:�\�g�C�5�%����TҾj��	 j��C(����]P����[�{������Y�5��aX�X�<��k::��:�� ;؟5;2R@;8uE;ϲG;�H;�H;��H;��H;#�H;G�H;	�H;D�H;N�H;9�H;n�H;7�H;O�H;A�H;�H;G�H;!�H;��H;��H;"�H;�H;ղG;6uE;4R@;ܟ5;�� ;2��: �k:X�<�^X�4����Y����{���[�]P����콪C(�	 j�j���TҾ��5�%�g�C�:�\�cm�      �ޞ�������_F�>�W�W�-���?Kɾ�G����O����ƽǸ��̈́-���ۼㄼ24�ǐ��ζ�4]:���:;��1;�c>;E�D;x\G;*sH;w�H;5�H;G�H; �H;M�H;�H;K�H;k�H;]�H;��H;^�H;k�H;H�H;
�H;M�H;��H;H�H;:�H;{�H;.sH;�\G;E�D;�c>;��1;;���:@]:�ζ�ǐ�24�ㄼ��ۼ̈́-�Ǹ��ƽ�����O��G��?Kɾ��W�-�>�W�_F�������      ��ſ���Lw���ޞ�����>�W�5�%�����hɰ��|x�e{+�ѱ����J��  �Ͷ��W�1�(���+�� 
9��:��;�-;��<;^�C;�G;�TH;#�H;��H;��H;��H;+�H;�H;h�H;��H;v�H;��H;r�H;��H;c�H;�H;+�H;��H;��H;��H;(�H;�TH;�G;]�C;��<;�-;��;��:� 
9+�%���W�1�Ͷ���  ��J���ѱ�e{+��|x�hɰ�����5�%�>�W������ޞ�Lw�����      ������Կp���ޞ�_F�g�C�-E�"�;�I��D���"��e�c�{��֯���J��ѻɢ)�PK�#��:�
;�M*;n�:;�C;ȸF;�8H;-�H;H�H;Z�H;��H;�H;�H;��H;��H;��H;��H;��H;��H;}�H;�H;�H;��H;a�H;M�H;.�H;�8H;ӸF;�C;n�:;�M*;�
;#��:K�ʢ)��ѻ��J��֯�{�e�c�"����D��I��"�;-E�g�C�`F��ޞ�p���Կ��      ����������ԿLw�����:�\�"����k��Y0X�����;����w����������]����F�����ɒ:��;�';��9;�oB;�zF;�!H;t�H;��H;�H;r�H;�H;�H;��H;��H;��H;��H;��H;��H;�H;�H;�H;n�H;	�H;��H;w�H;�!H;�zF;�oB;��9; �';��;�ɒ:����F��黨�]����������w��;�����Y0X�k�����"�:�\����Lw���Կ��𿝏�       $�������忇�����cm�U�-�����Ph��Vde�!-�֪ɽ�v��'�$�~�ɼxmj�4���X����ņ:jx;�%;4�8;HB; RF;�H;�H;�H;��H;E�H;�H;�H;v�H;��H;��H;�H;��H;��H;v�H;�H;�H;A�H;��H;�H;�H; H;.RF;EB;2�8;�%;hx;�ņ:���X�2���xmj�~�ɼ'�$��v��֪ɽ!-�Vde�Ph������U�-�cm��������忝����      �>���8���*�O������˿p��E�b�C\�4m־^��Q�:��J�(��D�B�;��������-/��F�����>:wt�:p ;�J6;�DA;^IF;�NH;��H;�!I;�I;�I;|I;NI;�I;I I;��H;	�H;��H;H I;�I;NI;|I;�I;�I;�!I;��H;�NH;kIF;�DA;�J6;p ;ut�:��>:<���-/���������;��D�B�(���J�Q�:�^��4m־C\�E�b�p���˿����O���*���8�      ��8��4��g&�6��<����<ƿ񲗿�>]����O�Ѿ�p���*7����$W��KR?��|�p8�������ʅ����G: �:�!;�6;�kA;iYF;�TH;G�H;�!I;�I;�I;eI;(I;�I;; I;��H;��H;��H;; I;�I;)I;gI;�I;�I;�!I;I�H;�TH;tYF;�kA;�6;�!;{ �:��G:�������p8���|�KR?�$W�����*7��p��O�Ѿ����>]�񲗿�<ƿ<���6���g&��4�      ��*��g&��#�t�T[�qL�������M�r5��>ľ����,��D�蒐��5�0�ݼ���q
��x�uk���b:3l�:�#;Ǘ7;X�A;��F;�dH;�I;%"I;�I;GI;I;�I;�I;��H;Y�H;��H;R�H;��H;�I;�I;I;AI;�I;&"I;�I;�dH;��F;W�A;×7;�#;1l�:��b:�tk��x��q
���0�ݼ�5�蒐��DὪ�,����>ľr5���M����qL��T[�t��#��g&�      O�6��t����˿@1��7�y�Î6��z �����2�l�+��ͽ"�����&���˼<�k������X�� �~��:<�;�&;�9;o�B;��F;�}H;�	I;2"I;I;�I;{I;UI;%I;��H;�H;a�H;��H;��H;"I;RI;{I;�I;I;5"I;�	I;�}H;��F;m�B;~9;�&;<�;|��:ԙ ���X����<�k���˼��&�"����ͽ+�2�l������z �Î6�7�y�@1���˿���t�6��      ����<���T[忶˿�T���{�R�����E۾җ����M���	������j��3�d����O�8�׻��/�0��G��:� 
;�*;S;;�jC;�'G;כH;�I;�!I;�I;wI;�
I;�I;�I;!�H;��H;��H;��H;"�H;�I;�I;�
I;sI;�I;�!I;�I;ڛH;�'G;�jC;N;;�*;� 
;E��:�����/�6�׻��O�d���3���j������	���M�җ���E۾���{�R���T���˿T[�<���      �˿�<ƿqL��@1����>]���)��$��ֳ���{���,�q��'��P`I��J���,���3/��+��� �0-69�4�:ք;�o.;.=;BaD;��G;T�H;�I;!I;AI;,I;�	I;�I;� I;��H;��H;C�H;��H;��H;� I;�I;�	I;)I;CI;!I;�I;S�H;��G;@aD;.=;�o.;Ԅ;�4�:`-69� ��+���3/��,���J��P`I�&��q�齤�,���{�ֳ��$����)��>]��@1��qL���<ƿ      p��񲗿���7�y�{�R���)�nv��>ľ^���I�Xl����������&�ҮҼ�}�0B�Ȯ�������!:�*�:&z;^3;Mj?;v\E;��G;��H;KI;I;mI;�I;XI;�I;��H;��H;C�H;��H;A�H;��H;��H;�I;WI;�I;pI;I;KI;��H;��G;v\E;Ij?;\3;&z;�*�:��!:���Ȯ��/B��}�ҮҼ��&��������Xl��I�^���>ľnv���)�{�R�7�y����񲗿      E�b��>]���M�Î6�����$���>ľ#q��y�Z�+�Q9ݽ W����L����!F���G�
�׻ ;�o칄Ȋ:�i;P$;��7;W�A;�IF;CH;��H;� I;EI;WI;�I;	I;�I;��H;��H;t�H;��H;r�H;��H;��H;I;I;�I;ZI;EI;� I;��H;CH;�IF;S�A;��7;P$;�i;�Ȋ:o��;��׻ �G� F�������L� W��P9ݽ+�y�Z�#q���>ľ�$�����Î6���M��>]�      C\����q5��z ��E۾ֳ�^��y�Z�K?#����A����j�$��Cϼ �����ǵ���lۺ�9�9h4�:D�;G�,;[�;; �C;�G;"�H;�I;�!I;�I;%I;I;sI;$I;��H;��H;��H;�H;��H;��H;��H;#I;sI;I;'I;�I;�!I;�I;"�H;�G;�C;\�;;J�,;A�;z4�:�9�9�lۺƵ����� ��Cϼ$����j��A�����K?#�y�Z�^��ֳ��E۾�z �q5����      4m־O�Ѿ�>ľ����җ����{��I�+����V���{�=�/�#���,��==�@�һg�@�8� ���k:��:�a;��3;j?;T2E;��G;C�H;I;P I;�I;�I; 	I;�I;��H;��H;��H;��H;9�H;��H;��H;��H;��H;�I; 	I;�I;�I;Q I;I;A�H;��G;P2E;j?;��3;�a;��:��k:,� �c�@�>�һ<=��,��#��=�/��{��V�����+��I���{�җ�������>ľO�Ѿ      ^���p����2�l���M���,�Xl�P9ݽ�A���{���5��J��;���T[� ?�����VP��(P�9��:��;*;�9;7kB;��F;WNH;X�H; I;iI;�I; I;�I;!I;F�H;��H;��H;��H;I�H;��H;��H;��H;D�H;!I;�I;I;�I;lI;�I;V�H;[NH;��F;8kB;�9;*;��;��:8P�9FP������ ?��T[�;���J����5��{��A��P9ݽXl���,���M�1�l����p��      P�:��*7���,�+���	�q�齁��� W����j�=�/��J���I���k�j�
.��_�� ���Ȋ:5o�:�;Fr3;�>;�D;P�G;$�H;�I;!I;�I;cI;b
I;�I;A I;��H;z�H;��H;��H;A�H;��H;��H;|�H;��H;? I;�I;g
I;mI;�I;!I;�I;(�H;O�G;	�D;�>;Gr3;�;7o�:�Ȋ:� ��[��	.��h��k��I���J��=�/���j� W������p�齂�	�+���,��*7�      �J�����D��ͽ���&�������L�$��"��;���k����gI����/��/�0�>:)��:�B;C�,;��:;�B;mxF;x<H;��H;�I;tI;�I;I;�I;�I;p�H;Z�H;�H;O�H;�H;N�H;�H;N�H;�H;W�H;n�H;�I;�I;I;�I;sI;�I;��H;v<H;nxF;�B;��:;N�,;�B;#��:L�>:x/���/�fI������k�;��#��$����L����&������ͽ�D����      '��$W��璐�"�����j�Q`I���&����Cϼ�,���T[�i�hI��];��nk��:�4�:�;�&;��6;�!@;2E;��G;��H;�I;� I;2I;�I;�
I;I;Q I;��H;��H;��H;@�H;v�H;'�H;v�H;@�H;��H;��H;��H;V I;I;�
I;�I;0I;� I;�I;�H;��G;2E;�!@;��6;�&;�;5�:�:�nk�Y;�gI��h��T[��,��Bϼ�����&�P`I���j�"���璐�$W��      C�B�KR?��5���&��3��J��ѮҼF�� ��<=�?�
.����/��nk� ��9*׳:��;$!;?3;��=;��C;��F;�cH;��H;oI;�I;�I;I;�I;�I;"�H;��H;r�H;`�H;!�H;g�H;�H;e�H; �H;b�H;u�H;��H;%�H;�I;�I;I;�I;�I;qI;��H;�cH;�F;��C;��=;C3; !;��;.׳: ��9�nk���/�
.��?�<=���� F��ѮҼ�J���3���&��5�KR?�      7���|�.�ݼ��˼d���,���}���G����>�һ����^���/��:0׳:��;Vb;��0;r<;��B;�IF;LH;�H;�I;P I;�I;I;9
I;�I; I;�H;8�H;��H;�H;�H;]�H;�H;\�H;�H;�H;��H;6�H;�H; I;�I;=
I;I;�I;Q I;�I;�H;OH;�IF;��B;u<;��0;Yb;�;4׳:�:�/�^������=�һ�����G��}��,��d����˼.�ݼ�|�      ~���n8����<�k���O��3/�-B��׻õ��\�@�>P��� ��L�>:5�:��;Zb;��/;;;!�A;j�E;��G;ҭH;�
I;H I;�I;�I;�I;�I;�I;f�H;�H;��H;}�H;��H;��H;Q�H;�H;M�H;��H;��H;x�H;��H;�H;i�H;�I;�I;�I;�I;�I;G I;�
I;խH;��G;q�E;$�A;;;��/;Zb;��;5�:D�>:� ��:P��\�@������׻.B��3/���O�=�k���m8��      ������q
����0�׻�+��®���;��lۺ� �HP�9�Ȋ:��:�;$!;��0;;;��A;�pE;S�G;��H;��H;�I;I;0I;I;�I;VI;��H;#�H;X�H;��H; �H;��H;��H;G�H;�H;D�H;��H;��H;��H;��H;[�H;(�H;��H;VI;�I;�I;3I;I;�I;��H;��H;X�G;�pE;��A;;;��0;"!;�;��:�Ȋ:�P�9� ��lۺ�;�Į���+��-�׻����q
���       /������x���X���/�� ������n��9�9ĩk:��:;o�:�B;�&;C3;u<;#�A;�pE;GtG;�|H;�H;I;UI;&I;�I;N
I;�I;3 I;-�H;�H;��H;`�H;��H;��H;��H;X�H;E�H;W�H;��H;��H;��H;]�H;��H;�H;-�H;5 I;�I;J
I;�I;&I;OI;	I;�H;�|H;GtG;�pE;%�A;r<;D3;�&;�B;;o�:��:��k:�9�9�n����� ���/���X��x����      <���ʅ���tk��� � ���-69��!:�Ȋ:z4�:��:��;�;H�,;��6;��=;��B;q�E;]�G;�|H;x�H;ZI;�I;eI;<I;�I;I;jI;*�H;��H;�H;��H;��H;��H;��H;��H;n�H;U�H;j�H;��H;��H;��H;��H;��H;�H;��H;-�H;fI;I;�I;9I;bI;�I;]I;x�H;�|H;W�G;o�E;��B;��=;��6;H�,;�;��;��:�4�:�Ȋ:��!:�-69���̙ �uk�䅍�      ��>:\�G:|�b:z��:1��:�4�:�*�:�i;A�;�a;*;Cr3;��:;�!@;��C;�IF;��G;��H;�H;WI;  I;"I;I;�I;�I;?I;�H;p�H;��H;[�H;*�H;��H;}�H;��H;��H;��H;c�H;��H;��H;��H;y�H;��H;-�H;^�H;��H;n�H;��H;:I;�I;�I;I;$I; I;WI;�H;��H;��G;�IF;��C;�!@;��:;Dr3;*;�a;A�;�i;�*�:�4�:G��:t��:��b:\�G:      qt�:� �:Ml�:P�;� 
;ڄ;(z;P$;P�,;��3;�9;�>;�B;2E;�F;VH;ۭH;��H;I;�I;&I;^I;I;�I;�I;��H;�H;3�H;��H;{�H;��H;��H;t�H;��H;�H;��H;��H;��H;�H;��H;o�H;��H;��H;{�H;��H;3�H;��H;��H;�I;�I;I;`I;&I;�I;I;��H;ۭH;RH;�F;2E;�B;�>;�9;��3;P�,;P$;,z;ք;� 
;F�;5l�:� �:      .p ;�!;�#;�&;�*;�o.;m3;��7;c�;;j?;@kB;�D;qxF;��G;�cH;�H;�
I;�I;UI;cI;I;I;�I;=I;�H;t�H;s�H;�H;��H;��H;��H;d�H;u�H;��H;9�H;�H;��H;��H;5�H;��H;q�H;c�H;��H;��H;��H;�H;n�H;t�H;�H;9I;�I;I;I;cI;SI;�I;�
I;
�H;�cH;��G;qxF;�D;CkB;j?;f�;;��7;j3;�o.;�*;�&;�#;�!;      �J6;�6;��7;~9;E;;.=;Mj?;T�A;�C;T2E;��F;S�G;x<H;��H;��H;�I;K I;I;(I;9I;�I;�I;=I;3�H;��H;��H;D�H;�H;!�H;��H;k�H;V�H;x�H;�H;��H;W�H;-�H;Q�H;��H;�H;v�H;T�H;k�H;��H;�H;�H;=�H;��H;��H;/�H;4I;�I;�I;6I;%I;I;G I;�I;��H;�H;u<H;Q�G;��F;Q2E;�C;[�A;Hj?;.=;S;;~9;��7;�6;      EA;�kA;O�A;k�B;�jC;PaD;~\E;�IF;�G;��G;bNH;0�H;��H;�I;xI;[ I;�I;<I;�I;�I;�I;�I;�H;��H;��H;d�H;�H;2�H;��H;|�H;O�H;h�H;��H;B�H;��H;��H;��H;��H;��H;E�H;��H;b�H;Q�H;{�H;��H;2�H;�H;c�H;��H;��H;�H;�I;�I;�I;�I;7I;�I;Z I;tI;�I;��H;0�H;dNH;��G;�G;�IF;~\E;FaD;�jC;m�B;M�A;�kA;      [IF;sYF;��F;��F;v'G;��G;��G;CH;#�H;I�H;]�H;�I;�I;� I;�I;�I;�I;I;M
I;I;=I;��H;r�H;��H;_�H;;�H;G�H;��H;�H;_�H;I�H;��H;�H;��H;9�H;�H;�H;�H;4�H;��H;�H;��H;I�H;\�H;{�H;��H;A�H;?�H;c�H;��H;q�H;��H;?I;I;M
I;�I;�I;�I;�I;� I;�I;�I;a�H;J�H;&�H;CH;��G;��G;�'G;��F;��F;pYF;      �NH;�TH;�dH;�}H;ϛH;T�H;��H;��H;�I;I; I;!I;qI;3I;�I;I;�I;�I;�I;jI;�H;�H;s�H;G�H;�H;C�H;��H;��H;Q�H;P�H;��H;��H;W�H;��H;��H;��H;z�H;��H;��H;��H;V�H;��H;��H;M�H;J�H;��H;��H;H�H;�H;C�H;p�H;�H;�H;hI;�I;�I;�I;I;�I;/I;qI;!I; I;I;�I;��H;��H;O�H;�H;�}H;�dH;{TH;      ��H;L�H;�I;�	I;�I;�I;VI;� I;�!I;X I;oI;�I;�I;�I;I;=
I;�I;SI;4 I;(�H;n�H;.�H;	�H;�H;+�H;��H;�H;`�H;G�H;w�H;��H;4�H;��H;t�H;6�H;�H;��H;�H;3�H;u�H;��H;2�H;��H;v�H;B�H;_�H;{�H;��H;/�H;�H;	�H;0�H;m�H;'�H;1 I;PI;�I;=
I;�I;�I;�I;�I;pI;U I;�!I;� I;WI;�I;�I;�	I;�I;@�H;      �!I;�!I;"I;D"I;�!I;!I;�I;II;�I;�I;�I;qI;"I;�
I;�I;�I;�I;��H;3�H;��H;��H;��H;��H;�H;��H;v�H;G�H;G�H;��H;��H;&�H;��H;D�H;��H;��H;��H;��H;��H;��H;��H;C�H;��H;%�H;��H;��H;F�H;C�H;v�H;��H;�H;��H;��H;��H;��H;1�H;��H;�I;�I;�I;�
I;I;mI;�I;�I;�I;II;�I;!I;�!I;D"I;!"I;�!I;      �I;I;�I;I;�I;?I;nI;]I;(I;�I;I;n
I;�I;!I;�I; I;o�H;"�H;�H;!�H;_�H;v�H;��H;��H;x�H;V�H;L�H;z�H;��H;�H;��H;?�H;��H;��H;c�H;C�H;2�H;C�H;_�H;��H;��H;=�H;��H;�H;��H;v�H;F�H;X�H;y�H;��H;��H;y�H;[�H;�H;�H;!�H;o�H; I;�I; I;�I;j
I;I;�I;'I;ZI;tI;?I;�I;I;�I;I;      �I;�I;LI;�I;vI;,I;�I;I;I;	I;�I;�I;�I;[ I;+�H;�H;%�H;`�H;��H;��H;3�H;��H;��H;k�H;N�H;I�H;��H;��H;,�H;��H;�H;��H;p�H;4�H;�H;��H;��H;��H;�H;6�H;p�H;��H;�H;��H;%�H;��H;��H;I�H;Q�H;j�H;��H;��H;0�H;��H;��H;^�H;'�H;�H;(�H;Z I;�I;�I;�I;	I;I;I;�I;%I;�I;�I;NI;�I;      }I;pI;I;vI;�
I;�	I;[I;I;zI;�I;%I;F I;t�H;��H;��H;<�H;��H;��H;e�H;��H;��H;��H;c�H;R�H;e�H;��H;��H;7�H;��H;A�H;��H;N�H;�H;��H;��H;��H;��H;��H;��H;��H;�H;M�H;��H;@�H;��H;2�H;��H;��H;h�H;N�H;g�H;��H;��H;��H;d�H;��H;��H;?�H;��H;��H;r�H;F I;(I;�I;xI;
I;bI;�	I;�
I;yI;I;oI;      YI;6I;�I;XI;�I;�I;�I;I;I;��H;H�H;��H;\�H;��H;w�H;��H;��H;�H;��H;��H;��H;u�H;t�H;v�H;��H;�H;W�H;��H;K�H;��H;m�H;�H;��H;��H;��H;g�H;`�H;g�H;��H;��H;��H;�H;l�H;��H;G�H;��H;U�H;�H;��H;v�H;z�H;u�H;��H;��H;��H;�H;��H;��H;y�H;��H;\�H;��H;K�H;��H;!I;~I;�I;�I;�I;RI;�I;6I;      �I;�I;�I;I;�I;� I;��H;��H;��H;��H;��H;��H; �H;��H;g�H;�H;��H;��H;��H;��H;��H;��H;��H;�H;<�H;{�H;��H;w�H;��H;��H;1�H;��H;��H;g�H;Q�H;B�H;4�H;C�H;P�H;i�H;��H;��H;2�H;��H;��H;r�H;��H;{�H;A�H;�H;��H;��H;��H;��H;��H;��H;��H;�H;g�H;��H;�H;��H;��H;��H;�H;��H; I;� I;�I; I;�I;�I;      B I;P I; I;��H;0�H;{�H;��H;��H;��H;��H;��H;��H;Z�H;K�H;-�H;�H;��H;��H;��H;��H;��H;�H;5�H;��H;��H;/�H;��H;5�H;��H;e�H; �H;��H;��H;P�H;.�H;�H;#�H; �H;*�H;S�H;��H;��H; �H;b�H;��H;2�H;��H;0�H;��H;��H;9�H;�H;��H;��H;��H;��H; �H;�H;+�H;K�H;Z�H;��H;��H;��H;��H;��H;��H;|�H;0�H;��H;  I;Q I;      ��H;��H;X�H;�H;��H;��H;M�H;{�H;��H;��H;��H;��H;��H;z�H;k�H;]�H;R�H;C�H;Z�H;n�H;��H;��H;��H;E�H;��H;�H;��H;�H;��H;I�H;��H;��H;l�H;B�H;#�H;�H;�H;�H; �H;H�H;n�H;��H;��H;D�H;��H;�H;��H;�H;��H;F�H;�H;��H;��H;j�H;[�H;J�H;V�H;a�H;i�H;}�H;��H;��H;��H;��H;��H;y�H;T�H;��H;��H;�H;T�H;��H;      �H;��H;��H;f�H;��H;>�H;��H;��H;�H;9�H;V�H;L�H;V�H;1�H;"�H;!�H;�H;�H;I�H;\�H;m�H;��H;��H;"�H;��H;��H;u�H;��H;��H;9�H;��H;��H;d�H;3�H;%�H;�H;�H;�H;"�H;4�H;h�H;��H;��H;4�H;��H;��H;u�H;�H;��H;#�H;��H;��H;g�H;W�H;I�H;$�H;�H;%�H; �H;4�H;Y�H;K�H;W�H;<�H;�H;��H;��H;?�H;��H;j�H;��H;��H;      ��H;��H;R�H;�H;��H;��H;L�H;x�H;��H;��H;��H;��H;��H;}�H;k�H;]�H;U�H;C�H;Z�H;n�H;��H;��H;��H;E�H;��H;�H;��H;�H;��H;I�H;��H;��H;n�H;C�H;#�H;�H;�H;�H; �H;F�H;n�H;��H;��H;B�H;��H;��H;��H;�H;��H;F�H;�H;��H;��H;j�H;[�H;L�H;U�H;c�H;i�H;}�H;��H;��H;��H;��H;��H;{�H;T�H;��H;��H;�H;Y�H;��H;      7 I;P I;��H;��H;/�H;x�H;��H;��H;��H;��H;��H;��H;\�H;K�H;.�H;�H;��H;��H;��H;��H; �H;�H;5�H;��H;��H;,�H;��H;5�H;��H;c�H;��H;��H;��H;P�H;-�H;�H;#�H;"�H;,�H;Q�H;��H;��H;��H;_�H;��H;/�H;��H;0�H;��H;��H;9�H;�H;��H;��H;��H;��H; �H;�H;*�H;M�H;\�H;��H;��H;��H;��H;��H;��H;w�H;4�H;��H; I;V I;      �I;�I;�I; I;�I;� I;��H;��H;��H;��H;��H;��H;�H;��H;i�H;�H;��H;��H;��H;��H;��H;��H;��H;�H;?�H;y�H;��H;w�H;��H;��H;/�H;��H;��H;h�H;Q�H;A�H;4�H;B�H;P�H;h�H;��H;��H;/�H;��H;��H;r�H;��H;|�H;A�H;�H;��H;��H;��H;��H;��H;��H;��H;�H;i�H;��H; �H;��H;��H;��H;�H;��H; I;� I;�I;"I;�I;�I;      VI;;I;�I;RI;�I;�I;�I;�I;!I;��H;H�H;��H;]�H;��H;z�H;��H;��H;�H;��H;��H;��H;v�H;t�H;v�H;��H;�H;U�H;��H;H�H;��H;i�H;�H;��H;��H;��H;g�H;`�H;g�H;��H;��H;��H;�H;j�H;��H;A�H;��H;V�H;�H;��H;s�H;{�H;u�H;~�H;��H;��H;�H;��H;��H;y�H;��H;^�H;��H;K�H;��H; I;�I;�I;�I;�I;]I;�I;6I;      rI;pI;I;rI;�
I;�	I;`I;I;wI;�I;(I;H I;t�H;��H;��H;=�H;��H;��H;d�H;��H;��H;��H;d�H;R�H;h�H;��H;��H;4�H;��H;?�H;��H;L�H;�H;��H;��H;��H;��H;��H;��H;��H;�H;M�H;��H;=�H;��H;2�H;��H;��H;e�H;K�H;k�H;��H;��H;��H;d�H;��H;��H;@�H;��H;��H;w�H;I I;)I;�I;{I;I;aI;�	I;�
I;xI;I;lI;      �I;�I;KI;�I;{I;,I;�I; I;I;	I;�I;�I;�I;] I;,�H;�H;'�H;`�H;��H;��H;4�H;��H;��H;k�H;R�H;C�H;��H;��H;*�H;��H;�H;��H;o�H;5�H;�H;��H;��H;��H;�H;6�H;p�H;��H;�H;��H;%�H;��H;��H;J�H;N�H;h�H;��H;��H;/�H;��H;��H;a�H;(�H;�H;,�H;] I;�I;�I;�I;	I;I;I;�I;*I;�I;�I;PI;�I;      �I;�I;�I;I;�I;MI;qI;bI;,I;�I;I;k
I;�I;!I;�I; I;o�H;#�H;�H;�H;a�H;x�H;��H;��H;{�H;R�H;I�H;w�H;��H;�H;��H;<�H;��H;��H;b�H;B�H;2�H;D�H;_�H;��H;��H;=�H;��H;�H;��H;v�H;I�H;Y�H;v�H;��H;��H;y�H;\�H;�H;�H;#�H;o�H; I;�I;#I;�I;j
I;I;�I;(I;`I;qI;?I;�I;'I; I;�I;      �!I;�!I;2"I;@"I;�!I;!I;�I;II;�I;�I;�I;oI; I;�
I;�I;�I;�I;��H;0�H;��H;��H;��H;��H; �H;��H;q�H;D�H;F�H;��H;��H;#�H;��H;C�H;��H;��H;��H;��H;��H;��H;��H;D�H;��H;%�H;��H;��H;C�H;F�H;x�H;��H;�H;��H;��H;��H;��H;4�H;��H;�I;�I;�I;�
I;!I;oI;�I;�I;�I;KI;�I;!I;�!I;C"I;2"I;�!I;      ��H;B�H;|I;�	I;�I;�I;WI;� I;�!I;X I;oI;�I;�I;�I;I;?
I;�I;SI;3 I;'�H;p�H;0�H;�H;�H;/�H;��H;{�H;]�H;G�H;u�H;��H;3�H;��H;t�H;3�H;�H;��H;�H;3�H;u�H;��H;3�H;��H;u�H;C�H;\�H;|�H;��H;+�H;�H;�H;0�H;k�H;(�H;5 I;RI;�I;?
I;I;�I;�I;�I;pI;X I;�!I;� I;YI;�I;�I;�	I;�I;B�H;      �NH;�TH;�dH;�}H;ߛH;[�H;��H;��H;�I;I; I;!I;qI;3I;�I;I;�I;�I;�I;hI;�H;�H;n�H;H�H;�H;@�H;��H;��H;O�H;L�H;��H;��H;V�H;��H;��H;��H;z�H;��H;��H;��H;W�H;��H;��H;M�H;K�H;�H;��H;J�H;�H;D�H;u�H;�H;�H;lI;�I;�I;�I;I;�I;2I;qI;!I; I;I;�I;��H;��H;W�H;�H;�}H;�dH;�TH;      OIF;sYF;��F;��F;}'G;ǈG;��G;CH;+�H;I�H;^�H;�I;�I;� I;�I;�I;�I;I;M
I;I;AI;��H;o�H;��H;b�H;8�H;D�H;��H;��H;\�H;I�H;��H;�H;}�H;9�H;�H;	�H;�H;6�H;��H;�H;��H;L�H;]�H;y�H;��H;D�H;A�H;_�H;��H;t�H;��H;?I;I;N
I;I;�I; I;�I;� I;�I;�I;a�H;J�H; �H;CH;��G;��G;�'G;��F;��F;dYF;      EA;�kA;M�A;g�B;�jC;RaD;�\E;�IF;�G;��G;dNH;3�H;��H;�I;{I;[ I;�I;<I;�I;�I;�I;�I;�H;��H;��H;[�H;�H;2�H;��H;y�H;O�H;f�H;��H;B�H;��H;��H;��H;��H;��H;C�H;��H;f�H;U�H;{�H;��H;/�H;�H;d�H;��H;��H;�H;�I;�I;�I;�I;:I;�I;^ I;{I;�I;��H;/�H;aNH;��G;�G;�IF;~\E;FaD;�jC;m�B;M�A;�kA;      �J6;�6;��7;�9;D;;".=;Kj?;Z�A;"�C;R2E;��F;T�G;v<H;��H;��H;�I;J I;I;&I;6I;�I;�I;6I;0�H;��H;��H;@�H;�H; �H;��H;k�H;U�H;w�H;�H;��H;S�H;.�H;T�H;��H;�H;{�H;V�H;o�H;��H;�H;�H;C�H;��H;��H;3�H;:I;�I;�I;9I;)I;I;L I;�I;��H;��H;u<H;P�G;��F;Q2E;�C;Q�A;Lj?;.=;Y;;�9;��7;�6;      p ;�!;�#;�&;�*;�o.;e3;��7;h�;;j?;>kB;�D;qxF;��G;�cH;�H;�
I;�I;UI;eI;I;I;�I;=I;�H;k�H;o�H;�H;��H;��H;��H;e�H;r�H;��H;8�H;�H;��H;�H;6�H;��H;w�H;g�H;��H;��H;��H;�H;r�H;t�H;�H;=I;�I;I;!I;hI;XI;�I;�
I;�H;�cH;��G;qxF;�D;>kB;j?;f�;;��7;e3;�o.;�*;�&;�#;�!;      ot�:� �:;l�:D�;� 
;�;,z;
P$;Q�,;��3;�9;
�>;�B;2E;�F;WH;ۭH;��H;I;�I;(I;`I;I;�I;�I;��H;�H;3�H;��H;y�H;��H;��H;o�H;��H;�H;��H;��H;��H;�H;��H;u�H;��H;��H;}�H;��H;1�H;�H;��H;�I;�I;I;cI;)I;�I;I;��H;٭H;UH;�F;2E;�B;�>;�9;��3;Q�,;
P$;$z;Ȅ;� 
;8�;;l�:� �:      P�>:��G:��b:~��:1��:�4�:�*�:�i;E�;�a;*;Fr3;��:;�!@;��C;�IF;��G;��H;�H;XI;  I;$I;I;�I;�I;6I;��H;m�H;��H;Z�H;,�H;��H;z�H;��H;��H;��H;d�H;��H;��H;��H;|�H;��H;0�H;^�H;��H;m�H;�H;=I;�I;�I;I;$I; I;[I;�H;��H;��G;�IF;��C;�!@;��:;Dr3;*;�a;D�;�i;�*�:�4�:S��:���:��b:x�G:      ��������tk��� � ��.69��!:�Ȋ:�4�:��:��;�;M�,;��6;��=;��B;r�E;[�G;�|H;z�H;]I;�I;cI;<I;�I;I;eI;*�H;��H;�H;��H;��H;��H;��H;��H;j�H;V�H;m�H;��H;��H;��H;��H;��H;�H;��H;*�H;iI;I;�I;@I;fI;�I;^I;{�H;�|H;Z�G;q�E;��B;��=;��6;J�,;�;��;��:�4�:�Ȋ:��!:�-69����� ��tk�����       /������x���X���/�� � ����n��9�9��k:��:7o�:�B;�&;H3;w<;$�A;�pE;GtG;�|H;�H;
I;UI;(I;�I;J
I;�I;4 I;.�H;�H;��H;^�H;��H;��H;��H;W�H;E�H;W�H;��H;��H;��H;^�H;��H;�H;-�H;4 I;�I;K
I;�I;*I;VI;I;�H;�|H;FtG;�pE;#�A;r<;F3;�&;�B;;o�:��:ĩk:�9�9�n����� ���/���X��x����      ������q
����,�׻�+��®���;��lۺ� �pP�9�Ȋ:��:�;&!;��0;;;��A;�pE;V�G;��H;��H;�I;I;6I;�I;�I;VI;��H;"�H;[�H;��H;��H;��H;��H;F�H;�H;G�H;��H;��H;��H;��H;]�H;#�H;��H;UI;�I;�I;0I;I;�I;��H;��H;X�G;�pE;��A;;;��0;$!;�;#��:�Ȋ:�P�9� ��lۺ�;�Į���+��.�׻����q
���      ~���n8����;�k���O��3/�-B��׻µ��\�@�8P��� ��L�>: 5�:��;[b;��/;;;!�A;n�E;��G;խH;�
I;H I;�I;�I;�I;�I;�I;e�H;�H;��H;z�H;��H;��H;O�H;�H;O�H;��H;��H;x�H;��H;�H;h�H;�I;�I;�I;�I;�I;H I;�
I;׭H;��G;q�E;!�A;;;��/;[b;��;5�:P�>:� ��>P��]�@������׻.B��3/���O�<�k���m8��      7���|�/�ݼ��˼d���,���}���G����>�һ����[���/��:6׳:��;Tb;��0;r<;��B;�IF;PH;
�H;�I;T I;�I;I;9
I;�I; I;�H;6�H;��H;�H;�H;\�H;�H;\�H;�H;�H;��H;4�H;�H; I;�I;:
I;I;�I;O I;�I;
�H;RH;�IF;��B;q<;��0;Wb;�;4׳:�:�/�_������>�һ�����G��}��,��d����˼0�ݼ�|�      D�B�KR?��5���&��3��J��ѮҼF�� ��<=�?�
.����/��nk� ��90׳:��;"!;A3;��=;��C;�F;�cH;��H;rI;�I;�I;I;�I;�I;%�H;��H;s�H;c�H;#�H;d�H;�H;e�H;!�H;b�H;s�H;��H;$�H;�I;�I;I;�I;�I;nI;��H;�cH;�F;��C;��=;?3;!;��;*׳:��9�nk���/�.��?�<=����F��ҮҼ�J���3���&��5�KR?�      '��$W��璐�"�����j�P`I���&����Bϼ�,���T[�h�gI��Y;��nk��:�4�:�;�&;��6;�!@;2E;��G;��H;�I;� I;0I;�I;�
I;I;V I;��H;��H;��H;A�H;t�H;'�H;w�H;?�H;��H;��H;��H;S I;I;�
I;�I;.I;� I;�I;��H;��G;2E;�!@;��6;�&;�;�4�:�:�nk�Z;�hI��i��T[��,��Bϼ�����&�P`I���j�"���璐�$W��      �J�����D��ͽ���&�������L�$��"��;���k����fI����/�x/�<�>:'��:�B;H�,;��:;�B;rxF;y<H;��H;�I;pI;�I; I;�I;�I;n�H;Y�H;�H;P�H;�H;N�H;�H;O�H;�H;V�H;m�H;�I;�I;!I;�I;oI;�I;��H;v<H;rxF;�B;��:;K�,;�B;#��:<�>:|/���/�gI������k�;��#��$����L����&������ͽ�D����      P�:��*7���,�+���	�p�齁��� W����j�=�/��J���I���k�i�	.��]�����Ȋ:5o�:�;Kr3;�>;�D;Q�G;)�H;�I;!I;�I;iI;b
I;�I;? I;��H;|�H;��H;��H;B�H;��H;��H;{�H;��H;> I;�I;d
I;mI;�I;!I;�I;$�H;P�G;�D;�>;Cr3;�;/o�:�Ȋ:� ��_��	.��j��k��I���J��=�/���j� W������p�齂�	�+���,��*7�      ^���p����1�l���M���,�Xl�P9ݽ�A���{���5��J��;���T[� ?�����LP�� P�9��:��;*;�9;<kB;��F;[NH;Z�H;�I;lI;�I; I;�I;"I;D�H;��H;��H;��H;J�H;��H;��H;��H;D�H; I;�I;I;�I;kI;�I;V�H;WNH;��F;>kB;�9;*;��;��:(P�9HP������ ?��T[�;���J����5��{��A��P9ݽXl���,���M�1�l����p��      4m־O�Ѿ�>ľ����җ����{��I�+����V���{�=�/�#���,��<=�>�һd�@�0� ���k:��:�a;��3;j?;T2E;��G;C�H;I;P I;�I;�I;	I;�I;��H;��H;��H;��H;9�H;��H;��H;��H;��H;�I; 	I;�I;�I;Q I;I;B�H;��G;R2E;j?;��3;�a;��:��k:0� �b�@�?�һ<=��,��#��=�/��{��V�����+��I���{�җ�������>ľO�Ѿ      C\����q5��z ��E۾ֳ�^��y�Z�K?#����A����j�$��Dϼ �����Ƶ���lۺ�9�9t4�:H�;H�,;[�;;�C;�G;"�H;�I;�!I;�I;%I;	I;sI;$I;��H;��H;��H;�H;��H;��H;��H;#I;sI;I;$I;�I;�!I;�I;"�H;�G;"�C;\�;;J�,;@�;v4�:x9�9�lۺƵ����� ��Cϼ$����j��A�����K?#�y�Z�^��ֳ��E۾�z �q5����      E�b��>]���M�Î6�����$���>ľ#q��y�Z�+�Q9ݽ W����L����!F�� �G�	�׻;� o칊Ȋ:�i;P$;��7;W�A;�IF;CH;��H;� I;BI;VI;�I;
I;�I;��H;��H;t�H;��H;r�H;��H;��H;I;I;�I;ZI;EI;� I;��H;CH;�IF;V�A;��7;P$;�i;�Ȋ:o��;��׻�G�!F�������L� W��P9ݽ+�y�Z�#q���>ľ�$�����Î6���M��>]�      p��񲗿���7�y�{�R���)�nv��>ľ^���I�Xl����������&�ҮҼ�}�/B�Ȯ�������!:�*�:&z;^3;Lj?;t\E;��G;��H;II;I;mI;�I;WI;�I;��H;��H;C�H;��H;C�H;��H;��H;�I;XI;�I;pI;�I;LI;��H;��G;t\E;Lj?;b3;&z;�*�:��!:���Ȯ��.B��}�ҮҼ��&��������Xl��I�^���>ľnv���)�{�R�7�y����񲗿      �˿�<ƿqL��@1����>]���)��$��ֳ���{���,�q��&��P`I��J���,���3/��+��� �`-69�4�:ք;�o.;.=;@aD;��G;Q�H;�I;!I;BI;,I;�	I;�I;� I;��H;��H;E�H;��H;��H;� I;�I;�	I;*I;BI;!I;�I;T�H;��G;@aD;.=;�o.;ք;�4�:p-69� ��+���3/��,���J��P`I�&��q�齤�,���{�ֳ��$����)��>]��@1��qL���<ƿ      ����<���T[忶˿�T���{�R�����E۾җ����M���	������j��3�d����O�8�׻��/���K��:� 
;�*;P;;�jC;�'G;ԛH;�I;�!I;�I;wI;�
I;�I;�I;�H;��H;��H;��H;"�H;�I;�I;�
I;vI;�I;�!I;�I;ۛH;�'G;�jC;R;;�*;� 
;C��:����/�6�׻��O�d���3���j������	���M�җ���E۾���{�R���T���˿T[�<���      O�6��t����˿@1��7�y�Î6��z �����2�l�+��ͽ"�����&���˼<�k������X�ؙ ����:<�;�&;�9;o�B;��F;�}H;�	I;1"I;I;�I;yI;TI;%I;��H;�H;c�H;�H;��H;"I;TI;|I;�I;I;3"I;�	I;�}H;��F;m�B;�9;�&;<�;|��:̙ ���X����<�k���˼��&�"����ͽ+�2�l������z �Î6�7�y�@1���˿���t�6��      ��*��g&��#�t�T[�qL�������M�r5��>ľ����,��D�蒐��5�0�ݼ���q
��x�uk���b:1l�:�#;ɗ7;Z�A;��F;�dH;�I;#"I;�I;HI;I;�I;�I;��H;Y�H;��H;T�H;��H;�I;�I;I;BI;�I;("I;�I;�dH;��F;T�A;ė7;�#;1l�:��b:�tk��x��q
���0�ݼ�5�蒐��DὪ�,����>ľr5���M����qL��T[�t��#��g&�      ��8��4��g&�6��<����<ƿ񲗿�>]����O�Ѿ�p���*7����$W��KR?��|�p8�������ȅ����G: �:�!;�6;�kA;hYF;�TH;F�H;�!I;�I;�I;eI;(I;�I;; I;��H;��H;��H;; I;�I;)I;hI;�I;�I;�!I;I�H;�TH;vYF;�kA;�6;�!;{ �:��G:���������p8���|�KR?�$W�����*7��p��O�Ѿ����>]�񲗿�<ƿ<���6���g&��4�      �Aq���i���U�F:�@�����<���u���{A�d5�� ��~^Z�����A���]�����d��I",��5����ѺX��9���:%�;aY4;M�@;RVF;��H;�GI;�bI;OI;:I;�)I;I;{I;�I;�I;�I;zI;�I;{I;I;�)I;:I;OI;�bI;�GI;��H;^VF;H�@;]Y4;�;���:P��9��Ѻ�5��H",��d������]��A�����~^Z�� ��d5�{A�u���<�������@�F:���U���i�      ��i���b�Z�O�.5�1i�������������q<�����e��`
V�GE	�!���IY�i9�B�����(��R����Ⱥt�:\��:�;D�4;C�@;#hF;��H;II;ybI;�NI;�9I;�)I;�I;[I;�I;]I;ZI;WI;�I;WI;�I;�)I;�9I;�NI;|bI;II;��H;.hF;B�@;A�4;�;V��:h�:��Ⱥ�R����(�B���i9��IY�!��GE	�`
V��e������q<������������1i�.5�Z�O���b�      ��U�Z�O�H-?�.�'���L�ῴ欿a�{�ea/���뾝���I����c���ZN�Z5������;H�` ��b�����":��:�;��5;�`A;��F;N�H;MI;�aI;�MI;�8I;�(I;BI;�I;:I;I;I;�I;9I;�I;BI;�(I;�8I;�MI;�aI;MI;O�H;��F;�`A;��5;{�;��:��":V���b ��:H�����Z5���ZN�c������I�������ea/�a�{��欿L����.�'�H-?�Z�O�      F:�.5�.�'��������jȿ���l$_���W�Ҿە���6�����*���`=�:�漬)��GG�$6�����<�Q:��:�/";�7;b&B;��F;��H;�RI;�`I;xKI;7I;�'I;>I;I;�I;qI;p
I;kI;�I;I;<I;�'I;7I;zKI;�`I;�RI;��H;��F;a&B;
�7;�/";��:0�Q:���$6��FG��)��:���`=��*������6�ە��W�Ҿ��l$_����jȿ�������.�'�.5�      @�1i�������I�ѿk��� ���q<��:��a����q����Wн潅���'�Sb̼�zl��.��F�X�H����:��;Ԏ&;ʫ9;'C;>MG;��H;:YI;�^I;�HI;�4I;�%I;�I;I;�I;�
I;�	I;�
I;�I;I;�I;�%I;�4I;�HI;�^I;:YI;��H;CMG;'C;ū9;ю&;��;��:4��G�X��.���zl�Sb̼��'�潅��Wн����q��a���:��q<� ��k���I�ѿ������1i�      �������L��jȿk���������O���{]׾z����I�����A��=�d�m�|֮�
RH��jλI�$�p(�z��:JN;��+;�<;�3D;��G;�I;�^I;l[I;�DI;"2I;�#I;CI;�I;]I;�	I;�I;�	I;]I;�I;CI;�#I; 2I;�DI;l[I;�^I;�I;��G;�3D;�<;��+;HN;n��:@(�I�$��jλ
RH�|֮�m�=�d��A������I�z���{]׾����O�����k���jȿL�Ῡ��      <��������欿��� ����O��x����� ���l���"��ܽ���`=����t���k"�*R��2ۺؓ�9�?�:_L;��0;��>;�ME;K#H;�%I;�aI;�VI;�@I;�.I;=!I;>I;I;
I;MI;�I;JI;
I;I;@I;=!I;�.I;�@I; WI;�aI;�%I;P#H;�ME;��>;��0;^L;�?�:���92ۺ*R���k"�t������`=����ܽ��"��l�� ����뾁x���O� ������欿����      u�������a�{�k$_��q<�������}��w��	�6�����!���h����᷾�� d�{.���^e��H[���Z:h��:�, ;��5;�A;�VF;��H;�@I;obI;�QI;�;I;=+I;mI;I;7I;}	I;�I;,I;�I;	I;7I;I;kI;;+I;�;I;�QI;ubI;�@I;��H;�VF;�A;��5;�, ;`��:��Z:�H[��^e�z.�� d�෾�����h�!������	�6�w���}��������q<�k$_�a�{�����      {A��q<�ea/����:�{]׾� ��w��>�CE	�����ٽ����3�\�꼘���",��W��Y�� 
Q����:�M
;�f);��:;'@C;�?G;R�H;HTI;�_I;$KI;�6I;N'I;eI;�I;;I;�I;oI;�I;lI;�I;;I;�I;jI;O'I;�6I;,KI;�_I;GTI;S�H;�?G;'@C;��:;�f);�M
;���: 
Q�Z���W��
",�����\�꼗�3�ٽ������CE	�>�w��� ��{]׾�:���ea/��q<�      d5�������W�Ҿ�a��z����l�	�6�CE	���Ƚk���aG����c֮��W����g�k�"���c,:���:��;��1;B�>;@E;"�G;I;&_I;AZI;3DI;�1I;0#I;EI; I;
I;I;�I;I;�I;I;
I;�I;CI;3#I;�1I;:DI;GZI;&_I;I;'�G;>E;D�>;��1;��;���:�c,: ��c�k�����W�b֮�����aG�k����ȽCE	��6��l�z����a��W�Ҿ������      � ���e�����ە����q��I���"���������k���ZN�Z� ¼M�y��$��Q���� � PX���:0;*�&;�w8;o B;��F;ԐH;W@I;�aI;jRI;=I;,I;�I;�I;\I;�I;4I;I;eI;I;8I;�I;^I;�I;�I;,I;=I;pRI;�aI;T@I;ڐH;��F;r B;�w8;(�&;(0;��: DX��� ��Q���$�K�y�¼Z��ZN�k������������"��I���q�ە������e��      }^Z�`
V��I��6�������ܽ!��ٽ���aG�Z�	�ȼ�)��{�(�c��DG5������Z:!�:S;'1;��=;��D;/�G;��H;�XI;^I;~II;�5I;�&I;�I;�I;�
I;�I;MI;a I;��H;a I;MI;�I;�
I;�I;�I;�&I;�5I;�II;^I;�XI;��H;1�G;��D;��=;'1;S;-�:��Z:���AG5�b��z�(��)��	�ȼY��aG�ٽ��!���ܽ������6��I�_
V�      ���FE	��������Wн�A�����h���3����¼�)��/x/��һl�X�f#����9Z��:�>;2f);i`9;_&B;��F;g}H;�6I;PaI;�UI;`@I;�.I;� I;GI;(I;�I;NI;Q I;��H;��H;��H;P I;NI;�I;(I;KI;!I;�.I;d@I;�UI;NaI;�6I;g}H;��F;d&B;g`9;=f);�>;Z��:��9`#��i�X�
�һ.x/�)��¼�����3��h��󑽠A���Wн��콹��FE	�      �A��!��b���*��潅�>�d��`=����\��b֮�K�y�z�(��һ�]e�܄���f9���:<�;G1";�4;�m?;�E;��G;h�H;�WI;�^I;KI;q7I;�'I;�I;$I;�
I;$I;I;m�H;��H;;�H;��H;k�H;I;!I;�
I;(I;�I;�'I;v7I;	KI;|^I;�WI;g�H;��G;�E;�m?;#�4;M1";:�;���:�f9ڄ���]e��һz�(�J�y�b֮�[�꼗���`=�=�d�潅��*��c��!��      �]��IY��ZN��`=���'�l����߷�������W��$�c��l�X������9���:e��:t�;��0;��<;T�C;"G;��H;�?I;&aI;�TI;>@I;/I;U!I;�I;I;yI;�I;��H;}�H;�H;��H;�H;|�H;��H;�I;vI;I;�I;Z!I;/I;>@I;�TI;)aI;�?I;��H;%G;U�C;��<;��0;r�;q��:���:�9ڄ��i�X�b���$��W�����෾����l���'��`=��ZN��IY�      ���h9�X5��8��Sb̼|֮�s��} d�
",�����Q��CG5�j#���f9���:��:�;��-;��:;�KB;>VF;KH;�I;�\I;\I;�HI;6I;'I;I;�I;
I;BI;��H;��H;��H;Z�H;��H;X�H;��H;��H;��H;AI;
I;�I;I;"'I;6I;�HI; \I;�\I;�I;KH;@VF;�KB;��:;��-;�;��:���:�f9l#��@G5��Q�����	",�~ d�s��z֮�Tb̼9��Y5��h9�      �d��@��������)���zl�	RH��k"�v.���W��\�k�~� ������9���:q��:�;�-;ѫ9;HaA;��E;*�G;x�H;SI;`I;�OI;�<I;�,I;�I;.I;I;zI;TI;��H;��H;��H;��H;a�H;��H;��H;��H;��H;TI;~I;I;1I;�I;�,I;�<I;�OI;`I;�RI;y�H;*�G;��E;IaA;̫9;�-;�;s��:���:��9���z� �\�k��W��u.���k"�RH��zl��)������@���      A",���(�9H�BG��.���jλ$R���^e�V���� 8X���Z:P��:8�;s�;��-;ʫ9;|A;�cE;!�G;��H;RGI;�`I;�UI;;BI;�1I;�#I;�I;�I;�I;�I;��H;H�H;��H;�H;�H;��H;�H;	�H;��H;E�H;��H;�I;�I;�I;�I;�#I;�1I;ABI;�UI;�`I;SGI;��H;%�G;�cE;zA;ͫ9;��-;s�;8�;N��:��Z:  X���Q���^e�&R���jλ�.��CG�7H���(�      �5���R��` ��6��J�X�:�$�ۺ�H[��Q��c,:��:)�:�>;M1";��0;��:;HaA;�cE;��G;w�H;�=I;.`I;tYI;�FI;�5I;�'I;�I;�I;�
I;�I;��H;�H;�H;��H;�H;��H;<�H;��H;}�H;��H;�H;�H;��H;�I;�
I;�I;�I;�'I;�5I;�FI;mYI;1`I;�=I;z�H;��G;�cE;LaA;��:;��0;K1";�>;)�:��:�c,:�Q��H[�$ۺ?�$�G�X�$6��_ ���R��      ��Ѻ��ȺH���|��D�� (�H��9��Z:���:���:*0;S;9f);!�4;��<;�KB;��E;+�G;|�H;`:I;R_I;�[I;%JI;9I;�*I;�I;�I; I;]I;I;��H;��H;�H;/�H;��H;7�H;��H;2�H;��H;.�H;�H;��H;��H;I;\I;I;�I;�I;�*I;9I;!JI;�[I;V_I;b:I;|�H;$�G;��E;�KB;��<;�4;7f);S;*0;���:���:��Z:0��9�'�(�����`����Ⱥ      ���90�:0�":,�Q:��:|��:�?�:f��:�M
;�;(�&;'1;g`9;�m?;U�C;BVF;,�G;��H;�=I;Q_I;\I;�KI;;I;�,I;� I;�I;�I;�I;HI;��H;5�H;x�H;5�H;��H;��H;��H;��H;��H;��H;��H;2�H;r�H;7�H;��H;GI;�I;�I;�I;� I;�,I;;I;�KI;\I;R_I;�=I;��H;,�G;BVF;U�C;�m?;i`9;'1;.�&;�;�M
;b��:�?�:r��:��:�Q:\�":0�:      ���:v��:��:��:��;LN;_L;�, ;�f);��1;�w8;��=;e&B;�E;)G;KH;}�H;YGI;6`I;�[I;�KI;�;I;�-I;3"I;0I;I;	I;dI;��H;��H;��H;j�H;y�H;�H;F�H;��H;e�H;��H;C�H;�H;x�H;f�H;��H;��H;��H;eI;	I;I;3I;2"I;�-I;�;I;�KI;�[I;3`I;UGI;}�H;KH;)G;�E;d&B;��=;�w8;��1;�f);�, ;eL;HN;��;��:��:^��:      :�;�;w�;�/";Ǝ&;��+;��0;��5;��:;I�>;| B;��D;��F;��G; �H;�I;SI; aI;tYI;$JI;;I;�-I;�"I;I;�I;�	I;.I;I�H;r�H;Z�H;��H;��H;��H;��H;��H;��H;a�H;��H;��H;��H;��H;��H;��H;X�H;m�H;N�H;'I;�	I;�I; I;�"I;�-I;;I;$JI;tYI;�`I;SI;�I; �H;��G;��F;��D; B;E�>;��:;��5;��0;��+;ێ&;�/";t�;̔;      [Y4;K�4;��5;
�7;��9;�<;��>;�A; @C;CE;��F;3�G;g}H;k�H;�?I;�\I;`I;�UI;�FI;9I;�,I;."I;I;&I;]
I;�I;��H;��H;��H;��H;��H;��H;��H;��H;��H;��H;i�H;��H;��H;��H;��H;��H;��H;��H;��H;��H;��H;�I;_
I;#I;�I;."I;�,I; 9I;�FI;�UI;`I;�\I;�?I;g�H;g}H;2�G;��F;AE;%@C;�A;��>;�<;ȫ9;�7;��5;A�4;      h�@;>�@;�`A;]&B;C;4D;�ME;�VF;�?G;*�G;ސH;��H;�6I;�WI;0aI;+\I;�OI;FBI;�5I;�*I;� I;5I;�I;d
I;�I; I;3�H;��H;'�H;��H;��H;��H;N�H;|�H;��H;��H;h�H;��H;��H;|�H;I�H;��H;�H;��H;�H;��H;-�H; I;�I;c
I;�I;7I;� I;�*I;�5I;BBI;�OI;-\I;-aI;�WI;�6I;��H;��H;*�G;�?G;�VF;�ME;�3D;*C;^&B;�`A;?�@;      NVF;.hF;��F;��F;1MG;��G;Q#H;��H;T�H;#I;]@I;�XI;VaI;�^I;�TI;�HI;�<I;�1I;�'I;�I;�I;I;�	I;�I; I;?�H;�H;[�H;��H;��H;z�H;K�H;@�H;{�H;	�H;��H;~�H;��H;�H;{�H;?�H;G�H;z�H;��H;��H;Y�H;�H;C�H; I;�I;�	I;I;�I;�I;�'I;�1I;�<I;�HI;�TI;�^I;VaI;�XI;b@I;!I;T�H;��H;R#H;��G;JMG;��F;��F;(hF;      ��H;��H;E�H;��H;��H;�I;�%I;�@I;KTI;*_I;�aI;^I;�UI;KI;A@I;	6I;�,I;�#I;�I;�I;�I;	I;-I;��H;-�H;�H;J�H;�H;0�H;p�H;)�H;�H;;�H;��H;:�H;��H;��H;��H;7�H;��H;9�H;�H;)�H;o�H;)�H;�H;C�H;�H;1�H;��H;,I;	I;�I;�I;�I;�#I;�,I;6I;<@I;KI;�UI;^I;�aI;)_I;JTI;�@I;�%I;�I;��H;��H;E�H;��H;      �GI;II;MI;�RI;.YI;�^I;�aI;sbI;�_I;JZI;qRI;�II;b@I;y7I;/I;"'I;�I;�I;�I;�I;�I;aI;G�H;��H;��H;T�H;�H;�H;~�H;)�H;�H;�H;h�H;��H;v�H;A�H;6�H;@�H;u�H;��H;g�H;	�H;�H;&�H;z�H;�H;
�H;Y�H;��H;��H;E�H;aI;�I;�I;�I;�I;�I;#'I;/I;u7I;a@I;�II;tRI;JZI;�_I;pbI;�aI;z^I;:YI;�RI;MI;II;      �bI;ubI;�aI;�`I;�^I;k[I;WI;�QI; KI;9DI;=I;�5I;�.I;�'I;\!I;I;6I;�I;�
I;`I;NI;��H;n�H;��H;�H;��H;%�H;}�H;#�H;��H;��H;;�H;��H;,�H;��H;��H;��H;��H;��H;-�H;��H;8�H;��H;��H;�H;|�H;"�H;��H;�H;��H;n�H;��H;JI;\I;�
I;�I;5I;I;Z!I;�'I;�.I;�5I;=I;<DI;)KI;�QI;WI;g[I;�^I;�`I;�aI;sbI;      OI;�NI;�MI;sKI;�HI;�DI;�@I;�;I;�6I;�1I;,I;�&I;!I;�I;�I;�I;I;�I;�I;I;��H;��H;V�H;��H;��H;��H;n�H;*�H;�H; �H;&�H;�H;��H;��H;G�H;!�H;�H;!�H;C�H;��H;��H;}�H;&�H;��H;��H;(�H;g�H;��H;��H;��H;X�H;��H;��H;I;�I;�I;I;�I;�I;�I;!I;�&I;,I;�1I;�6I;�;I;�@I;�DI;�HI;yKI;�MI;�NI;       :I;�9I;�8I;&7I;�4I;!2I;�.I;K+I;S'I;9#I;�I;�I;QI;/I;I;"
I;�I;�I;��H;��H;=�H;��H;��H;��H;��H;v�H;)�H;�H;��H;-�H;��H;��H;_�H;�H;��H;��H;��H;��H;��H;�H;_�H;��H;��H;)�H;��H;�H;#�H;w�H;��H;��H;��H;��H;9�H;��H;��H;�I;�I;$
I;I;.I;RI;�I;�I;:#I;V'I;I+I; /I;2I;�4I;(7I;�8I;�9I;      �)I;�)I;�(I;�'I;�%I;�#I;@!I;pI;mI;HI;�I;�I;.I;�
I;}I;HI;\I;��H;�H;��H;}�H;i�H;��H;��H;��H;B�H;�H;�H;>�H;��H;��H;w�H;��H;��H;w�H;N�H;9�H;Q�H;s�H;��H;��H;w�H;��H;�H;8�H;�H;	�H;B�H;��H;��H;��H;l�H;x�H;��H;�H;��H;^I;JI;}I;�
I;+I;�I;�I;HI;kI;mI;I!I;�#I;�%I;�'I;�(I;�)I;      %I;�I;MI;AI;�I;<I;>I;I;�I;�I;_I;�
I;�I;(I;�I;  I;��H;K�H;#�H;�H;?�H;{�H;��H;��H;K�H;<�H;9�H;l�H;��H;��H;Y�H;��H;��H;U�H;�H;�H;�H;�H;�H;X�H;��H;��H;[�H;��H;��H;i�H;5�H;9�H;N�H;��H;��H;{�H;9�H;�H;#�H;N�H;��H; I;�I;(I;�I;�
I;bI;�I;�I;I;@I;6I;�I;;I;WI;�I;      vI;\I;�I;I;I;�I;I;=I;>I;
I;�I;�I;VI;$I;��H;��H;��H;��H;��H;5�H;��H;�H;��H;��H;r�H;t�H;��H;��H;0�H;��H;	�H;��H;X�H;�H;��H;��H;��H;��H;��H;�H;Z�H;��H;�H;��H;*�H;��H;��H;t�H;x�H;��H;��H;�H;��H;.�H;��H;��H;��H;��H;��H;$I;UI;�I;�I;
I;AI;:I;I;�I;	I;I;�I;eI;      �I;�I;@I;�I;�I;WI;I;�	I;�I;I;AI;[I;] I;x�H;��H;��H;��H;�H;��H;��H;��H;B�H;��H;��H;��H;��H;1�H;u�H;��H;H�H;��H;v�H;�H;��H;��H;��H;��H;��H;��H;��H;�H;z�H;��H;C�H;��H;t�H;1�H;��H;��H;��H;��H;B�H;��H;��H;��H;�H;��H;��H;��H;x�H;^ I;YI;BI;I;�I;�	I;I;ZI;�I;�I;@I;�I;      ~I;dI;I;nI;�
I;�	I;VI;�I;oI;�I;%I;h I;��H;��H;�H;Z�H;��H;�H;��H;6�H;��H;��H;��H;u�H;��H;��H;��H;A�H;��H;'�H;��H;P�H;�H;��H;��H;}�H;|�H;��H;��H;��H;	�H;S�H;��H;!�H;��H;@�H;��H;��H;��H;z�H;��H;��H;��H;3�H;��H;�H;��H;^�H;�H;��H;��H;g I;(I;�I;qI;�I;]I;�	I;�
I;oI; I;rI;      �I;WI;I;t
I;�	I;�I;�I;5I;�I;"I;pI;��H;�H;E�H;��H;��H;m�H;��H;A�H;��H;��H;h�H;]�H;[�H;b�H;u�H;��H;:�H;��H;$�H;��H;;�H;�H;��H;��H;w�H;��H;z�H;��H;��H;�H;=�H;��H;�H;��H;6�H;��H;w�H;f�H;]�H;d�H;h�H;��H;��H;A�H;��H;m�H;��H;��H;H�H;�H;��H;sI;%I;�I;5I;�I;�I;�	I;x
I;I;dI;      ~I;eI; I;nI;�
I;�	I;TI;�I;oI;�I;$I;i I;��H;��H;�H;Z�H;��H;�H;��H;6�H;��H;��H;��H;w�H;��H;��H;��H;A�H;��H;$�H;��H;P�H;	�H;��H;��H;}�H;|�H;��H;��H;��H;	�H;S�H;��H;�H;��H;=�H;��H;��H;��H;x�H;��H;��H;��H;3�H;��H;�H;��H;_�H;�H;��H;��H;h I;(I;�I;sI;�I;[I;�	I;�
I;uI;I;lI;      �I;�I;;I;�I;�I;VI;I;�	I;�I;I;BI;[I;] I;x�H;��H;��H;��H;�H;��H;��H;��H;D�H;��H;��H;��H;��H;0�H;t�H;��H;G�H;��H;v�H;�H;��H;��H;��H;��H;��H;��H;��H;�H;x�H;��H;@�H;��H;q�H;1�H;�H;��H;��H;��H;C�H;��H;��H;��H;�H;��H;��H;��H;z�H;` I;\I;CI;I;�I;�	I;I;VI;�I;�I;AI;�I;      vI;[I;�I;I;I;�I;I;@I;AI;
I;�I;�I;UI;$I;��H;��H;��H;��H;��H;4�H;��H;�H;��H;��H;w�H;t�H;��H;��H;0�H;��H;�H;��H;X�H;�H;��H;��H;��H;��H;��H;�H;Z�H;��H;�H;��H;)�H;��H;��H;w�H;w�H;��H;��H;�H;��H;/�H;��H;��H;��H;��H;��H;&I;VI;�I;�I;
I;BI;?I;I;�I;I;I;�I;\I;      "I;�I;PI;:I;�I;?I;=I;I;�I;�I;aI;�
I;�I;(I;�I; I;��H;L�H;!�H;�H;?�H;|�H;��H;��H;N�H;6�H;5�H;k�H;��H;��H;X�H;��H;��H;U�H;�H;�H;�H;�H;�H;W�H;��H;��H;Y�H;��H;��H;h�H;6�H;:�H;K�H;��H;��H;|�H;8�H;�H;#�H;N�H;��H; I;�I;*I;�I;�
I;bI;�I;�I;I;DI;;I;�I;EI;XI;�I;      �)I;�)I;�(I;�'I;�%I;�#I;D!I;nI;jI;HI;�I;�I;+I;�
I;�I;HI;\I;��H;
�H;��H;�H;l�H;��H;��H;��H;A�H;	�H;�H;?�H;�H;��H;t�H;��H;��H;w�H;J�H;9�H;N�H;s�H;��H;��H;w�H;��H;}�H;8�H;�H;�H;D�H;��H;��H;��H;l�H;y�H;��H;
�H;��H;^I;JI;I;�
I;/I;�I;�I;JI;mI;nI;F!I;�#I;�%I;�'I;�(I;�)I;      :I;�9I;�8I;7I;�4I;$2I;�.I;I+I;U'I;7#I;�I;�I;QI;0I;I;"
I;�I;�I;��H;��H;@�H;��H;��H;��H;��H;s�H;%�H;�H;��H;*�H;��H;��H;]�H;�H;��H;��H;��H;��H;��H;�H;_�H;��H;��H;'�H;��H;�H;&�H;y�H;��H;��H;��H;��H;9�H;��H;��H;�I;�I;$
I;I;0I;RI;�I;�I;:#I;U'I;I+I;�.I;!2I;�4I;*7I;�8I;�9I;      'OI;�NI;�MI;}KI;|HI;�DI;�@I;�;I;�6I;�1I;,I;�&I;!I;�I;�I;�I;I;�I;�I;I;��H;��H;V�H;��H;��H;��H;k�H;(�H;�H; �H;&�H;}�H;��H;��H;F�H; �H;�H;!�H;C�H;��H;��H;�H;&�H;��H;��H;(�H;k�H;��H;��H;��H;Z�H;��H;��H;I;�I;�I;I;�I;�I;�I;!I;�&I;,I;�1I;�6I;�;I;�@I;�DI;�HI;�KI;�MI;�NI;      �bI;sbI;�aI;�`I;~^I;q[I;WI;�QI;,KI;7DI;=I;�5I;�.I;�'I;_!I;I;5I;�I;�
I;]I;OI;��H;m�H;��H;�H;��H;$�H;}�H;#�H;��H;��H;:�H;��H;,�H;��H;��H;��H;��H;��H;,�H;��H;:�H;��H;��H;�H;z�H;$�H;��H;�H;��H;o�H;��H;KI;\I;�
I;�I;5I;I;^!I;�'I;�.I;�5I;=I;9DI;)KI;�QI;WI;l[I;�^I;�`I;�aI;obI;      �GI;II;MI;�RI;*YI;�^I;�aI;wbI;�_I;KZI;qRI;�II;a@I;{7I;/I;%'I;�I;�I;�I;�I;�I;dI;E�H;��H;��H;O�H;�H;�H;~�H;&�H;�H;�H;e�H;��H;u�H;>�H;7�H;A�H;t�H;��H;h�H;�H;�H;(�H;z�H;�H;�H;X�H;��H;��H;H�H;cI;�I;�I;�I;�I;�I;%'I;/I;x7I;b@I;�II;sRI;JZI;�_I;pbI;�aI;�^I;9YI;�RI;MI;II;      ��H;ȗH;G�H;��H;��H;�I;�%I;�@I;NTI;*_I;�aI;#^I;�UI;KI;C@I;6I;�,I;�#I;�I;�I;�I;	I;)I;��H;0�H;�H;G�H;�H;/�H;l�H;(�H;�H;8�H;��H;8�H;��H;��H;��H;7�H;��H;9�H;�H;*�H;n�H;+�H;�H;G�H;�H;.�H;��H;.I;	I;�I;�I;�I;�#I;�,I;6I;B@I;KI;�UI;^I;�aI;)_I;KTI;�@I;�%I;�I;��H;��H;J�H;��H;      BVF;.hF;��F;��F;7MG;��G;K#H;��H;[�H;!I;^@I;�XI;VaI;�^I;�TI;�HI;�<I;�1I;�'I;�I;�I;I;�	I;�I; I;<�H;�H;]�H;��H;��H;y�H;H�H;=�H;{�H;�H;��H;��H;��H;�H;{�H;@�H;I�H;}�H;��H;��H;[�H;�H;E�H; I;�I;�	I;I;�I;�I;�'I;�1I;�<I;�HI;�TI;�^I;VaI;�XI;`@I;!I;R�H;��H;M#H;��G;FMG;��F;��F;hF;      f�@;?�@;�`A;X&B;C;
4D;�ME;�VF;�?G;*�G;��H;��H;�6I;�WI;3aI;.\I;�OI;HBI;�5I;�*I;� I;7I;�I;d
I;�I; I;.�H;��H;$�H;��H;��H;��H;I�H;{�H;��H;��H;f�H;��H;��H;~�H;L�H;��H;�H;��H;!�H;��H;0�H; I;�I;c
I;�I;8I;� I;�*I;�5I;EBI;�OI;0\I;3aI;�WI;�6I;��H;ܐH;*�G;�?G;�VF;�ME;�3D;&C;^&B;�`A;>�@;      9Y4;5�4;��5;�7;��9;�<;��>;�A;(@C;@E;��F;3�G;g}H;h�H;�?I;�\I;`I;�UI;�FI;9I;�,I;,"I;�I;&I;_
I;�I;��H;��H;��H;��H;��H;��H;��H;��H;��H;��H;g�H;��H;��H;��H;��H;��H;��H;��H;��H;��H;��H;�I;\
I;'I;�I;."I;�,I;9I;�FI;�UI;`I;�\I;�?I;h�H;g}H;3�G;��F;>E;$@C;�A;��>;�<;Ы9;+�7;��5;�4;      '�;�;q�;�/";Ď&;��+;��0;��5;��:;I�>;x B;��D;��F;��G;�H;�I;SI;�`I;tYI;$JI;;I;�-I;�"I;I;�I;�	I;)I;L�H;r�H;V�H;��H;��H;��H;��H;��H;��H;d�H;��H;��H;��H;��H;��H;��H;[�H;n�H;K�H;,I;�	I;�I;I;�"I;�-I;;I;%JI;uYI;�`I;SI;�I;�H;��G;��F;��D;x B;H�>;��:;��5;��0;��+;Ǝ&;�/";o�;ʔ;      ���:x��:��:��:��;TN;fL;�, ;�f);��1;�w8;��=;d&B;�E;,G;KH;|�H;XGI;3`I;�[I;�KI;�;I;�-I;2"I;5I;I;	I;eI;��H;��H;��H;i�H;x�H;�H;B�H;��H;g�H;��H;B�H;�H;{�H;j�H;��H;��H;��H;dI;	I;I;1I;6"I;�-I;�;I;�KI;�[I;5`I;XGI;}�H;KH;*G;�E;d&B;��=;�w8;��1;�f);�, ;_L;;N;��;��:��:d��:      ��9��:��":4�Q:��:���:�?�:f��:�M
;�;,�&;'1;j`9;�m?;Y�C;DVF;*�G;��H;�=I;R_I;\I;�KI;;I;�,I;� I;�I;�I;�I;HI;��H;5�H;v�H;4�H;��H;��H;��H;��H;��H;��H;��H;5�H;u�H;9�H;��H;GI;�I;�I;�I;� I;�,I;;I;�KI;\I;U_I;�=I;��H;,�G;DVF;Y�C;�m?;j`9;'1;.�&;�;�M
;n��:�?�:|��:��:<�Q:��":L�:      r�Ѻ��ȺR���~��@���'�H��9�Z:���:���:,0;S;:f); �4;��<;�KB;��E;(�G;z�H;b:I;X_I;�[I;$JI;9I;�*I;�I;�I; I;_I;I;��H;��H;�H;1�H;��H;3�H;��H;6�H;��H;-�H;�H;��H;��H;I;]I; I;�I;�I;�*I;9I;%JI;�[I;V_I;c:I;|�H;'�G;��E;�KB;��<;!�4;:f);S;-0;���:���:��Z:0��90(�4�����T�����Ⱥ      �5���R��_ �� 6��K�X�:�$�"ۺ�H[� Q��c,:��:-�:�>;M1";��0;��:;IaA;�cE;��G;y�H;�=I;1`I;tYI;�FI;�5I;�'I;�I;�I;�
I;�I;��H;�H;�H;��H;~�H;��H;<�H;��H;{�H;��H;�H;�H;��H;�I;�
I;�I;�I;�'I;�5I;�FI;tYI;1`I;�=I;|�H;��G;�cE;IaA;��:;��0;K1";�>;-�:��:�c,:�Q��H[�"ۺ<�$�K�X�6��b ���R��      D",���(�:H�CG��.���jλ$R��~^e�O���� ,X���Z:T��:<�;w�;��-;ͫ9;{A;�cE;%�G;��H;UGI;�`I;�UI;BBI;�1I;�#I;�I;�I;�I;�I;��H;G�H;��H;
�H;�H;��H;�H;�H;��H;H�H;�H;�I;�I;�I;�I;�#I;�1I;9BI;�UI;�`I;VGI;��H;'�G;�cE;{A;̫9;��-;v�;:�;T��:��Z: (X���Q���^e�$R���jλ�.��CG�<H���(�      �d��@��������)���zl�RH��k"�t.���W��^�k�}� �����9���:y��:�;�-;Ы9;HaA;��E;/�G;{�H;SI;`I;�OI;�<I;�,I;�I;4I;I;|I;TI;��H;��H;��H;��H;c�H;��H;��H;��H;��H;QI;~I;I;/I;�I;�,I;�<I;�OI;`I;SI;{�H;(�G;��E;HaA;Ы9;�-;�;y��:���:�9���{� �^�k��W��u.���k"�RH��zl��)������@���      ���h9�Y5��8��Sb̼z֮�s��} d�	",�����Q��@G5�l#���f9���:��:�;��-;��:;�KB;BVF;KH;�I;�\I;#\I;�HI;6I;'I;I;�I;
I;BI;��H;��H;��H;X�H;��H;X�H;��H;��H;��H;?I;
I;�I;I;'I;6I;�HI;\I;�\I;�I;KH;<VF;�KB;��:;��-;�;��:���:�f9j#��DG5��Q�����
",�~ d�t��{֮�Tb̼8��Z5��h9�      �]��IY��ZN��`=���'�l����෾������W��$�b��k�X�܄���9���:m��:s�;��0;��<;Y�C;&G;�H;�?I;,aI;�TI;<@I;/I;[!I;�I;I;yI;�I;��H;}�H;�H;��H;�H;z�H;��H;�I;uI;I;�I;[!I;/I;<@I;�TI;&aI;�?I;�H;'G;R�C;��<;��0;p�;q��:���:�9܄��l�X�c���$��W�����෾����l���'��`=��ZN��IY�      �A��!��c���*��潅�=�d��`=����\��b֮�J�y�y�(��һ�]e�؄��@�f9���::�;K1";�4;�m?;�E;��G;k�H;�WI;�^I;
KI;t7I;�'I;�I;(I;�
I;!I;I;m�H;��H;;�H;��H;j�H;I;!I;�
I;%I;�I;�'I;r7I;
KI;}^I;�WI;j�H;��G;�E;�m?;!�4;H1";:�;���:�f9ڄ���]e��һz�(�J�y�b֮�\�꼖���`=�=�d�潅��*��b��!��      ���FE	��������Wн�A�����h���3����¼�)��.x/��һh�X�d#����9V��:�>;7f);m`9;b&B;��F;k}H;�6I;PaI;�UI;a@I;�.I;� I;JI;(I;�I;PI;Q I;��H;��H;��H;P I;NI;�I;%I;HI; !I;�.I;`@I;�UI;NaI;�6I;g}H;��F;b&B;f`9;:f);�>;P��:��9f#��h�X��һ/x/��)��¼�����3��h��󑽠A���Wн��콺��FE	�      }^Z�`
V��I��6�������ܽ!��ٽ���aG�Z�	�ȼ�)��z�(�b��CG5������Z:)�:S;'1;��=;��D;3�G;��H;�XI;^I;~II;�5I;�&I;�I;�I;�
I;�I;MI;` I;��H;a I;KI;�I;�
I;�I;�I;�&I;�5I;~II;^I;�XI;��H;1�G;��D;��=;'1;S;%�:��Z:���EG5�b��{�(��)��	�ȼZ��aG�ٽ��!���ܽ������6��I�_
V�      � ���e�����ە����q��I���"���������k���ZN�Z�¼L�y��$��Q���� � PX���:#0;/�&;�w8;u B;��F;ڐH;Z@I;�aI;oRI;=I;,I;�I;�I;\I;�I;4I;I;eI;I;4I;�I;\I;�I;�I;,I;=I;oRI;�aI;V@I;ԐH;��F;v B;�w8;#�&;#0;��: PX��� ��Q���$�L�y� ¼Z��ZN�k������������"��I���q�ە������e��      d5�������W�Ҿ�a��z����l��6�CE	���Ƚk���aG����c֮��W����c�k�$���c,:���:�;��1;D�>;CE;'�G;I;&_I;CZI;9DI;�1I;4#I;EI; I;
I;	I;�I;I;�I;	I;
I;�I;BI;2#I;�1I;:DI;EZI;$_I;I;"�G;@E;I�>;��1;��;���:�c,:"��b�k�����W�c֮�����aG�k����ȽCE	�	�6��l�z����a��W�Ҿ������      {A��q<�ea/����:�{]׾� ��w��>�CE	�����ٽ����3�\�꼘���
",��W��]��@
Q����:�M
;�f);��:;(@C;�?G;P�H;HTI;�_I;*KI;�6I;P'I;hI;�I;>I;�I;oI;�I;mI;�I;<I;�I;gI;O'I;�6I;*KI;�_I;GTI;S�H;�?G;*@C;��:;�f);�M
;���: Q�Z���W��
",�����\�꼗�3�ٽ������CE	�>�w��� ��{]׾�:���ea/��q<�      u�������a�{�k$_��q<�������}��w��	�6�����!���h����᷾� d�z.���^e��H[���Z:l��:�, ;��5;�A;�VF;��H;�@I;pbI;�QI;�;I;>+I;kI;I;9I;~	I;�I;.I;�I;	I;7I;I;kI;>+I;�;I;�QI;rbI;�@I;��H;�VF;�A;��5;�, ;`��:��Z:�H[��^e�y.��� d�᷾�����h�!������	�6�w���}��������q<�k$_�a�{�����      <��������欿��� ����O��x����� ���l���"��ܽ���`=����t���k"�,R��6ۺ���9�?�:_L;��0;��>;�ME;K#H;�%I;�aI; WI;�@I;�.I;<!I;@I;I;
I;MI;�I;LI;I;I;@I;=!I;�.I;�@I; WI;�aI;�%I;Q#H;�ME;��>;��0;_L;�?�:��96ۺ*R���k"�t������`=����ܽ��"��l�� ����뾁x���O� ������欿����      �������L��jȿk���������O���{]׾z����I�����A��=�d�m�|֮�	RH��jλI�$� (�|��:FN;��+;�<;�3D;��G;�I;�^I;l[I;�DI;%2I;�#I;BI;�I;^I;�	I;�I;�	I;^I;�I;CI;�#I;!2I;�DI;l[I;�^I;�I;��G;�3D;�<;��+;IN;t��: (�J�$��jλ
RH�|֮�m�=�d��A������I�z���{]׾����O�����k���jȿL�Ῡ��      @�1i�������I�ѿk��� ���q<��:��a����q����Wн潅���'�Sb̼�zl��.��G�X�8����:��;Ҏ&;ȫ9;'C;8MG;��H;8YI;�^I;�HI;�4I;�%I;�I;
I;�I;�
I;�	I;�
I;�I;I;�I;�%I;�4I;�HI;�^I;:YI;��H;CMG;$C;ɫ9;Ԏ&;��;��:4��G�X��.���zl�Sb̼��'�潅��Wн����q��a���:��q<� ��k���I�ѿ������1i�      F:�.5�.�'��������jȿ���l$_���W�Ҿە���6�����*���`=�;�漬)��GG�$6�����@�Q:��:�/";	�7;b&B;��F;��H;�RI;�`I;vKI;7I;�'I;;I;I;�I;oI;q
I;mI;�I;I;>I;�'I;7I;|KI;�`I;�RI;��H;��F;^&B;�7;�/";��:,�Q:���$6��EG��)��:���`=��*������6�ە��W�Ҿ��l$_����jȿ�������.�'�.5�      ��U�Z�O�H-?�.�'���L�ῴ欿a�{�ea/���뾝���I����c���ZN�Z5������:H�a ��`�����":��:~�;��5;�`A;��F;K�H;MI;�aI;�MI;�8I;�(I;@I;�I;7I;I;	I;I;9I;�I;BI;�(I;�8I;�MI;�aI;MI;Q�H;��F;�`A;��5;{�;��:��":T���b ��:H�����Z5���ZN�c������I�������ea/�a�{��欿L����.�'�H-?�Z�O�      ��i���b�Z�O�.5�1i�������������q<�����e��`
V�GE	�!���IY�i9�B�����(��R����Ⱥt�:\��:�;D�4;C�@;!hF;��H;II;xbI;�NI;�9I;�)I;�I;[I;�I;[I;\I;ZI;�I;[I;�I;�)I;�9I;�NI;|bI;II;��H;-hF;>�@;A�4;�;V��:h�:��Ⱥ�R����(�B���i9��IY�!��GE	�`
V��e������q<������������1i�.5�Z�O���b�      ඕ�S���Ѭ��.�_���7�{�}߿����,b��V�,l¾Hx�c.���Ž��t�)��d����?�N������x9���:T�;��2;9@@;bfF;9�H;��I;R�I;|I;�[I;�CI;2I;�%I;[I;�I;2I;�I;ZI;�%I;2I;�CI;�[I;"|I;R�I;��I;?�H;pfF;5@@;��2;P�;���:��x9��N����?�d��)����t���Žc.�Hx�,l¾�V��,b����}߿{���7�.�_�Ѭ��S���      S���D���#}��+Y��3�����$ڿ$��ý\����(���s��3�5����p�b�R���<<�7���������9U��:ջ;S%3;Kp@;�yF;��H;��I;�I;�{I;K[I;LCI;�1I;P%I;I;WI;I;QI;I;N%I;�1I;NCI;H[I;�{I;�I;��I;��H;�yF;Jp@;R%3;л;K��:���9����7���<<�R��b��p�5����3��s�(�����ý\�$���$ڿ����3��+Y�#}�D���      Ѭ��#}�>tf��lG�ע%��p�.�ʿZ����>M����T�����d�Ȥ�̷�-�d��
��I���1�b���R��Ь�9���: ;�U4;��@;ձF;4�H;܎I;��I;�yI;�YI;6BI;�0I;�$I;�I;�I;I;�I;�I;�$I;�0I;7BI;�YI;�yI;��I;ގI;6�H;�F;��@;�U4;;���:Ь�9J��d����1��I���
�-�d�̷�Ȥ���d�T�������>M�Z���.�ʿ�p�ע%��lG�>tf�#}�      .�_��+Y��lG�f.�{���꿲���M䂿��5���󾍰��N�N�V��Q�� �Q����{����h!��g��`񳺀	:c
�:��;_16;��A;<G;I;8�I;x�I;lvI;KWI;h@I;k/I;�#I;�I;
I;�I;I;�I;�#I;k/I;k@I;HWI;ovI;z�I;8�I;I;DG;��A;]16;��;[
�:t	:V񳺆g���h!�{������ �Q�Q��V��N�N���������5�M䂿�������{�f.��lG��+Y�      ��7��3�֢%�{��<����ſ	���½\�<����Ͼ����`�3��轻z��|�9�\�Ἑ���z��7}�|dt�(�^:g+�:��#;��8;��B;sG;q%I;��I;�I;	rI;TI;�=I;p-I;"I;HI;�I;zI;�I;JI;"I;p-I;�=I;TI;rI;�I;��I;t%I;sG;��B;��8;��#;e+�:�^:ldt��7}��z����\��|�9��z����`�3�������Ͼ<��½\�	�����ſ�<��{�֢%��3�      {�����p������ſ$���Ps���1�1r���d���d�|I�ΈŽ��}�^*�IC���^��B�v�D��F๘ �:��;r); 7;;*D;4�G;UHI;��I;��I;�lI;�OI;�:I;+I; I;�I;yI;,I;uI;�I; I;+I;�:I;�OI;�lI;��I;��I;UHI;=�G;,D;7;;p);��;� �:�F�v�D��B��^�IC��^*���}�ΈŽ|I��d��d��1r����1��Ps�$����ſ��꿃p����      }߿�$ڿ.�ʿ����	����Ps�QX:����%l¾�ǆ���7����75���Q�����t���75�i����� �8�ɼ:��;��.;��=;�EE;�YH;�hI;$�I;��I;%fI;KI;#7I;E(I;�I;�I;�I;wI;�I;�I;�I;E(I;#7I;KI;+fI;��I;&�I;�hI;�YH;�EE;��=;��.;��;�ɼ:��8���j���75��t������Q�75�������7��ǆ�%l¾���QX:��Ps�	�������.�ʿ�$ڿ      ���$��Z���M䂿½\���1�����J˾蝒�C�N�x��H������U�'�c�Ҽ��|��z��n��Bx����&:�P�:��;�W4;Ҡ@;#gF;a�H;�I; �I;0�I;_I;�EI;3I; %I;BI;�I;�I;�I;�I;�I;BI;!%I;3I;�EI;!_I;2�I;"�I;�I;e�H;)gF;͠@;�W4;��;�P�:��&:>x���n���z���|�b�ҼU�'����H���x��C�N�蝒��J˾�����1�½\�M䂿Z���$��      �,b�ý\��>M���5�<��0r��%l¾蝒�"&W��3�7Sؽ�z��YG����{I����?���̻��-��
����:��;��&;|9;�C;�dG;KI;@�I;P�I;MvI;{WI;)@I;�.I;�!I;�I;UI;�I;�I;�I;VI;�I;�!I;�.I;,@I;WI;RvI;T�I;@�I;NI;�dG;�C;|9;��&;��;"��:x
����-���̻��?�{I�����YG��z��7Sؽ�3�"&W�蝒�%l¾0r��<����5��>M�ý\�      �V������������Ͼ�d���ǆ�C�N��3��c�[����\�2��(C���o���	��눻L𳺸��9��:�h;P�/;7�=;HE;�2H;�WI;��I;��I;�kI;�OI;!:I;�)I;"I;�I;�I;�I;xI;�I;�I;�I;$I;�)I;$:I;�OI;�kI;��I;��I;�WI;�2H;HE;:�=;T�/;�h;)��:���9H��눻��	��o�'C��2����\�[���c཰3�C�N��ǆ��d����Ͼ���������      ,l¾(��T������������d���7�x��8Sؽ[���d�C*�bkּ+\����'�)���R�0~��|�:�Z;ӣ#;:=7;*�A;�F;T�H;o�I;�I;��I;�`I;�GI;�3I;'%I;rI;�I;SI;K
I;J	I;M
I;TI;�I;tI;'%I;�3I;�GI;�`I;��I;�I;n�I;[�H;�F;+�A;?=7;ԣ#;�Z;��:~���R�(����'�+\��bkּB*��d�[��7Sؽx����7��d���������T���(��      Gx��s���d�M�N�_�3�|I����H����z����\�B*�	�ݼH���-<<��ڻ�V�4dt�4�&:���:=C;�</;OD=;ԈD;��G;�8I;ǘI;��I;tI;$VI;Z?I;�-I;d I;�I;ZI;�
I;�I;I;�I;�
I;]I;�I;b I;�-I;`?I;.VI;tI;��I;ǘI;�8I;��G;ڈD;TD=;�</;IC;���:8�&:dt��V��ڻ,<<�G���	�ݼB*���\��z��G������|I�`�3�M�N���d��s�      c.��3�Ȥ�V����͈Ž75�����YG�2��bkּG����xC��>�c6}���� �x9p��:
	;.�&;�;8;��A;��F;��H;0yI;��I;��I;0fI;�KI;K7I;|'I;�I;�I;XI;I;�I;�I;�I;I;XI;�I;�I;�'I;R7I;�KI;4fI;��I;��I;7yI;��H;��F;��A;�;8;:�&;	;l��:`�x9 ���_6}��>��xC�G���akּ2��YG����75��͈Ž��V��Ȥ��3�      ��Ž4���̷�Q���z����}��Q�T�'����'C��+\��,<<��>n��8��@�8��:6��:�;�'3;��>;�E;gH;_<I;˗I;��I;�vI;�XI;�AI;u/I;�!I;�I;�I;S	I;cI;%I;tI;#I;bI;T	I;�I;�I;�!I;}/I;�AI;�XI;�vI;��I;җI;a<I;jH;�E;��>;�'3;�;8��:F��:@�2�ກn���>�,<<�*\��'C�����T�'��Q���}��z��Q��̷�4���      ��t��p�-�d��Q�|�9�^*����a�ҼzI���o���'��ڻc6}�8�� 9���:Zm�:��;��.;<;�oC;=7G;��H;ӁI;ӜI;ԅI; fI;<LI;�7I;�'I;�I;uI;LI;HI;�I;� I;Q I;� I;�I;JI;OI;rI;�I;�'I;�7I;ELI;fI;ЅI;ٜI;ՁI;��H;A7G;�oC;<;��.;��;lm�:��:09�6��a6}��ڻ��'��o�zI��a�Ҽ���^*�|�9� �Q�-�d��p�      '��a��
����\��IC���t����|���?���	�(���V����@���:��:�h;#�+;��9;��A;|fF;X�H;u_I;��I;��I;sI;�VI;s@I;�.I;� I;TI;I;�I;jI;O I;�H;�H;~�H;L I;jI;�I;I;YI;� I;�.I;y@I;�VI;�rI;��I;��I;u_I;[�H;~fF;��A;��9;!�+;�h;��:��:������V�$����	���?���|��t��HC��]������
�a�      a��Q���I��{�������^��75��z���̻�눻�R�dt�`�x9F��:hm�:�h;_�*;��8;��@;�E;:(H;h8I;��I;�I;J~I;�`I;�HI;�5I;[&I;tI;2I;�	I;�I;� I;��H;W�H;��H;S�H;��H;� I;�I;�	I;6I;uI;_&I;�5I;�HI;�`I;Q~I;�I;��I;i8I;<(H;�E;��@;ٍ8;c�*;�h;lm�:D��:P�x9dt��R��눻��̻�z��75��^����|����I��O��      ��?��<<��1��h!��z��B�b���n����-�>��}��8�&:f��:6��:��; �+;؍8;B�@;�]E;h�G;GI;�I;R�I;8�I;liI;;PI;<I;�+I;�I;nI;PI;+I;sI;��H;��H;R�H;��H;O�H;��H;��H;pI;)I;TI;rI;�I;�+I;<I;4PI;riI;6�I;L�I;�I;II;m�G;�]E;>�@;ۍ8;�+;��;4��:d��:8�&:�}��>𳺀�-��n��d���B黳z��h!� �1��<<�      N��<��a����g���7}�e�D����*x��0
�����9��:���:	;�;��.;��9;��@;�]E;n�G;?I;�I;�I;N�I;�pI;�VI;�AI;~0I;�"I;�I;�I;�I;�I;��H;^�H;w�H;a�H;��H;^�H;t�H;\�H;��H;�I;�I;�I;�I;�"I;z0I;�AI;�VI;�pI;H�I;�I;�I;AI;m�G;�]E;��@;��9;��.;�;	;���:��:���98
��.x�����l�D��7}��g��a���<��      ������>��>񳺈dt��Fเ�8��&:"��:+��:�Z;EC;5�&;�'3;<;��A;�E;q�G;AI;[|I;ĜI;��I;�uI;r[I;FI;�4I;,&I;�I;II;�	I;�I;9�H;��H;6�H;u�H;�H;�H;z�H;q�H;5�H;��H;7�H;�I;�	I;II;�I;(&I;�4I;FI;r[I;{uI;��I;ȜI;[|I;AI;k�G;�E;��A;<;�'3;3�&;HC;�Z;%��:(��:��&: �8�F�pdt�V�X�຺���       �x9��9��9p	:��^:� �:�ɼ:�P�:��;�h;ԣ#;�</;�;8;��>;�oC;�fF;=(H;PI;�I;ĜI;��I;�wI;q^I;;II;�7I;	)I;I;�I;�I;GI;L I;I�H;S�H;:�H;��H;��H;��H;��H;��H;9�H;Q�H;C�H;O I;II;�I;�I;I;)I;�7I;8II;k^I;�wI;��I;ÜI;�I;II;<(H;fF;�oC;��>;�;8;�</;أ#;�h;��;�P�:�ɼ:� �:(�^:d	:h��9��9      ���:m��:���:�
�:Y+�:��;��;��;��&;W�/;C=7;TD=;��A;�E;D7G;_�H;n8I;�I;�I;��I;�wI;�_I;�JI;�9I;�*I;�I;6I;<I;I;9I;��H;��H;�H;=�H;��H;�H;��H;�H;��H;<�H;�H;��H;�H;;I;I;=I;1I;�I;�*I;�9I;�JI;�_I;�wI;��I;	�I;�I;l8I;[�H;C7G;�E;��A;VD=;D=7;S�/;��&;��;��;��;�+�:k
�:���:Q��:      h�;һ;;��;��#;z);��.;�W4;(|9;@�=;4�A;�D;��F;tH;��H;|_I;ƓI;X�I;P�I;�uI;p^I;�JI;):I;#,I;8 I;�I;QI;�I;$I;��H;��H;4�H;�H;k�H;d�H;��H;T�H;��H;`�H;m�H;�H;3�H;�H;��H;I;�I;MI;�I;< I;,I;":I;�JI;r^I;�uI;P�I;Q�I;ÓI;y_I;��H;nH;��F;��D;8�A;<�=;(|9;�W4;��.;t);��#; �;;��;      ��2;\%3;�U4;Y16;��8;$7;;��=;Ϡ@;�C;JE;�F;��G;��H;d<I;ՁI;��I;�I;<�I;�pI;n[I;9II;�9I;",I;� I;I;I;VI;�I;K�H;f�H;]�H;+�H;=�H;��H;��H;a�H;�H;]�H;��H;��H;:�H;*�H;`�H;c�H;G�H;�I;OI;I;I;� I;,I;�9I;8II;m[I;�pI;5�I;�I;��I;ӁI;^<I;��H;��G;�F;IE;�C;Ԡ@;��=;7;;��8;V16;�U4;S%3;      U@@;Gp@;��@;��A;��B;7D;�EE;&gF;�dG;�2H;_�H;�8I;6yI;ٗI;ߜI;��I;V~I;viI;�VI;FI;�7I;�*I;A I;%I;`I;�I;@I;��H;��H;��H;�H;#�H;��H;p�H;��H;&�H;��H;!�H;��H;r�H;��H;�H; �H;��H;��H;��H;9I;�I;aI;!I;; I;�*I;�7I;FI;�VI;siI;V~I;��I;ܜI;՗I;6yI;�8I;a�H;�2H;�dG;&gF;�EE;,D;��B;��A;��@;Hp@;      bfF;�yF;ӱF;=G;sG;A�G;�YH;q�H;QI;�WI;v�I;јI;��I;��I;ׅI;
sI;�`I;:PI;�AI;�4I;	)I;�I;�I;I;�I;UI;��H;�H;��H;W�H;0�H;f�H;�H;-�H;u�H;�H;�H;�H;q�H;-�H;�H;c�H;0�H;T�H;��H;�H;��H;WI;�I;I;~I;�I;	)I;�4I;�AI;5PI;�`I;sI;ԅI;��I;��I;ϘI;{�I;�WI;RI;o�H;�YH;4�G;sG;GG;ӱF;�yF;      M�H;��H;,�H;I;h%I;UHI;�hI;�I;D�I;��I;�I;��I;�I;�vI;"fI;�VI;�HI;<I;�0I;.&I;I;2I;QI;VI;;I;��H;�H;��H;l�H;4�H;o�H;��H;��H;	�H;l�H;�H;�H;�H;i�H;�H;��H;��H;o�H;2�H;f�H;��H;��H;��H;@I;TI;QI;6I;I;)&I;~0I;<I;�HI;�VI;fI;�vI;�I;��I;�I;��I;A�I;�I;�hI;SHI;%I;�I;+�H;��H;      ��I;�I;َI;?�I;��I;��I;/�I;"�I;S�I;��I;��I;tI;2fI;�XI;>LI;w@I;�5I;�+I;�"I;�I;�I;8I;�I;�I;��H;��H;��H;a�H;I�H;_�H;��H;��H;��H;��H;��H;B�H;'�H;?�H;��H; �H;��H;��H;��H;^�H;E�H;_�H;��H;��H;��H;�I;�I;;I;�I;�I;�"I;�+I;�5I;y@I;<LI;�XI;1fI;tI;��I;��I;S�I;�I;.�I;��I;��I;@�I;َI;��I;      R�I;ޛI;��I;��I;ܔI;��I;��I;7�I;KvI;�kI;�`I;/VI;�KI;�AI;�7I;�.I;c&I;�I;�I;LI;�I;{I; I;G�H;��H;��H;c�H;H�H;c�H;��H;��H;��H;��H;&�H;��H;��H;R�H;��H;��H;)�H;��H;��H;��H;��H;_�H;H�H;_�H;��H;��H;C�H; I;{I;�I;II;�I;�I;c&I;�.I;�7I;�AI;�KI;.VI;�`I;�kI;OvI;7�I;��I;��I;�I;��I;��I;ۛI;      "|I;�{I;�yI;hvI;rI;�lI;)fI;#_I;}WI;�OI;�GI;g?I;R7I;�/I;�'I;� I;|I;nI;�I;�	I;NI;6I;��H;b�H;��H;M�H;0�H;a�H;��H;��H;��H;��H; �H;��H;�H;��H;��H;��H;�H;��H;��H;��H;��H;��H;��H;a�H;,�H;P�H;��H;_�H;��H;8I;II;�	I;�I;lI;{I;� I;�'I;}/I;R7I;c?I;�GI;�OI;WI;_I;/fI;�lI;	rI;ovI;�yI;�{I;      �[I;e[I;�YI;UWI;TI;�OI;KI;�EI;0@I;):I;�3I;�-I;�'I;�!I;�I;\I;=I;VI;�I;�I;V I;�H;�H;]�H;�H;,�H;m�H;��H;��H;��H;��H;��H;Y�H;��H;z�H;\�H;U�H;[�H;u�H;��H;Z�H;��H;��H;��H;��H;��H;i�H;-�H; �H;\�H;�H; �H;P I;�I;�I;VI;=I;]I;�I;�!I;�'I;�-I;�3I;+:I;0@I;�EI;(KI;�OI;TI;VWI;�YI;c[I;      �CI;WCI;6BI;b@I;�=I;�:I;&7I;	3I;�.I;�)I;*%I;k I;�I;�I;xI;I;
I;.I;�I;>�H;P�H;��H;2�H;'�H;!�H;^�H;��H;��H;��H;��H;��H;D�H;��H;O�H;�H;��H;��H;��H;�H;R�H;��H;B�H;��H;��H;��H;��H;��H;_�H;#�H;!�H;7�H;��H;J�H;:�H;�I;0I;
I;I;xI;�I;�I;h I;+%I;�)I;�.I;3I;,7I;�:I;�=I;i@I;=BI;ZCI;      2I;�1I;�0I;n/I;s-I;+I;B(I;!%I;�!I;!I;wI;�I;�I;�I;SI;�I;�I;wI;��H;��H;^�H;�H;�H;4�H;��H;�H;��H;��H;��H;�H;V�H;��H;5�H;��H;��H;��H;p�H;��H;��H;��H;3�H;��H;U�H;��H;��H;��H;��H;�H;��H;7�H;�H;�H;W�H;��H;��H;wI;�I;�I;SI;�I;�I;�I;zI;"I;�!I;%I;E(I;	+I;x-I;k/I;�0I;�1I;      �%I;S%I;�$I;�#I;"I; I;�I;KI;�I;�I;�I;eI;bI;\	I;QI;qI;� I;��H;a�H;;�H;A�H;<�H;g�H;��H;i�H;%�H;�H;�H;*�H;��H;��H;Q�H;��H;��H;^�H;;�H;'�H;;�H;^�H;��H;��H;R�H;��H;��H;%�H;��H;�H;%�H;n�H;��H;n�H;<�H;;�H;5�H;a�H;��H;� I;rI;OI;\	I;`I;cI;�I;�I;�I;HI;�I; I;"I;�#I;�$I;\%I;      QI;6I;�I;�I;VI;�I;�I;�I;]I;�I;aI;�
I;I;mI;�I;T I;��H;��H;x�H;v�H;��H;��H;]�H;��H;��H;g�H;b�H;��H;��H;�H;q�H;�H;��H;\�H;�H;�H;�H;�H;�H;_�H;��H;�H;q�H;
�H;��H;��H;b�H;i�H;��H;��H;c�H;��H;��H;r�H;x�H;��H;��H;X I;�I;oI;I;�
I;cI;�I;_I;�I;�I;�I;TI;�I;�I;8I;      �I;`I;�I;I;�I;vI;�I;�I;�I;�I;U
I;I;�I;*I;� I;�H;Z�H;N�H;b�H;|�H;��H;�H;��H;O�H;�H;�H;�H;A�H;��H;��H;Y�H;��H;��H;9�H;	�H;��H;��H;��H;�H;?�H;��H;��H;Y�H;��H;��H;A�H;�H;�H;�H;Q�H;��H;�H;��H;z�H;b�H;U�H;]�H;��H;� I;,I;�I;I;V
I;�I;�I;�I;�I;vI;�I;
I;�I;nI;      :I;I;�I;�I;vI;(I;}I;�I;�I;{I;X	I;I;�I;I;[ I;	�H;��H;��H;��H; �H;��H;��H;S�H;��H;��H;�H;�H;,�H;Y�H;��H;O�H;��H;s�H;#�H;�H;��H;��H;��H;�H;$�H;t�H;��H;Q�H;��H;S�H;)�H;�H;	�H;��H;��H;W�H;��H;��H;�H;��H;��H;��H;�H;[ I;�I;�I;I;[	I;|I;�I;�I;�I;(I;vI;�I;�I;I;      �I;aI;�I;I;�I;yI;�I;�I;�I;�I;T
I;I;�I;,I;� I;�H;Z�H;N�H;b�H;|�H;��H;�H;��H;O�H;�H;�H;�H;A�H;��H;��H;Y�H;��H;��H;;�H;	�H;��H;��H;��H;�H;=�H;��H;��H;Y�H;��H;��H;?�H;�H;�H;�H;P�H;��H;�H;��H;z�H;b�H;U�H;[�H;��H;� I;,I;�I;I;X
I;�I;�I;�I;�I;wI;�I;I;�I;hI;      GI;6I;�I;�I;VI;�I;�I;�I;]I;�I;bI;�
I;I;oI;�I;T I;��H;��H;z�H;v�H;��H;��H;_�H;��H;��H;f�H;b�H;��H;��H;�H;p�H;�H;��H;\�H;�H;�H;�H;�H;�H;_�H;��H;�H;q�H;	�H;��H;��H;b�H;j�H;��H;��H;c�H;��H;��H;r�H;z�H;��H;��H;X I;�I;pI;I;�
I;cI;�I;_I;�I;�I;�I;XI;�I;�I;=I;      �%I;S%I;�$I;�#I;"I; I;�I;NI;�I;�I;�I;dI;`I;\	I;RI;qI;� I;��H;c�H;9�H;A�H;?�H;j�H;��H;l�H;%�H;�H;�H;,�H;��H;��H;Q�H;��H;��H;_�H;9�H;'�H;;�H;\�H;��H;��H;R�H;��H;��H;%�H;��H;�H;(�H;o�H;��H;n�H;=�H;;�H;6�H;d�H;��H;� I;tI;TI;^	I;aI;dI;�I;�I;�I;KI;�I; I;"I;�#I;�$I;T%I;      	2I;�1I;�0I;h/I;p-I;+I;B(I;&%I;�!I;!I;wI;�I;�I;�I;VI;�I;�I;wI;��H;��H;\�H;�H;�H;7�H;��H;�H;��H;��H;��H;�H;U�H;��H;3�H;��H;��H;��H;p�H;��H;��H;��H;2�H;��H;U�H;��H;��H;��H;��H;�H;��H;4�H;�H;�H;U�H;��H;��H;wI;�I;�I;SI;�I;�I;�I;xI;"I;�!I;#%I;I(I;+I;w-I;u/I;�0I;�1I;      �CI;YCI;,BI;b@I;�=I;�:I;*7I;3I;�.I;�)I;.%I;k I;�I;�I;{I;I;
I;0I;�I;>�H;Q�H;��H;4�H;&�H;#�H;^�H;��H;��H;��H;��H;��H;A�H;��H;N�H;�H;��H;��H;��H;�H;O�H;��H;B�H;��H;��H;��H;��H;��H;a�H;!�H;�H;9�H;��H;I�H;:�H;�I;0I;
I;I;zI;�I;�I;l I;-%I;�)I;�.I;3I;*7I;�:I;�=I;i@I;/BI;VCI;      �[I;h[I;�YI;OWI;TI;�OI;KI;�EI;0@I;):I;�3I;�-I;�'I;�!I;�I;]I;?I;VI;�I;�I;W I;�H;�H;]�H; �H;)�H;j�H;��H;��H;��H;~�H;��H;Y�H;��H;z�H;[�H;T�H;\�H;u�H;��H;Z�H;��H;��H;��H;��H;��H;j�H;/�H;�H;Y�H;�H;�H;P I;�I;�I;VI;@I;_I;�I;�!I;�'I;�-I;�3I;+:I;1@I;�EI;%KI;�OI;TI;\WI;�YI;g[I;      +|I;�{I;�yI;svI;�qI;�lI;)fI;&_I;�WI;�OI;�GI;g?I;S7I;�/I;�'I;� I;|I;oI;�I;�	I;PI;9I;��H;`�H;��H;L�H;0�H;b�H;��H;��H;��H;��H;��H;��H;�H;��H;��H;��H;�H;��H;��H;��H;��H;��H;��H;_�H;/�H;Q�H;��H;\�H;��H;9I;JI;�	I;�I;nI;{I;� I;�'I;�/I;R7I;d?I;�GI;�OI;|WI;#_I;+fI;�lI;rI;yvI;�yI;�{I;      Y�I;ޛI;��I;��I;ΔI;��I;��I;5�I;TvI;�kI;�`I;0VI;�KI;�AI;�7I;�.I;c&I;�I;�I;JI;�I;|I;I;H�H;��H;��H;b�H;I�H;c�H;��H;��H;��H;��H;&�H;��H;��H;P�H;��H;��H;&�H;��H;��H;��H;��H;^�H;D�H;a�H;��H;��H;@�H;!I;|I;�I;JI;�I;�I;b&I;�.I;�7I;�AI;�KI;,VI;�`I;�kI;PvI;7�I;��I;��I;��I;��I;��I;؛I;      ��I;��I;ώI;?�I;��I;��I;/�I;'�I;U�I; �I;��I;tI;1fI;�XI;BLI;y@I;�5I;�+I;�"I;�I;�I;<I;�I;�I;��H;��H;��H;a�H;K�H;\�H;��H;��H;��H;��H;��H;?�H;)�H;A�H;��H; �H;��H;��H;��H;^�H;E�H;\�H;��H; �H;��H;�I;�I;;I;�I;�I;�"I;�+I;�5I;y@I;ALI;�XI;2fI;tI;��I;��I;T�I; �I;/�I;��I;��I;@�I;ڎI;��I;      =�H;��H;,�H;I;v%I;\HI;�hI;�I;F�I;��I;�I;��I;�I;�vI;#fI;�VI;�HI;<I;�0I;+&I;I;6I;NI;ZI;>I;��H;�H;��H;j�H;0�H;l�H;��H;��H;�H;j�H;�H;�H;�H;h�H;	�H;��H;��H;o�H;2�H;h�H;��H;�H;��H;=I;TI;TI;6I;I;,&I;�0I;<I;�HI;�VI; fI;�vI;�I;��I;�I;��I;C�I;�I;�hI;WHI;|%I;I;/�H;��H;      [fF;�yF;�F;6G;sG;F�G;�YH;s�H;WI;�WI;v�I;ҘI;��I;��I;؅I;sI;�`I;<PI;�AI;�4I;)I;�I;~I;!I;�I;PI;��H;�H;��H;S�H;/�H;e�H;�H;-�H;t�H;�H;�H;�H;q�H;-�H;�H;f�H;3�H;T�H;��H; �H;��H;YI;�I;I;�I;�I;)I;�4I;�AI;:PI;�`I;sI;مI;��I;��I;ΘI;y�I;�WI;MI;k�H;�YH;6�G;sG;<G;ȱF;�yF;      R@@;Gp@;��@;��A;��B;:D;�EE;(gF;�dG;�2H;a�H;�8I;5yI;֗I;��I;��I;V~I;xiI;�VI;FI;�7I;�*I;; I;#I;`I;�I;;I;��H;��H;��H;�H;"�H;��H;p�H;��H;"�H;��H;"�H;��H;r�H;��H;"�H;!�H;��H;��H;��H;=I;�I;]I;!I;> I;�*I;�7I;FI;�VI;uiI;X~I;��I;��I;֗I;7yI;�8I;]�H;�2H;�dG;(gF;�EE;.D;��B;��A;��@;Ep@;      ��2;G%3;�U4;`16;��8;*7;;��=;Р@;�C;IE;�F;��G;��H;_<I;ցI;��I;�I;:�I;�pI;n[I;;II;�9I;,I;� I;I;I;QI;�I;J�H;b�H;^�H;+�H;;�H;��H;��H;^�H;�H;`�H;��H;��H;>�H;+�H;c�H;d�H;H�H;�I;SI;I;I;� I;,I;�9I;;II;o[I;�pI;9�I;�I;��I;ՁI;_<I;��H;��G;�F;HE;�C;ˠ@;��=; 7;;��8;{16;�U4;0%3;      Z�;ӻ;;�;��#;x);��.;�W4;+|9;A�=;1�A;�D;��F;rH;��H;~_I;œI;V�I;N�I;�uI;q^I;�JI;%:I;#,I;< I;zI;NI;�I;%I;��H;�H;6�H;�H;k�H;c�H;��H;U�H;��H;`�H;k�H;�H;6�H;�H;��H;!I;�I;QI;�I;8 I;",I;%:I;�JI;t^I;�uI;R�I;R�I;ƓI;~_I;��H;pH;��F;ވD;2�A;A�=;)|9;�W4;��.;v);��#;	�;;��;      ���:k��:���:c
�:Y+�:��;��;��;��&;V�/;D=7;ZD=;��A;�E;H7G;_�H;l8I;��I;	�I;��I;�wI;�_I;�JI;�9I;�*I;�I;4I;=I;�I;9I; �H;��H;�H;<�H;��H;�H;��H;�H;��H;;�H;�H;��H;�H;=I;I;<I;6I;�I;�*I;�9I;�JI;�_I; xI;��I;�I;�I;l8I;_�H;D7G;�E;��A;VD=;F=7;V�/;��&;��;��;��;�+�:Q
�:���:Y��:      0�x9З�9���9p	:��^:� �:�ɼ:�P�:��;�h;أ#;�</;�;8;��>;�oC;�fF;=(H;NI;�I;ĜI;��I;�wI;n^I;;II;�7I;)I;I;�I;�I;GI;M I;H�H;Q�H;=�H;��H;��H;��H;��H;��H;9�H;S�H;F�H;O I;LI;�I;�I;I;)I;�7I;<II;p^I;�wI;��I;ŜI;�I;LI;>(H;�fF;�oC;��>;�;8;�</;ڣ#;�h;��;�P�:�ɼ:� �:@�^:|	:��9H��9      ������D��>񳺈dt��F� �8��&:.��:%��:�Z;IC;7�&;�'3;!<;��A;�E;p�G;AI;\|I;ȜI;��I;�uI;r[I;FI;�4I;'&I;�I;LI;�	I;�I;9�H;��H;6�H;t�H;z�H;�H;{�H;q�H;2�H;��H;7�H;�I;�	I;JI;�I;+&I;�4I;FI;u[I;�uI;��I;ȜI;\|I;CI;n�G;�E;��A;<;�'3;6�&;FC;�Z;��:(��:��&: �8�Fเdt�P�J�ຖ���      N��;��`����g���7}�e�D����*x��(
�����9��:���:	;�;��.;��9;��@;�]E;n�G;AI;�I;�I;N�I;�pI;�VI;�AI;z0I;�"I;�I;�I;�I;�I;��H;]�H;w�H;`�H;��H;`�H;t�H;\�H;��H;�I;�I;�I;�I;�"I;}0I;�AI;�VI;�pI;P�I;	�I;�I;CI;m�G;�]E;��@;��9;��.;�;	;���:��:���9(
��*x�����g�D��7}��g��c���7��      ��?��<<��1��h!��z��B�b���n����-�:��}��8�&:d��:6��:��;#�+;ۍ8;A�@;�]E;m�G;JI;�I;U�I;9�I;riI;7PI;<I;�+I;�I;nI;SI;+I;qI;��H;��H;O�H;��H;Q�H;��H;��H;sI;(I;TI;nI;�I;�+I;<I;7PI;kiI;9�I;S�I;�I;GI;n�G;�]E;B�@;ۍ8;!�+;��;4��:d��:4�&:�}��>𳺀�-��n��b���B黴z��h!��1��<<�      a��P���I��z�������^��75��z���̻�눻�R�dt�P�x9D��:nm�:�h;c�*;ލ8;��@;�E;>(H;k8I;I;�I;R~I;�`I;�HI;�5I;b&I;qI;5I;�	I;�I;� I;��H;V�H;��H;V�H;��H;� I;�I;�	I;6I;tI;]&I;�5I;�HI;�`I;K~I;�I;I;k8I;9(H;�E;��@;܍8;b�*;�h;lm�:D��:P�x9dt��R��눻��̻�z��75��^����|����I��O��      '��b��
����\��HC���t����|���?���	�&���V�
���@���:��:�h;!�+;��9;��A;�fF;]�H;{_I;��I;��I;sI;�VI;u@I;�.I;� I;XI;I;�I;mI;Q I;~�H;�H;~�H;L I;hI;�I;	I;VI;� I;�.I;u@I;�VI;�rI;��I;��I;{_I;]�H;zfF;��A;��9; �+;�h;��:��:������V�&����	���?���|��t��HC��]������
�a�      ��t��p�-�d��Q�|�9�^*����a�ҼzI���o���'��ڻa6}�2���8���:hm�:��;��.;<;�oC;C7G;��H;ցI;ۜI;ԅI;fI;?LI;�7I;�'I;�I;tI;NI;KI;�I;� I;P I;� I;�I;JI;NI;qI;�I;�'I;�7I;?LI;fI;хI;ӜI;؁I;��H;C7G;�oC;<;��.;��;hm�:��:09�6��b6}��ڻ��'��o�zI��a�Ҽ���^*�|�9� �Q�-�d��p�      ��Ž4���̷�Q���z����}��Q�T�'����'C��*\��,<<��>n��,��@�>��:6��:�;�'3;��>;�E;kH;d<I;՗I;��I;�vI;�XI;�AI;y/I;�!I;�I;�I;T	I;cI;"I;tI;%I;aI;T	I;�I;�I;�!I;y/I;�AI;�XI;�vI;��I;˗I;d<I;pH;�E;��>;�'3;�;6��:B��:��8�຀n���>�,<<�*\��'C�����T�'��Q���}��z��Q��̷�4���      c.��3�Ȥ�V����͈Ž75�����YG�2��akּG����xC��>�^6}�����0�x9l��:	;5�&;�;8;��A;��F;��H;6yI;��I;�I;0fI;�KI;O7I;'I;�I;�I;[I;I;�I;�I;�I;I;XI;�I;�I;}'I;N7I;�KI;1fI;�I;��I;0yI;��H;��F;��A;�;8;7�&;	;f��:0�x9���_6}��>��xC�G���akּ2��YG����75��͈Ž��V��Ȥ��3�      Gx��s���d�M�N�_�3�|I����G����z����\�B*�	�ݼH���,<<��ڻ�V� dt�(�&:���:DC;�</;TD=;ۈD;��G;�8I;ȘI;��I;tI;+VI;\?I;�-I;b I;�I;]I;�
I;�I;I;�I;�
I;\I;�I;a I;�-I;\?I;+VI;tI;��I;ĘI;�8I;��G;ވD;SD=;�</;FC;���:0�&:(dt��V��ڻ,<<�H���	�ݼB*���\��z��G������|I�`�3�M�N���d��s�      ,l¾(��T������������d���7�x��8Sؽ[���d�C*�bkּ+\����'�(���R�0~��~�:�Z;ڣ#;@=7;/�A;�F;Z�H;q�I;�I;��I;�`I;�GI;�3I;'%I;tI;�I;TI;M
I;L	I;M
I;TI;�I;rI;$%I;�3I;�GI;�`I;��I;�I;n�I;V�H;�F;1�A;==7;ͣ#;�Z;x�:0~���R�(����'�+\��bkּC*��d�[��7Sؽx����7��d���������T���(��      �V������������Ͼ�d���ǆ�C�N��3��c�[����\�2��(C���o���	��눻L����9!��:�h;T�/;<�=;LE;�2H;�WI;��I;��I;�kI;�OI;%:I;�)I;"I;�I;�I;�I;xI;�I;�I;�I;"I;�)I;":I;�OI;�kI;��I;��I;�WI;�2H;IE;>�=;S�/;�h;#��:���9L��눻��	��o�(C��2����\�[���c཰3�C�N��ǆ��d����Ͼ���������      �,b�ý\��>M���5�<��0r��%l¾蝒�"&W��3�7Sؽ�z��YG����{I����?���̻��-�x
����:��;��&;|9;�C;�dG;NI;?�I;Q�I;SvI;}WI;,@I;�.I;�!I;�I;UI;�I;�I;�I;VI;�I;�!I;�.I;)@I;yWI;RvI;S�I;@�I;MI;�dG;�C;"|9;��&;��;&��:�
����-���̻��?�{I�����YG��z��7Sؽ�3�"&W�蝒�%l¾0r��<����5��>M�ý\�      ���$��Z���M䂿½\���1�����J˾蝒�C�N�x��H������U�'�b�Ҽ��|��z��n��>x����&:�P�:��;�W4;Ӡ@;(gF;c�H;�I;�I;2�I;_I;�EI;3I;!%I;DI;�I;�I;�I;�I;�I;DI; %I;3I;�EI;_I;1�I; �I;�I;c�H;#gF;Ҡ@;�W4;��;�P�:��&:Bx���n���z���|�b�ҼU�'����H���x��C�N�蝒��J˾�����1�½\�M䂿Z���$��      }߿�$ڿ.�ʿ����	����Ps�QX:����%l¾�ǆ���7����75���Q�����t���75�j�����`�8�ɼ:��;��.;��=;�EE;�YH;�hI;#�I;��I;(fI;KI;#7I;E(I;�I;�I;�I;wI;�I;�I;�I;E(I;%7I;KI;(fI;��I;&�I;�hI;�YH;�EE;��=;��.;��;�ɼ:��8���h���75��t������Q�75�������7��ǆ�%l¾���QX:��Ps�	�������.�ʿ�$ڿ      {�����p������ſ$���Ps���1�1r���d���d�|I�ΈŽ��}�^*�IC���^��B�u�D��F๚ �:��;p);7;;,D;3�G;THI;��I;��I;�lI;�OI;�:I;+I; I;�I;yI;-I;yI;�I; I;+I;�:I;�OI;�lI;��I;��I;WHI;;�G;*D; 7;;t);��;� �:�F�w�D��B��^�IC��^*���}�ΈŽ|I��d��d��1r����1��Ps�$����ſ��꿃p����      ��7��3�֢%�{��<����ſ	���½\�<����Ͼ����`�3��轻z��|�9�\�Ἑ���z��7}�pdt�0�^:e+�:��#;��8;��B;sG;o%I;��I;�I;rI;TI;�=I;p-I;"I;GI;�I;zI;�I;JI;"I;p-I;�=I;TI;	rI;�I;��I;v%I;sG;��B;��8;��#;g+�:�^:ldt��7}��z����\��|�9��z����`�3�������Ͼ<��½\�	�����ſ�<��{�֢%��3�      .�_��+Y��lG�f.�{���꿲���M䂿��5���󾍰��N�N�V��Q�� �Q����{����h!��g��V񳺌	:]
�:��;\16;��A;9G;�I;6�I;x�I;kvI;LWI;i@I;j/I;�#I;�I;	I;�I;I;�I;�#I;m/I;k@I;KWI;qvI;z�I;9�I;I;DG;��A;`16;��;]
�:t	:V񳺆g���h!�{������ �Q�Q��V��N�N���������5�M䂿�������{�f.��lG��+Y�      Ѭ��#}�>tf��lG�ע%��p�.�ʿZ����>M����T�����d�Ȥ�̷�-�d��
��I���1�c���P����9���:;�U4;��@;ӱF;2�H;܎I;��I;�yI;�YI;6BI;�0I;�$I;�I;�I;�I;�I;�I;�$I;�0I;7BI;�YI;�yI;��I;��I;8�H;�F;��@;�U4;;���:���9H��b����1��I���
�-�d�̷�Ȥ���d�T�������>M�Z���.�ʿ�p�ע%��lG�>tf�#}�      S���D���#}��+Y��3�����$ڿ$��ý\����(���s��3�5����p�b�R���<<�6���������9U��:ӻ;R%3;Kp@;�yF;��H;��I;�I;�{I;L[I;LCI;�1I;Q%I;I;TI;I;QI;I;P%I;�1I;OCI;H[I;�{I;�I;��I;��H;�yF;Hp@;S%3;л;O��:���9����7���<<�R��b��p�5����3��s�(�����ý\�$���$ڿ����3��+Y�#}�D���      ����,������T���J�Q�ř$�4�����<�}�H(�?�׾�T���L+���սj��
��L���iO���ͻ��� #m8vo�:`�;X�1;��?;�uF;j I;i�I;��I;��I;YvI;�WI;�AI;�1I;�'I;�!I;�I;�!I;�'I;�1I;�AI;�WI;XvI;��I;��I;l�I;m I;�uF;��?;V�1;^�;po�:�!m8�����ͻ�iO�L��
��j����ս�L+��T��?�׾H(�<�}���4���ř$�J�Q�T��������,��      �,��a��#P���{���K��x �����p�����w��$���Ҿf���  (���ѽѷ��&������K�Aɻ#��`��8���:~�;��1;�@;p�F;!I;߿I;�I;��I;�uI;%WI;hAI;�1I;�'I;�!I;�I;�!I;�'I;�1I;hAI;&WI;�uI;��I;�I;�I;%I;|�F;�@;��1;~�;~��:���8 ��Aɻ��K����&�ѷ����ѽ  (�f�����Ҿ�$���w�p��������x ���K��{�#P��a��      ����#P�������d���;�#���㿲���#f�d��ž��z���;�ƽ$0v�S5�0����o@�����vi� au9KK�:];�73;&�@;��F;JI;��I;P�I;V�I;�sI;�UI;B@I;�0I;�&I;!I;0I;!I;�&I;�0I;A@I;�UI;�sI;Y�I;P�I;��I;MI;��F;%�@;�73;];EK�: au9ri������o@�0���S5�$0v�;�ƽ����z�žd��#f�������#����;���d����#P��      T����{���d��F�ř$�:����ɿ.蒿��K�P���j���Yb�F�0���r�a����>�����.��d��b�غ ��9�Y�:2X;�25;'�A;\!G;L7I;v�I;D�I;S�I;�pI;�SI;�>I;{/I;�%I;" I;/I; I;�%I;v/I;>I;�SI;�pI;T�I;D�I;v�I;L7I;f!G;$�A;�25;2X;�Y�:��9\�غ�d����.�>������r�a�0���F��Yb��j��P����K�.蒿��ɿ:��ř$��F���d��{�      J�Q���K���;�ř$��;
��޿�����w�r,���澝���&�D������I��#�G�����N��������H�����9:d��:�n!;��7;��B;M�G;�YI;,�I;Z�I;��I;�lI;uPI;<I;�-I;$I;�I;�I;�I;$I;�-I;<I;uPI;�lI;��I;Z�I;/�I;�YI;U�G;��B;��7;�n!;d��:��9:B����������N�����#�G��I������&�D��������r,���w�����޿�;
�ř$���;���K�      ř$��x �"��9���޿o���Ʌ���F�}�
��~����z��$���ս���@2+���ϼPp�����F�]� �*�"��:�;�8';��:;��C; H;�}I;�I;q�I;ًI;mgI;�LI; 9I;9+I;""I;�I;)I;�I; "I;4+I;9I;�LI;hgI;ۋI;s�I;"�I;�}I;H;��C;��:;�8';�;��:�*�F�]�����Pp���ϼ@2+������ս�$���z��~��}�
��F�Ʌ��o����޿9��"���x �      4��������㿊�ɿ���Ʌ����P�c��;�׾�`��S�H����@��Q�a���ˡ���D��ɻ� ��׭��W�:�;fI-;;|=;!CE;��H;�I;��I;u�I;��I;iaI;#HI;�5I;p(I;�I;�I;QI;�I;�I;p(I;�5I;"HI;faI;��I;v�I;��I;�I;��H;&CE;;|=;dI-;�;�W�: ׭�� ��ɻ�D�ˡ����Q�a��@����S�H��`��;�׾d����P�Ʌ�������ɿ�㿳���      ��p�������.蒿��w��F�c��ʰ� ����Yb�)����ѽ�%��D4�ן�X����� H���潺��9Pr�:��;�93;*Q@;~vF;�H;�I;��I;��I;�zI;�ZI;CI;�1I;b%I;?I;�I;"I;�I;BI;c%I;�1I;CI;�ZI;�zI;��I;��I;�I;�H;�vF;'Q@;�93;��;Jr�:��9�潺�G�����X��֟�D4��%����ѽ)���Yb� ���ʰ�c���F���w�.蒿����p���      <�}���w�#f���K�q,�}�
�;�׾ �����k���'�dz꽝I���;V�<M�����iO�fG�ioE����D��:I� ;��$;��8;_�B;��G;/KI;�I;�I;A�I;	qI;�SI;�=I;�-I;"I;jI;I;�I;I;mI;"I;�-I;�=I;�SI;qI;D�I;�I;�I;/KI; �G;_�B;��8;��$;G� ;R��:���hoE�eG໨iO����;M��;V��I��dz���'���k� ���;�׾}�
�r,���K�#f���w�      G(��$�d��P������~���`���Yb���'��U�F$��C�m�%����ϼ�/��;��������غp8�9D��:�F;�G.;|=;KE;�\H;�I;v�I;z�I;��I;gI; LI;�7I;)I;pI;rI;rI;'I;qI;rI;pI;)I;�7I;LI;gI;��I;�I;u�I;�I;�\H;KE;|=;�G.;�F;V��:�8�9��غ����;���/����ϼ%��C�m�F$���U���'��Yb��`���~�����P��d���$�      ?�׾��Ҿž�j��������z�S�H�)��dz�F$���/v�2+�ݐ�����5��ɻ24� (�����:f��:<o!;P6;
lA;��F;t�H;��I;��I;�I;G}I;�\I;[DI;	2I;r$I;�I;HI;�I;�I;�I;II;�I;r$I;2I;^DI;�\I;M}I;�I;��I;��I;z�H;��F;lA;P6;=o!;|��:���:�'��+4��ɻ��5���ܐ�2+��/v�F$��dz�)��S�H���z������j��ž��Ҿ      �T��f�����z��Yb�&�D��$�����ѽ�I��C�m�2+�������I�K��ﻎ�p�<������91T�:�/;v�-;j�<;FzD;_H;�mI;��I;}�I;��I;�oI;�RI;�<I;,I;�I;I;/I;�I;�I;�I;.I;I;�I;,I;�<I;�RI;�oI;��I;}�I;��I;�mI;_H;LzD;q�<;x�-;�/;;T�:��9.�����p���H�K�������2+�C�m��I����ѽ���$�&�D��Yb���z�f���      �L+�  (���F�������ս�@���%���;V�$��ܐ�����~MS�J��!��fD���n8q�:�;h�$;_7;.�A;h�F;��H;b�I;d�I;��I;�I;QbI;�HI;5I;(&I;/I;>I;�I;�
I;
I;�
I;�I;>I;/I;%&I;5I;�HI;XbI;�I;��I;b�I;i�I;��H;k�F;5�A;_7;s�$;�;q�: �n8`D� ��I��}MS�����ܐ�$���;V��%���@����ս����F�����'�      ��ս��ѽ;�ƽ0����I�����Q�a�D4�;M���ϼ��H�K�L��HG��Wf�0�o���:�B�:�Y;��1;Ul>;�E;�/H;#qI;��I;��I;ܘI; sI;�UI;�>I;�-I;b I;�I;�I;�
I;I;0I;I;�
I;�I;�I;` I;�-I;�>I;�UI;sI;ژI;��I;�I;#qI;�/H;�E;Wl>;��1;�Y;�B�:��:P�o�Tf�FG��K��H�K�����ϼ;M�D4�P�a�����I��0���;�ƽ��ѽ      i��ѷ��$0v�q�a�#�G�?2+���՟�����/����5���"��Vf�xج��g:E�:�;I-;g;;OC;SG;�I;ͶI;�I; �I;
�I;
cI;~II;�5I;n&I;�I;7I;�I;�I;PI;XI;NI;�I;�I;9I;�I;t&I;�5I;�II;cI;
�I;��I; �I;ͶI;�I;SG;OC;"g;;I-;�;O�:�g:xج�Sf�!������5��/�����՟���?2+�$�G�q�a�$0v�ѷ��      	��&�S5���������ϼʡ��X���iO�;���ɻ��p�tD�0�o��g:`�:JG;v*;v9;��A;�uF; �H;ƔI;��I;��I;I�I;�pI;4TI;M>I;-I;�I;}I;�I;VI;�I;�I;�I;�I;�I;VI;�I;zI;�I;-I;R>I;:TI;�pI;D�I;��I;��I;ƔI;%�H;�uF;��A;y9;t*;LG;`�:�g:P�o�tD⺎�p��ɻ:���iO�X��ˡ����ϼ������S5�%�      L�����0���>����N��Pp��D����bG�����+4�.��� �n8��:M�:QG;
�(;��7;`�@;��E;QQH;mI;��I;��I;��I;&}I;�^I;�FI;�3I;�$I;\I;�I;�	I;I;�I;��H;O�H;��H;�I;I;�	I;�I;aI;�$I;�3I;�FI;�^I;!}I;��I;��I;��I;mI;UQH;��E;c�@;��7;�(;OG;S�:��:��n8.���'4�����bGໄ���D�Pp��N��?���2������      �iO�ޔK��o@���.���������ɻ�G��coE���غ�'����9q�:�B�:�;t*;��7;�P@;�\E;�H;�II;��I;m�I;�I;Y�I;?hI;�NI;c:I;9*I;xI;�I;�I;I;I;2�H;a�H;��H;\�H;/�H;I;I;�I;�I;{I;:*I;f:I;�NI;;hI;a�I;�I;g�I;��I;�II;�H;�\E;�P@;��7;r*;�;�B�:q�:��9�'����غ_oE��G���ɻ����~����.��o@�ޔK�      ��ͻFɻ�����d�����5�]�� ��潺����8�9���:=T�:�;�Y;"I-;}9;a�@;�\E;��G;55I;��I;G�I;ߵI;V�I;epI;�UI;V@I;4/I;}!I;�I;@I;�I;�I;"�H;��H;�H;��H;�H;��H;!�H;�I;�I;CI;�I;}!I;9/I;S@I;�UI;npI;Y�I;صI;J�I;��I;95I;��G;�\E;d�@;w9; I-;�Y;�;=T�:���:�8�9����潺� �=�]�����d������Fɻ      ���%��ni�H�غT����*� ֭�В�9N��:V��:z��:�/;p�$;��1;"g;;��A;��E;�H;75I;=�I;��I;P�I;��I;�vI;O[I;aEI;�3I;6%I;�I;�I;P	I;�I;}�H;a�H;'�H;��H;n�H;��H;"�H;`�H;}�H;�I;Q	I;�I;�I;9%I;�3I;^EI;W[I;�vI;��I;P�I;��I;?�I;:5I;�H;��E;��A; g;;��1;l�$;�/;~��:R��:R��: ��9`֭�Ї*�F���b�غyi�3��      �+m8 ��8�_u9Ȱ�9x�9:$��:�W�:Xr�:G� ;�F;=o!;y�-;_7;Yl>;OC;�uF;UQH;�II;��I;��I;��I;��I;�zI;�_I;?II;N7I;d(I;aI;�I;I;�I;, I;u�H;��H;�H;��H;u�H;��H;�H;��H;p�H;& I;�I;I;�I;dI;a(I;K7I;DII;�_I;{zI;��I;��I;��I;��I;�II;UQH;�uF;OC;Rl>;_7;v�-;Bo!;�F;D� ;Nr�:�W�:��:��9:���9@`u9���8      ho�:���:aK�:�Y�:R��: �;�;��;��$;�G.;P6;q�<;1�A;�E;SG;'�H;mI;��I;L�I;T�I;��I;�{I;zaI;�KI;�9I;�*I;�I;�I;�I;'I;� I;��H;��H;k�H;��H;�H;��H;�H;��H;j�H;��H;��H;� I;(I;�I;�I;�I;�*I;�9I;�KI;saI;�{I;��I;Q�I;L�I;��I;mI;$�H;SG;�E;2�A;q�<;P6;�G.;��$;��;�;�;���:�Y�:OK�:���:      u�;~�;];@X;�n!;�8';rI-;�93;��8;|=;lA;TzD;n�F;�/H;�I;ΔI;��I;o�I;ߵI;��I;�zI;waI;zLI;!;I;a,I;3 I;!I;�I;=I;�I;w�H;��H;g�H;o�H;
�H;U�H;"�H;O�H;�H;p�H;e�H;��H;z�H;�I;9I;�I;I;3 I;g,I;;I;sLI;xaI;�zI;��I;ߵI;j�I;��I;˔I;�I;�/H;l�F;SzD;lA;|=;��8;�93;pI-;�8';�n!;@X;];b�;      U�1;��1;�73;�25;��7;��:;7|=;(Q@;X�B;NE;��F;`H;��H;&qI;ͶI;��I;��I;�I;V�I;�vI;�_I;�KI;;I;�,I;� I;I;�I;I;uI;��H;r�H;n�H;#�H;��H;q�H;��H;��H;��H;n�H;��H;!�H;m�H;w�H;��H;qI;I;�I;I;� I;�,I;;I;�KI;�_I;�vI;S�I;�I;��I;��I;̶I; qI;��H;`H;��F;KE;\�B;.Q@;5|=;��:;��7;�25;�73;��1;      ��?;�@;�@; �A;��B;�C;(CE;�vF;��G;�\H;~�H;�mI;f�I;
�I;#�I;��I;��I;f�I;spI;\[I;JII;�9I;h,I;� I;rI;aI;�I;�I;j�H;��H;��H;.�H;W�H;��H;��H;^�H;3�H;X�H;��H;��H;U�H;(�H;��H;��H;f�H;�I;�I;aI;uI;� I;d,I;�9I;LII;W[I;rpI;a�I;��I;��I;#�I;�I;f�I;�mI;|�H;�\H;��G;~vF;*CE;��C;��B;�A;�@;�@;      �uF;|�F;��F;]!G;C�G;H;��H;#�H;5KI;+�I;��I;��I;f�I;��I;�I;M�I;+}I;AhI;�UI;^EI;O7I;�*I;0 I;I;]I;�I;HI;��H;��H;��H;'�H;@�H;��H;^�H;��H;�H;��H;�H;��H;`�H;��H;;�H;'�H;��H;��H;��H;BI;�I;aI;I;. I;�*I;N7I;\EI;�UI;>hI;*}I;O�I; �I;��I;f�I;��I;��I;(�I;5KI; �H;��H; H;Z�G;j!G;��F;{�F;      x I;-I;BI;P7I;�YI;�}I;�I;�I;�I;z�I;��I;��I;��I;��I;
�I;�pI;�^I;�NI;Z@I;�3I;k(I;�I;$I;�I;�I;GI;��H;%�H;��H;2�H;#�H;j�H;�H;�H;��H;	�H;��H;�H;�H;�H;�H;f�H;#�H;1�H;��H;#�H;��H;II;�I;�I;"I;�I;i(I;�3I;W@I;�NI;�^I;�pI;�I;ژI;��I;��I;��I;v�I;�I;�I;�I;�}I; ZI;E7I;BI;I;      e�I;�I;��I;{�I;�I; �I;��I;��I;�I;��I;�I;��I;�I;sI;cI;7TI;�FI;`:I;6/I;5%I;eI;�I;�I;I;�I;��H;%�H;��H;F�H;"�H;Z�H;��H;��H;�H;[�H;�H;��H;��H;Z�H;�H;��H;��H;Z�H;!�H;B�H;��H;�H;��H;�I;I;�I;�I;dI;4%I;4/I;]:I;�FI;:TI;cI;sI;�I;��I;�I;��I;�I;��I;��I;�I;(�I;}�I;��I;ۿI;      ��I;��I;H�I;T�I;P�I;s�I;y�I;��I;=�I;��I;P}I;�oI;XbI;�UI;�II;T>I;�3I;?*I;�!I;�I;�I;�I;7I;pI;c�H;��H;��H;D�H;3�H;W�H;��H;��H;��H;��H;|�H;5�H;.�H;1�H;z�H;��H;��H;��H;��H;U�H;-�H;C�H;��H;��H;g�H;nI;:I;�I;�I;�I;�!I;<*I;�3I;U>I;�II;�UI;UbI;�oI;S}I;��I;A�I;��I;|�I;m�I;Z�I;X�I;L�I;��I;      ��I;��I;a�I;P�I;��I;ًI;��I;�zI;qI;gI;�\I;�RI;�HI;�>I;�5I;-I;�$I;wI;�I;�I;#I;"I;�I;��H;��H;��H;2�H;%�H;\�H;��H;��H;��H;��H;�H;��H;|�H;]�H;{�H;��H;�H;��H;��H;��H;��H;X�H;%�H;-�H;��H;��H;��H;�I;%I;I;�I;�I;vI;�$I;!-I;�5I;�>I;�HI;�RI;�\I;gI;qI;�zI;��I;ڋI;��I;Y�I;`�I;��I;      YvI;�uI;�sI;�pI;�lI;mgI;jaI;�ZI;�SI;
LI;dDI;�<I;5I;�-I;x&I;�I;fI;�I;FI;W	I;�I;� I;v�H;r�H;��H;#�H;"�H;^�H;��H;��H;��H;��H;��H;\�H;�H;��H;��H;��H;
�H;^�H;��H;��H;��H;��H;��H;[�H;!�H;&�H;��H;r�H;z�H;� I;�I;T	I;GI;�I;fI;�I;w&I;�-I;5I;�<I;bDI;LI;�SI;�ZI;saI;egI;�lI;�pI;�sI;�uI;      �WI;/WI;�UI;�SI;gPI;�LI;#HI;CI;�=I;�7I;2I;,I;+&I;i I;�I;~I;�I;�I;�I;�I;3 I;��H;��H;j�H;+�H;6�H;e�H;��H;��H;��H;��H;��H;E�H;��H;|�H;A�H;K�H;C�H;z�H;��H;H�H;��H;��H;��H;��H;��H;c�H;7�H;.�H;d�H;�H;��H;, I;�I;�I;�I;�I;�I;�I;i I;+&I;
,I;2I;�7I;�=I;CI;)HI;�LI;rPI;�SI;�UI;2WI;      �AI;wAI;F@I;�>I;<I;9I;�5I;�1I;�-I;	)I;u$I;�I;2I;�I;<I;�I;�	I;I;�I;��H;}�H;��H;d�H;�H;U�H;��H;�H;��H;��H;��H;��H;D�H;��H;]�H;�H;��H;��H;��H;�H;`�H;��H;H�H;��H;��H;��H;��H;�H;��H;Y�H;�H;h�H;��H;w�H;��H;�I;I;�	I;�I;=I;�I;3I;�I;y$I;)I;�-I;�1I;�5I;9I;<I;�>I;S@I;wAI;      �1I;�1I;�0I;r/I;�-I;,+I;s(I;j%I;"I;{I;�I;I;GI;�I;�I;[I;I;I;%�H;e�H;��H;j�H;l�H;��H;��H;T�H;�H;�H; �H; �H;Y�H;��H;_�H;��H;��H;��H;~�H;��H;��H;��H;`�H;��H;Y�H;�H;��H;�H;�H;V�H;��H;��H;q�H;h�H;��H;`�H;%�H;I;I;]I;�I;�I;EI;I;�I;{I;"I;h%I;y(I;-+I;�-I;v/I;�0I;�1I;      �'I;�'I;�&I;�%I;$I;"I;�I;NI;tI;�I;VI;@I;�I;�
I;�I;�I;�I;2�H;��H;(�H;�H;��H;�H;b�H;��H;��H;x�H;^�H;��H;��H;	�H;|�H;�H;��H;��H;\�H;X�H;a�H;~�H;��H;�H;�H;�H;��H;z�H;Z�H;z�H;��H;��H;c�H;
�H;��H;�H;"�H;��H;4�H;�I;�I;�I;�
I;�I;@I;XI;�I;tI;MI;�I;"I;$I;�%I;�&I;�'I;      �!I;�!I;!I;" I;�I;�I;�I;�I;I;}I;�I;�I;�
I;I;UI;�I;��H;^�H;�H;��H;��H;�H;N�H;��H;T�H;�H;�H;�H;<�H;��H;��H;D�H;��H;��H;a�H;+�H;.�H;/�H;_�H;��H;��H;G�H;��H;{�H;8�H;�H;�H;�H;W�H;��H;R�H;�H;��H;��H;�H;c�H;��H;�I;XI;"I;�
I;�I;�I;}I;I;�I;�I;�I;�I;% I;!I;�!I;      �I;�I;BI;.I;�I;%I;XI;,I;�I;,I;�I;�I;
I;=I;dI;�I;Z�H;��H;��H;s�H;��H;��H;�H;��H;-�H;��H;��H;��H;3�H;a�H;��H;K�H;��H;{�H;W�H;(�H;�H;-�H;T�H;~�H;��H;N�H;��H;\�H;.�H;��H;��H;��H;.�H;��H;"�H;��H;x�H;p�H;��H;��H;Z�H;�I;dI;@I;
I;�I;�I;.I;�I;*I;\I;%I;�I;3I;@I;�I;      �!I;�!I;!I; I;�I;�I;�I;�I;I;|I;�I;�I;�
I;I;UI;�I;��H;^�H;�H;��H;��H;�H;N�H;��H;T�H;�H;�H;�H;>�H;�H;��H;G�H;��H;��H;b�H;+�H;.�H;.�H;_�H;��H;��H;G�H;��H;y�H;8�H; �H;�H;�H;W�H;��H;R�H;�H;��H;��H;�H;c�H;��H;�I;WI;I;�
I;�I;�I;{I; I;�I;�I;�I;�I;) I;!I;�!I;      �'I;�'I;�&I;�%I;$I;"I;�I;QI;tI;�I;WI;BI;�I;�
I;�I;�I;�I;3�H;��H;(�H;�H;��H;�H;`�H;��H;��H;x�H;^�H;��H;��H;�H;|�H;�H;��H;��H;^�H;X�H;a�H;�H;��H;�H;~�H;�H;��H;z�H;X�H;z�H;��H;��H;b�H;
�H;��H;�H;$�H;��H;6�H;�I;�I;�I;�
I;�I;BI;XI;�I;uI;QI;�I;"I;$I;�%I;�&I;�'I;      �1I;�1I;�0I;u/I;�-I;3+I;r(I;m%I;"I;zI;�I;I;EI;�I;�I;[I;I;I;&�H;d�H;��H;k�H;l�H;��H;��H;V�H;�H;�H;�H;�H;W�H;��H;_�H;��H;��H;��H;~�H;��H;��H;��H;`�H;��H;W�H;�H;��H;�H;�H;W�H;��H;��H;q�H;k�H;��H;a�H;(�H;I;I;`I;�I;�I;GI;I;�I;{I;"I;i%I;|(I;0+I;�-I;y/I;�0I;�1I;      �AI;}AI;J@I;~>I;<I;9I;�5I;�1I;�-I;	)I;v$I;�I;3I;�I;?I;�I;�	I;I;�I;��H;}�H;��H;c�H;�H;V�H;��H;�H;��H;��H;��H;��H;D�H;��H;\�H;�H;��H;��H;��H;�H;]�H;��H;G�H;��H;��H;��H;��H;�H;��H;V�H;�H;j�H;��H;v�H;��H;�I;I;�	I;�I;?I;�I;4I;�I;w$I;)I;�-I;�1I;�5I;9I;<I;�>I;W@I;xAI;      �WI;2WI;�UI;�SI;hPI;�LI;'HI;CI;�=I;�7I;2I;,I;,&I;i I;�I;�I;�I;�I;�I;�I;4 I;��H;��H;g�H;.�H;7�H;e�H;��H;��H;��H;��H;��H;E�H;��H;~�H;A�H;K�H;D�H;z�H;��H;G�H;��H;��H;��H;��H;��H;b�H;9�H;+�H;a�H;�H;��H;, I;�I;�I;�I;�I;�I;�I;k I;.&I;,I;2I;�7I;�=I;CI;*HI;�LI;iPI;�SI;�UI;/WI;      OvI;�uI;�sI;�pI;�lI;ngI;maI;�ZI;�SI;
LI;eDI;�<I;5I;�-I;z&I;�I;iI;�I;GI;U	I;�I;� I;w�H;r�H;��H;!�H;!�H;^�H;��H;��H;��H;��H;��H;\�H;�H;��H;��H;��H;
�H;^�H;��H;��H;��H;��H;��H;[�H;!�H;'�H;��H;n�H;{�H;� I;�I;U	I;HI;�I;iI;�I;{&I;�-I;5I;�<I;eDI;
LI;�SI;�ZI;saI;jgI;�lI;�pI;�sI;�uI;      ��I;��I;\�I;Y�I;��I;�I;��I;�zI;qI;gI;�\I;�RI;�HI;�>I;�5I; -I;�$I;xI;�I;�I;%I;'I;�I;��H;��H;��H;1�H;&�H;^�H;��H;��H;��H;��H;�H;��H;{�H;]�H;|�H;��H;�H;��H;��H;��H;��H;X�H;"�H;.�H;��H;��H;��H;�I;'I;!I;�I;�I;wI;�$I;!-I;�5I;�>I;�HI;�RI;�\I;gI;qI;�zI;��I;׋I;��I;b�I;f�I;��I;      ��I;��I;Z�I;P�I;A�I;z�I;w�I;��I;G�I;��I;P}I;�oI;VbI;�UI;�II;V>I;�3I;@*I;!I;�I;�I;�I;9I;rI;g�H;��H;��H;D�H;2�H;T�H;��H;��H;��H;��H;|�H;4�H;-�H;4�H;z�H;��H;��H;��H;��H;U�H;,�H;@�H;��H;��H;d�H;jI;;I;�I;�I;�I;�!I;<*I;�3I;Y>I;�II;�UI;XbI;�oI;P}I;��I;B�I;��I;}�I;t�I;P�I;Q�I;Z�I;��I;      r�I;ۿI;��I;{�I;�I;-�I;��I;��I;�I;��I;�I;��I;�I;sI;cI;:TI;�FI;b:I;6/I;5%I;gI;�I;�I;I;�I;��H;!�H;��H;F�H;�H;X�H;��H;��H;�H;\�H;��H;��H; �H;[�H;�H;��H;��H;Z�H;�H;B�H;��H;!�H;��H;�I;I;�I;�I;bI;5%I;7/I;_:I;�FI;;TI;cI;sI;�I;��I;�I;��I;�I;��I;��I;�I;'�I;}�I;��I;ۿI;      g I;6I;BI;W7I;�YI;�}I;�I;�I;�I;y�I;��I;��I;��I;ޘI;�I;�pI;�^I;�NI;X@I;�3I;l(I;�I;!I;�I;�I;BI;��H;%�H;��H;/�H;"�H;i�H;�H;�H;��H;�H;��H;�H;~�H;�H;�H;i�H;%�H;1�H;��H;"�H;��H;LI;�I;�I;%I;�I;i(I;�3I;Z@I;�NI;�^I;�pI;
�I;ܘI;��I;~�I;��I;v�I;�I;�I;�I;�}I;�YI;Z7I;CI;I;      �uF;|�F;��F;X!G;I�G;H;��H;$�H;9KI;'�I;��I;��I;f�I;��I;�I;P�I;*}I;ChI;�UI;^EI;S7I;�*I;. I;I;`I;�I;EI;��H;��H;��H;&�H;>�H;��H;]�H;��H;�H;��H;�H;��H;]�H;��H;>�H;(�H;��H;��H;��H;GI;�I;^I;I;0 I;�*I;O7I;_EI;�UI;>hI;-}I;P�I;�I;��I;f�I;��I;��I;+�I;/KI;�H;��H;H;T�G;]!G;��F;n�F;      ��?;�@;�@;�A;��B;
�C;*CE;�vF;�G;�\H;~�H;�mI;f�I;	�I;'�I;��I;��I;f�I;spI;Y[I;LII;�9I;g,I;� I;uI;ZI;�I;�I;j�H;��H;��H;-�H;U�H;��H;��H;[�H;3�H;[�H;��H;��H;W�H;-�H;��H;��H;f�H;�I;�I;cI;rI;� I;i,I;�9I;LII;Z[I;vpI;c�I;��I;��I;&�I;	�I;h�I;�mI;{�H;�\H;��G;~vF;*CE;��C;��B;�A;�@;�@;      6�1;��1;�73;�25;�7;��:;5|=;(Q@;`�B;IE;��F;cH;��H;"qI;жI;��I;��I;�I;U�I;�vI;�_I;�KI;;I;�,I;� I;I;�I;I;uI;��H;t�H;o�H;!�H;��H;m�H;��H;��H;��H;m�H;��H;&�H;o�H;x�H;��H;tI;I;�I;I;� I;�,I;;I;�KI;�_I;�vI;X�I;�I;��I;��I;ͶI;"qI;��H;`H;��F;IE;[�B;$Q@;7|=;��:;��7;�25;�73;��1;      l�;��;];HX;�n!;�8';nI-;�93;��8;|=;lA;SzD;l�F;�/H;�I;ΔI;��I;r�I;�I;��I;�zI;xaI;vLI;";I;g,I;* I;I;�I;>I;�I;x�H;��H;e�H;m�H;
�H;U�H;%�H;S�H;�H;l�H;e�H;��H;}�H;�I;:I;�I;"I;1 I;d,I;";I;wLI;xaI;�zI;��I;�I;m�I;��I;ΔI;�I;�/H;n�F;PzD;lA;|=;��8;�93;jI-;�8';�n!;JX;];j�;      jo�:���:WK�:�Y�:V��:(�;�;��;��$;�G.;P6;u�<;2�A;�E;SG;(�H;mI;��I;L�I;V�I;��I;�{I;vaI;�KI;�9I;�*I;�I;�I;�I;%I;� I;��H;��H;k�H;��H;�H;��H;�H;��H;h�H;��H;��H;� I;)I;�I;�I;�I;�*I;�9I;�KI;waI;�{I;��I;V�I;N�I;��I;mI;'�H;SG;�E;2�A;q�<;P6;�G.;��$;��;�;�;~��:�Y�:OK�:���:      @(m8���8�`u9ذ�9h�9:*��:�W�:Pr�:I� ;�F;Bo!;y�-;_7;Vl>;OC;�uF;UQH;�II;��I;��I;��I;��I;~zI;�_I;DII;H7I;a(I;bI;�I;I;�I;* I;s�H;��H;�H;��H;u�H;��H; �H;��H;s�H;) I;�I;I;�I;bI;b(I;L7I;BII;�_I;~zI;��I;��I;��I;��I;�II;UQH;�uF;OC;Wl>;_7;v�-;Co!;�F;E� ;Vr�:�W�:"��:��9:��9Pau9���8      q����oi�B�غT���܇*��֭�@��9Z��:P��:~��:�/;p�$;��1;%g;;��A;��E;�H;95I;?�I;��I;S�I;��I;�vI;V[I;[EI;�3I;5%I;�I;�I;Q	I;�I;}�H;b�H;'�H;��H;n�H;��H;"�H;]�H;|�H;�I;U	I;�I;�I;5%I;�3I;_EI;R[I;�vI;��I;Q�I;��I;?�I;:5I;�H;��E;��A;"g;;��1;o�$;�/;~��:L��:X��:��9`֭���*�J���\�غri� ��      ��ͻFɻ�����d�����5�]�� ��潺x���8�9���:=T�:�;�Y;&I-;}9;c�@;�\E;��G;95I;��I;K�I;ߵI;V�I;npI;�UI;S@I;6/I;!I;�I;AI;�I;�I;!�H;��H;�H;��H;�H;��H;�H;�I;�I;DI;�I;}!I;6/I;T@I;�UI;hpI;Z�I;ݵI;K�I;��I;95I;��G;�\E;c�@;y9;"I-;�Y;�;=T�:���:�8�9����潺� �8�]�����d������Bɻ      �iO�ܔK��o@���.��������ɻ�G��_oE���غ�'����9q�:�B�:�;t*;��7;�P@;�\E;�H;�II;��I;o�I;�I;a�I;<hI;�NI;d:I;=*I;wI;�I;�I;I;I;0�H;_�H;��H;a�H;-�H;I;I;�I;�I;zI;<*I;d:I;�NI;>hI;Z�I;�I;k�I;��I;�II;�H;�\E;�P@;��7;t*;�;�B�:q�:��9�'����غ_oE��G���ɻ��������.��o@�ܔK�      L�����0���=����N��Pp��D����bG�����(4�*�����n8��:U�:QG;�(;��7;`�@;��E;WQH;mI;��I;��I;��I;$}I;�^I;�FI;�3I;�$I;_I;�I;�	I;I;�I;��H;O�H;��H;�I;I;�	I;�I;aI;�$I;�3I;�FI;�^I;#}I;��I;��I;��I;mI;PQH;��E;a�@;��7;�(;OG;S�:��:��n80���'4�����bGໄ���D�Pp��N��>���2������      	��&�S5���������ϼˡ��X���iO�;���ɻ��p�pD� �o��g:`�:JG;t*;y9;��A;�uF;'�H;˔I;��I;��I;I�I;�pI;5TI;T>I;-I;�I;}I;�I;[I;�I;�I;�I;�I;�I;TI;�I;xI;�I;-I;R>I;5TI;�pI;E�I;��I;��I;˔I;%�H;�uF;��A;w9;r*;KG;`�:�g:0�o�pD⺎�p��ɻ;���iO�X��̡����ϼ������T5�%�      j��ѷ��$0v�q�a�#�G�?2+���՟�����/����5���!��Tf�Xج��g:M�:�; I-;g;;OC;SG;�I;϶I;!�I; �I;�I;cI;�II;�5I;r&I;�I;7I;�I;�I;MI;WI;NI;�I;�I;6I;�I;q&I;�5I;�II;cI;	�I;��I;�I;жI;�I;SG;�NC;"g;;I-;�;M�:�g:xج�Tf�"������5��/�����֟���?2+�$�G�r�a�$0v�ѷ��      ��ս��ѽ;�ƽ0����I�����P�a�D4�;M���ϼ��H�K�K��FG��Qf���o���:�B�:�Y;��1;\l>;�E;�/H;&qI;�I;��I;ژI;sI;�UI;�>I;�-I;b I;�I;�I;�
I;I;/I;I;�
I;�I;�I;^ I;�-I;�>I;�UI;sI;٘I;��I;��I;&qI;�/H;�E;Pl>;��1;�Y;�B�:��:0�o�Wf�FG��K��H�K�����ϼ;M�D4�Q�a�����I��0���;�ƽ��ѽ      �L+���'���F�������ս�@���%���;V�$��ܐ�����}MS�J�� ��bD�@�n8q�:�;o�$;_7;2�A;o�F;�H;i�I;d�I;��I;�I;YbI;�HI;5I;'&I;/I;AI;�I;�
I;
I;�
I;�I;>I;/I;"&I;5I;�HI;YbI;�I;��I;`�I;c�I;��H;o�F;2�A;�^7;r�$;�;q�:��n8fD� ��J��~MS�����ܐ�$���;V��%���@����ս����F�����'�      �T��f�����z��Yb�&�D��$�����ѽ�I��C�m�2+�������H�K��ﻋ�p�6���В�9;T�:�/;}�-;n�<;MzD;aH;�mI;��I;z�I;��I;�oI;�RI;�<I;,I;�I;I;/I;�I;�I;�I;/I;I;�I; ,I;�<I;�RI;�oI;��I;z�I;��I;�mI;`H;PzD;n�<;r�-;�/;5T�:В�94�����p���H�K�������2+�C�m��I����ѽ���$�&�D��Yb���z�f���      ?�׾��Ҿž�j��������z�S�H�)��dz�G$���/v�2+�ܐ�����5��ɻ/4�(�����:p��:Do!;P6;lA;��F;x�H;��I;��I;�I;M}I;�\I;`DI;	2I;r$I;�I;HI;�I;�I;�I;HI;�I;r$I;2I;]DI;�\I;M}I;�I;��I;��I;u�H;��F;lA;P6;8o!;p��:���: (��.4��ɻ��5���ݐ�2+��/v�G$��dz�)��S�H���z������j��ž��Ҿ      G(��$�d��P������~���`���Yb���'��U�F$��C�m�%����ϼ�/��:��������غ�8�9P��:�F;�G.;|=;NE;�\H;!�I;u�I;z�I;��I;gI;LI;�7I;)I;qI;rI;rI;'I;qI;rI;pI;)I;�7I;LI;gI;��I;|�I;u�I;�I;�\H;NE;|=;�G.;�F;P��:�8�9��غ����;���/����ϼ%��C�m�F$���U���'��Yb��`���~�����P��d���$�      <�}���w�#f���K�q,�}�
�;�׾ �����k���'�dz꽝I���;V�<M�����iO�fG�joE����N��:L� ;��$;��8;_�B;�G;0KI;�I;�I;D�I;	qI;�SI;�=I;�-I;"I;kI;I;�I;I;kI;"I;�-I;�=I;�SI;qI;B�I;�I;�I;0KI;��G;d�B;��8;��$;D� ;R��:���hoE�fG໨iO����;M��;V��I��dz���'���k� ���;�׾}�
�r,���K�#f���w�      ��p�������.蒿��w��F�c��ʰ� ����Yb�)����ѽ�%��D4�ן�X����� H���潺��9Xr�:��;�93;,Q@;�vF;�H;	�I;��I;��I;�zI;�ZI;CI;�1I;c%I;?I;�I;"I;�I;BI;b%I;�1I;CI;�ZI;�zI;��I;��I;�I;�H;�vF;,Q@;�93;��;Hr�:��9�潺�G�����X��ן�D4��%����ѽ)���Yb� ���ʰ�c���F���w�.蒿����p���      4��������㿊�ɿ���Ʌ����P�c��;�׾�`��S�H����@��Q�a���ˡ���D��ɻ� � ׭��W�:�;dI-;;|=;#CE;��H;�I;��I;v�I;��I;iaI;"HI;�5I;r(I;�I;�I;SI;�I;�I;p(I;�5I;"HI;haI;��I;v�I;��I;�I;��H;#CE;>|=;jI-;�;�W�:�֭�� ��ɻ�D�ˡ����Q�a��@����S�H��`��;�׾d����P�Ʌ�������ɿ�㿳���      ř$��x �"��9���޿o���Ʌ���F�}�
��~����z��$���ս���@2+���ϼPp�����F�]��*�&��:�;�8';��:;��C;�H;�}I;�I;t�I;ڋI;ngI;�LI;9I;9+I;!"I;�I;*I;�I;""I;7+I;9I;�LI;jgI;ڋI;t�I;#�I;�}I;H;��C;��:;�8';�;��:�*�F�]�����Pp���ϼ@2+������ս�$���z��~��}�
��F�Ʌ��o����޿9��"���x �      J�Q���K���;�ř$��;
��޿�����w�r,���澝���&�D������I��#�G�����N��������B�����9:d��:�n!;��7;¹B;J�G;�YI;+�I;Z�I;��I;�lI;sPI;<I;�-I;
$I;�I;�I;�I;$I;�-I;<I;uPI;�lI;��I;\�I;/�I;�YI;T�G;��B;��7;�n!;b��:��9:B����������N�����#�G��I������&�D��������r,���w�����޿�;
�ř$���;���K�      T����{���d��F�ř$�:����ɿ.蒿��K�P���j���Yb�F�0���r�a����>�����.��d��\�غ��9�Y�:2X;�25;&�A;Y!G;I7I;t�I;D�I;R�I;�pI;�SI;>I;y/I;�%I;" I;0I; I;�%I;v/I;�>I;�SI;�pI;V�I;D�I;w�I;M7I;f!G;$�A;�25;2X;�Y�:��9V�غ�d����.�>������r�a�0���F��Yb��j��P����K�.蒿��ɿ:��ř$��F���d��{�      ����#P�������d���;�#���㿲���#f�d��ž��z���;�ƽ$0v�S5�0����o@�����si�@au9IK�:];�73;(�@;��F;GI;��I;R�I;U�I;�sI;�UI;A@I;�0I;�&I;!I;0I;!I;�&I;�0I;B@I;�UI;�sI;Y�I;P�I;��I;MI;��F;%�@;�73;];EK�: au9qi������o@�0���S5�$0v�;�ƽ����z�žd��#f�������#����;���d����#P��      �,��a��#P���{���K��x �����p�����w��$���Ҿf���  (���ѽѷ��&�����K�@ɻ �����8���:~�;��1;�@;m�F;"I;߿I;�I;��I;�uI;&WI;hAI;�1I;�'I;�!I;�I;�!I;�'I;�1I;iAI;(WI;�uI;��I;�I;�I;&I;|�F;�@;��1;~�;~��:���8��Bɻ��K����&�ѷ����ѽ  (�f�����Ҿ�$���w�p��������x ���K��{�#P��a��      D(��q'���o��N�d��X1�~x�	Ŀ����3�v���x����4�j��Y+���'���ü7yY��kٻp&���p�V��:?;��0;��?;F;k I;�I;��I;,�I;j�I;MdI;�KI;�9I;n.I;�'I;�%I;�'I;k.I;�9I;�KI;OdI;h�I;0�I;��I;�I;m I;ЀF;��?;��0;;;N��: �p�p&��kٻ7yY���ü�'�Y+��j�ཽ�4��x��v���3����	Ŀ~x��X1�d�N��o��q'��      q'���X��f^�������]]���,�P9�6g��T�����/����o��f1��hܽ���-$�]l���|U�`�Իz!� �,���:�;�51;��?;8�F;C'I;c�I;�I;?�I;��I;�cI;@KI;z9I; .I;{'I;�%I;v'I;!.I;w9I;AKI;�cI;��I;A�I;�I;f�I;D'I;C�F;��?;�51;�;�: �,�u!�`�Ի�|U�]l���-$����hܽf1��o���ྚ�/�T���6g��P9���,��]]�����f^���X��      �o��f^���ē��4z�5K�h��R��&ﱿT�v��X#���Ѿń��&�o�нb̀�^��t���I�I��ǻ�4� #9��::�;$�2;��@;��F;�:I;��I;��I;��I;w�I;MbI;�II;�8I;[-I;�&I;�$I;�&I;[-I;�8I;JI;MbI;s�I;��I;��I;��I;�:I;��F;��@;!�2;:�;��:�"9�4��ǻJ�I�t���^��b̀�o�н�&�ń���Ѿ�X#�T�v�&ﱿR��h��5K��4z��ē�f^��      N������4z���V��X1��<�sؿ����RZ��	�(���IUo����]y��,l�X��R��?�7������ Ƴ9��:��;\�4;ntA;`2G;�XI;��I;M�I;�I;��I;�_I;�GI;#7I;�+I;�%I;�#I;�%I;�+I;!7I;�GI;�_I;�I;�I;N�I;��I;�XI;j2G;mtA;\�4;��;��:�ų9������?�7��R��X�,l�]y�����IUo�(����	��RZ����sؿ�<��X1���V��4z�����      d��]]�4K��X1�Zf��nQ��S���[58��A���נ���O���_什�Q����>ߓ��� ��V��x氺 �":��: ;�07;�B;3�G;�{I;��I;��I;��I;;|I;8\I;MEI;5I;5*I;1$I;)"I;-$I;5*I;5I;MEI;8\I;7|I;��I;��I;��I;�{I;<�G;�B;�07; ;��:�":r氺�V���� �>ߓ�����Q�_什����O��נ��A��[58�S���nQ���Zf��X1�4K��]]�      �X1���,�h���<��5g��e_���U�͂�֌Ⱦń�*�-�h��O ��%�2�	?ټ_�{� "��n��O���u:�P ;�&;0#:;A�C;�%H;�I;$�I;��I;�I;_vI;�WI;�AI;{2I;(I;D"I;^ I;@"I;(I;w2I;�AI;�WI;\vI;�I;��I;(�I;�I;�%H;C�C;+#:;�&;�P ;��u:��O��n� "�_�{�	?ټ%�2�O ��h��*�-�ń�֌Ⱦ͂��U�e_��5g��<�h����,�      ~x�O9�R��sؿnQ��e_��6�_��X#�p���f��9�S�{�����l�A�w���M���Ի��+��<T���:�e;�\,;�/=;�BE;V�H;}�I;��I;��I;��I;�oI;�RI;>I;]/I;}%I;�I;FI;�I;~%I;]/I;>I;�RI;�oI;��I;��I;��I;z�I;]�H;�BE;�/=;�\,;�e;��:`<T���+���Ի�M�w��A�l�����{�9�S��f��p���X#�6�_�e_��nQ��sؿR��O9�      	Ŀ6g��&ﱿ���S����U��X#�t��d���HUo��#��hܽ����n<����:����� ��᝻2�Ժ�t�9n��:�V;Ї2;� @;X�F;�I;��I;E�I;+�I;k�I; hI;MI;�9I;�+I;�"I;jI;�I;iI;�"I;�+I;�9I;MI;�gI;o�I;,�I;H�I;��I;�I;\�F;� @;ԇ2;�V;h��:�t�92�Ժ�᝻�� �:�������n<�����hܽ�#�HUo�d���s���X#��U�S������&ﱿ6g��      ���T���T�v��RZ�[58�͂�p��d���foy�]1�_O��[什�`�L�����myY��컏�T��1���u:
��:L#;98;�B;j�G;�lI;�I;�I;.�I;v�I;�_I;GI;�4I;%(I;�I;�I;I;�I;�I;%(I;�4I;GI;�_I;z�I;/�I;�I;�I;�lI;p�G;�B;98;O#;��:��u:�1���T���myY����L���`�[什_O��]1�foy�d���p��͂�[58��RZ�T�v�T���      �3���/��X#��	��A��֌Ⱦ�f��HUo�]1�ʰ��{n��мx��'��>ټ�@���k�ʼ����P�39�#�:4R;e-;�/=;�	E;`xH;��I;�I;q�I; �I;vI;aWI;�@I;�/I;#$I;;I;�I;6I;�I;<I;#$I;�/I;�@I;dWI;vI;�I;v�I;�I;��I;fxH;�	E;�/=;e-;4R;�#�:`�39��ȼ���k��@���>ټ�'�мx�{n��ʰ��]1�HUo��f��ՌȾ�A���	��X#���/�      v���ྃ�Ѿ(����נ�ń�9�S��#�_O��{n��Ì���2���𛼀�>���Ի��B��#�Tm:�G�:e ;��5;�FA;��F;�I;Q�I;T�I;��I;k�I;njI;�NI;:I;�*I;�I;�I;�I;KI;�I;�I;�I;�*I;:I;�NI;qjI;o�I;��I;U�I;N�I;�I;��F;�FA;��5;c ;�G�:`m:�#���B���Ի��>�������2�Ì�{n��_O���#�9�S�ń��נ�(�����Ѿ��      �x���o��
ń�IUo���O�*�-�{��hܽ[什мx���2�rb��TR��T|U�T2��4��갺�u�9��:D;��,;�h<;grD;S%H;ďI;j�I;��I;�I;�I;�^I;FI;V3I;�%I;�I;^I;hI;4I;hI;^I;�I;�%I;S3I;FI;�^I;�I;�I;��I;g�I;ˏI;T%H;krD;�h<;��,;D;��:�u�9갺4��T2��S|U�SR��rb����2�мx�[什�hܽ{�*�-���O�IUo�
ń��o��      ��4�f1��&������h�ང�������`��'���SR��B�]�|��V���X���Fo����:p�;,#;�6;VtA;W�F;�	I;u�I;��I;q�I;�I;�pI;�SI;�=I;�,I;w I;�I;�I;GI;9I;FI;�I;�I;y I;�,I;�=I;�SI;�pI;�I;q�I;��I;}�I;�	I;X�F;\tA;�6;8#;v�;���:�Do��X��V��{��B�]�SR����'��`��������h��������&�f1�      j�ྲྀhܽo�н]y��^什O ��l��n<�L���>ټ��T|U�~�������1�H�����u:gl�:�;i71;Y)>;W	E;JH;X�I;��I;��I;�I;׃I;YbI;�HI;&5I;c&I;gI;qI;<I;%I;
I;%I;:I;rI;gI;`&I;+5I;�HI;bbI;��I;�I;��I;��I;X�I;JH;^	E;Y)>;s71;�;al�:�u:H����1�����|��S|U��𛼿>ټL���n<�l�O ��^什]y��o�н�hܽ      X+����b̀�,l��Q�%�2�A��������@����>�T2��V���1�X�� $R:���:�;{\,;8;;�;C;�eG;Y9I;��I;1�I;��I;D�I;�qI;�TI;b>I;8-I;3 I;zI;rI;�
I;I;I;I;�
I;tI;|I;. I;;-I;d>I;�TI;�qI;D�I;��I;8�I;��I;[9I;�eG;�;C;B;;�\,;�;���: $R:X��1�V��R2��~�>��@��������A�$�2��Q�,l�b̀���      �'�-$�^��X����	?ټw��9���myY��k���Ի4���X��H���$R:���:�R;�);�8;��A;��F;7�H;-�I;��I;��I;��I;�I;�`I;�GI;�4I;�%I;JI;�I;�I;oI;I;EI;I;kI;�I;�I;GI;�%I;�4I;�GI;�`I;�I;��I;��I;��I;-�I;>�H;��F;��A;�8;�);�R;���:($R:H����X��4����Ի�k�lyY�9���w��?ټ���X�^��~-$�      ��ü\l��u����R��=ߓ�^�{��M��� ���ļ����B�갺 Fo��u:���:�R;7�';!17;Å@;��E;�lH;2�I;l�I;��I;�I;z�I;�lI;�QI;&<I;�+I;�I;�I;eI;�I;BI;/I;�I;+I;AI;�I;eI;�I;�I;�+I;*<I;�QI;�lI;t�I;�I;��I;k�I;6�I;�lH;�E;ą@;17;:�';�R;���:�u: Fo�갺~�B�ż���컈� ��M�^�{�>ߓ��R��v���Zl��      0yY��|U�I�I�<�7��� ��!���Ի�᝻��T� ��#��u�9���:al�:�;�);17;6 @;A]E;�$H;hkI;�I;Y�I;��I;*�I;�wI;�ZI;�CI;w1I;N#I;%I;�I;-	I;rI;9I;k�H;��H;h�H;6I;pI;-	I;�I;*I;R#I;z1I;�CI;�ZI;�wI;1�I;��I;U�I;�I;lkI;�$H;C]E;3 @;17;�);�;al�:���:�u�9|#�����T��᝻��Ի�!��� �>�7�H�I��|U�      �kٻf�Ի�ǻ����V���n���+�"�ԺԷ1���39xm:��:t�;�;�\,;�8;ą@;H]E;�
H;QVI;u�I;��I;��I;f�I;��I;�bI;cJI;&7I;�'I;�I;.I;�
I;8I;;I;i�H;��H;y�H;��H;f�H;9I;8I;�
I;2I;�I;�'I;*7I;bJI;�bI;�I;j�I;��I;��I;{�I;TVI;�
H;B]E;ǅ@;�8;�\,;�;t�;��:�m:��39�1�"�Ժ��+��n��V������ǻf�Ի      p&�{!��4���氺��O� <T��t�9��u:�#�:�G�:D;3#;r71;D;;��A;�E;�$H;SVI;�I;��I;�I;��I;��I;iI;*PI;<I;�+I;I;�I;�I;�I;�I;5�H;��H;��H;�H;��H;��H;2�H;�I;�I;�I;�I;I;�+I;<I;'PI;iI;�I;��I;�I;��I;�I;TVI;�$H;�E;��A;B;;l71;0#;D;�G�:�#�:��u:�t�9 <T�ܬO�t氺���4��!�      ��p� �,��!9�ų9�":��u:��:p��:��:8R;e ;��,;�6;Z)>;�;C;��F;�lH;rkI;y�I;��I;��I;�I;u�I;�mI;zTI;'@I;�/I;$"I;YI;�I;�I;�I;u�H;u�H;��H;W�H;��H;P�H;��H;t�H;t�H;�I;�I;�I;WI;'"I;�/I;&@I;�TI;�mI;p�I;�I;��I;��I;{�I;mkI;�lH;��F;�;C;V)>;�6;��,;g ;6R; ��:l��:��:��u:�":�ų9�!9 �,�      F��:��:�:#��:̸�:�P ;�e;�V;Q#;e-;��5;�h<;YtA;`	E;�eG;?�H;8�I;�I;��I;�I;�I;��I;pI;OWI;�BI;C2I;�$I;tI;pI;C	I;tI;��H;��H;�H;Z�H;5�H;��H;/�H;W�H;�H;��H;��H;xI;D	I;oI;wI;�$I;C2I;�BI;NWI;pI;��I;�I;�I;��I;�I;8�I;=�H;�eG;Z	E;YtA;�h<;��5;e-;S#;�V;�e;�P ;��:��:��:��:      P;�;6�;��;� ;�&;�\,;�2; 98;�/=;�FA;urD;[�F;JH;`9I;4�I;s�I;_�I;��I;��I;u�I;pI;MXI;�DI;�3I;`&I;"I;�I;�
I;pI;��H;��H;��H;��H;;�H;I�H;�H;C�H;8�H;��H;��H;��H;��H;oI;~
I;�I;I;`&I;�3I;�DI;HXI;
pI;v�I;��I;��I;W�I;r�I;3�I;_9I;JH;Y�F;srD;�FA;�/=;98;އ2;�\,;�&; ;��;0�;�;      ��0;�51;�2;W�4;�07;3#:;�/=;� @;�B;�	E;��F;U%H;�	I;[�I;��I;��I;��I;��I;g�I;��I;�mI;HWI;�DI;�4I;@'I;0I;I;}I;<I;0 I;-�H;��H;{�H;��H;d�H;��H;j�H;��H;a�H;��H;|�H;��H;1�H;. I;8I;I;�I;3I;D'I;�4I;�DI;KWI;�mI;��I;f�I;��I;��I;��I;��I;U�I;�	I;U%H;��F;�	E;�B;� @;�/=;##:;�07;T�4;�2;�51;      ��?;��?;��@;dtA;��B;K�C;�BE;[�F;p�G;dxH;�I;ϏI;y�I;��I;;�I;��I;�I;5�I;�I;iI;�TI;�BI;�3I;I'I;�I;I;I;�I;� I;��H;�H;m�H;b�H;��H;��H;/�H;��H;*�H;��H;��H;a�H;i�H;�H;��H;� I;�I;I;�I;�I;G'I;�3I;�BI;�TI;iI;�I;1�I;�I;��I;8�I;��I;{�I;ϏI;�I;dxH;l�G;X�F;�BE;?�C;�B;ctA;��@;��?;      F;F�F;��F;b2G;*�G;&H;]�H;�I;�lI;��I;X�I;t�I;��I;��I;��I;��I;}�I;�wI;�bI;)PI;*@I;=2I;_&I;3I;|I;;I; I;I;��H;G�H;z�H;W�H;~�H;(�H;^�H;��H;��H;��H;[�H;(�H;~�H;S�H;z�H;F�H;��H;I;I;>I;�I;1I;\&I;C2I;*@I;'PI;�bI;�wI;~�I;��I;��I;��I;��I;s�I;\�I;��I;�lI;�I;^�H;�%H;?�G;p2G;��F;F�F;      y I;N'I;�:I;�XI;�{I;�I;��I;�I;�I;�I;Z�I;��I;q�I;�I;F�I;	�I;�lI;�ZI;fJI;"<I;�/I;�$I;#I;I;I;I;I;��H;w�H;��H;M�H;U�H;��H;��H;�H;��H;q�H;��H;�H;��H;��H;R�H;P�H;��H;q�H;��H;I;!I;I; I;#I;�$I;�/I;<I;fJI;�ZI;�lI;�I;C�I;�I;p�I;��I;Z�I;�I;�I;�I;z�I;�I;�{I;�XI;�:I;8'I;      ��I;i�I;��I;��I;��I;%�I;��I;E�I;�I;z�I;��I;�I;�I;�I;�qI;�`I;�QI;�CI;&7I;�+I;("I;pI;�I;I;�I;� I;��H;m�H;��H;W�H;U�H;��H;��H;��H;��H;��H;q�H;��H;��H;��H;��H;��H;U�H;V�H;��H;m�H;��H; I;�I;}I;�I;sI;'"I;�+I;%7I;�CI;�QI;�`I;�qI;��I;�I;�I;��I;x�I;�I;D�I;��I;�I;��I;��I;��I;_�I;      ��I;�I;��I;]�I;��I;��I;��I;0�I;*�I;�I;q�I;�I;�pI;cbI;�TI;�GI;-<I;}1I;�'I;I;`I;iI;
I;8I;� I;��H;o�H;��H;Q�H;Q�H;��H;R�H;A�H;��H;��H;��H;��H;��H;��H;��H;C�H;N�H;��H;O�H;O�H;��H;j�H;��H;� I;4I;~
I;kI;\I;I;�'I;z1I;,<I;�GI;�TI;bbI;�pI;�I;u�I;�I;-�I;0�I;��I;��I;��I;`�I;��I;��I;      0�I;=�I;��I;�I;��I;�I;��I;u�I;z�I;vI;wjI;�^I;�SI;�HI;f>I;�4I;�+I;O#I;�I;�I;�I;?	I;lI;, I;��H;@�H;��H;Z�H;V�H;��H;,�H;�H;9�H;��H;�H;��H;��H;��H;�H;��H;8�H;�H;,�H;��H;R�H;Z�H;��H;B�H;��H;* I;pI;B	I;�I;�I;�I;N#I;�+I;�4I;d>I;�HI;�SI;�^I;wjI; vI;z�I;o�I;��I;�I;��I;�I;��I;:�I;      g�I;��I;z�I; �I;7|I;`vI;�oI;hI;�_I;kWI;�NI;FI;�=I;/5I;@-I;�%I;�I;,I;2I;�I;�I;vI;��H;-�H;�H;w�H;O�H;[�H;��H;/�H;�H;�H;V�H;��H;v�H;/�H;��H;-�H;u�H;��H;X�H;�H;�H;,�H;��H;X�H;L�H;x�H;�H;-�H;��H;xI;�I;�I;5I;*I;�I;�%I;@-I;.5I;�=I;FI;�NI;nWI;�_I;hI;�oI;[vI;A|I;�I;y�I;��I;      MdI;�cI;FbI;�_I;*\I;�WI;�RI;MI;
GI;�@I;:I;^3I;�,I;j&I;5 I;MI;�I;�I;�
I;�I;�I;��H;��H;��H;k�H;O�H;R�H;��H;V�H;�H;�H;O�H;��H;&�H;��H;��H;��H;��H;��H;(�H;��H;O�H;�H;�H;P�H;��H;Q�H;P�H;p�H;��H;��H;��H;�I;�I;�
I;�I;�I;QI;5 I;j&I;�,I;]3I;:I;�@I;	GI;MI;�RI;�WI;4\I;�_I;QbI;�cI;      �KI;OKI;JI;�GI;LEI;�AI;>I;�9I;�4I;�/I;�*I;�%I;| I;mI;~I;�I;jI;/	I;=I;�I;~�H;��H;��H;u�H;a�H;u�H;��H;��H;J�H;<�H;S�H;��H;�H;��H;K�H;�H;/�H;�H;H�H;��H;�H;��H;Q�H;6�H;F�H;��H;��H;w�H;e�H;w�H;��H;��H;z�H;�I;?I;/	I;lI;�I;�I;mI;} I;�%I;�*I;�/I;�4I;�9I;>I;�AI;PEI;�GI;JI;OKI;      �9I;{9I;�8I;7I;5I;n2I;^/I;�+I;)(I;.$I; I;�I;�I;yI;|I;�I;�I;rI;?I;7�H;|�H;�H;��H;��H;��H;�H;��H;��H;��H;��H;��H;&�H;��H;6�H;��H;��H;��H;��H;��H;9�H;��H;(�H;��H;��H;��H;��H;��H; �H;��H;��H;��H;�H;v�H;0�H;?I;vI;�I;�I;|I;{I;�I;�I;
 I;1$I;,(I;�+I;g/I;p2I;5I;7I;�8I;�9I;      b.I;=.I;c-I;�+I;A*I;(I;�%I;�"I;�I;LI;�I;pI;�I;GI;�
I;uI;LI;9I;k�H;��H;��H;U�H;5�H;U�H;��H;P�H;�H;��H;��H;�H;q�H;��H;K�H;��H;��H;��H;}�H;��H;��H;��H;K�H;��H;o�H;�H;��H;��H;�H;Q�H;��H;V�H;8�H;U�H;��H;��H;k�H;<I;MI;xI;�
I;JI;�I;oI;�I;OI;�I;�"I;�%I;(I;=*I;,I;a-I;?.I;      �'I;�'I;�&I;�%I;&$I;A"I;�I;tI;�I;�I;�I;tI;MI;*I;I;I;3I;j�H;��H;��H;^�H;.�H;B�H;��H;&�H;��H;��H;��H;��H;��H;-�H;��H; �H;��H;��H;c�H;q�H;f�H;��H;��H; �H;��H;,�H;��H;��H;��H;��H;��H;'�H;��H;F�H;/�H;X�H;��H;��H;o�H;6I;I;I;/I;MI;qI;�I;�I;�I;qI; I;A"I;*$I;�%I;�&I;�'I;      �%I;�%I;�$I;�#I;%"I;[ I;MI;�I;I;<I;WI;AI;CI;(
I;I;LI;�I; �H;~�H;	�H;��H;��H;�H;[�H;��H;��H;j�H;t�H;��H;��H;��H;��H;0�H;��H;}�H;m�H;v�H;o�H;z�H;��H;2�H;��H;��H;��H;��H;q�H;k�H;��H;��H;\�H;�H;��H;��H;�H;~�H;�H;�I;OI;I;+
I;DI;?I;]I;?I;I;�I;RI;[ I;""I;�#I;�$I;�%I;      �'I;�'I;�&I;�%I;'$I;D"I;�I;sI;�I;�I;�I;tI;MI;-I;I;I;3I;h�H;��H;��H;`�H;/�H;B�H;��H;&�H;��H;��H;��H;��H;��H;-�H;��H;!�H;��H;��H;c�H;q�H;f�H;��H;��H; �H;��H;,�H;��H;��H;��H;��H;��H;'�H;��H;F�H;.�H;X�H;��H;��H;o�H;5I;I;I;,I;MI;qI;�I;�I;�I;sI; I;D"I;*$I;�%I;�&I;�'I;      X.I;?.I;^-I;�+I;A*I;(I;�%I;�"I;�I;MI;�I;qI;�I;GI;�
I;uI;LI;;I;m�H;��H;��H;W�H;5�H;S�H;��H;O�H;�H;��H;��H;�H;o�H;��H;J�H;��H;��H;��H;}�H;��H;��H;��H;M�H;��H;o�H;�H;��H;��H;�H;S�H;��H;S�H;9�H;V�H;��H;��H;k�H;<I;OI;xI;�
I;JI;�I;pI;�I;MI;�I;�"I;�%I;(I;@*I;,I;a-I;C.I;      �9I;{9I;�8I;7I;5I;w2I;`/I;�+I;,(I;0$I; I;�I;�I;yI;}I;�I;�I;uI;?I;6�H;}�H;�H;��H;��H;��H; �H;��H;��H;��H;��H;��H;&�H;��H;6�H;��H;��H;��H;��H;��H;6�H;��H;&�H;��H;��H;��H;��H;��H;#�H;��H;��H;��H;�H;r�H;5�H;@I;vI;�I;�I;}I;|I;�I;�I; I;1$I;-(I;�+I;j/I;r2I; 5I;!7I;�8I;9I;      �KI;VKI;JI;�GI;JEI;�AI;>I;�9I;�4I;�/I;�*I;�%I;} I;kI;�I;�I;jI;1	I;?I;�I;�H;��H;��H;w�H;e�H;t�H;��H;��H;K�H;<�H;Q�H;��H;�H;��H;K�H;�H;/�H;�H;J�H;��H;�H;��H;Q�H;5�H;D�H;��H;��H;w�H;b�H;t�H;��H;��H;x�H;�I;?I;/	I;jI;�I;�I;mI;~ I;�%I;�*I;�/I;�4I;�9I;>I;�AI;NEI;HI;JI;RKI;      FdI;�cI;<bI;�_I;-\I;�WI;�RI;MI;	GI;�@I;:I;`3I;�,I;j&I;8 I;NI;�I;�I;�
I;�I;�I;��H;��H;��H;p�H;P�H;R�H;��H;Y�H;�H;	�H;O�H;��H;#�H;��H;��H;��H;��H;��H;&�H;��H;O�H;	�H;�H;P�H;��H;O�H;Q�H;m�H;��H;��H;��H;�I;�I;�
I;�I;�I;QI;8 I;j&I;�,I;`3I;:I;�@I;
GI;MI;�RI;�WI;,\I;�_I;AbI;�cI;      ^�I;��I;}�I;��I;<|I;bvI;�oI;hI;�_I;mWI;�NI;FI;�=I;25I;B-I;�%I;�I;*I;5I;�I;�I;yI;��H;-�H;�H;t�H;L�H;[�H;��H;/�H;	�H;�H;V�H;��H;x�H;-�H;��H;/�H;t�H;��H;V�H;�H;	�H;,�H;��H;U�H;L�H;z�H;�H;*�H;��H;yI;�I;�I;6I;*I;�I;�%I;@-I;25I;�=I;FI;�NI;mWI;�_I;hI;�oI;_vI;F|I;�I;��I;��I;      7�I;C�I;��I;�I;��I;�I;��I;w�I;}�I;!vI;rjI;�^I;�SI;�HI;j>I;�4I;�+I;P#I;�I;�I;�I;C	I;nI;, I;��H;=�H;��H;[�H;X�H;��H;,�H;�H;6�H;��H;�H;��H;��H;��H;�H;��H;9�H;�H;,�H;��H;Q�H;X�H;��H;C�H;��H;' I;rI;B	I;�I;�I;�I;N#I;�+I;�4I;g>I;�HI;�SI;�^I;tjI;!vI;x�I;s�I;��I;�I;��I;�I;��I;<�I;      ��I;�I;��I;V�I;��I;��I;��I;0�I;4�I;�I;q�I;�I;�pI;cbI;�TI;�GI;-<I;~1I;�'I;I;aI;lI;~
I;8I;� I;��H;m�H;��H;S�H;M�H;��H;R�H;A�H;��H;��H;��H;��H;��H;��H;��H;C�H;P�H;��H;N�H;M�H;��H;l�H;��H;� I;1I;�
I;lI;\I;I;�'I;z1I;,<I;�GI;�TI;cbI;�pI;�I;r�I;�I;.�I;2�I;��I;��I;��I;[�I;��I;��I;      	�I;`�I;��I;��I;��I;2�I;��I;K�I;�I;x�I;��I;�I;�I;�I;�qI;�`I;�QI;�CI;&7I;�+I;)"I;sI;�I;�I;�I;� I;��H;m�H;��H;S�H;V�H;��H;��H;��H;��H;��H;s�H;��H;��H;��H;��H;��H;V�H;T�H;��H;i�H;��H;� I;�I;{I;�I;qI;%"I;�+I;(7I;�CI;�QI;�`I;�qI;��I;�I;�I;��I;z�I;�I;D�I;��I;"�I;��I;��I;��I;`�I;      g I;U'I;�:I;�XI;�{I;"�I;~�I;�I;�I;�I;X�I;��I;m�I;�I;F�I;�I;�lI;�ZI;fJI;<I;�/I;�$I;!I;I;I;I;I;��H;w�H;��H;L�H;U�H;��H;��H;�H;��H;q�H;��H;�H;��H;��H;V�H;O�H;��H;s�H;��H;I;!I;I; I;%I;�$I;�/I; <I;iJI;�ZI;�lI;�I;F�I;�I;n�I;��I;Z�I;�I;�I;�I;��I;�I;�{I;�XI;�:I;@'I;      ��F;E�F;��F;^2G;.�G;&H;Y�H;�I;�lI;��I;X�I;u�I;��I;��I;��I;��I;{�I;�wI;�bI;)PI;.@I;@2I;]&I;5I;�I;8I;I;I;��H;C�H;z�H;W�H;|�H;(�H;^�H;��H;��H;��H;[�H;(�H;~�H;W�H;|�H;D�H;��H;I;I;>I;}I;3I;_&I;A2I;,@I;*PI;�bI;�wI;~�I;��I;��I;��I;��I;q�I;\�I;��I;�lI;�I;]�H;�%H;8�G;c2G;��F;8�F;      ��?;��?;��@;ctA;��B;N�C;�BE;[�F;r�G;fxH;�I;ԏI;{�I;��I;>�I;��I;�I;5�I;�I;iI;�TI;�BI;�3I;K'I;�I;{I;I;�I;� I;}�H;�H;n�H;`�H;��H;��H;*�H;��H;+�H;��H;��H;b�H;m�H;�H;��H;� I;�I;I;�I;�I;H'I;�3I;�BI;�TI;iI;�I;1�I;�I;��I;>�I;��I;|�I;ϏI;�I;gxH;n�G;W�F;�BE;@�C;�B;dtA;��@;��?;      ��0;~51;�2;\�4;�07;:#:;�/=;� @;�B;�	E;��F;W%H;�	I;X�I;��I;��I;��I;�I;g�I;��I;�mI;IWI;�DI;�4I;E'I;,I;�I;I;;I;- I;.�H;��H;|�H;��H;d�H;��H;k�H;��H;a�H;��H;�H;��H;3�H;1 I;9I;}I; I;3I;B'I;�4I;�DI;IWI;�mI;��I;j�I;��I;��I;��I;��I;W�I;�	I;T%H;��F;�	E;�B;� @;�/=;0#:;�07;u�4;�2;g51;      K;�;*�;��;� ;�&;�\,;އ2;#98;�/=;�FA;urD;X�F;JH;c9I;5�I;r�I;_�I;��I;��I;v�I;
pI;IXI;�DI;�3I;Y&I;I;�I;�
I;lI;��H;��H;��H;��H;;�H;I�H;�H;H�H;8�H;��H;��H;��H;��H;pI;
I;�I;"I;_&I;�3I;�DI;IXI;
pI;w�I;��I;��I;Y�I;s�I;4�I;c9I;JH;[�F;rrD;�FA;�/=; 98;ڇ2;�\,;�&;� ;��;(�;�;      J��:��: �:��:и�:�P ;�e;�V;S#;e-;��5;�h<;YtA;]	E;�eG;?�H;6�I;�I;��I;�I; �I;��I;pI;NWI;�BI;?2I;�$I;vI;pI;B	I;vI;��H;��H;�H;W�H;0�H;��H;3�H;V�H;�H;��H;��H;|I;F	I;nI;tI;�$I;D2I;�BI;RWI;pI;��I;�I;�I;��I;�I;6�I;>�H;�eG;^	E;ZtA;�h<;��5;e-;S#;�V;�e;�P ;���:���:��:��:      ��p� �,��"9�ų9��":��u:��:l��:
��:2R;f ;��,;�6;Z)>;�;C;��F;�lH;pkI;y�I;��I;��I;�I;s�I;�mI;�TI;#@I;�/I;%"I;YI;�I;�I;�I;t�H;t�H;��H;S�H;��H;T�H;��H;o�H;u�H;�I;�I;�I;WI;%"I;�/I;&@I;}TI;�mI;r�I;�I;��I;��I;{�I;mkI;�lH;��F;�;C;Z)>;�6;��,;i ;6R;��:p��:��:��u:(�": Ƴ9 #9 �,�      �o&�t!��4���氺�O� <T�u�9��u:�#�:�G�:D;3#;p71;F;;��A;�E;�$H;QVI;�I;��I;�I;��I; �I;iI;'PI;<I;�+I;I;�I;�I;�I;�I;5�H;��H;��H;�H;��H;��H;0�H;�I;�I;�I;�I;I;�+I;<I;)PI;iI;�I;��I;�I;��I;�I;TVI;�$H;�E;��A;D;;o71;1#;D;�G�:�#�:��u:�t�9 <T� �O�x氺����4�z!�      �kٻf�Ի�ǻ����V���n���+�"�Ժȷ1���39|m:��:v�;�;�\,;�8;Ņ@;F]E;�
H;SVI;{�I;��I;��I;g�I;�I;�bI;`JI;(7I;�'I;�I;/I;�
I;8I;;I;j�H;��H;y�H;��H;d�H;8I;8I;�
I;2I;�I;�'I;&7I;cJI;�bI; �I;m�I;��I;��I;y�I;TVI;�
H;C]E;Ņ@;�8;�\,;�;t�;��:xm:��39Է1�"�Ժ��+��n��V��
����ǻb�Ի      3yY��|U�J�I�<�7��� ��!���Ի�᝻��T� ��#��u�9���:al�:�;�);17;6 @;C]E;�$H;mkI;�I;\�I;��I;2�I;�wI;�ZI;�CI;}1I;L#I;'I;�I;-	I;sI;8I;k�H;��H;m�H;5I;pI;-	I;�I;)I;P#I;z1I;�CI;�ZI;�wI;*�I;��I;Y�I;�I;ikI;�$H;B]E;5 @;17;�);�;al�:���:�u�9�#� ���T��᝻��Ի�!��� �=�7�M�I��|U�      ��ü\l��u����R��=ߓ�^�{��M��� ���ż��~�B�갺 Fo��u:���:�R;:�';17;ą@;�E;�lH;8�I;p�I;��I;�I;x�I;�lI;�QI;,<I;�+I;�I;�I;eI;�I;EI;.I;�I;.I;AI;�I;bI;�I;�I;�+I;*<I;�QI;�lI;v�I;�I;��I;o�I;6�I;�lH;�E;ą@;17;9�';�R;���:�u: Fo�갺}�B�Ƽ���컈� ��M�]�{�>ߓ��R��v���[l��      �'�-$�^��W����?ټw��9���lyY��k���Ի2���X��X���,$R:���:�R;�);�8;��A;��F;>�H;3�I;��I;��I;��I;�I;�`I;�GI;�4I;�%I;JI;�I;�I;qI;I;CI;I;mI;�I;�I;FI;�%I;�4I;�GI;�`I;�I;��I;��I;��I;1�I;=�H;��F;��A;�8;�);�R;���: $R:H����X��5����Ի�k�myY�9���w��?ټ���X�^��-$�      X+����c̀�,l��Q�$�2�A��������@���>�T2��V���1�0��,$R:���:�;�\,;?;;�;C;�eG;c9I;��I;8�I;��I;B�I;�qI;�TI;b>I;;-I;1 I;zI;uI;�
I;I;I;I;�
I;rI;zI;- I;9-I;`>I;�TI;�qI;B�I;��I;3�I;��I;`9I;�eG;�;C;A;;}\,;�;���:$R:`��1�V��T2���>��@��������A�$�2��Q�,l�c̀���      j�ཱུhܽo�н]y��^什O ��l��n<�L���>ټ��R|U�|������~1�(����u:al�:�;o71;^)>;]	E;JH;Z�I;��I;��I;�I;ڃI;_bI;�HI;+5I;c&I;eI;rI;<I;"I;
I;&I;9I;qI;gI;_&I;(5I;�HI;]bI;ۃI;�I;��I;��I;\�I;JH;]	E;S)>;r71;�;_l�:�u:H����1�����}��T|U��𛼿>ټL���n<�l�O ��^什]y��o�н�hܽ      ��4�f1��&������h�ང�������`��'���SR��B�]�|��V���X�� Fo����:r�;3#;$�6;\tA;\�F;�	I;}�I;��I;n�I;�I;�pI;�SI;�=I;�,I;w I;�I;�I;FI;9I;FI;�I;�I;y I;�,I;�=I;�SI;�pI;�I;p�I;��I;v�I;�	I;\�F;YtA;�6;5#;p�;���:�Eo��X��V��|��B�]�SR����'��`��������h��������&�f1�      �x���o��
ń�IUo���O�*�-�{��hܽ[什мx���2�rb��SR��S|U�S2��3��
갺�u�9��:D;��,;�h<;orD;W%H;͏I;j�I;��I;�I;
�I;�^I;FI;U3I;�%I;�I;^I;hI;5I;iI;\I;�I;�%I;R3I;FI;�^I;�I;�I;��I;g�I;ƏI;U%H;qrD;�h<;��,;D;��:�u�9
갺4��T2��T|U�TR��rb����2�мx�[什�hܽ{�*�-���O�IUo�
ń��o��      v���ྃ�Ѿ(����נ�ń�9�S��#�_O��{n��Ì���2�����>���Ի��B��#�\m:�G�:j ;��5;�FA;��F;�I;R�I;S�I;��I;o�I;njI;�NI;:I;�*I;�I;�I;�I;LI;�I;�I;�I;�*I;:I;�NI;njI;o�I;��I;S�I;N�I;�I;��F;�FA;��5;_ ;�G�:Pm:�#���B���Ի��>�������2�Ì�{n��_O���#�9�S�ń��נ�(�����Ѿ��      �3���/��X#��	��A��ՌȾ�f��HUo�]1�ʰ��{n��мx��'��>ټ�@���k�ȼ����`�39�#�:8R;e-;�/=;�	E;dxH;��I;�I;q�I;�I;vI;eWI;�@I;�/I;&$I;;I;�I;6I;�I;<I;#$I;�/I;�@I;cWI;vI;�I;s�I;�I;��I;axH;�	E;�/=;e-;.R;�#�:P�39��Ǽ���k��@���>ټ�'�мx�{n��ʰ��]1�HUo��f��ՌȾ�A���	��X#���/�      ���T���T�v��RZ�[58�͂�p��d���foy�]1�_O��[什�`�L�����lyY��컐�T��1���u:��:P#;98;�B;p�G;�lI;�I;�I;2�I;w�I;�_I;GI;�4I;&(I;�I;�I;I;�I;�I;%(I;�4I;GI;�_I;s�I;/�I;�I;�I;�lI;n�G;�B;98;L#; ��:��u:��1���T���myY����L���`�[什_O��]1�foy�d���p��͂�[58��RZ�T�v�T���      	Ŀ6g��&ﱿ���S����U��X#�s��d���HUo��#��hܽ����n<����:����� ��᝻2�Ժ�t�9z��:�V;ԇ2;� @;\�F;�I;��I;D�I;,�I;i�I; hI;MI;�9I;�+I;�"I;iI;�I;iI;�"I;�+I;�9I;MI; hI;k�I;+�I;E�I;��I;�I;Y�F;� @;ׇ2;�V;f��:�t�92�Ժ�᝻�� �:�������n<�����hܽ�#�HUo�d���s���X#��U�S������&ﱿ6g��      ~x�O9�R��sؿnQ��e_��6�_��X#�p���f��9�S�{�����l�A�w���M���Ի��+�`<T���:�e;�\,;�/=;�BE;V�H;z�I;��I;��I;��I;�oI;�RI;>I;]/I;}%I;�I;FI;�I;%I;]/I;>I;�RI;�oI;��I;��I;��I;}�I;Z�H;�BE;0=;�\,;�e;��:0<T���+���Ի�M�w��A�l�����{�9�S��f��p���X#�6�_�e_��nQ��sؿR��O9�      �X1���,�h���<��5g��e_���U�͂�֌Ⱦń�*�-�h��O ��%�2�	?ټ^�{� "��n���O���u:�P ;�&;0#:;A�C;�%H;�I;$�I;��I;�I;`vI;�WI;�AI;z2I;(I;C"I;` I;C"I;(I;x2I;�AI;�WI;]vI;�I;��I;)�I;�I;�%H;A�C;3#:;�&;�P ;��u:�O��n� "�^�{�?ټ%�2�O ��h��*�-�ń�֌Ⱦ͂��U�e_��5g��<�h����,�      d��]]�4K��X1�Zf��nQ��S���[58��A���נ���O���_什�Q����>ߓ��� ��V��n氺$�":��: ;�07;�B;0�G;�{I;��I;��I;��I;;|I;5\I;LEI;5I;0*I;1$I;+"I;-$I;5*I;5I;MEI;7\I;8|I;��I;��I;��I;�{I;:�G;�B;�07;	 ;��:�":n氺�V���� �>ߓ�����Q�_什����O��נ��A��[58�S���nQ���Zf��X1�4K��]]�      N������4z���V��X1��<�sؿ����RZ��	�(���IUo����]y��,l�X��R��?�7�������0Ƴ9��:��;\�4;ntA;^2G;�XI;��I;N�I;�I;��I;�_I;�GI;"7I;�+I;�%I;�#I;�%I;�+I;7I;�GI;�_I;�I;�I;N�I;��I;�XI;i2G;mtA;^�4;��;��:�ų9������>�7��R��X�,l�]y�����IUo�(����	��RZ����sؿ�<��X1���V��4z�����      �o��f^���ē��4z�5K�h��R��&ﱿT�v��X#���Ѿń��&�o�нc̀�^��t���J�I��ǻ�4� #9��::�;$�2;��@;��F;�:I;��I;��I;��I;y�I;MbI;�II;�8I;X-I;�&I;�$I;�&I;\-I;�8I;�II;MbI;u�I;��I;��I;��I;�:I;��F;��@;$�2;:�;��:�"9�4��ǻI�I�t���^��b̀�o�н�&�ń���Ѿ�X#�T�v�&ﱿR��h��5K��4z��ē�f^��      q'���X��f^�������]]���,�P9�6g��T�����/����o��f1��hܽ���-$�]l���|U�`�Իw!� �,���:�;�51;��?;7�F;C'I;c�I;�I;?�I;��I;�cI;@KI;z9I;!.I;y'I;�%I;v'I;!.I;x9I;AKI;�cI;��I;A�I;�I;f�I;D'I;E�F;��?;�51;�;��: �,�t!�a�Ի�|U�]l���-$����hܽf1��o���ྚ�/�T���6g��P9���,��]]�����f^���X��   