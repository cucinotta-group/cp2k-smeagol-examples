H   �V�\V�/@                        �V�\V�/@                        �V�\V�/@H      H   H   H            m����������Ѣ��1�j��5���	��ȿ(8����7�E�꾃S���7�
3�}L���)���Ƽ��\�܉ݻ8+��Nɸ*�:sx;��0;�?;��F;$,I;��I;'�I;�I;f�I;iI;;OI;�<I;1I;�)I;�'I;�)I;1I;�<I;:OI;iI;f�I;�I;$�I;��I;$,I;��F;�?;��0;vx;*�:`Nɸ:+�܉ݻ��\���Ƽ�)�}L��
3��7��S��E�꾪�7�(8���ȿ��	��5�1�j�Ѣ����������      ��������B��^�����c�721�&X��ÿjڇ�t�3��s��7��}74�`�=ى���&��Mü�X���ػ;�%���J�;��:c;��0;��?;^�F;3I;'�I;��I;)�I;��I;�hI;�NI;r<I;�0I;�)I;�'I;�)I;�0I;r<I;�NI;�hI;��I;&�I;��I;'�I;3I;^�F;��?;��0;c;;��:��J�=�%���ػ�X� Nü��&�=ى�`�}74��7���s�t�3�jڇ��ÿ&X�721���c�^����B�����      �����B����F��y�P���#�N�������x|��'�ZD־�X��p�)�Խ�Ă�F<�2_��l-M���ʻ���-�8=��:�;NK2;^v@;��F;�FI;��I;Q�I;f�I;C�I;gI;MI;�;I;�/I;�(I;'I;�(I;�/I;�;I;~MI;gI;C�I;a�I;O�I;��I;�FI;��F;^v@;HK2;�;=��:�-�8
����ʻk-M�2_��F<��Ă�Խp�)��X��ZD־�'��x|����N�����#�y�P�F�����B��      Ѣ��^���F���/]��5�N���,ݿ-8��sm_��K��t��Y�s�$>����7�o��3��۩���:�LT��p����)�9g�:�<;�_4;UhA;a8G;�dI;G�I;w�I;��I;��I;ndI;]KI;�9I;�.I;�'I;�%I;�'I;�.I;�9I;\KI;ldI;��I;��I;t�I;G�I;�dI;^8G;ThA;�_4;�<;g�:*�9r���LT����:��۩��3�7�o����$>�Y�s��t���K�sm_�-8���,ݿN���5��/]�F��^���      1�j���c�y�P��5���t��J���jڇ�Iv<�*���r���_S��������	+T��� �$$���G#������0�� �:3��:��;f7;��B;ѮG;��I;Z�I;��I;�I;́I;�`I;�HI;�7I;�,I;H&I;B$I;H&I;�,I;�7I;�HI;�`I;́I;�I;��I;Z�I;��I;ϮG;��B;b7;��;3��:�:�0�������G#�$$���� �	+T���������_S�r��*���Iv<�jڇ�J���t�����5�y�P���c�      �5�721���#�N��u���ÿ�ҕ�Z������̾�X����0�3�/W����5�|zܼ/��H���s�hT\�h�n:a��:*�%;��9;��C;2/H;W�I;V�I;O�I;¦I;�{I;O\I;EI;5I;n*I;W$I;Y"I;W$I;n*I;5I;EI;P\I;�{I;��I;J�I;V�I;V�I;0/H;��C;��9;*�%;a��:p�n:lT\��s�H��0��|zܼ��5�/W��3佀�0��X����̾���Z��ҕ��ÿu��N����#�721�      ��	�&X�N����,ݿJ����ҕ��d��'�A��%���z�W����k���0�o��G��*���Q�z�ػ��0�p�~�j�:��;~,;�=;�BE;٬H;��I;��I;��I;*�I;�tI;WI;AI;�1I;�'I;�!I; I;�!I;�'I;�1I; AI;	WI;�tI;(�I;��I;��I;��I;٬H;�BE;�=;~,;��;p�:��~���0�y�ػ�Q��*���G�0�o�k������z�W�%���A�꾍'��d��ҕ�J����,ݿN���&X�      �ȿ�ÿ���-8��jڇ�Z��'�����n8��Y�s�-�&�W�/g??��V�琼GG#�>7���Sܺ��9�W�:��;hL2;�@;*�F;EI;��I;��I;��I;��I;�lI;QI;�<I;=.I;�$I;dI;�I;dI;�$I;=.I;�<I;QI;�lI;��I;��I;��I;��I;EI;*�F;�@;hL2;��;�W�:��9�Sܺ=7��GG#�琼�V�g??�/W�-�&�Y�s�n8�������'�Z�jڇ�-8������ÿ      (8��jڇ��x|�sm_�Iv<����A��n8��$6~�p74��l��{���5nc�2���^����\��9� Z���=��n:���:;#;�8;	�B;��G;�xI;��I;��I;ϵI;�I;ydI;�JI;�7I;[*I;z!I;�I;�I;�I;z!I;[*I;�7I;�JI;ydI;�I;̵I;��I;��I;�xI;��G;�B;�8;<#;���:�n:��=��Z��9���\��^��2��5nc�{����l��p74�$6~�n8��A�꾐��Iv<�sm_��x|�jڇ�      ��7�t�3��'��K�*�����̾%���Y�s�p74����!N��̇|�ށ)�4zܼ�Y��0 �h������pX9m��:f�;G-;T=;�E;K�H;��I;s�I;�I;�I;Z{I;�[I;�CI;�2I;V&I;I;lI;�I;lI;I;V&I;�2I;�CI;�[I;\{I;�I;�I;r�I;��I;H�H;�E;S=;G-;h�;k��:pX9����i��0 ��Y��4zܼށ)�̇|�!N�����p74�Y�s�%�����̾*����K��'�t�3�      E���s�ZD־�t��r���X��z�W�-�&��l��!N���Ă�h�5�����vQ����A�$�ػo�G�� /�<f:�b�:��;��5;�9A;��F;&+I;�I;�I;M�I;��I;ooI;�RI;�<I;\-I;�!I;�I;AI;�I;CI;�I;�!I;[-I;�<I;�RI;qoI;��I;N�I;�I;�I;#+I;��F;�9A;��5;��;�b�:<f:� /�p�G�$�ػ��A�vQ������h�5��Ă�!N���l��-�&�z�W��X��r���t��ZD־�s�      �S���7���X��Y�s��_S���0����W�{���̇|�h�5�d���ک�(�X�c �V�J3�� �9���:4�;F�,;�L<;�oD;P.H;�I;��I;��I;��I;��I;xcI;�II;6I;(I;�I;�I;�I;�I;�I;�I;�I;(I;6I;�II;xcI;��I;��I;��I;��I;�I;M.H;�oD;�L<;G�,;3�;���: �9L3��V�c �(�X��ک�e��h�5�̇|�{���Wལ����0��_S�Y�s��X���7��      �7�}74�p�)�$>����3�k���/5nc�ށ)������ک�fa��Q�1����M�`�ȸ���:2�;�#;��6;HhA;��F;�I;��I;��I;V�I;��I;�uI;�WI;�@I;I/I;�"I;XI;AI;�I;�I;�I;BI;ZI;�"I;K/I;�@I;�WI;�uI;��I;S�I;��I;�I;�I;��F;JhA;��6;�#;2�;���:��ȸ�M�1����Q�fa��ک�����ށ)�5nc�/k���3����$>�p�)�}74�      
3�`�Խ�������/W��0�o�f??�1��4zܼuQ��(�X��Q��6��n����Ϲ��n:n�:W>;��0;�>;uE;�SH;��I;�I;��I;��I;��I;gI;eLI;8I;�(I;MI;5I;�I;^I;�I;^I;�I;4I;NI;�(I;8I;gLI;gI;��I;��I;��I;�I;��I;�SH;uE;�>;��0;W>;n�:��n:��Ϲl���6���Q�(�X�uQ��3zܼ1��f??�0�o�.W���������Խ`�      }L��=ى��Ă�7�o�
+T���5��G��V��^���Y����A�c �1���n�����@�J:�l�:-f;d,;�:;P5C;UlG;,EI;A�I;��I;��I;ӝI;�vI;�XI;�AI;�/I;O"I;'I;�I;�I;<	I;�I;<	I;�I;�I;)I;T"I;�/I;�AI;�XI;�vI;ӝI;��I;��I;>�I;(EI;VlG;N5C;�:;e,;0f;�l�:@�J:���n��2���c ���A��Y���^���V��G���5�
+T�7�o��Ă�=ى�      �)���&�F<��3��� �|zܼ�*��琼��\�0 �"�ػV��M���ϹL�J:�j�:��;��(;�e8;�A;V�F;�H;f�I;��I;G�I;=�I;��I;�eI;�KI;Z7I;(I;%I;PI;I;�I;I;lI;I;�I;I;OI;)I;(I;\7I;�KI;�eI;��I;@�I;G�I;��I;a�I;�H;U�F;�A;�e8;��(;��;�j�:L�J:��Ϲ�M�V�"�ػ0 ���\�琼�*��{zܼ�� ��3�F<���&�      ��Ƽ�Mü2_���۩�$$��/���Q�FG#��9�g��n�G�J3����ȸ��n:�l�:��;]�';�7;�v@;j�E;XvH;:�I;��I;�I;��I;ƕI;�qI;�UI;r?I;".I;� I;RI;�I;#	I;�I;,I;dI;,I;�I;&	I;�I;TI;� I;".I;q?I;�UI;�qI;ɕI;��I;�I;��I;:�I;WvH;k�E;�v@;�7;_�';��;�l�:��n:��ȸJ3��o�G�g���9�FG#��Q�.��$$���۩�2_���Mü      ��\��X�k-M���:��G#�J��z�ػ>7���Z������ /���9���:n�:0f;��(;�7;�@;h]E;�-H;xwI;��I;	�I;�I; �I;}I;_I;#GI;04I;�%I;�I;I;�
I;~I;bI;k I;��H;k I;bI;~I;�
I; I;�I;�%I;-4I;%GI;_I;}I;�I;�I;�I;��I;uwI;�-H;h]E;�@;�7;��(;0f;n�:���:��9� /������Z�?7��z�ػI���G#���:�k-M��X�      ׉ݻ��ػ��ʻJT�������s���0��Sܺ��=��X9Df:���:2�;Z>;f,;�e8;�v@;f]E;sH;GbI;T�I;��I;��I;׭I;��I;BgI;CNI;:I;,*I;�I;�I;:I;uI;FI;��H;��H;��H;��H;��H;GI;wI;<I;�I;�I;)*I;:I;@NI;EgI;��I;ԭI;~�I;��I;Q�I;IbI;sH;i]E;�v@;�e8;h,;Z>;2�;���:Df:�X9��=��Sܺ��0��s�����JT����ʻ��ػ      8+�)�%�	��t����0��xT\���~���9�n:g��:�b�:1�;�#;��0;�:;ەA;f�E;�-H;CbI;��I;��I;��I;H�I;��I;nI;ATI;K?I;u.I;-!I;�I;?I;�I;�I;:�H;��H;I�H;��H;K�H;��H;:�H;�I;�I;@I;�I;'!I;w.I;H?I;BTI;nI;�I;F�I;��I;��I;��I;EbI;�-H;g�E;ەA;�:;��0;�#;1�;�b�:e��: �n:��9��~�lT\��0��x���	��3�%�      �Mɸ@�J��.�8�)�9�:t�n:p�:�W�:���:h�;��;C�,;��6;�>;N5C;R�F;XvH;wwI;T�I;��I;y�I;�I;��I;�rI;�XI;yCI;.2I;i$I;I;.I;#	I;�I;��H;l�H;�H;��H;��H;��H;�H;l�H;��H;�I;#	I;-I;I;l$I;,2I;yCI;�XI;�rI;��I;�I;w�I;��I;T�I;xwI;WvH;R�F;P5C;�>;��6;C�,;��;f�;���:�W�:n�:��n:��:�)�9`.�8��J�      8�:u��:[��:�f�:+��:q��:ĭ;��;A#;D-;��5;�L<;FhA;tE;UlG;�H;8�I;��I;��I;��I;�I;1�I;2uI;�[I;�FI;5I;�&I;rI;�I;�
I;�I;��H;O�H;��H;��H;��H;��H;��H;��H;��H;L�H;��H;�I;�
I;�I;tI;�&I;5I;�FI;�[I;1uI;3�I;�I;��I;��I;��I;5�I;�H;VlG;tE;GhA;�L<;��5;D-;A#;��;ĭ;w��:U��:�f�:[��:g��:      zx;c;�;�<;{�;)�%;�,;dL2;�8;T=;�9A;�oD;��F;�SH;+EI;a�I;��I;	�I;��I;H�I;��I;5uI;�\I;�GI;�6I;�(I; I;�I;�I;�I;� I;��H;��H;B�H;��H;	�H;��H;	�H;��H;D�H;��H;��H;� I;�I;�I;�I;I;�(I;�6I;�GI;�\I;5uI;��I;M�I;��I;�I;��I;`�I;+EI;�SH;��F;�oD;�9A;S=;�8;dL2;�,;*�%;��;�<;�;�b;      0;��0;VK2;�_4;d7;��9;�=;�@;�B;�E;��F;M.H;�I;��I;@�I;��I;�I;�I;֭I;��I;�rI;�[I;�GI;a7I;�)I;@I;�I;�I;pI;-I;�H;��H;:�H;/�H;�H;D�H;��H;D�H;�H;1�H;9�H;��H;�H;-I;pI;�I;�I;@I;�)I;^7I;�GI;�[I;�rI;��I;׭I;�I;�I;��I;@�I;��I;�I;M.H;��F;�E;	�B;�@;�=;��9;j7;�_4;RK2;��0;      ��?;��?;Jv@;YhA;��B;��C;�BE;#�F;��G;D�H;!+I;�I;{�I;�I;��I;E�I;��I; �I;��I;nI;�XI;�FI;�6I;�)I;�I;I;wI;�I;�I;x�H;��H;�H;��H;j�H;T�H;��H;p�H;��H;T�H;h�H;��H;�H;��H;x�H;�I;�I;wI;I;�I;�)I;�6I;�FI;�XI;nI;��I;�I;��I;D�I;��I;�I;y�I;�I;!+I;C�H;��G;%�F;�BE;��C;��B;XhA;Iv@;��?;      ��F;r�F;��F;d8G;ήG;+/H;֬H;;I;�xI;��I;�I;��I;��I;��I;��I;:�I;ƕI;}I;>gI;>TI;uCI; 5I;�(I;<I;I;�I;uI;�I;��H;!�H;;�H;��H;�H;��H;��H;7�H;.�H;7�H;��H;��H;
�H;��H;;�H;!�H;��H;�I;uI;�I;I;<I;�(I;5I;qCI;?TI;AgI;}I;ĕI;9�I;��I;��I;��I;��I;�I;��I;�xI;=I;֬H;)/H;ҮG;b8G;��F;g�F;      2,I;3I;�FI;�dI;��I;Y�I;��I;��I;��I;p�I;�I;��I;P�I;��I;ѝI;��I;�qI;_I;ANI;K?I;.2I;�&I;I;�I;sI;vI;.I;��H;R�H;@�H;��H;��H;x�H;a�H;m�H;��H;��H;��H;k�H;`�H;w�H;��H;��H;@�H;R�H;��H;,I;vI;wI;�I;I;�&I;+2I;K?I;ANI;_I;�qI;��I;ԝI;��I;S�I;��I;�I;o�I;��I;��I;��I;T�I;��I;�dI;�FI;�2I;      ��I;)�I;��I;C�I;U�I;R�I;��I;��I;��I;�I;P�I;��I;��I;��I;�vI;�eI;�UI;GI;:I;w.I;k$I;rI;�I;�I;�I;�I;��H;r�H;]�H;��H;��H;?�H;��H;��H;b�H;�H;��H;�H;b�H;��H;��H;@�H;��H;��H;]�H;t�H;��H;�I;�I;�I;�I;tI;h$I;w.I;:I;GI;�UI;�eI;�vI;��I;��I;��I;P�I;�I;��I;��I;��I;R�I;_�I;A�I;��I;5�I;      8�I;��I;H�I;z�I;��I;F�I;��I;��I;͵I;�I;��I;��I;�uI;gI;�XI;�KI;t?I;,4I;,*I;*!I;I;�I;�I;rI;�I;��H;Q�H;]�H;��H;��H; �H;��H;��H;��H;z�H;�H;��H;	�H;{�H;��H;��H;��H;!�H;��H;��H;]�H;T�H;��H;�I;rI;�I;�I;I;+!I;,*I;-4I;r?I;�KI;�XI;gI;�uI;��I;��I;�I;͵I;��I;��I;H�I;��I;z�I;H�I;v�I;      �I;,�I;g�I;��I;�I;ƦI;*�I;��I;"�I;^{I;uoI;�cI;�WI;kLI;�AI;Z7I;(.I;�%I;�I;�I;.I;�
I;�I;-I;s�H; �H;@�H;��H;��H;(�H;��H;��H;��H;��H;a�H;4�H;5�H;4�H;a�H;��H;��H;��H;��H;(�H;��H;��H;>�H;�H;v�H;.I;�I;�
I;-I;�I;�I;�%I;'.I;Z7I;�AI;kLI;�WI;�cI;toI;^{I;"�I;��I;+�I;ƦI;�I;��I;c�I;)�I;      e�I;��I;F�I;��I;ԁI;�{I;�tI;�lI;~dI;�[I;�RI;�II;�@I;8I;�/I;(I;� I;�I;�I;CI;(	I;�I;� I;�H;��H;=�H;��H;��H;�H;��H;|�H;x�H;��H;%�H;��H;��H;m�H;��H;��H;%�H;��H;z�H;|�H;��H; �H;��H;��H;;�H;��H;�H;� I;�I;&	I;CI;�I;�I;� I;(I;�/I;8I;�@I;�II;�RI;�[I;}dI;�lI;�tI;�{I;ҁI;��I;F�I;��I;      !iI;�hI;gI;rdI;�`I;L\I;WI;QI;�JI;�CI;�<I; 6I;I/I;�(I;U"I;*I;[I;I;?I;�I;�I;��H;��H;��H;�H;��H;��H;?�H;��H;��H;v�H;��H;�H;u�H;)�H;��H;��H;��H;)�H;u�H; �H;��H;w�H;��H;��H;?�H;��H;��H;�H;��H;��H;��H;�I;�I;?I;I;[I;*I;U"I;�(I;I/I; 6I;�<I;�CI;�JI;QI;WI;O\I;�`I;rdI;gI;�hI;      :OI;�NI;�MI;aKI;�HI;EI;AI;�<I;�7I;�2I;\-I;(I;�"I;NI;)I;PI;�I;�
I;xI;�I;��H;M�H;��H;=�H;��H;�H;x�H;��H;��H;��H;��H;�H;U�H;�H;��H;w�H;k�H;w�H;��H;�H;R�H;�H;��H;��H;��H;��H;v�H;�H;��H;>�H;��H;M�H;��H;�I;xI;�
I;�I;RI;'I;NI;�"I;(I;\-I;�2I;�7I;�<I;AI;EI;�HI;aKI;�MI;�NI;      �<I;w<I;x;I;�9I;�7I;�4I;�1I;@.I;]*I;U&I;�!I;�I;XI;8I;�I;I;+	I;{I;KI;@�H;s�H;��H;B�H;4�H;e�H;��H;[�H;��H;��H;��H;"�H;t�H;��H;��H;K�H;2�H;	�H;2�H;M�H;��H;��H;v�H;"�H;��H;��H;��H;]�H;��H;g�H;2�H;B�H;��H;r�H;@�H;KI;}I;*	I;I;�I;9I;XI;�I;�!I;U&I;_*I;C.I;�1I; 5I;�7I;�9I;y;I;p<I;      1I;�0I;�/I;�.I;�,I;f*I;�'I;�$I;~!I;I;�I;�I;DI;�I;�I;�I;�I;\I;��H;��H;�H;��H;��H;�H;N�H;��H;g�H;_�H;z�H;a�H;��H;*�H;��H;O�H;��H;��H;��H;��H;��H;O�H;��H;-�H;��H;d�H;}�H;_�H;g�H;��H;N�H;�H;��H;��H;�H;��H;��H;]I;�I;�I;�I;�I;DI;�I;�I;I;~!I;�$I;�'I;j*I;�,I;�.I;�/I;�0I;      �)I;�)I;�(I;�'I;U&I;P$I;�!I;jI;�I;lI;FI;I;�I;gI;@	I;!I;3I;d I;��H;O�H;��H;��H;�H;G�H;��H;4�H;��H;��H;�H;4�H;��H;��H;u�H;6�H;��H;��H;��H;��H;��H;3�H;t�H;��H;��H;4�H;�H;��H;��H;3�H;��H;G�H;�H;��H;��H;P�H;��H;e I;2I;"I;@	I;eI;�I;I;DI;mI;�I;jI;�!I;T$I;K&I;�'I;�(I;�)I;      �'I;�'I;
'I;�%I;F$I;U"I; I;�I;�I;�I;�I;�I;�I;�I;�I;oI;iI;��H; �H;��H;��H;��H;��H;��H;m�H;*�H;��H;��H;��H;:�H;q�H;��H;m�H;�H;��H;��H;��H;��H;��H;�H;j�H;��H;q�H;;�H;��H;��H;��H;,�H;m�H;��H;��H;��H;��H;��H; �H;��H;gI;oI;�I;�I;�I;�I;�I;�I;�I;�I; I;Y"I;;$I;�%I;'I;�'I;      �)I;�)I;�(I;�'I;U&I;P$I;�!I;jI;�I;jI;FI;I;�I;gI;@	I;"I;3I;d I;��H;O�H; �H;��H;�H;G�H;��H;4�H;��H;��H;�H;3�H;��H;��H;u�H;6�H;��H;��H;��H;��H;��H;3�H;t�H;��H;��H;5�H;�H;��H;��H;3�H;��H;G�H;�H;��H;��H;P�H;��H;e I;2I;!I;@	I;eI;�I;I;FI;lI;�I;jI;�!I;T$I;K&I;�'I;�(I;�)I;      1I;�0I;�/I;�.I;�,I;f*I;�'I;�$I;~!I;I;�I;�I;DI;�I;�I;�I;�I;\I;��H;��H;�H;��H;��H;�H;N�H;��H;h�H;_�H;{�H;a�H;��H;,�H;��H;O�H;��H;��H;��H;��H;��H;O�H;��H;/�H;��H;d�H;}�H;_�H;e�H;��H;N�H;�H;��H;��H;�H;��H;��H;]I;�I;�I;�I;�I;DI;�I;�I;I;~!I;�$I;�'I;j*I;�,I;�.I;�/I;�0I;      �<I;w<I;x;I;�9I;�7I;�4I;�1I;@.I;]*I;U&I;�!I;�I;XI;8I;�I;I;-	I;{I;KI;@�H;v�H;��H;B�H;4�H;g�H;��H;]�H;��H;��H;��H;"�H;t�H;��H;��H;M�H;2�H;	�H;2�H;K�H;��H;��H;v�H;"�H;��H;��H;��H;[�H;��H;e�H;2�H;B�H;��H;r�H;@�H;KI;}I;(	I;I;�I;9I;XI;�I;�!I;U&I;_*I;C.I;�1I;5I;�7I;�9I;y;I;p<I;      =OI;�NI;�MI;cKI;�HI;EI;AI;�<I;�7I;�2I;\-I;(I;�"I;NI;'I;RI;�I;�
I;xI;�I;��H;M�H;��H;>�H;��H;�H;x�H;��H;��H;��H;��H;�H;S�H;�H;��H;w�H;k�H;w�H;��H;�H;R�H;�H;��H;��H;��H;��H;v�H;�H;��H;=�H;��H;M�H;��H;�I;xI;�
I;�I;PI;)I;PI;�"I;(I;[-I;�2I;�7I;�<I;AI;EI;�HI;dKI;MI;�NI;      !iI;�hI;gI;rdI;�`I;L\I;WI;QI;�JI;�CI;�<I; 6I;I/I;�(I;U"I;*I;\I;I;?I;�I;�I;��H;��H;��H;�H;��H;��H;?�H;��H;��H;w�H;��H;�H;u�H;)�H;��H;��H;��H;)�H;u�H; �H;��H;v�H;��H;��H;?�H;��H;��H;�H;��H;��H;��H;�I;�I;?I;I;YI;*I;U"I;�(I;I/I; 6I;�<I;�CI;�JI;QI;WI;M\I;�`I;rdI;gI;�hI;      e�I;��I;F�I;��I;ԁI;�{I;�tI;�lI;~dI;�[I;�RI;�II;�@I;8I;�/I;(I;� I;�I;�I;AI;*	I;�I;� I;�H;��H;=�H;��H;��H;�H;��H;|�H;x�H;��H;%�H;��H;��H;m�H;��H;��H;%�H;��H;z�H;|�H;��H; �H;��H;��H;;�H;��H;�H;� I;�I;$	I;CI;�I;�I;� I;(I;�/I;8I;�@I;�II;�RI;�[I;}dI;�lI;�tI;�{I;ҁI;��I;F�I;��I;      �I;,�I;f�I;��I;
�I;��I;*�I;��I;#�I;]{I;uoI;�cI;�WI;lLI;�AI;Z7I;(.I;�%I;�I;�I;1I;�
I;�I;-I;v�H; �H;@�H;��H;��H;*�H;��H;��H;��H;��H;a�H;4�H;5�H;4�H;a�H;��H;��H;��H;��H;'�H;��H;��H;>�H;�H;s�H;.I;�I;�
I;-I;�I;�I;�%I;'.I;\7I;�AI;iLI;�WI;�cI;uoI;^{I;#�I;��I;+�I;æI;�I;��I;f�I;-�I;      2�I;~�I;O�I;x�I;��I;C�I;��I;��I;̵I;�I;��I;��I;�uI;gI;�XI;�KI;t?I;,4I;,*I;+!I;I;�I;�I;rI;�I;��H;Q�H;]�H;��H;��H;!�H;��H;��H;��H;z�H;�H;��H;	�H;z�H;��H;��H;��H; �H;��H;��H;]�H;R�H;��H;�I;rI;�I;�I;I;+!I;,*I;-4I;r?I;�KI;�XI;gI;�uI;��I;��I;�I;͵I;��I;��I;E�I;��I;u�I;N�I;~�I;      ��I;)�I;��I;A�I;U�I;R�I;��I;��I;��I;�I;Q�I;��I;��I;��I;�vI;�eI;�UI;GI;:I;w.I;n$I;tI;�I;�I;�I;�I;��H;t�H;]�H;��H;��H;@�H;��H;��H;`�H;�H;��H;�H;b�H;��H;��H;@�H;��H;��H;\�H;r�H;��H;�I;�I;�I;�I;rI;h$I;w.I;:I;GI;�UI;�eI;�vI;��I;��I;��I;N�I;�I;��I;��I;��I;O�I;a�I;C�I;��I;5�I;      ,,I;3I;�FI;�dI;��I;S�I;��I;��I;��I;p�I;�I;��I;S�I;��I;ӝI;��I;�qI;_I;ANI;L?I;02I;�&I; I;�I;wI;yI;.I;��H;T�H;A�H;��H;��H;w�H;`�H;k�H;��H;��H;��H;m�H;`�H;x�H;��H;��H;@�H;R�H;��H;,I;vI;sI;�I;I;�&I;)2I;K?I;ANI;_I;�qI;��I;ѝI;��I;P�I;��I;�I;p�I;��I;��I;��I;R�I;��I;�dI;�FI;�2I;      ��F;k�F;��F;d8G;ήG;,/H;֬H;=I;�xI;��I;�I;��I;��I;��I;��I;:�I;ƕI;}I;AgI;?TI;vCI;5I;�(I;=I;I;�I;uI;�I;��H;"�H;;�H;��H;�H;��H;��H;7�H;.�H;7�H;��H;��H;
�H;��H;;�H; �H;��H;�I;rI;�I;I;:I;�(I; 5I;oCI;>TI;>gI;}I;ĕI;:�I;��I;��I;��I;��I;�I;��I;�xI;=I;׬H;+/H;ҮG;d8G;��F;b�F;      ��?;��?;Jv@;XhA;��B;��C;�BE;#�F;��G;D�H;#+I;�I;y�I;�I;��I;E�I;��I; �I;��I;nI;�XI;�FI;�6I;�)I;�I;I;xI;�I;�I;x�H;��H;�H;��H;h�H;R�H;��H;p�H;��H;T�H;h�H;��H;�H;��H;w�H;�I;�I;vI;I;�I;�)I;�6I;�FI;�XI;nI;��I;�I;��I;E�I;��I;�I;{�I;�I;!+I;C�H;��G;%�F;�BE;��C;��B;YhA;Iv@;��?;      ȁ0;��0;XK2;�_4;^7;��9;�=;�@;�B;�E;��F;M.H;�I;��I;@�I;��I;�I;�I;׭I;��I;�rI;�[I;�GI;a7I;�)I;@I;�I;�I;qI;.I;�H;��H;9�H;/�H;�H;D�H;��H;D�H;�H;/�H;9�H;��H;�H;*I;mI;�I;�I;@I;�)I;`7I;�GI;�[I;�rI;��I;֭I;�I;�I;��I;>�I;��I;�I;M.H;��F;�E;�B;�@;�=;��9;n7;�_4;VK2;��0;      wx;c;�;�<;{�;,�%;�,;dL2;�8;T=;�9A;�oD;��F;�SH;+EI;a�I;��I;�I;��I;K�I;��I;5uI;�\I;�GI;�6I;�(I; I;�I;�I;�I;� I;��H;��H;D�H;��H;	�H;��H;	�H;��H;B�H;��H;��H;� I;�I;�I;�I;I;�(I;�6I;�GI;�\I;5uI;��I;K�I;��I;�I;��I;a�I;,EI;�SH;��F;�oD;�9A;R=;�8;fL2;�,;.�%;��;�<;�;c;      8�:s��:[��:�f�:+��:u��:ĭ;��;A#;D-;��5;�L<;GhA;tE;UlG;�H;7�I;��I;��I;��I;�I;3�I;5uI;�[I;�FI;5I;�&I;tI;�I;�
I;�I;��H;M�H;��H;��H;��H;��H;��H;��H;��H;M�H;��H;�I;�
I;�I;rI;�&I;5I;�FI;�[I;/uI;1�I;�I;��I;��I;��I;7�I;�H;VlG;tE;FhA;�L<;��5;D-;A#;��;ĭ;q��:W��:�f�:Y��:i��:      `Nɸ��J� /�8�)�9�:X�n:r�:�W�:���:f�;��;C�,;��6;�>;N5C;R�F;XvH;wwI;T�I;��I;z�I;�I;��I;�rI;�XI;yCI;,2I;l$I;I;.I;#	I;�I;��H;k�H;�H;��H;��H;��H;�H;l�H;��H;�I;#	I;,I;I;i$I;+2I;yCI;�XI;�rI;��I;�I;t�I;��I;T�I;xwI;WvH;R�F;M5C;�>;��6;A�,;��;d�;���:�W�:v�:|�n:�:�)�9 /�8��J�      :+�(�%���z����0��xT\���~���9�n:g��:�b�:1�;�#;��0;�:;ەA;g�E;�-H;EbI;��I;��I;��I;J�I;��I;nI;BTI;K?I;w.I;-!I;�I;@I;�I;�I;:�H;��H;K�H;��H;K�H;��H;:�H;�I;�I;?I;�I;'!I;u.I;H?I;ATI;nI;�I;F�I;��I;��I;��I;CbI;�-H;f�E;ەA;�:;��0;�#;0�;�b�:e��:�n:��9��~�hT\��0��x�����3�%�      ׉ݻ��ػ��ʻJT�������s���0��Sܺ��=��X9@f:���:2�;Z>;f,;�e8;�v@;i]E;sH;GbI;T�I;��I;��I;׭I;��I;DgI;CNI;:I;,*I;�I;�I;;I;wI;GI;��H;��H;��H;��H;��H;FI;tI;;I;�I;�I;)*I;:I;?NI;DgI;��I;ӭI;}�I;��I;P�I;IbI;sH;i]E;�v@;�e8;h,;Z>;2�;���:Df:�X9��=��Sܺ��0��s�����JT����ʻ��ػ      ��\��X�k-M���:��G#�J��z�ػ@7���Z������ /���9���:n�:/f;��(;�7;�@;h]E;�-H;wwI;��I;�I;�I;�I;}I;_I;%GI;04I;�%I;�I;I;�
I;~I;bI;k I;��H;k I;bI;~I;�
I; I;�I;�%I;-4I;#GI;_I;}I; �I;	�I;�I;��I;twI;�-H;h]E;�@;�7;��(;0f;n�:���:��9� /������Z�@7��z�ػI���G#���:�k-M��X�      ��Ƽ�Mü2_���۩�$$��/���Q�FG#��9�g��n�G�J3����ȸ��n:�l�:��;`�';�7;�v@;j�E;XvH;:�I;��I;�I;��I;ǕI;�qI;�UI;t?I;".I;� I;TI;�I;&	I;�I;,I;dI;,I;�I;$	I;�I;TI;� I;$.I;o?I;�UI;�qI;ǕI;��I;�I;��I;:�I;WvH;k�E;�v@;�7;]�';��;�l�:��n:��ȸJ3��l�G�h���9�FG#��Q�.��$$���۩�2_���Mü      �)���&�F<��3��� �|zܼ�*��琼��\�0 �#�ػX��M���ϹL�J:�j�:��;��(;�e8;�A;U�F;�H;d�I;��I;G�I;?�I;��I;�eI;�KI;Z7I;(I;&I;PI;I;�I;I;lI;I;�I;I;OI;&I;(I;Z7I;�KI;�eI;��I;?�I;H�I;��I;a�I;�H;T�F;�A;�e8;��(;��;�j�:L�J:��Ϲ�M�V�"�ػ0 ���\�琼�*��{zܼ�� ��3�F<���&�      }L��=ى��Ă�7�o�	+T���5��G��V��^���Y����A�c �1���n�����@�J:�l�:/f;e,;�:;N5C;VlG;.EI;C�I;��I;��I;֝I;�vI;�XI;�AI;�/I;Q"I;*I;�I;�I;<	I;�I;<	I;�I;�I;'I;Q"I;�/I;�AI;�XI;�vI;ѝI;��I;��I;=�I;(EI;UlG;N5C;�:;d,;2f;�l�:@�J:���n��1���c ���A��Y���^���V��G���5�
+T�7�o��Ă�=ى�      
3�`�Խ�������/W��0�o�f??�1��4zܼuQ��(�X��Q��6��l����Ϲ��n:n�:W>;��0;�>;uE;�SH;��I;�I;��I;��I;��I;gI;eLI;8I;�(I;PI;5I;�I;^I;�I;^I;�I;4I;LI;�(I;8I;eLI;gI;��I;��I;��I;�I;��I;�SH;uE;�>;��0;W>;n�:��n:��Ϲn���6���Q�(�X�uQ��3zܼ1��g??�0�o�.W���������Խ`�      �7�}74�p�)�$>����3�k���/5nc�ށ)������ک�fa��Q�1����M�`�ȸ���:2�;�#;��6;JhA;��F;�I;�I;��I;V�I;��I;�uI;�WI;�@I;I/I;�"I;ZI;BI;�I;�I;�I;AI;XI;�"I;H/I;�@I;�WI;�uI;��I;S�I;��I;��I;�I;��F;HhA;��6;�#;2�;���:��ȸ�M�1����Q�fa��ک�����ށ)�5nc�/k���3����$>�p�)�}74�      �S���7���X��Y�s��_S���0����W�{���̇|�h�5�e���ک�(�X�c �V�J3�� �9���:3�;C�,;�L<;�oD;P.H;�I;��I;��I;��I;��I;xcI;�II;6I;(I;�I;�I;�I;�I;�I;�I;�I;(I;6I;�II;xcI;��I;��I;��I;��I;�I;M.H;�oD;�L<;F�,;3�;���:( �9L3��X�c �(�X��ک�e��h�5�̇|�{���Wལ����0��_S�Y�s��X���7��      E���s�ZD־�t��r���X��z�W�-�&��l��!N���Ă�h�5�����vQ����A�$�ػo�G�� /�<f:�b�:��;��5;�9A;��F;#+I;�I;�I;N�I;��I;qoI;�RI;�<I;\-I;�!I;�I;CI;�I;AI;�I;�!I;[-I;�<I;�RI;ooI;��I;M�I;�I;�I;&+I;��F;�9A;��5;��;�b�:<f:� /�p�G�$�ػ��A�vQ������h�5��Ă�!N���l��-�&�z�W��X��r���t��ZD־�s�      ��7�t�3��'��K�*�����̾%���Y�s�p74����!N��̇|�ށ)�4zܼ�Y��0 �h������pX9m��:d�;G-;T=;�E;H�H;��I;s�I;�I;�I;Z{I;�[I;�CI;�2I;V&I;I;mI;�I;lI;I;V&I;�2I;�CI;�[I;Z{I;�I;�I;r�I;��I;K�H;�E;S=;G-;f�;k��:pX9����h��0 ��Y��4zܼށ)�̇|�!N�����p74�Y�s�%�����̾*����K��'�t�3�      (8��jڇ��x|�sm_�Iv<����A��n8��$6~�p74��l��{���5nc�2���^����\��9� Z���=��n:���:<#;�8;	�B;��G;�xI;��I;��I;еI;�I;ydI;�JI;�7I;[*I;z!I;�I;�I;�I;z!I;[*I;�7I;�JI;ydI;�I;̵I;��I;��I;�xI;��G;�B;�8;;#;���:�n:��=��Z��9���\��^��2��5nc�{����l��p74�$6~�n8��A�꾐��Iv<�sm_��x|�jڇ�      �ȿ�ÿ���-8��jڇ�Z��'�����n8��Y�s�-�&�W�/g??��V�琼FG#�>7���Sܺ��9�W�:��;hL2;�@;*�F;EI;��I;��I;��I;��I;�lI;QI;�<I;?.I;�$I;dI;�I;eI;�$I;?.I;�<I;QI;�lI;��I;��I;��I;��I;DI;*�F;�@;hL2;��;�W�:��9�Sܺ=7��GG#�琼�V�g??�/W�-�&�Y�s�n8�������'�Z�jڇ�-8������ÿ      ��	�&X�N����,ݿJ����ҕ��d��'�A��%���z�W����k���0�o��G��*���Q�z�ػ��0�p�~�j�:��;�,;�=;�BE;٬H;��I;��I;��I;*�I;�tI;WI; AI;�1I;�'I;�!I; I;�!I;�'I;�1I;AI;WI;�tI;(�I;��I;��I;��I;٬H;�BE;�=;},;��;n�:��~���0�y�ػ�Q��*���G�0�o�k������z�W�%���A�꾍'��d��ҕ�J����,ݿN���&X�      �5�721���#�N��t���ÿ�ҕ�Z������̾�X����0�3�/W����5�|zܼ/��H���s�lT\�`�n:a��:)�%;��9;��C;2/H;W�I;V�I;O�I;¦I;�{I;O\I;EI;5I;n*I;W$I;Y"I;X$I;m*I;5I;EI;P\I;�{I;��I;J�I;V�I;V�I;0/H;��C;��9;*�%;a��:p�n:lT\��s�G��0��|zܼ��5�/W��3佀�0��X����̾���Z��ҕ��ÿu��N����#�721�      1�j���c�y�P��5���t��J���jڇ�Iv<�*���r���_S��������	+T��� �$$���G#������0����:3��:��;f7;��B;ѮG;��I;Z�I;��I;�I;́I;�`I;�HI;�7I;�,I;J&I;B$I;H&I;�,I;�7I;�HI;�`I;́I;�I;��I;Z�I;��I;ϮG;��B;b7;��;3��:�:�0�������G#�$$���� �	+T���������_S�r��*���Iv<�jڇ�J���t�����5�y�P���c�      Ѣ��^���F���/]��5�N���,ݿ-8��sm_��K��t��Y�s�$>����7�o��3��۩���:�LT��p����)�9g�:�<;�_4;ThA;^8G;�dI;G�I;w�I;��I;��I;ndI;]KI;�9I;�.I;�'I;�%I;�'I;�.I;�9I;\KI;kdI;��I;��I;t�I;G�I;�dI;a8G;UhA;�_4;�<;g�:*�9r���LT����:��۩��3�7�o����$>�Y�s��t���K�sm_�-8���,ݿN���5��/]�F��^���      �����B����F��y�P���#�N�������x|��'�ZD־�X��p�)�Խ�Ă�F<�2_��k-M���ʻ
���-�8=��:�;NK2;^v@;��F;�FI;��I;Q�I;d�I;C�I;gI;MI;�;I;�/I;�(I;'I;�(I;�/I;�;I;~MI;gI;C�I;c�I;O�I;��I;�FI;��F;^v@;HK2;�;=��:�-�8	����ʻk-M�2_��F<��Ă�Խp�)��X��ZD־�'��x|����N�����#�y�P�F�����B��      ��������B��^�����c�721�&X��ÿjڇ�t�3��s��7��}74�`�=ى���&��Mü�X���ػ;�%���J�;��:c;��0;��?;^�F;3I;'�I;��I;)�I;��I;�hI;�NI;r<I;�0I;�)I;�'I;�)I;�0I;r<I;�NI;�hI;��I;&�I;��I;'�I;�2I;^�F;��?;��0;c;;��:��J�=�%���ػ�X� Nü��&�=ى�`�}74��7���s�t�3�jڇ��ÿ&X�721���c�^����B�����      F(��r'���o��O�d��X1�x�Ŀ����3�y���x����4�l��Y+���'���ü)yY��kٻ�o&� �p����:�;�0;Ͷ?;�F;� I;B�I;�I;e�I;��I;�dI;�KI;:I;�.I;�'I;&I;�'I;�.I;:I;�KI;�dI;��I;e�I;	�I;B�I;� I;�F;Ͷ?;�0;�;���:��p��o&��kٻ(yY���ü�'�Y+��l�ཾ�4��x��y���3����Ŀx��X1�d�O��o��r'��      r'���X��f^�������]]���,�Q9�8g��V�����/����o��h1��hܽ��~-$�Yl���|U�F�Ի1!� �,���:2;�51;�?;��F;q'I;��I;[�I;w�I;�I;dI;�KI;�9I;f.I;�'I;�%I;�'I;g.I;�9I;KI;dI;�I;t�I;X�I;��I;q'I;��F;�?;�51;6;��: �,�1!�D�Ի�|U�Yl��~-$����hܽh1��o���ྚ�/�V���8g��Q9���,��]]�����f^���X��      �o��f^���ē��4z�6K�i��T��'ﱿV�v��X#���Ѿń��&�p�нb̀�]��o���=�I�lǻz4��%9]�:��;O�2;Յ@;(�F;';I;4�I;A�I;ײI;��I;�bI;?JI;�8I;�-I;�&I;%I;�&I;�-I;�8I;?JI;�bI;��I;ԲI;?�I;4�I;&;I;(�F;Յ@;I�2;��;]�:&9{4�lǻ=�I�p���]��b̀�p�н�&�ń���Ѿ�X#�V�v�'ﱿT��i��6K��4z��ē�f^��      O������4z���V��X1��<�uؿ����RZ��	�*���KUo����^y��,l�W��R��2�7�𻱻r���ǳ9x��:)�;��4;�tA;�2G;�XI;��I;��I;E�I;8�I;`I;>HI;c7I;>,I;�%I;�#I;�%I;>,I;d7I;<HI;`I;8�I;D�I;��I;��I;�XI;�2G;�tA;��4;,�;x��:�ǳ9r��𻱻2�7��R��W�,l�^y�����KUo�*����	��RZ����uؿ�<��X1���V��4z�����      d��]]�6K��X1�[f��oQ��V���]58��A���נ���O���_什�Q����8ߓ��� �rV���尺��":S��:T ;&17;N�B;��G;*|I;(�I;��I;�I;}|I;|\I;�EI;\5I;z*I;o$I;m"I;o$I;x*I;\5I;�EI;|\I;}|I;�I;��I;(�I;+|I;��G;M�B; 17;V ;W��:��":�尺rV���� �8ߓ�����Q�_什����O��נ��A��]58�V���oQ���[f��X1�6K��]]�      �X1���,�i���<��8g��f_���U�΂�،Ⱦ
ń�+�-�j��P ��$�2�?ټQ�{��!�sn��O���u:0Q ;&;c#:;��C;H&H;T�I;g�I;�I;�I;�vI;XI;0BI;�2I;T(I;�"I;� I;�"I;V(I;�2I;0BI;XI;�vI;�I;�I;g�I;S�I;F&H;��C;_#:;&;0Q ;��u:�O�sn��!�Q�{�?ټ$�2�P ��i��+�-�
ń�،Ⱦ΂��U�f_��7g��<�i����,�      x�Q9�T��uؿoQ��f_��8�_��X#�t���f��;�S�{�����l�@�w���M�x�Ի��+�8T��:�e;],;40=;�BE;��H;��I;!�I;��I;��I;�oI;
SI;R>I;�/I;�%I;4 I;�I;4 I;�%I;�/I;T>I;SI;�oI;��I;��I;!�I;��I;��H;�BE;00=;],;�e; �:@8T���+�x�Ի�M�w��@�l�����{�;�S��f��t���X#�8�_�f_��oQ��uؿT��Q9�      Ŀ8g��'ﱿ���V����U��X#�v��f���JUo��#��hܽ����n<����5���}� ��᝻��Ժ w�9��:�V;�2;!@;��F;#I;<�I;��I;o�I;��I;ChI;QMI;�9I;0,I;�"I;�I;I;�I;�"I;0,I;�9I;SMI;ChI;��I;l�I;��I;:�I;#I;��F;!@;�2;�V;��:�v�9��Ժ�᝻}� �5�������n<�����hܽ�#�JUo�f���v���X#��U�V������'ﱿ8g��      ���V���V�v��RZ�]58�΂�t��f���hoy�_1�`O��[什�`�J�����ayY���Q�T���1���u:���:�#;_98;K�B;��G;:mI;R�I;A�I;q�I;��I;`I;DGI;55I;h(I;�I;�I;NI;�I;�I;h(I;55I;GGI;`I;��I;o�I;C�I;M�I;<mI;��G;F�B;]98;�#;���:��u:��1�O�T���`yY����K���`�[什`O��_1�hoy�f���t��΂�]58��RZ�V�v�V���      �3���/��X#��	��A��،Ⱦ�f��JUo�_1�̰��|n��Լx��'��>ټ�@���k��������P�39?$�:sR;Pe-;0=;
E;�xH;ͯI;S�I;��I;F�I;TvI;�WI;�@I;50I;g$I;�I;�I;zI;�I;�I;g$I;50I;�@I;�WI;UvI;C�I;��I;Q�I;ͯI;�xH;
E;0=;Pe-;sR;=$�:P�39��𺪼���k��@���>ټ�'�Լx�|n��̰��_1�JUo��f��،Ⱦ�A���	��X#���/�      y���྅�Ѿ*����נ�
ń�;�S��#�`O��|n��Ì���2����s�>�߾ԻF�B��#�Pm:fH�:� ;޼5;�FA;��F;�I;��I;��I;�I;��I;�jI;�NI;O:I;!+I;> I;I;�I;�I;�I;I;> I;+I;R:I;�NI;�jI;��I;�I;��I;��I;�I;��F;�FA;�5;� ;bH�:Pm:�#�H�B�޾Իs�>�������2�Ì�|n��`O���#�;�S�
ń��נ�*�����Ѿ��      �x���o��ń�KUo���O�+�-�{��hܽ[什Լx���2�nb��NR��G|U�<2�����鰺�w�9?�:YD;��,;i<;�rD;�%H;�I;��I;#�I;I�I;M�I;_I;KFI;�3I;�%I;I;�I;�I;yI;�I;�I;I;�%I;�3I;KFI;_I;L�I;I�I;"�I;��I;�I;�%H;�rD;i<; �,;XD;?�:�w�9�鰺��:2��G|U�NR��nb����2�Լx�[什�hܽ{�+�-���O�KUo�ń��o��      ��4�h1��&������i�ཅ�������`��'���NR��6�]�p���U��pX���6o�.��:��;t#;^�6;�tA;��F;�	I;��I;�I;��I;\�I; qI;�SI;�=I;	-I;� I;�I;I;�I;I;�I;I;�I;� I;-I;�=I;�SI; qI;\�I;��I;�I;��I;�	I;��F;�tA;^�6;r#;��;4��:�6o�lX���U��p��6�]�NR����'��`��������i��������&�h1�      k�ླྀhܽp�н^y��_什P ��l��n<�J���>ټ��F|U�p������E1�������u:�l�:L�;�71;�)>;�	E;SJH;��I;��I;��I;+�I;�I;�bI;�HI;j5I;�&I;�I;�I;I;cI;`
I;cI;I;�I;�I;�&I;m5I;�HI;�bI; �I;*�I;��I;��I;��I;QJH;�	E;�)>;�71;M�;�l�:��u:����D1�����p��G|U��𛼺>ټJ���n<�l�P ��_什^y��p�н�hܽ      X+����b̀�,l��Q�$�2�@��������@��s�>�<2���U��G1�x��%R:1��:(;�\,;�;;0<C;�eG;�9I;��I;y�I;�I;��I;�qI;�TI;�>I;z-I;n I;�I;�I;I;SI;RI;SI;I;�I;�I;r I;}-I;�>I;�TI;�qI;��I;�I;y�I;��I;�9I;�eG;0<C;�;;�\,;*;/��:%R:x��G1� V��<2��s�>��@��������@�$�2��Q�,l�b̀���      �'�~-$�]��W����?ټw��5���_yY��k�޾Ի��nX������%R:��:�R;�);"�8;͡A;ҀF;y�H;p�I;��I;��I;�I;L�I;aI;7HI;�4I;�%I;�I;I;�I;�I;TI;�I;TI;�I;�I;I;�I;�%I;�4I;3HI;aI;I�I;�I;��I;��I;l�I;z�H;πF;͡A;"�8;�);�R;��:%R:����pX����޾Ի�k�_yY�5���w��?ټ���W�\��~-$�      ��üWl��o����R��8ߓ�P�{��M�|� � �컨���D�B��鰺�6o���u:7��:�R;u�';Y17;�@;F�E;�lH;v�I;��I;��I;N�I;��I;mI;�QI;l<I;�+I;�I;I;�I;&I;�I;kI;�I;kI;�I;'I;�I;I;�I;�+I;k<I;�QI;	mI;��I;O�I;��I;��I;v�I;�lH;H�E;�@;[17;v�';�R;7��:��u:�6o��鰺F�B����� ��|� ��M�P�{�8ߓ��R��o���Xl��      *yY��|U�<�I�1�7��� ��!�x�Ի�᝻N�T����#��w�9,��:�l�:*;�);W17;p @;]E;%H;�kI;O�I;��I;;�I;r�I;�wI;�ZI;�CI;�1I;�#I;kI;�I;q	I;�I;wI;��H;A�H;��H;xI;�I;p	I;�I;kI;�#I;�1I;�CI;�ZI;�wI;r�I;8�I;��I;Q�I;�kI;	%H;]E;s @;V17;�);*;�l�:,��:�w�9�#����N�T��᝻x�Ի�!��� �1�7�<�I��|U�      �kٻD�Իfǻ𻱻tV��ln���+���Ժ�1�P�39Xm:E�:��;O�;�\,;"�8; �@;�]E;�
H;�VI;��I;1�I;5�I;��I;I�I;�bI;�JI;h7I;(I;�I;pI;I;{I;xI;��H;&�H;��H;&�H;��H;xI;zI;I;rI;�I;(I;h7I;�JI;�bI;I�I;��I;1�I;1�I;��I;�VI;�
H;�]E;��@;"�8;�\,;P�;��;E�:Xm:P�39ض1���Ժ��+�gn�rV��𻱻fǻD�Ի      �o&�!�x4�r���尺�O�`8T��v�9��u:9$�:fH�:WD;p#;�71;;;ǡA;B�E;%H;�VI;U�I;��I;W�I;ǭI;A�I;QiI;oPI;b<I;;,I;aI;I;I;�I;�I;q�H;�H;��H;H�H;��H;�H;q�H;�I;�I;I;I;^I;;,I;`<I;nPI;SiI;;�I;­I;Y�I;��I;W�I;�VI;%H;C�E;ǡA;;;�71;p#;UD;bH�:9$�:��u:�v�9`8T��O��尺r��w4�)!�      ��p� ,�`&9�ǳ9܍":��u: �:��:���:sR;� ;��,;\�6;�)>;/<C;̀F;�lH;�kI;��I;��I;��I;^�I;��I;�mI;�TI;l@I;�/I;f"I;�I;�I;I;�I;��H;��H;��H;��H;�H;��H;��H;��H;��H;�I;I;�I;�I;g"I;�/I;l@I;�TI;�mI;��I;^�I;��I;��I;��I;�kI;�lH;̀F;0<C;�)>;\�6;��,;� ;qR;���:��:�:��u:��":�ǳ9`&9 �,�      ɳ�:%�:}�:j��:O��::Q ;�e;�V;�#;Me-;�5;i<;�tA;�	E;�eG;v�H;u�I;O�I;0�I;W�I;\�I;:�I;JpI;�WI;4CI;�2I;�$I;�I;�I;�	I;�I;:�H;��H;B�H;��H;p�H;�H;p�H;��H;C�H;��H;:�H;�I;�	I;�I;�I;�$I;�2I;6CI;�WI;HpI;<�I;Z�I;Z�I;1�I;Q�I;s�I;u�H;�eG;�	E;�tA;i<;�5;Me-;�#;�V;�e;<Q ;u��:j��:}�:�:      �;6;��;%�;L ;&;],;�2;b98;0=;�FA;�rD;��F;SJH;�9I;l�I;��I;��I;5�I;ǭI;��I;MpI;�XI;�DI;-4I;�&I;gI;+I;�
I;�I;��H;��H;-�H;�H;x�H;��H;L�H;��H;x�H;�H;-�H;��H;��H;�I;�
I;+I;dI;�&I;04I;�DI;�XI;MpI;��I;ɭI;5�I;��I;��I;k�I;�9I;SJH;��F;�rD;�FA;0=;`98;�2;],;&;V ;#�;��;(;      #�0;�51;U�2;��4;%17;b#:;;0=;!@;L�B;
E;��F;�%H;�	I;��I;��I;��I;��I;;�I;��I;<�I;�mI;�WI;�DI;�4I;�'I;vI;DI;�I;xI;r I;p�H;!�H;��H;��H;��H;��H;��H;��H;��H;��H;��H;#�H;r�H;o I;xI;�I;DI;vI;�'I;�4I;�DI;�WI;�mI;>�I;��I;>�I;��I;��I;��I;��I;�	I;�%H;��F;
E;K�B;!@;:0=;c#:;*17;��4;U�2;�51;      ٶ?;�?;��@;�tA;M�B;��C;�BE;��F;��G;�xH;�I;�I;��I;��I;y�I;��I;R�I;q�I;M�I;UiI;�TI;6CI;34I;�'I;�I;�I;WI;"I;� I;��H;X�H;��H;��H;�H;�H;h�H;5�H;h�H;�H;�H;��H;��H;Z�H;��H;� I;$I;WI;�I;�I;�'I;04I;9CI;�TI;WiI;M�I;t�I;O�I;��I;y�I;��I;��I;�I;�I;�xH;��G;��F;�BE;��C;N�B;�tA;��@;�?;      &�F;��F;�F;�2G;��G;?&H;��H;I;;mI;ʯI;��I;��I;�I;��I;
�I;�I;��I;�wI;�bI;kPI;h@I;�2I;�&I;sI;�I;�I;cI;BI;�H;��H;��H;��H;��H;h�H;��H;�H;��H;�H;��H;i�H;��H;��H;��H;��H;�H;CI;cI;�I;�I;sI;�&I;�2I;d@I;lPI;�bI;�wI;��I;�I;�I;��I;�I;��I;��I;ǯI;:mI;I;��H;A&H;��G;�2G;�F;��F;      � I;r'I;$;I;�XI;(|I;W�I;��I;7�I;R�I;Q�I;��I;#�I;��I;*�I;��I;I�I;mI;�ZI;�JI;b<I;�/I;�$I;eI;GI;SI;dI;JI;.�H;��H;��H;��H;��H;�H;�H;W�H;��H;��H;��H;V�H;�H;�H;��H;��H;��H;��H;/�H;II;dI;XI;GI;dI;�$I;�/I;b<I;�JI;�ZI;mI;G�I;��I;*�I;��I;#�I;��I;N�I;S�I;8�I;��I;T�I;.|I;�XI;$;I;p'I;      4�I;��I;:�I;��I;#�I;d�I;�I;��I;D�I;��I;�I;K�I;Z�I; �I;�qI;aI;�QI;�CI;g7I;;,I;f"I;�I;,I;�I; I;DI;.�H;��H;��H;��H;��H;��H;��H;��H;�H;��H;��H;��H;�H;��H;��H;��H;��H;��H;��H;��H;.�H;DI;!I;�I;+I;�I;c"I;<,I;g7I;�CI;�QI;aI;�qI;�I;Y�I;K�I;�I;��I;D�I;��I;�I;d�I;-�I;��I;8�I;��I;      �I;X�I;9�I;��I;��I;	�I;��I;l�I;o�I;C�I;��I;M�I;qI;�bI;�TI;3HI;n<I;�1I;(I;`I;�I;�I;�
I;{I;� I;�H;��H;��H;��H;��H;��H;��H;��H;��H;*�H;��H;��H;��H;*�H;��H;��H;��H;��H;��H;��H;��H;��H;�H;� I;}I;�
I;�I;�I;aI;(I;�1I;l<I;3HI;�TI;�bI;qI;L�I;��I;B�I;q�I;l�I;��I;	�I;��I;��I;8�I;J�I;      l�I;{�I;ڲI;E�I;��I;"�I;��I;��I;��I;XvI;�jI;%_I;�SI;�HI;�>I;�4I;�+I;�#I;�I;I;�I;�	I;�I;r I;��H;��H;��H;��H;��H;��H;n�H;T�H;w�H;��H;Q�H;�H;��H;�H;Q�H;��H;v�H;U�H;n�H;��H;��H;��H;��H;��H;��H;r I;�I;�	I;�I;	I;�I;�#I;�+I;�4I;�>I;�HI;�SI;%_I;�jI;XvI;��I;��I;��I;"�I;��I;D�I;ԲI;x�I;      ��I;�I;��I;@�I;�|I;�vI;�oI;ChI;#`I;�WI;OI;RFI;�=I;p5I;~-I;�%I;�I;hI;tI;I;I;�I;��H;s�H;T�H;��H;��H;��H;��H;q�H;N�H;Q�H;��H;
�H;��H;r�H;4�H;r�H;��H;
�H;��H;S�H;N�H;o�H;��H;��H;��H;��H;W�H;s�H;��H;�I;I;I;tI;kI;�I;�%I;~-I;o5I;�=I;RFI;OI;�WI;"`I;EhI;�oI;�vI;�|I;?�I;��I;�I;      �dI;&dI;�bI;`I;z\I;XI;SI;TMI;GGI;�@I;R:I;�3I;-I;�&I;u I;�I;I;�I;#I;�I;�I;=�H; �H;&�H;��H;��H;��H;��H;��H;U�H;N�H;��H;��H;h�H;�H;��H;��H;��H;�H;h�H;��H;��H;P�H;V�H;��H;��H;��H;��H;��H;&�H;��H;>�H;�I;�I;#I;�I;I;�I;u I;�&I;-I;�3I;R:I;�@I;GGI;TMI;SI;XI;y\I;`I;�bI; dI;      �KI;�KI;AJI;CHI;�EI;,BI;N>I;�9I;85I;10I;!+I;�%I;� I;�I;�I;I;�I;i	I;}I;�I;��H;��H;+�H;��H;��H;��H;�H;��H;��H;{�H;��H;��H;S�H;��H;��H;]�H;m�H;]�H;��H;��H;P�H;��H;��H;}�H;��H;��H;�H;��H;��H;��H;*�H;��H;��H;�I;}I;j	I;�I;I;�I;�I;� I;�%I;!+I;30I;65I;�9I;N>I;/BI;�EI;CHI;CJI;�KI;      :I;�9I;�8I;j7I;a5I;�2I;�/I;4,I;i(I;e$I;A I;I;�I;�I;�I;�I;-I;�I;~I;w�H;��H;C�H;�H;��H;�H;e�H;��H;��H;��H;��H;�H;g�H;��H;{�H;7�H;�H;��H;�H;7�H;{�H;��H;j�H;�H;��H;��H;��H;��H;e�H;�H;��H;�H;C�H;��H;w�H;~I;�I;-I;�I;�I;�I;�I;I;? I;e$I;l(I;5,I;�/I;�2I;W5I;j7I;�8I;�9I;      �.I;t.I;�-I;C,I;�*I;M(I;�%I;�"I;�I;�I;I;�I;I;�I;I;�I;�I;sI;��H;�H;��H;��H;z�H;��H;�H;��H;S�H;�H;(�H;Q�H;��H;�H;��H;<�H;��H;��H;��H;��H;��H;<�H;��H;�H;��H;T�H;+�H;�H;R�H;��H;�H;��H;x�H;��H;��H;�H;��H;tI;�I;�I;I;�I;I;�I;I;�I;�I;�"I;�%I;P(I;�*I;C,I;�-I;k.I;      �'I;�'I;�&I;�%I;|$I;{"I;5 I;�I;�I;�I;�I;�I;�I;kI;WI;XI;rI;��H;*�H;��H;��H;p�H;��H;��H;e�H;�H;��H;��H;��H;�H;r�H;��H;[�H;�H;��H;��H;��H;��H;��H;�H;[�H;��H;r�H;�H;��H;��H;��H;�H;f�H;��H;��H;p�H;��H;��H;*�H;��H;qI;XI;WI;jI;�I;�I;�I;�I;�I;�I;5 I;"I;r$I;�%I; 'I;�'I;      &I;�%I;%I;�#I;q"I;� I;�I;I;PI;tI;�I;}I;I;f
I;SI;�I;�I;7�H;��H;M�H;�H;�H;M�H;��H;1�H;��H;��H;��H;��H;��H;9�H;��H;m�H;��H;��H;��H;��H;��H;��H;��H;k�H;��H;9�H;��H;��H;��H;��H;��H;1�H;��H;M�H;�H;�H;M�H;��H;9�H;�I;�I;SI;f
I;I;}I;�I;wI;QI;I;�I;� I;g"I;�#I;%I;�%I;      �'I;�'I;�&I;�%I;|$I;{"I;5 I;�I;�I;�I;�I;�I;�I;kI;WI;XI;rI;��H;*�H;��H;��H;p�H;��H;��H;f�H;�H;��H;��H;��H;�H;r�H;��H;[�H;�H;��H;��H;��H;��H;��H;�H;[�H;��H;r�H;�H;��H;��H;��H;�H;e�H;��H;��H;p�H;��H;��H;*�H;��H;qI;XI;WI;jI;�I;�I;�I;�I;�I;�I;5 I;"I;r$I;�%I;�&I;�'I;      �.I;t.I;�-I;C,I;�*I;M(I;�%I;�"I;�I;�I;I;�I;I;�I;I;�I;�I;sI;��H;�H;��H;��H;z�H;��H;�H;��H;S�H;�H;*�H;Q�H;��H;�H;��H;<�H;��H;��H;��H;��H;��H;<�H;��H;�H;��H;S�H;+�H;�H;R�H;��H;�H;��H;x�H;��H;��H;�H;��H;tI;�I;�I;I;�I;I;�I;I;�I;�I;�"I;�%I;Q(I;�*I;C,I;�-I;k.I;      :I;�9I;�8I;j7I;_5I;�2I;�/I;4,I;k(I;e$I;A I;I;�I;�I;�I;�I;.I;�I;~I;w�H;��H;C�H;�H;��H;�H;h�H;��H;��H;��H;��H;�H;g�H;��H;{�H;7�H;�H;��H;�H;7�H;{�H;��H;j�H;�H;��H;��H;��H;��H;e�H;�H;��H;�H;C�H;��H;w�H;~I;�I;,I;�I;�I;�I;�I;I;A I;e$I;l(I;5,I;�/I;�2I;U5I;j7I;�8I;�9I;      �KI;�KI;DJI;FHI;�EI;,BI;N>I;�9I;85I;10I;!+I;�%I;� I;�I;�I;I;�I;j	I;}I;�I;��H;��H;+�H;��H;��H;��H;�H;��H;��H;{�H;��H;��H;R�H;��H;��H;]�H;m�H;]�H;��H;��H;P�H;��H;��H;}�H;��H;��H;�H;��H;��H;��H;*�H;��H;��H;�I;}I;i	I;�I;I;�I;�I;� I;�%I;!+I;30I;85I;�9I;N>I;.BI;�EI;EHI;@JI;�KI;      �dI;&dI;�bI;
`I;|\I;XI;	SI;TMI;GGI;�@I;R:I;�3I;-I;�&I;u I;�I;I;�I;#I;�I;�I;>�H; �H;&�H;��H;��H;��H;��H;��H;U�H;P�H;��H;��H;h�H;�H;��H;��H;��H;�H;h�H;��H;��H;N�H;V�H;��H;��H;��H;��H;��H;&�H;��H;=�H;�I;�I;#I;�I;I;�I;u I;�&I;-I;�3I;R:I;�@I;HGI;TMI;SI;XI;y\I;
`I;�bI;"dI;      ��I;�I;��I;?�I;�|I;�vI;�oI;ChI;"`I;�WI;OI;RFI;�=I;p5I;~-I;�%I;�I;iI;tI;I;I;�I;��H;u�H;W�H;��H;��H;��H;��H;q�H;N�H;Q�H;��H;
�H;��H;r�H;4�H;r�H;��H;
�H;��H;Q�H;N�H;o�H;��H;��H;��H;��H;T�H;u�H;��H;�I;I;I;tI;iI;�I;�%I;~-I;q5I;�=I;RFI;OI;�WI;"`I;EhI;�oI;�vI;�|I;@�I;��I;�I;      e�I;y�I;ٲI;D�I;��I;�I;��I;��I;��I;VvI;�jI;%_I;�SI;�HI;�>I;�4I;�+I;�#I;�I;I;�I;�	I;�I;r I;��H;��H;��H;��H;��H;��H;n�H;T�H;w�H;��H;Q�H;�H;��H;�H;Q�H;��H;w�H;U�H;n�H;��H;��H;��H;��H;��H;��H;r I;�I;�	I;�I;I;�I;�#I;�+I;�4I;�>I;�HI;�SI;%_I;�jI;XvI;��I;��I;��I;!�I;��I;D�I;ٲI;|�I;      �I;T�I;=�I;��I;��I;�I;��I;l�I;q�I;B�I;��I;M�I;qI;�bI;�TI;3HI;n<I;�1I;(I;cI;�I;�I;�
I;{I;� I;�H;��H;��H;��H;��H;��H;��H;��H;��H;(�H;��H;��H;��H;*�H;��H;�H;��H;��H;��H;��H;��H;��H;�H;� I;}I;�
I;�I;�I;`I;(I;�1I;l<I;4HI;�TI;�bI;qI;M�I;��I;C�I;o�I;o�I;��I;	�I;��I;��I;=�I;T�I;      4�I;��I;:�I;��I;#�I;d�I;�I;��I;D�I;��I;�I;K�I;Y�I; �I;�qI;aI;�QI;�CI;g7I;<,I;i"I;�I;.I;�I;!I;DI;.�H;��H;��H;��H;��H;��H;��H;��H;�H;��H;��H;��H;�H;��H;��H;��H;��H;��H;��H;��H;.�H;DI; I;�I;)I;�I;c"I;<,I;g7I;�CI;�QI;aI;�qI;�I;Z�I;K�I;�I;��I;F�I;��I;�I;a�I;0�I;��I;8�I;��I;      � I;q'I;$;I;�XI;&|I;S�I;��I;7�I;R�I;P�I;��I;#�I;��I;*�I;��I;I�I;mI;�ZI;�JI;d<I;�/I;�$I;gI;GI;XI;gI;JI;/�H;��H;��H;��H;��H;�H;�H;V�H;��H;��H;��H;W�H;�H;�H;��H;��H;��H;��H;.�H;II;dI;SI;DI;cI;�$I;�/I;b<I;�JI;�ZI;mI;G�I;��I;*�I;��I;#�I;��I;P�I;R�I;8�I;��I;R�I;(|I;�XI;!;I;f'I;      *�F;��F;%�F;�2G;��G;B&H;��H;I;:mI;ʯI;��I;��I;�I;��I;
�I;�I;��I;�wI;�bI;lPI;i@I;�2I;�&I;uI;�I;�I;dI;CI;�H;��H;��H;��H;��H;i�H;��H;�H;��H;�H;��H;h�H;��H;��H;��H;��H;�H;BI;bI;�I;�I;pI;�&I;�2I;d@I;kPI;�bI;�wI;��I;�I;
�I;��I;�I;��I;��I;ȯI;8mI;I;��H;?&H;��G;�2G;"�F;��F;      ٶ?;�?;��@;�tA;M�B;��C;�BE;��F;��G;�xH;�I;�I;��I;��I;y�I;��I;Q�I;r�I;M�I;WiI;�TI;9CI;34I;�'I;�I;�I;XI;$I;� I;��H;Z�H;��H;��H;�H;�H;h�H;5�H;h�H;�H;�H;��H;��H;X�H;��H;� I;"I;VI;�I;�I;�'I;04I;6CI;�TI;WiI;M�I;t�I;O�I;��I;y�I;��I;��I;�I;�I;�xH;��G;��F;�BE;��C;K�B;�tA;��@;�?;      *�0;�51;Z�2;��4;17;g#:;50=;!@;M�B;
E;��F;�%H;�	I;��I;��I;��I;��I;=�I;��I;>�I;�mI;�WI;�DI;�4I;�'I;wI;EI;�I;{I;r I;r�H;!�H;��H;��H;��H;��H;��H;��H;��H;��H;��H;#�H;p�H;o I;wI;�I;BI;vI;�'I;�4I;�DI;�WI;�mI;>�I;��I;=�I;��I;��I;��I;��I;�	I;�%H;��F;
E;L�B;!@;50=;g#:;.17;��4;X�2;�51;      �;@;��;#�;N ;&;	],;�2;b98;0=;�FA;�rD;��F;SJH;�9I;l�I;��I;��I;5�I;ȭI;��I;MpI;�XI;�DI;04I;�&I;gI;+I;�
I;�I;��H;��H;.�H;�H;x�H;��H;L�H;��H;x�H;�H;+�H;��H;��H;�I;�
I;+I;dI;�&I;-4I;�DI;�XI;MpI;��I;ȭI;5�I;��I;��I;l�I;�9I;SJH;��F;�rD;�FA;0=;`98;�2;],;&;R ;%�;��;2;      ɳ�:%�:}�:j��:O��::Q ;�e;�V;�#;Me-;�5;i<;�tA;�	E;�eG;v�H;s�I;O�I;1�I;Y�I;]�I;<�I;LpI;�WI;6CI;�2I;�$I;�I;�I;�	I;�I;:�H;��H;C�H;��H;p�H;�H;p�H;��H;B�H;��H;:�H;�I;�	I;�I;�I;�$I;�2I;4CI;�WI;HpI;:�I;Z�I;Z�I;0�I;Q�I;s�I;v�H;�eG;�	E;�tA;i<;�5;Me-;�#;�V;�e;:Q ;{��:j��:}�:�:      ��p� �,��&9�ǳ9܍":��u:"�:��:���:qR;� ;��,;\�6;�)>;0<C;̀F;�lH;�kI;��I;��I;��I;^�I;��I;�mI;�TI;n@I;�/I;g"I;�I;�I;I;�I;��H;��H;��H;��H;�H;��H;��H;��H;��H;�I;I;�I;�I;f"I;�/I;l@I;�TI;�mI;��I;^�I;��I;��I;��I;�kI;�lH;̀F;/<C;�)>;\�6;��,;� ;pR;���:��:&�:��u:��":�ǳ9�&9 �,�      �o&�!�s4�v���尺�O�@8T��v�9��u:=$�:bH�:UD;p#;�71;;;ǡA;C�E;%H;�VI;U�I;��I;Y�I;ǭI;?�I;SiI;oPI;b<I;;,I;cI;I;I;�I;�I;q�H;�H;��H;H�H;��H;�H;q�H;�I;�I;I;I;\I;;,I;`<I;nPI;QiI;;�I;­I;W�I;��I;W�I;�VI;%H;B�E;ǡA;;;�71;p#;TD;bH�:7$�:��u: w�9@8T��O��尺r��x4�*!�      �kٻD�Իfǻ𻱻tV��mn���+���Ժ�1�P�39Xm:E�:��;P�;�\,;"�8; �@;�]E;�
H;�VI;��I;1�I;7�I;��I;I�I;�bI;�JI;h7I;(I;�I;rI;I;{I;xI;��H;&�H;��H;&�H;��H;xI;zI;I;pI;�I;(I;h7I;�JI;�bI;I�I;��I;0�I;1�I;��I;�VI;�
H;�]E;��@;"�8;�\,;O�;��;E�:Xm:P�39�1���Ժ��+�in�qV��𻱻fǻD�Ի      )yY��|U�<�I�2�7��� ��!�x�Ի�᝻N�T����#��w�9,��:�l�:(;�);Y17;r @;]E;%H;�kI;Q�I;��I;;�I;r�I;�wI;�ZI;�CI;�1I;�#I;kI;�I;q	I;�I;xI;��H;A�H;��H;wI;�I;p	I;�I;kI;�#I;�1I;�CI;�ZI;�wI;r�I;6�I;��I;O�I;�kI;	%H;]E;r @;W17;�);*;�l�:,��:�w�9�#����N�T��᝻x�Ի�!��� �1�7�<�I��|U�      ��üWl��o����R��8ߓ�P�{��M�|� � �컨���E�B��鰺�6o���u:7��:�R;x�';Y17;�@;F�E;�lH;v�I;��I;��I;O�I;��I;mI;�QI;n<I;�+I;�I;I;�I;'I;�I;kI;�I;kI;�I;'I;�I;I;�I;�+I;i<I;�QI;mI;��I;N�I;��I;��I;v�I;�lH;H�E;�@;[17;u�';�R;7��:��u:�6o��鰺D�B����� ��|� ��M�P�{�8ߓ��R��o���Xl��      �'�~-$�]��W� ���?ټw��5���_yY��k�޾Ի��pX������%R:��:�R;�);"�8;͡A;рF;z�H;o�I;��I;��I;�I;L�I;aI;7HI;�4I;�%I;�I;I;�I;�I;TI;�I;TI;�I;�I;I;�I;�%I;�4I;3HI;aI;G�I;�I;��I;��I;l�I;y�H;΀F;͡A;"�8;�);�R;��:%R:����nX����޾Ի�k�_yY�5���w��?ټ���W�]��~-$�      X+����b̀�,l��Q�$�2�@��������@��t�>�<2�� V��G1�x��%R:1��:(;�\,;�;;/<C;�eG;�9I;��I;y�I;�I;��I;�qI;�TI;�>I;}-I;o I;�I;�I;I;SI;RI;SI;I;�I;�I;p I;z-I;�>I;�TI;�qI;��I;�I;y�I;��I;�9I;�eG;/<C;�;;�\,;*;/��:%R:x��G1��U��<2��s�>��@��������@�#�2��Q�,l�b̀���      k�ླྀhܽp�н^y��_什P ��l��n<�J���>ټ��G|U�p������D1�������u:�l�:M�;�71;�)>;�	E;UJH;��I;��I;��I;-�I; �I;�bI;�HI;m5I;�&I;�I;�I;I;cI;`
I;cI;I;�I;�I;�&I;j5I;�HI;�bI;�I;*�I;��I;��I;��I;OJH;�	E;�)>;�71;L�;�l�:��u:����E1�����p��F|U��𛼺>ټJ���n<�l�P ��_什^y��p�н�hܽ      ��4�h1��&������i�ཅ�������`��'���NR��6�]�p���U��nX��@6o�0��:��;r#;\�6;�tA;��F;�	I;��I;�I;��I;\�I;!qI;�SI;�=I;	-I;� I;�I;I;�I;I;�I;I;�I;� I;	-I;�=I;�SI;qI;\�I;��I; �I;��I;�	I;��F;�tA;^�6;r#;��;4��:�6o�pX���U��p��6�]�NR����'��`��������i��������&�h1�      �x���o��ń�KUo���O�+�-�{��hܽ[什Լx���2�nb��NR��G|U�:2�����鰺�w�9?�:XD;��,;i<;�rD;�%H;�I;��I;#�I;I�I;M�I;_I;KFI;�3I;�%I;I;�I;�I;yI;�I;�I;I;�%I;�3I;KFI;_I;L�I;I�I; �I;��I;�I;�%H;�rD;i<;��,;XD;?�:�w�9�鰺��<2��G|U�NR��nb����2�Լx�[什�hܽ{�+�-���O�KUo�ń��o��      y���྅�Ѿ*����נ�
ń�;�S��#�`O��|n��Ì���2����s�>�޾ԻE�B��#�Pm:hH�:� ;�5;�FA;��F;�I;��I;��I;�I;��I;�jI;�NI;O:I;!+I;> I;I;�I;�I;�I;I;> I;+I;Q:I;�NI;�jI;��I;�I;��I;��I;�I;��F;�FA;޼5;� ;fH�:Pm:�#�H�B��Իs�>�������2�Ì�|n��`O���#�;�S�
ń��נ�*�����Ѿ��      �3���/��X#��	��A��،Ⱦ�f��JUo�_1�̰��|n��Լx��'��>ټ�@���k��������P�39?$�:qR;Pe-;0=;
E;�xH;ͯI;S�I;��I;F�I;TvI;�WI;�@I;50I;g$I;�I;�I;zI;�I;�I;g$I;40I;�@I;�WI;TvI;C�I;��I;Q�I;ίI;�xH;
E;0=;Pe-;sR;=$�:P�39��𺪼���k��@���>ټ�'�Լx�|n��̰��_1�JUo��f��،Ⱦ�A���	��X#���/�      ���V���V�v��RZ�]58�΂�t��f���hoy�_1�`O��[什�`�K�����`yY���Q�T���1���u:���:�#;_98;I�B;��G;;mI;R�I;C�I;r�I;��I;`I;EGI;65I;h(I;�I;�I;NI;�I;�I;h(I;45I;BGI;`I;��I;o�I;A�I;M�I;:mI;��G;F�B;]98;�#;���:��u:��1�O�T���ayY����J���`�[什`O��_1�hoy�f���t��΂�]58��RZ�V�v�V���      Ŀ8g��'ﱿ���V����U��X#�v��f���JUo��#��hܽ����n<����5���|� ��᝻��Ժ w�9��:�V;�2;!@;��F;#I;<�I;��I;o�I;��I;ChI;QMI;�9I;1,I;�"I;�I;I;�I;�"I;1,I;�9I;QMI;ChI;��I;l�I;��I;:�I;"I;��F;!@;�2;�V;��:�v�9��Ժ�᝻}� �5�������n<�����hܽ�#�JUo�f���v���X#��U�V������'ﱿ8g��      x�Q9�T��uؿoQ��f_��8�_��X#�t���f��;�S�{�����l�@�w���M�x�Ի��+�08T��:�e;],;40=;�BE;��H;��I;!�I;��I;��I;�oI;
SI;U>I;�/I;�%I;4 I;�I;4 I;�%I;�/I;Q>I;
SI;�oI;�I;��I;!�I;��I;��H;�BE;10=;],;�e; �:@8T���+�v�Ի�M�w��@�l�����{�;�S��f��t���X#�8�_�f_��oQ��uؿT��Q9�      �X1���,�i���<��7g��f_���U�΂�،Ⱦ
ń�+�-�i��P ��$�2�?ټQ�{��!�sn��O���u:0Q ;&;c#:;��C;H&H;T�I;g�I;�I;�I;�vI;XI;2BI;�2I;V(I;�"I;� I;�"I;T(I;�2I;/BI;XI;�vI;�I;�I;g�I;S�I;F&H;��C;_#:;&;0Q ;��u:�O�sn��!�Q�{�?ټ$�2�P ��j��+�-�
ń�،Ⱦ΂��U�f_��7g��<�i����,�      d��]]�6K��X1�[f��oQ��V���]58��A���נ���O���_什�Q����8ߓ��� �rV���尺�":W��:T ;%17;M�B;��G;*|I;(�I;��I;�I;}|I;z\I;�EI;\5I;z*I;o$I;m"I;o$I;x*I;\5I;�EI;|\I;}|I;�I;��I;(�I;+|I;��G;N�B;"17;V ;S��:��":�尺rV���� �8ߓ�����Q�_什����O��נ��A��]58�V���oQ���[f��X1�6K��]]�      O������4z���V��X1��<�uؿ����RZ��	�*���KUo����^y��,l�W��R��2�7�𻱻r��ǳ9x��:)�;��4;�tA;�2G;�XI;��I;��I;G�I;8�I;`I;>HI;d7I;>,I;�%I;�#I;�%I;>,I;c7I;<HI;`I;8�I;D�I;��I;��I;�XI;�2G;�tA;��4;,�;x��:�ǳ9r��𻱻2�7��R��W�,l�^y�����KUo�*����	��RZ����uؿ�<��X1���V��4z�����      �o��f^���ē��4z�6K�i��T��'ﱿV�v��X#���Ѿń��&�p�нb̀�]��o���=�I�lǻ{4��%9]�:��;O�2;Յ@;(�F;&;I;4�I;A�I;ײI;��I;�bI;?JI;�8I;�-I;�&I;%I;�&I;�-I;�8I;?JI;�bI;��I;ԲI;?�I;4�I;&;I;(�F;Յ@;I�2;��;]�:�%9{4�lǻ<�I�p���]��b̀�p�н�&�ń���Ѿ�X#�V�v�'ﱿT��i��6K��4z��ē�f^��      r'���X��f^�������]]���,�Q9�8g��V�����/����o��h1��hܽ��~-$�Yl���|U�D�Ի1!� �,���:2;�51;�?;��F;q'I;��I;[�I;w�I;�I;dI;�KI;�9I;f.I;�'I;�%I;�'I;g.I;�9I;KI;dI;�I;t�I;X�I;��I;p'I;��F;�?;�51;6;��: �,�1!�F�Ի�|U�Yl��~-$����hܽh1��o���ྚ�/�V���8g��Q9���,��]]�����f^���X��      ����,������U���L�Q�Ǚ$�5�����=�}�I(�C�׾�T���L+���սj��	��L���iO���ͻ>���-m8�o�:��;|�1;��?;/vF;� I;��I;��I;��I;�vI;�WI;BI;22I;(I;"I;. I;"I;(I;22I;BI;�WI;�vI;��I;��I;��I;� I;/vF;��?;z�1;��;�o�: .m8?����ͻ�iO�L��	��j����ս�L+��T��C�׾I(�=�}���5���Ǚ$�L�Q�U��������,��      �,��b��$P���{���K��x �����r�����w��$���Ҿh��� (���ѽѷ��%����ՔK�(ɻݟ����8��:��;��1;7@;ʊF;NI;"�I;X�I;�I;�uI;nWI;�AI;�1I;�'I;�!I; I;�!I;�'I;�1I;�AI;oWI;�uI;��I;U�I;"�I;NI;ɊF;7@;��1;��;��:���8ݟ�(ɻԔK����%�ѷ����ѽ (�h�����Ҿ�$���w�r��������x ���K��{�$P��b��      ����$P�������d���;�$���㿴���#f�f�� ž��z���=�ƽ$0v�R5�*����o@�f���-i�0du9�K�:j];83;h�@;?�F;xI;��I;��I;��I;tI;VI;�@I;#1I;('I;L!I;qI;L!I;&'I;#1I;�@I;VI;tI;��I;��I;��I;xI;?�F;h�@;83;m];�K�:0du9.i�g����o@�*���R5�$0v�=�ƽ����z� žf��#f�������$����;���d����$P��      U����{���d��F�Ǚ$�<����ɿ0蒿��K�R���j�� Zb�G�2���q�a����9�����.��d����غ���9+Z�:�X;�25;j�A;�!G;{7I;��I;��I;��I;�pI;�SI;�>I;�/I;�%I;a I;qI;a I;�%I;�/I;�>I;�SI;�pI;��I;��I;��I;{7I;�!G;h�A;�25;�X;+Z�:���9��غ�d����.�:������q�a�2���G� Zb��j��R����K�0蒿��ɿ<��Ǚ$��F���d��{�      L�Q���K���;�Ǚ$��;
��޿�����w�r,���澞���(�D������I��"�G����N��v���������x�9:ڨ�:o!;��7;�B;��G;(ZI;l�I;��I;��I;�lI;�PI;W<I;�-I;T$I; I;I; I;S$I;�-I;V<I;�PI;�lI;��I;��I;l�I;*ZI;��G;�B;��7;o!;ڨ�:��9:�������v���N�����"�G��I������(�D��������r,���w�����޿�;
�Ǚ$���;���K�      Ǚ$��x �$��<���޿q���˅���F�~�
��~����z��$���ս���>2+���ϼPp�q����]��*����:Y�;*9';ތ:;@�C;QH;�}I;b�I;��I;�I;�gI;�LI;\9I;x+I;d"I;6I;jI;5I;d"I;y+I;\9I;�LI;�gI;�I;��I;b�I;�}I;PH;?�C;ڌ:;)9';W�;���:�*��]�p���Pp���ϼ>2+������ս�$���z��~��~�
��F�˅��q����޿<��$���x �      5��������㿌�ɿ���˅����P�e��>�׾�`��U�H����@��Q�a���ơ���D��ɻ� ��έ�SX�:�;�I-;o|=;lCE;�H;K�I;!�I;��I;��I;�aI;eHI;�5I;�(I; I;I;�I;I; I;�(I;�5I;gHI;�aI;�I;��I;!�I;G�I;�H;iCE;j|=;�I-;�;SX�: ϭ�� ��ɻ�D�ơ����Q�a��@����U�H��`��>�׾e����P�˅�������ɿ�㿵���      ��r�������/蒿��w��F�e��̰�!����Yb�*����ѽ�%��D4�ԟ�X��y���G��:潺0��9�r�:1 ;+:3;bQ@;�vF;_�H;H�I;��I;ΤI;�zI;
[I;SCI;�1I;�%I;�I;�I;dI;�I;�I;�%I;�1I;UCI;
[I;�zI;ˤI;��I;E�I;_�H;�vF;]Q@;*:3;1 ;�r�: ��9:潺�G��z��X��ԟ�D4��%����ѽ*���Yb�!���̰�e���F���w�/蒿����r���      =�}���w�#f���K�r,�~�
�>�׾!�����k���'�fz꽝I���;V�:M�����iO�HG�,oE�������:�� ;�$;��8;��B;D�G;|KI;U�I;Z�I;��I;IqI;�SI;�=I;�-I;H"I;�I;YI;�I;YI;�I;H"I;�-I;�=I;�SI;GqI;��I;Z�I;R�I;|KI;A�G;��B;�8;�$;�� ;���:���+oE�HGໜiO����:M��;V��I��fz���'���k�!���>�׾~�
�r,���K�#f���w�      I(��$�f��R������~���`���Yb���'��U�H$��D�m�#����ϼ�/��.�������غ�:�9���:1G; H.;\|=;�E; ]H;h�I;��I;��I;=�I;BgI;ELI;'8I;I)I;�I;�I;�I;jI;�I;�I;�I;G)I;)8I;ELI;DgI;:�I;��I;��I;g�I;�\H;�E;Y|=; H.;3G;���:p:�9�غ����.���/����ϼ#��D�m�H$���U���'��Yb��`���~�����R��f���$�      C�׾��Ҿ ž�j��������z�U�H�*��fz�H$���/v�2+�ؐ�����5��ɻ�4�0&��:���:�o!;TP6;QlA;$�F;��H;ַI;��I;!�I;�}I;�\I;�DI;F2I;�$I;I;�I;�I;�I;�I;�I;I;�$I;H2I;�DI;�\I;�}I;!�I;��I;طI;��H; �F;MlA;TP6;|o!;���::&���4��ɻ��5���ؐ�2+��/v�H$��fz�*��U�H���z������j�� ž��Ҿ      �T��h�����z� Zb�(�D��$�����ѽ�I��C�m�2+�������>�K���Z�p���Ȕ�9�T�:0;��-;��<;�zD;�H;�mI;,�I;��I;ҕI;�oI;�RI;�<I;B,I; I;PI;tI;�I;I;�I;vI;PI; I;E,I;�<I;�RI;�oI;ҕI;��I;,�I;�mI;�H;�zD;��<;��-;0;�T�:���9Ɩ��W�p���>�K�������2+�C�m��I����ѽ���$�(�D� Zb���z�h���      �L+� (���G�������ս�@���%���;V�#��ؐ�����pMS�>�����C� 
o8�q�:;��$;B_7;t�A;��F;<�H;��I;��I;ɭI;#�I;�bI;�HI;Q5I;f&I;oI;�I;/I;I;H
I;I;0I;�I;oI;g&I;Q5I;�HI;�bI;#�I;ƭI;��I;��I;8�H;��F;u�A;B_7;��$;;�q�:�	o8�C���>��pMS�����ؐ�#���;V��%���@����ս����G��� (�      ��ս��ѽ=�ƽ2����I�����P�a�D4�:M���ϼ��>�K�>��-G��f���o�$��:bC�:�Y;)�1;�l>;#E;10H;_qI;D�I;/�I;�I;DsI;�UI;0?I;�-I;� I;�I;�I;I;TI;uI;TI;I;�I;�I;� I;�-I;2?I;�UI;DsI;�I;0�I;D�I;\qI;-0H;#E;�l>;)�1;�Y;fC�: ��:��o�f�,G��>��>�K�����ϼ9M�D4�P�a�����I��2���=�ƽ��ѽ      j��ѷ��#0v�q�a�"�G�>2+���ԟ�����/����5�����f��֬��g:��:J�;[I-;`g;;COC;NSG;�I;�I;d�I;C�I;H�I;NcI;�II;6I;�&I;I;xI;#I;�I;�I;�I;�I;�I;%I;xI;I;�&I;6I;�II;NcI;F�I;F�I;c�I;�I;�I;OSG;COC;cg;;[I-;N�;��:�g:�֬�f�������5��/�����ԟ���>2+�"�G�q�a�#0v�ѷ��      ��$�R5���������ϼš��X���iO�/���ɻX�p��C���o���g:u`�:�G;�*;�9;	�A;�uF;a�H;	�I;��I;�I;��I;�pI;yTI;�>I;^-I;�I;�I;:I;�I;�I;�I;I;�I;�I;�I;9I;�I;�I;^-I;�>I;yTI;�pI;��I;�I;��I;�I;c�H;�uF;	�A;�9;�*;�G;u`�:��g:��o��C�X�p��ɻ/���iO�X��š����ϼ������R5�%�      L�����*���9����N��Pp��D�x��GG໾����4����� 	o8$��:��:�G;H�(;�7;��@;�E;�QH;[mI;��I;=�I;ߢI;j}I;�^I;�FI;4I;&%I;�I;�I;3
I;PI; I;) I;��H;) I; I;QI;2
I;�I;�I;$%I;4I;�FI;�^I;l}I;ߢI;7�I;��I;]mI;�QH;
�E;��@;�7;I�(;�G;��:$��: 	o8�����4�����GG�x���D�Pp��N��9���*������      �iO�ԔK��o@���.�v��u����ɻ�G��+oE��غ&��Ȕ�9~q�:^C�:M�;�*;޶7;�P@; ]E;7H;JI;ýI;��I;O�I;��I;�hI;�NI;�:I;*I;�I;�I;I;XI;OI;o�H;��H;�H;��H;o�H;OI;XI;"I;�I;�I;|*I;�:I;�NI;�hI;��I;K�I;��I;ŽI;JI;8H;]E;�P@;ݶ7;�*;M�;bC�:�q�:Ȕ�9&���غ*oE��G���ɻs���u����.��o@�֔K�      ��ͻ(ɻa���~d������]�� �>潺����:�9:�T�:;�Y;^I-;�9;��@;]E;��G;y5I;��I;��I;�I;��I;�pI;�UI;�@I;v/I;�!I;�I;�I;�I;�I;`�H;��H;W�H;��H;W�H;��H;`�H;�I;�I;�I;�I;�!I;x/I;�@I;�UI;�pI;��I;�I;��I;��I;z5I;��G;]E;��@;�9;`I-;�Y;;�T�::�:�9���>潺� ��]�����d��a���(ɻ      >��ʟ�-i���غ������*�@ϭ� ��9���:���:���:0;��$;"�1;^g;;�A;�E;4H;u5I;�I;��I;��I;ۗI;�vI;�[I;�EI;�3I;v%I;�I;�I;�	I;�I;��H;��H;f�H;(�H;��H;*�H;f�H;��H;��H;�I;�	I;�I;�I;w%I;�3I;�EI;�[I;�vI;חI;��I;��I;��I;v5I;5H;�E;�A;^g;;"�1;��$;0;���:���:���:��9@ϭ��*�������غ,i�֟�      �/m8���8pdu9X��9d�9:���:WX�:�r�:�� ;3G;|o!;��-;@_7;�l>;BOC;�uF;�QH;JI;��I;��I;��I;��I;�zI;�_I;�II;�7I;�(I;�I;I;`I;'I;h I;��H;��H;B�H;#�H;��H;#�H;B�H;��H;��H;i I;(I;]I;I;�I;�(I;�7I;�II;�_I;�zI;��I;�I;��I;��I;JI;�QH;�uF;COC;�l>;@_7;��-;|o!;1G;�� ;�r�:SX�:���:h�9:h��9�du9@��8      �o�:%��:�K�:Z�:Ҩ�:a�;�;6 ;�$;H.;VP6;��<;o�A;!E;OSG;]�H;[mI;½I;��I;��I;��I;'|I;�aI;�KI;�9I;#+I;�I;�I;�I;jI;/I;4�H;�H;��H;/�H;M�H;�H;M�H;/�H;��H;�H;5�H;1I;fI;�I;�I;�I;%+I;�9I;�KI;�aI;)|I;��I;��I;��I;ŽI;XmI;\�H;QSG;!E;q�A;��<;TP6;H.;�$;6 ;�;c�;���:Z�:�K�:��:      ��;��;n];|X;o!;)9';�I-;(:3;��8;[|=;NlA;�zD;��F;00H;�I;�I;��I;��I;�I;ڗI;�zI;�aI;�LI;`;I;�,I;u I;fI;7I;|I;I;��H;<�H;��H;��H;H�H;��H;c�H;��H;H�H;��H;��H;=�H;��H;I;{I;:I;cI;v I;�,I;^;I;�LI;�aI;�zI;ޗI;�I;��I;��I;�I;�I;00H;��F;�zD;MlA;Y|=;��8;(:3;�I-;*9';o!;|X;p];��;      ��1;��1;83;�25;��7;ی:;v|=;]Q@;��B;�E;$�F;�H;6�H;_qI;�I;��I;;�I;P�I;��I;�vI;�_I;�KI;^;I;-I;.!I;]I;I;XI;�I;9�H;��H;��H;f�H;��H;��H;�H;��H;�H;��H;��H;c�H;��H;��H;6�H;�I;ZI;I;]I;/!I;-I;^;I;�KI;�_I;�vI;��I;R�I;:�I;��I;�I;_qI;6�H;�H;#�F;�E;��B;`Q@;t|=;݌:;ƶ7;�25;83;��1;      �?;A@;U�@;n�A;�B;B�C;fCE;�vF;C�G;�\H;��H;�mI;��I;F�I;d�I;�I;�I;��I;�pI;�[I;�II;�9I;�,I;5!I;�I;�I;�I;7I;��H;��H;��H;j�H;��H;0�H;.�H;��H;p�H;��H;/�H;/�H;��H;l�H;��H;��H;��H;9I;�I;�I;�I;1!I;�,I;�9I;�II;�[I;�pI;��I;�I;�I;d�I;D�I;��I;�mI;��H;�\H;A�G;�vF;fCE;@�C;�B;n�A;U�@;A@;      <vF;݊F;2�F;�!G;��G;KH;�H;U�H;zKI;d�I;ҷI;)�I;��I;.�I;@�I;��I;i}I;�hI;�UI;�EI;�7I;"+I;r I;\I;�I;	I;�I;��H;0�H;
�H;i�H;|�H;��H;��H;��H;Y�H;*�H;Y�H;��H;��H;��H;�H;i�H;
�H;/�H;��H;�I;	I;�I;ZI;r I;"+I;�7I;�EI;�UI;�hI;h}I;��I;C�I;.�I;��I;)�I;ѷI;a�I;yKI;W�H;�H;JH;��G;�!G;1�F;ъF;      � I;PI;wI;7I;*ZI;�}I;L�I;D�I;U�I;��I;��I;��I;ŭI;�I;H�I;�pI;�^I;�NI;�@I;�3I;�(I;�I;dI;I;�I;�I;�H;d�H;�H;w�H;e�H;��H;Z�H;Z�H;��H;G�H;�H;G�H;��H;Y�H;W�H;��H;g�H;v�H;�H;e�H;�H;�I;�I;I;dI;�I;�(I;�3I;�@I;�NI;�^I;�pI;H�I;�I;ƭI;��I;��I;��I;U�I;D�I;L�I;�}I;/ZI;�7I;uI;MI;      ��I;%�I;��I;��I;j�I;_�I;!�I;��I;]�I;��I;$�I;ՕI; �I;GsI;NcI;vTI;�FI;�:I;u/I;x%I;�I;�I;:I;[I;4I;��H;d�H;;�H;��H;d�H;��H;�H;�H;D�H;��H;@�H;.�H;@�H;��H;F�H;�H;"�H;��H;d�H;��H;;�H;d�H;��H;7I;]I;:I;�I;�I;x%I;u/I;�:I;�FI;wTI;NcI;GsI; �I;ՕI;"�I;��I;]�I;��I;!�I;_�I;u�I;��I;��I;2�I;      �I;U�I;��I;��I;��I;��I;��I;̤I;��I;:�I;�}I;�oI;�bI;�UI;�II;�>I; 4I;{*I;�!I;�I;I;�I;{I;�I;��H;2�H;�H;��H;m�H;��H;�H;��H;��H;;�H;��H;v�H;l�H;v�H;��H;;�H;��H;��H;�H;��H;n�H;��H;�H;0�H;��H;�I;{I;�I;I;�I;�!I;|*I;4I;�>I;�II;�UI;�bI;�oI;�}I;7�I;��I;̤I;��I;��I;��I;��I;��I;H�I;      ȟI;�I;��I;��I; �I;�I;��I;�zI;MqI;HgI;]I;�RI;�HI;6?I;6I;_-I;(%I;�I;�I;�I;`I;fI;	I;:�H;��H;�H;t�H;c�H;��H;�H;��H;��H;��H;^�H;��H;��H;��H;��H;��H;^�H;��H;��H;��H;�H;��H;e�H;t�H;�H;��H;9�H;I;gI;^I;�I;�I;�I;'%I;^-I;6I;6?I;�HI;�RI; ]I;HgI;MqI;�zI;��I;�I;��I;��I;��I;�I;      �vI;vI;tI;qI;�lI;�gI;�aI;
[I;�SI;HLI;�DI;�<I;S5I;�-I;�&I;�I;�I;�I;�I;�	I;-I;/I;��H;��H;��H;j�H;c�H;��H;�H;��H;��H;��H;*�H;��H;L�H;�H;��H;�H;L�H;��H;'�H;��H;��H;��H;�H;��H;d�H;h�H;��H;��H;��H;/I;*I;�	I;�I;�I;�I;�I;�&I;�-I;S5I;�<I;�DI;HLI;�SI;[I;�aI;�gI;�lI;qI;tI;vI;      �WI;|WI;VI;�SI;�PI;�LI;aHI;YCI;�=I;'8I;J2I;I,I;g&I;� I;I;�I;�I;I;�I;�I;o I;8�H;?�H;��H;i�H;|�H;��H; �H;��H;��H;��H;#�H;��H;�H;��H;��H;��H;��H;��H;�H;��H;&�H;��H;��H;��H;"�H;��H;{�H;m�H;��H;=�H;8�H;n I;�I;�I;I;�I;�I;I;� I;g&I;I,I;J2I;)8I;�=I;YCI;aHI;�LI;�PI;�SI;VI;vWI;      BI;�AI;�@I;�>I;[<I;Z9I;�5I;�1I;�-I;F)I;�$I; I;oI;�I;xI;:I;6
I;RI;�I;��H;��H;�H;��H;i�H;��H;��H;Z�H;�H;��H;��H;,�H;��H;��H;��H;M�H;!�H;)�H;!�H;M�H;��H;��H;��H;,�H;��H;��H;�H;W�H;��H;��H;i�H;��H;�H;��H;��H;�I;TI;6
I;:I;xI;�I;oI; I;�$I;G)I;�-I;�1I;�5I;[9I;V<I;�>I;�@I;�AI;      =2I;�1I;1I;�/I;�-I;q+I;�(I;�%I;K"I;�I;I;SI;�I;�I;'I;�I;WI;MI;d�H;��H;��H;��H;��H;��H;)�H;��H;V�H;C�H;9�H;]�H;��H;�H;��H;2�H;�H;��H;��H;��H;�H;2�H;��H;�H;��H;^�H;=�H;C�H;V�H;��H;,�H;��H;��H;��H;��H;��H;d�H;NI;UI;�I;'I;�I;�I;SI;I;�I;M"I;�%I;�(I;u+I;�-I;�/I;1I;�1I;      (I;�'I;)'I;�%I;e$I;\"I; I;�I;�I;�I;�I;}I;3I;	I;I;�I;'I;k�H;��H;j�H;I�H;0�H;H�H;��H;'�H;��H;��H;��H;��H;��H;K�H;��H;K�H;	�H;��H;��H;��H;��H;��H;	�H;H�H;��H;L�H;��H;��H;��H;��H;��H;(�H;��H;H�H;0�H;H�H;j�H;��H;m�H;%I;�I;I;
I;3I;}I;�I;�I;�I;�I; I;`"I;]$I;�%I;)'I;�'I;      "I;�!I;Q!I;b I;I;.I;"I;�I;cI;�I;�I;�I;"I;]I;�I;�I;0 I;��H;\�H;/�H;,�H;P�H;��H;�H;��H;S�H;D�H;@�H;w�H;��H;�H;��H; �H;��H;��H;p�H;j�H;p�H;��H;��H;�H;��H;�H;��H;z�H;@�H;C�H;R�H;��H;�H;��H;P�H;*�H;/�H;\�H;��H;. I;�I;�I;[I;"I;�I;�I;�I;cI;�I;"I;4I;I;b I;Q!I;�!I;      * I; I;yI;qI;I;dI;�I;eI;�I;dI;�I;I;H
I;{I;�I;I;��H;�H;��H;��H;��H;�H;c�H;��H;l�H;#�H;	�H;2�H;n�H;��H;��H;��H;)�H;��H;��H;l�H;P�H;l�H;��H;��H;(�H;��H;��H;��H;p�H;2�H;�H;%�H;l�H;��H;c�H;�H;��H;��H;��H;�H;��H;I;�I;{I;H
I;I;�I;gI;�I;eI;�I;hI;I;qI;yI;
 I;      "I;�!I;Q!I;b I;I;/I;"I;�I;cI;�I;�I;�I;"I;]I;�I;�I;0 I;��H;\�H;/�H;-�H;P�H;��H;�H;��H;S�H;D�H;@�H;w�H;��H;�H;��H; �H;��H;��H;p�H;j�H;p�H;��H;��H;�H;��H;�H;��H;z�H;@�H;C�H;R�H;��H;�H;��H;P�H;*�H;/�H;\�H;��H;. I;�I;�I;[I;"I;�I;�I;�I;cI;�I;"I;2I;I;b I;N!I;�!I;      (I;�'I;('I;�%I;e$I;\"I; I;�I;�I;�I;�I;}I;3I;	I;I;�I;'I;k�H;��H;j�H;J�H;0�H;H�H;��H;(�H;��H;��H;��H;��H;��H;L�H;��H;K�H;	�H;��H;��H;��H;��H;��H;	�H;H�H;��H;K�H;��H;��H;��H;��H;��H;'�H;��H;H�H;0�H;H�H;j�H;��H;m�H;%I;�I;I;
I;3I;}I;�I;�I;�I;�I; I;`"I;]$I;�%I;('I;�'I;      ?2I;�1I;1I;�/I;�-I;q+I;�(I;�%I;K"I;�I;I;SI;�I;�I;'I;�I;WI;MI;d�H;��H;�H;��H;��H;��H;,�H;��H;V�H;C�H;9�H;]�H;��H;�H;��H;2�H;�H;��H;��H;��H;�H;2�H;��H;�H;��H;^�H;<�H;C�H;V�H;��H;)�H;��H;��H;��H;��H;��H;d�H;NI;UI;�I;'I;�I;�I;SI;I;�I;M"I;�%I;�(I;u+I;�-I;�/I;1I;�1I;      BI;�AI;�@I;�>I;[<I;Z9I;�5I;�1I;�-I;F)I;�$I; I;oI;�I;xI;:I;7
I;RI;�I;��H;��H;�H;��H;i�H;��H;��H;Z�H;�H;��H;��H;,�H;��H;��H;��H;M�H;!�H;)�H;!�H;K�H;��H;��H;��H;,�H;��H;��H;�H;W�H;��H;��H;h�H;��H;�H;��H;��H;�I;RI;5
I;:I;xI;�I;nI; I;�$I;G)I;�-I;�1I;�5I;[9I;T<I;�>I;�@I;�AI;      �WI;|WI;VI;�SI;�PI;�LI;dHI;YCI;�=I;)8I;J2I;I,I;g&I;� I;I;�I;�I;I;�I;�I;r I;8�H;?�H;��H;m�H;|�H;��H;"�H;��H;��H;��H;#�H;��H;�H;��H;��H;��H;��H;��H;�H;��H;%�H;��H;��H;��H; �H;��H;{�H;i�H;��H;=�H;8�H;n I;�I;�I;I;�I;�I;I;� I;g&I;I,I;J2I;*8I;�=I;YCI;dHI;�LI;�PI;�SI;VI;xWI;      �vI;vI;tI;qI;�lI;�gI;�aI;
[I;�SI;FLI;�DI;�<I;S5I;�-I;�&I;�I;�I;�I;�I;�	I;.I;/I;��H;��H;��H;j�H;d�H;��H;�H;��H;��H;��H;)�H;��H;L�H;�H;��H;�H;L�H;��H;'�H;��H;��H;��H;�H;��H;c�H;h�H;��H;��H;��H;/I;*I;�	I;�I;�I;�I;�I;�&I;�-I;S5I;�<I;�DI;ILI;�SI;[I;�aI;�gI;�lI;qI;tI;vI;      I;�I;��I;��I;��I;�I;��I;�zI;NqI;GgI;]I;�RI;�HI;6?I;6I;^-I;(%I;�I;�I;�I;aI;gI;	I;:�H;��H;�H;v�H;e�H;��H;�H;��H;��H;��H;]�H;��H;��H;��H;��H;��H;^�H;��H;��H;��H;�H;��H;c�H;s�H;�H;��H;<�H;I;fI;^I;�I;�I;�I;'%I;a-I;6I;6?I;�HI;�RI;]I;GgI;PqI;�zI;��I;�I;��I;��I;��I;�I;      �I;Q�I;��I;��I;��I;��I;��I;̤I;��I;8�I;�}I;�oI;�bI;�UI;�II;�>I; 4I;{*I;�!I;�I;I;�I;|I;�I;��H;2�H;�H;��H;n�H;��H;�H;��H;��H;;�H;��H;v�H;l�H;v�H;��H;;�H;��H;��H;�H;��H;m�H;��H;�H;0�H;��H;�I;yI;�I;I;�I;�!I;|*I;4I;�>I;�II;�UI;�bI;�oI;�}I;:�I;��I;ΤI;��I;��I;��I;��I;��I;Q�I;      ��I;&�I;��I;��I;k�I;_�I;!�I;��I;]�I;��I;$�I;ՕI; �I;GsI;NcI;wTI;�FI;�:I;u/I;x%I;�I;�I;<I;]I;7I;��H;d�H;;�H;��H;g�H;��H; �H;�H;D�H;��H;@�H;.�H;@�H;��H;D�H;�H; �H;��H;c�H;��H;;�H;d�H;��H;4I;[I;9I;�I;�I;x%I;u/I;�:I;�FI;wTI;NcI;GsI; �I;ՕI;"�I;��I;^�I;��I;!�I;\�I;v�I;��I;��I;0�I;      � I;PI;uI;{7I;'ZI;�}I;K�I;D�I;U�I;��I;��I;��I;ƭI;�I;F�I;�pI;�^I;�NI;�@I;�3I;�(I;�I;fI;I;�I;�I;�H;e�H;�H;w�H;g�H;��H;X�H;Y�H;��H;G�H;�H;F�H;��H;Y�H;X�H;��H;e�H;v�H;�H;d�H;�H;�I;�I;I;cI;�I;�(I;�3I;�@I;�NI;�^I;�pI;F�I;�I;ŭI;��I;��I;��I;U�I;E�I;K�I;�}I;(ZI;z7I;rI;DI;      AvF;ԊF;<�F;�!G;��G;MH;�H;X�H;yKI;c�I;ҷI;'�I;��I;.�I;@�I;��I;i}I;�hI;�UI;�EI;�7I;"+I;r I;\I;�I;	I;�I;��H;0�H;�H;i�H;|�H;��H;��H;��H;Y�H;*�H;Y�H;��H;��H;��H;}�H;i�H;�H;/�H;��H;�I;	I;�I;YI;r I;"+I;�7I;�EI;�UI;�hI;h}I;��I;@�I;.�I;��I;)�I;ҷI;c�I;yKI;X�H;�H;KH;��G;�!G;9�F;̊F;      �?;A@;U�@;n�A;�B;B�C;fCE;�vF;A�G;�\H;��H;�mI;��I;D�I;d�I;�I;�I;��I;�pI;�[I;�II;�9I;�,I;5!I;�I;�I;�I;9I;��H;��H;��H;j�H;��H;/�H;.�H;��H;p�H;��H;.�H;/�H;��H;m�H;��H;��H;��H;7I;�I;�I;�I;2!I;�,I;�9I;�II;�[I;�pI;��I;�I;�I;d�I;D�I;��I;�mI;��H;�\H;A�G;�vF;fCE;B�C;�B;n�A;U�@;?@;      ��1;��1;83;�25;��7;�:;p|=;`Q@;��B;�E;#�F;�H;9�H;_qI;�I;��I;;�I;P�I;��I;�vI;�_I;�KI;`;I;-I;/!I;]I;I;ZI;�I;9�H;��H;��H;c�H;��H;��H;�H;��H;�H;��H;��H;e�H;��H;��H;6�H;�I;XI;I;]I;.!I;-I;];I;�KI;�_I;�vI;��I;R�I;:�I;��I;�I;_qI;8�H;�H;#�F;�E;��B;`Q@;p|=;�:;ɶ7;�25;83;��1;      ��;��;|];|X;o!;+9';�I-;(:3;��8;[|=;MlA;�zD;��F;00H;�I;�I;��I;��I;�I;ݗI;�zI;�aI;�LI;a;I;�,I;u I;fI;:I;}I;I;��H;=�H;��H;��H;H�H;��H;c�H;��H;H�H;��H;��H;<�H;��H;	I;yI;7I;dI;v I;�,I;];I;�LI;�aI;�zI;ݗI;�I;��I;��I;�I;�I;00H;��F;�zD;NlA;Y|=;��8;*:3;�I-;.9';o!;|X;r];��;      �o�:%��:�K�:Z�:Ԩ�:a�;�;5 ;�$;H.;TP6;��<;q�A;!E;OSG;]�H;ZmI;ýI;��I;��I;��I;)|I;�aI;�KI;�9I;%+I;�I;�I;�I;jI;1I;5�H;�H;��H;/�H;N�H;�H;M�H;/�H;��H;�H;2�H;/I;fI;�I;�I;�I;%+I;�9I;�KI;�aI;'|I;��I;��I;��I;ýI;ZmI;]�H;QSG;!E;o�A;��<;TP6;H.;�$;6 ;�;a�;���:Z�:�K�:��:       .m8���8�du9h��9d�9:���:YX�:�r�:�� ;1G;|o!;��-;@_7;�l>;COC;�uF;�QH;JI;��I;��I;��I;��I;�zI;�_I;�II;�7I;�(I;�I;I;`I;(I;h I;��H;��H;B�H;#�H;��H;#�H;B�H;��H;��H;i I;'I;]I;I;�I;�(I;�7I;�II;�_I;�zI;��I;�I;��I;��I;JI;�QH;�uF;BOC;�l>;@_7;��-;|o!;0G;�� ;�r�:YX�:���:x�9:h��9�du9`��8      >��̟�'i���غ������*� ϭ���9���:���:���:0;��$;"�1;^g;;�A;�E;4H;v5I;�I;��I;��I;ۗI;�vI;�[I;�EI;�3I;w%I;�I;�I;�	I;�I;��H;��H;f�H;+�H;��H;*�H;f�H;��H;��H;�I;�	I;�I;�I;v%I;�3I;�EI;�[I;�vI;חI;��I;��I;��I;u5I;5H;�E;�A;^g;;"�1;��$;0;���:���:���: ��9 ϭ��*�������غ*i�ן�      ��ͻ(ɻb����d������]�� �>潺����:�9:�T�:;�Y;^I-;�9;��@;]E;��G;z5I;��I;��I; �I;��I;�pI;�UI;�@I;x/I;�!I;�I;�I;�I;�I;`�H;��H;W�H;��H;W�H;��H;`�H;�I;�I;�I;�I;�!I;v/I;�@I;�UI;�pI;��I;�I;��I;��I;|5I;��G;]E;��@;�9;`I-;�Y;;�T�::�:�9���:潺� ��]����~d��a���(ɻ      �iO�ԔK��o@���.�v��u����ɻ�G��+oE��غ&��Ȕ�9�q�:^C�:M�;�*;޶7;�P@;]E;7H;JI;ŽI;��I;O�I;��I;�hI;�NI;�:I;*I;�I;�I; I;YI;OI;o�H;��H;�H;��H;o�H;OI;VI;I;�I;�I;|*I;�:I;�NI;�hI;��I;K�I;��I;ýI;JI;8H; ]E;�P@;޶7;�*;M�;^C�:~q�:Ȕ�9&���غ*oE��G���ɻs���u����.��o@�֔K�      L�����*���9����N��Pp��D�x��GG໾����4����� 	o8$��:��:�G;J�(;�7;��@;�E;�QH;]mI;��I;;�I;ߢI;j}I;�^I;�FI;4I;&%I;�I;�I;3
I;QI;!I;) I;��H;) I; I;QI;2
I;�I;�I;$%I;4I;�FI;�^I;l}I;ߢI;7�I;��I;[mI;�QH;
�E;��@;�7;H�(;�G;��:$��: 	o8�����4�����GG�x���D�Pp��N��9���*������      ��$�R5���������ϼš��X���iO�/���ɻX�p��C���o���g:u`�:�G;�*;�9;	�A;�uF;c�H;	�I;��I;�I;��I;�pI;yTI;�>I;^-I;�I;�I;:I;�I;�I;�I;I;�I;�I;�I;9I;�I;�I;^-I;�>I;yTI;�pI;��I;�I;��I;�I;a�H;�uF;	�A;�9;�*;�G;u`�:��g:��o��C�X�p��ɻ/���iO�X��š����ϼ������R5�%�      j��ѷ��#0v�q�a�"�G�>2+���ԟ�����/����5�����f��֬��g:��:K�;[I-;bg;;BOC;OSG;�I;�I;c�I;E�I;I�I;NcI;�II;6I;�&I;I;xI;%I;�I;�I;�I;�I;�I;%I;xI;I;�&I;6I;�II;NcI;F�I;E�I;d�I;�I;�I;NSG;BOC;cg;;[I-;M�;��:�g:�֬�f�������5��/�����ԟ���>2+�"�G�q�a�#0v�ѷ��      ��ս��ѽ=�ƽ2����I�����P�a�D4�9M���ϼ��>�K�>��-G��f���o�&��:dC�:�Y;(�1;�l>;#E;10H;_qI;D�I;/�I;�I;DsI;�UI;0?I;�-I;� I;�I;�I;I;TI;uI;TI;I;�I;�I;� I;�-I;2?I;�UI;DsI;�I;0�I;D�I;\qI;,0H;#E;�l>;(�1;�Y;fC�: ��:��o�f�-G��>��>�K�����ϼ9M�D4�P�a�����I��2���=�ƽ��ѽ      �L+� (���G�������ս�@���%���;V�#��ؐ�����pMS�>�����C� 
o8�q�:;��$;A_7;u�A;��F;<�H;��I;��I;ɭI;#�I;�bI;�HI;Q5I;f&I;oI;�I;0I;I;H
I;I;/I;�I;nI;d&I;Q5I;�HI;�bI;#�I;ƭI;��I;��I;6�H;��F;t�A;B_7;��$;;�q�:�	o8�C���>��pMS�����ؐ�#���;V��%���@����ս����G��� (�      �T��h�����z� Zb�(�D��$�����ѽ�I��C�m�2+�������>�K���W�p�����Д�9�T�:0;��-;��<;�zD;�H;�mI;,�I;��I;ҕI;�oI;�RI;�<I;B,I; I;RI;wI;�I;I;�I;vI;PI; I;C,I;�<I;�RI;�oI;ҕI;��I;,�I;�mI;�H;�zD;��<;��-;0;�T�:��9Ɩ��[�p���>�K�������2+�C�m��I����ѽ���$�(�D� Zb���z�h���      C�׾��Ҿ ž�j��������z�U�H�*��fz�H$���/v�2+�ؐ�����5��ɻ�4�(&��:���:|o!;TP6;QlA;$�F;��H;ַI;��I;!�I;�}I;�\I;�DI;F2I;�$I;I;�I;�I;�I;�I;�I;I;�$I;G2I;�DI;�\I;�}I;!�I;��I;طI;��H; �F;MlA;TP6;~o!;���::&���4��ɻ��5���ؐ�2+��/v�H$��fz�*��U�H���z������j�� ž��Ҿ      I(��$�f��R������~���`���Yb���'��U�H$��D�m�#����ϼ�/��.�������غp:�9���:0G; H.;\|=;�E;�\H;g�I;��I;��I;=�I;BgI;ELI;'8I;I)I;�I;�I;�I;jI;�I;�I;�I;G)I;'8I;ELI;DgI;:�I;��I;��I;h�I; ]H;�E;Y|=; H.;1G;���:�:�9�غ����.���/����ϼ#��D�m�H$���U���'��Yb��`���~�����R��f���$�      =�}���w�#f���K�r,�~�
�>�׾!�����k���'�fz꽝I���;V�:M�����iO�HG�,oE�������:�� ;�$;��8;��B;A�G;zKI;U�I;Z�I;��I;FqI;�SI;�=I;�-I;H"I;�I;YI;�I;YI;�I;H"I;�-I;�=I;�SI;GqI;��I;Z�I;R�I;|KI;D�G;��B;�8;�$;�� ;���:���+oE�IGໜiO����:M��;V��I��fz���'���k�!���>�׾~�
�r,���K�#f���w�      ��r�������/蒿��w��F�e��̰�!����Yb�*����ѽ�%��D4�ԟ�X��y���G��:潺0��9�r�:1 ;+:3;`Q@;�vF;_�H;H�I;��I;ΤI;�zI;
[I;SCI;�1I;�%I;�I;�I;dI;�I;�I;�%I;�1I;SCI;
[I;�zI;ˤI;��I;G�I;^�H;�vF;]Q@;*:3;1 ;�r�: ��9:潺�G��z��X��ԟ�D4��%����ѽ*���Yb�!���̰�e���F���w�/蒿����r���      5��������㿌�ɿ���˅����P�e��>�׾�`��U�H����@��Q�a���ơ���D��ɻ� ��έ�MX�:�;�I-;o|=;iCE;�H;I�I;!�I;��I;�I;�aI;eHI;�5I;�(I; I;I;�I;I; I;�(I;�5I;eHI;�aI;�I;��I;!�I;I�I;�H;lCE;l|=;�I-;�;SX�: ϭ�� ��ɻ�D�ơ����Q�a��@����U�H��`��>�׾e����P�˅�������ɿ�㿵���      Ǚ$��x �$��<���޿q���˅���F�~�
��~����z��$���ս���>2+���ϼPp�q����]��*����:W�;)9';ތ:;?�C;QH;�}I;b�I;��I;�I;�gI;�LI;^9I;y+I;d"I;6I;jI;6I;d"I;x+I;[9I;�LI;�gI;�I;��I;b�I;�}I;PH;@�C;ڌ:;)9';Y�;���:�*��]�p���Pp���ϼ>2+������ս�$���z��~��~�
��F�˅��q����޿<��$���x �      L�Q���K���;�Ǚ$��;
��޿�����w�r,���澞���(�D������I��"�G����N��v���������t�9:ڨ�:o!;��7;�B;��G;(ZI;l�I;��I;��I;�lI;�PI;W<I;�-I;T$I; I;I; I;S$I;�-I;V<I;�PI;�lI;��I;��I;l�I;*ZI;��G;�B;��7;o!;ڨ�:��9:�������v���N�����"�G��I������(�D��������r,���w�����޿�;
�Ǚ$���;���K�      U����{���d��F�Ǚ$�<����ɿ0蒿��K�R���j�� Zb�G�2���q�a����9�����.��d����غx��9+Z�:�X;�25;h�A;�!G;{7I;��I;��I;��I;�pI;�SI;�>I;�/I;�%I;a I;qI;a I;�%I;�/I;�>I;�SI;�pI;��I;��I;��I;{7I;�!G;j�A;�25;�X;+Z�:���9��غ�d����.�:������q�a�2���G� Zb��j��R����K�0蒿��ɿ<��Ǚ$��F���d��{�      ����$P�������d���;�$���㿴���#f�f�� ž��z���=�ƽ$0v�R5�*����o@�g���.i� du9�K�:j];83;h�@;?�F;xI;��I;��I;��I;tI;VI;�@I;#1I;('I;L!I;qI;L!I;('I;#1I;�@I;VI;tI;��I;��I;��I;xI;?�F;h�@;83;m];�K�:0du9.i�g����o@�*���R5�$0v�=�ƽ����z� žf��#f�������$����;���d����$P��      �,��b��$P���{���K��x �����r�����w��$���Ҿg��� (���ѽѷ��%����ՔK�(ɻݟ����8��:��;��1;7@;ʊF;NI;"�I;X�I;�I;�uI;nWI;�AI;�1I;�'I;�!I; I;�!I;�'I;�1I;�AI;oWI;�uI;��I;U�I;"�I;MI;ɊF;7@;��1;��;��:���8ݟ�(ɻԔK����%�ѷ����ѽ (�g�����Ҿ�$���w�r��������x ���K��{�$P��b��      ᶕ�T���Ҭ��/�_���7�{�!}߿����,b��V�.l¾Jx�d.���Ž��t�'��_����?��M��ٯ�P�x9���:��;ȼ2;w@@;�fF;_�H;ĉI;��I;T|I;\I;�CI;F2I;�%I;�I;�I;oI;�I;�I;�%I;D2I;�CI;\I;T|I;��I;ĉI;_�H;�fF;w@@;Ƽ2;��;���:`�x9ٯ��M����?�_��'����t���Žd.�Jx�.l¾�V��,b����!}߿{���7�/�_�Ҭ��T���      T���E���%}��+Y��3�����$ڿ&��ƽ\����(���s��3�6����p�a�N���<<������ؘ�9���:'�;v%3;�p@;zF;��H;=�I;6�I;�{I;�[I;�CI;�1I;�%I;cI;�I;DI;�I;fI;�%I;�1I;�CI;�[I;�{I;3�I;=�I;��H;zF;�p@;r%3;,�;���:ؘ�9������<<�N��a��p�6����3��s�(�����ƽ\�&���$ڿ����3��+Y�%}�E���      Ҭ��%}�?tf��lG�آ%��p�0�ʿ\����>M����V�����d�ɤ�̷�-�d��
�I����1�H������ ��9���:p;�U4;��@;0�F;^�H; �I;��I;�yI;�YI;�BI;1I;�$I;�I;I;�I;I;�I;�$I;1I;�BI;�YI;�yI;��I; �I;^�H;0�F;��@;�U4;s;���:��9���H�����1��I���
�-�d�̷�ɤ���d�V�������>M�\���0�ʿ�p�آ%��lG�?tf�%}�      /�_��+Y��lG�f.�{���꿲���O䂿��5���󾏰��O�N�W��S�� �Q����v����h!�kg����,
:�
�:A�;�16;��A;�G;.I;y�I;ƘI;�vI;�WI;�@I;�/I;�#I;�I;HI;�I;HI;�I;�#I;�/I;�@I;�WI;�vI;ØI;y�I;.I;�G;��A;�16;D�;�
�:0
:��kg���h!�v������ �Q�S��W��O�N���������5�O䂿�������{�f.��lG��+Y�      ��7��3�آ%�{��<����ſ
���Ľ\�=����Ͼ����a�3��轻z��{�9�Y�ἔ���z�_7}�hct���^:�+�:�#;ڍ8;��B;bsG;�%I;�I;1�I;?rI;STI;$>I;�-I;O"I;�I;$I;�I;$I;�I;Q"I;�-I;%>I;STI;<rI;/�I;�I;�%I;`sG;��B;֍8;��#;�+�:��^:hct�_7}��z����Y��{�9��z����a�3�������Ͼ=��Ľ\�
�����ſ�<��{�آ%��3�      {�����p������ſ&���Ps���1�3r���d���d�}I�ψŽ��}�]*�EC���^��B�@�D��D�� �:��;�);Q7;;oD;��G;�HI;�I;�I;�lI;1PI;
;I;U+I;[ I;�I;�I;kI;�I;�I;[ I;U+I;;I;1PI;�lI;�I;�I;�HI;��G;mD;L7;;�);��; �:�D�@�D��B��^�EC��]*���}�ψŽ}I��d��d��3r����1��Ps�&����ſ��꿄p����      !}߿�$ڿ0�ʿ����
����Ps�RX:����'l¾�ǆ���7����85���Q�����t���75�N��b���$�8Qʼ:��;�.;��=;�EE;ZH;�hI;f�I;��I;cfI;]KI;e7I;�(I;I;/I; I;�I; I;/I;I;�(I;g7I;\KI;bfI;��I;f�I;�hI;ZH;�EE;��=; �.;��;Sʼ:`$�8b��L���75��t������Q�85�������7��ǆ�'l¾���RX:��Ps�
�������0�ʿ�$ڿ      ���&��\���N䂿Ľ\���1�����J˾Ꝓ�F�N�y��I������T�'�_�Ҽ��|��z��n���w����&:Q�:�;�W4;	�@;kgF;��H;N�I;`�I;u�I;W_I;FI;H3I;_%I;�I;�I; I;�I; I;�I;�I;\%I;H3I;FI;W_I;r�I;`�I;K�I;��H;hgF;�@;�W4;�;Q�:��&:�w���n���z���|�_�ҼT�'����I���y��F�N�Ꝓ��J˾�����1�Ľ\�N䂿\���&��      �,b�ƽ\��>M���5�=��3r��'l¾Ꝓ�$&W��3�9Sؽ�z��XG����wI����?�u�̻Q�-�������:��;��&;g|9;C;�dG;�I;}�I;��I;�vI;�WI;l@I;�.I;�!I;�I;�I;I;�I;I;�I;�I;�!I;�.I;l@I;�WI;�vI;��I;z�I;�I;�dG;C;d|9;��&;��;���:���P�-�u�̻��?�wI�����XG��z��9Sؽ�3�$&W�Ꝓ�'l¾3r��=����5��>M�ƽ\�      �V������������Ͼ�d���ǆ�F�N��3��c�[����\�1��$C���o���	��눻�ﳺ���9���:�h;��/;��=;�E;=3H;�WI;��I;9�I; lI;�OI;d:I;(*I;_I;�I;1I;�I;�I;�I;1I;�I;]I;)*I;c:I;�OI;�kI;9�I;��I;�WI;93H;~E;}�=;��/;�h;���:���9�ﳺ�눻��	��o�$C��0����\�[���cི3�F�N��ǆ��d����Ͼ���������      .l¾(��V������������d���7�y��9Sؽ[���d�A*�_kּ&\����'���lR�`|����:�Z;�#;z=7;r�A;T�F;��H;��I;(�I;�I;-aI;�GI;34I;c%I;�I;�I;�I;�
I;�	I;�
I;�I;�I;�I;f%I;34I;�GI;*aI;�I;'�I;��I;��H;Q�F;n�A;z=7;�#;�Z;��:H|��mR�����'�&\��^kּA*��d�[��9Sؽy����7��d���������V���(��      Jx��s���d�O�N�a�3�}I����I����z����\�A*��ݼB���#<<��ڻЗV�Hct��&:��:�C;�</;�D=;�D;��G;79I;�I;�I;TtI;mVI;�?I;�-I;� I;�I;�I;�
I;7I;SI;7I;�
I;�I;�I;� I;�-I;�?I;kVI;TtI;�I;�I;59I;��G;�D;�D=;�</;�C;��:$�&:Lct�ЗV��ڻ#<<�B����ݼA*���\��z��I������}I�b�3�O�N���d��s�      d.��3�ɤ�W����ψŽ85�����XG�1��^kּB����xC�{>�+6}����� �x9؏�:L	;w�&;�;8;��A;�F;�H;yyI;ԝI;5�I;pfI;LI;�7I;�'I;�I;	I;�I;QI;�I;�I;�I;QI;�I;	I;�I;�'I;�7I;LI;qfI;1�I;֝I;vyI;�H;��F;��A;�;8;v�&;L	;܏�:��x9����+6}�{>��xC�B���^kּ1��XG����85��ψŽ��W��ɤ��3�      ��Ž6���̷�S���z����}��Q�T�'����$C��&\��#<<�|>�hn����� ����:���:P�;�'3;��>;�E;�H;�<I;�I;�I;�vI;YI;�AI;�/I;�!I;!I;/I;�	I;�I;aI;�I;aI;�I;�	I;/I;#I;�!I;�/I;�AI;YI;�vI;�I;�I;�<I;�H;�E;��>;�'3;P�;���:���: ����hn��|>�#<<�&\��$C�����T�'��Q���}��z��S��̷�6���      ��t��p�-�d� �Q�|�9�]*����`�ҼwI��	�o���'��ڻ,6}�����5�0�:�m�:��;+�.;^<;�oC;�7G;��H;�I;�I;�I;_fI;�LI;88I; (I;I;�I;�I;�I;�I;	I;� I;	I;�I;�I;�I;�I;I;(I;58I;�LI;]fI;�I;�I;�I;��H;�7G;�oC;^<;,�.;��;�m�:0�:�5����,6}��ڻ��'��o�wI��`�Ҽ���]*�|�9� �Q�-�d��p�      '��a��
�
���Y��EC���t����|���?���	���ЗV�����@�8�:C�:i;]�+;5�9;��A;�fF;��H;�_I;̛I;ّI;FsI;�VI;�@I;/I;-!I;�I;KI;I;�I;� I;��H;G�H;��H;� I;�I;I;MI;�I;-!I;/I;�@I;�VI;FsI;ؑI;țI;�_I;��H;�fF;��A;5�9;`�+;i;C�:8�: �����ЗV�����	���?���|��t��EC��Z��
����
�a�      _��L���I��v�������^��75��z�t�̻�눻kR�Hct���x9���:�m�:i;��*;�8;+�@;#�E;|(H;�8I;�I;W�I;�~I;�`I;�HI;�5I;�&I;�I;wI;:
I;�I;� I;0�H;��H;#�H;��H;0�H;� I;�I;<
I;wI;�I;�&I;�5I;�HI;�`I;�~I;S�I;��I;�8I;z(H;&�E;+�@;�8;��*;i;�m�:���:��x9Hct�lR��눻t�̻�z��75��^����v����I��N��      ��?��<<���1��h!��z��B�N���n��P�-��ﳺH|���&:֏�:���:��;Z�+;�8;z�@;/^E;��G;�I;-�I;��I;u�I;�iI;|PI;H<I;�+I;�I;�I;�I;jI;�I;�H;��H;��H;�H;��H;��H;�H;�I;kI;�I;�I;�I;�+I;E<I;}PI;�iI;q�I;��I;-�I;�I;��G;0^E;{�@;�8;Z�+;��;���:֏�:�&:H|���ﳺO�-��n��N���B黬z��h!���1��<<�      �M����D���jg��c7}�=�D�[���w��������9��:��:J	;Q�;/�.;2�9;)�@;/^E;��G;�I;�I;G�I;��I;�pI;�VI;�AI;�0I;�"I;�I;,I;.I;�I;��H;��H;��H;��H;�H;��H;��H;��H;��H;�I;.I;)I;�I;�"I;�0I;�AI;�VI;�pI;��I;I�I;�I;�I;��G;2^E;(�@;2�9;/�.;S�;J	;��:��:���9x���w��]��7�D�]7}�jg��D�����      ׯ���������tct��D�@$�8��&:���:���:�Z;�C;r�&;�'3;Z<;��A;!�E;��G;I;�|I;�I;�I;�uI;�[I;MFI;�4I;n&I;�I;�I;"
I;3I;x�H;�H;v�H;��H;��H;_�H;��H;��H;v�H;�H;y�H;3I; 
I;�I;�I;k&I;�4I;NFI;�[I;�uI;�I;�I;�|I;�I;��G;!�E;��A;X<;�'3;r�&;�C;�Z;���:���:��&:@$�8�D�Tct��𳺾�����      ��x9H��98��9
:��^: �:Sʼ:Q�:��;�h;�#;�</;�;8;��>;�oC;�fF;z(H;�I;�I;�I;�I;>xI;�^I;}II;�7I;L)I;MI;�I;�I;�I;� I;��H;��H;x�H;��H;��H;��H;��H;��H;x�H;��H;��H;� I;�I;�I;�I;JI;L)I;�7I;xII;�^I;?xI;�I;�I;�I;�I;z(H;�fF;�oC;��>;�;8;�</;�#;�h;��;Q�:Sʼ:�:��^:
:@��9���9      	��:���:��:�
�:�+�:��;�;�;��&;��/;}=7;�D=;��A;�E;�7G;��H;�8I;+�I;F�I;�I;;xI;�_I;%KI;�9I;7+I;@I;zI;{I;�I;}I;@�H;��H;Z�H;{�H;�H;L�H;(�H;L�H;�H;{�H;W�H;��H;B�H;zI;�I;}I;vI;@I;;+I;�9I;"KI;�_I;;xI;�I;G�I;-�I;�8I;��H;�7G;�E;��A;�D=;|=7;��/;��&;�;�;��;�+�:�
�:��:���:      ��;+�;s;;�;�#;�);�.;�W4;i|9;~�=;o�A;�D;��F;�H;��H;�_I;�I;��I;��I;�uI;�^I;&KI;f:I;a,I;| I;�I;�I;�I;cI;��H;C�H;r�H;J�H;��H;��H;��H;��H;��H;��H;��H;I�H;r�H;C�H;��H;bI;�I;�I;�I;} I;^,I;f:I;&KI;�^I;�uI;��I;��I;�I;�_I;��H;�H;�F;�D;n�A;}�=;h|9;�W4;�.;�);�#;:�;u; �;      ݼ2;�%3;�U4;�16;ٍ8;O7;;��=;�@;C;�E;T�F;��G;�H;�<I;�I;țI;V�I;u�I;�pI;�[I;xII;�9I;^,I;� I;^I;aI;�I;I;��H;��H;��H;h�H;}�H;�H;+�H;��H;A�H;��H;-�H;�H;{�H;j�H;��H;��H;��H;I;�I;aI;`I;� I;^,I;�9I;vII;�[I;�pI;x�I;T�I;țI;�I;�<I;�H;��G;S�F;~E;C;�@;��=;Q7;;��8;�16;�U4;|%3;      �@@;�p@;��@;��A;��B;oD;�EE;egF;�dG;93H;��H;69I;uyI;�I;�I;ّI;�~I;�iI;�VI;QFI;�7I;;+I;� I;dI;�I;�I;�I;��H;�H; �H;_�H;]�H;��H;��H;��H;]�H;;�H;^�H;��H;��H;��H;a�H;a�H;��H;�H;��H;I;�I;�I;aI;� I;=+I;�7I;TFI;�VI;�iI;�~I;ّI;�I;�I;syI;79I;��H;63H;�dG;egF;�EE;pD;��B;��A;��@;�p@;      �fF;0zF;$�F;�G;_sG;��G;ZH;��H;�I;�WI;��I;�I;НI;�I;�I;BsI;�`I;yPI;�AI;�4I;I)I;>I;�I;`I;�I;�I;-�H;B�H;
�H;��H;o�H;��H;V�H;k�H;��H;M�H;Q�H;M�H;��H;k�H;T�H;��H;r�H;��H;
�H;B�H;,�H;�I;�I;`I;�I;>I;D)I;�4I;�AI;zPI;�`I;@sI;�I;�I;НI;�I;��I;�WI;�I;��H;ZH;�G;dsG;�G;#�F;%zF;      p�H;��H;^�H;3I;�%I;�HI;�hI;K�I;�I;��I;(�I;�I;1�I;�vI;]fI;�VI;�HI;E<I;�0I;n&I;MI;zI;�I;�I;{I;0�H;G�H;)�H;��H;t�H;��H;4�H;#�H;H�H;��H;Q�H;Q�H;Q�H;��H;G�H;!�H;5�H;��H;u�H;��H;*�H;E�H;-�H;I;�I;�I;zI;LI;n&I;�0I;E<I;�HI;�VI;]fI;�vI;1�I;�I;'�I;��I;�I;K�I;�hI;�HI;�%I;5I;]�H;��H;      ��I;@�I;%�I;s�I;�I;�I;f�I;c�I;��I;>�I;��I;VtI;pfI;YI;�LI;�@I;�5I;�+I;�"I;�I;�I;{I;�I;I;��H;D�H;)�H;��H;��H;��H;&�H;��H;�H;?�H;��H;��H;g�H;��H;��H;?�H;��H;��H;'�H;��H;��H;��H;)�H;D�H;��H;I;�I;}I;�I;�I;�"I;�+I;�5I;�@I;�LI;YI;pfI;VtI;�I;=�I;��I;f�I;f�I;�I;��I;u�I;%�I;L�I;      ��I;3�I;��I;ɘI;+�I;�I;��I;u�I;�vI; lI;*aI;nVI;LI;�AI;78I;/I;�&I;�I;�I;�I;�I;�I;bI;��H;�H;�H;��H;��H;��H;�H;��H;��H;��H;e�H;�H;��H;��H;��H;�H;e�H;��H;��H;��H;�H;��H;��H;��H;
�H;�H;��H;bI;�I;�I;�I;�I;�I;�&I;/I;78I;�AI; LI;mVI;(aI;�kI;�vI;u�I;��I;�I;2�I;ɘI;��I;)�I;      ^|I;�{I;�yI;�vI;LrI;�lI;dfI;Z_I;�WI;�OI;�GI;�?I;�7I;�/I;"(I;.!I;�I;�I;)I;$
I;�I;zI;��H;��H;��H;��H;t�H;��H;�H;��H;��H;��H;<�H;��H;L�H;�H;�H;�H;L�H;��H;;�H;��H;��H;��H;�H;��H;r�H;��H;��H;��H;��H;{I;�I;%
I;*I;�I;�I;-!I;"(I;�/I;�7I;�?I;�GI;�OI;�WI;]_I;dfI;�lI;IrI;�vI;�yI;�{I;      \I;�[I;ZI;�WI;]TI;.PI;aKI;FI;r@I;i:I;74I;�-I;�'I;�!I;"I;�I;{I;�I;1I;5I;� I;B�H;D�H;��H;[�H;t�H;��H;)�H;��H;��H;��H;�H;��H;�H;��H;��H;��H;��H;��H;�H;��H;�H;��H;��H;��H;*�H;��H;r�H;^�H;��H;A�H;B�H;� I;5I;1I;�I;{I;�I;"I;�!I;�'I;�-I;74I;i:I;r@I; FI;aKI;.PI;ZTI;�WI;ZI;�[I;      �CI;�CI;�BI;�@I;%>I;
;I;e7I;K3I;�.I;(*I;h%I;� I;�I;(I;�I;OI;A
I;jI;�I;}�H;��H;��H;u�H;m�H;^�H;��H;3�H; �H;��H;��H;�H;��H;��H;��H;T�H;!�H;�H;!�H;T�H;��H;��H;��H;�H;��H;��H; �H;4�H;��H;a�H;m�H;t�H;��H;��H;}�H;�I;kI;@
I;QI;�I;(I;�I;� I;h%I;)*I;�.I;K3I;d7I;;I;%>I;�@I;�BI;�CI;      G2I;2I;1I;�/I;�-I;R+I;�(I;_%I;"I;]I;�I;�I;
I;3I;�I;I;�I;�I;��H;�H;��H;Z�H;L�H;��H;��H;T�H;%�H;�H;��H;A�H;��H;��H;r�H;,�H;��H;��H;��H;��H;��H;,�H;p�H;��H;��H;B�H;��H;�H;"�H;T�H;��H;��H;J�H;Z�H;��H;�H;��H;�I;�I;I;�I;3I;	I;�I;�I;_I;"I;a%I;�(I;S+I;�-I;�/I;1I;�1I;      �%I;�%I;�$I;�#I;X"I;S I;I;�I;�I;�I;�I;�I;�I;�	I;�I;�I;� I;�H;��H;z�H;�H;}�H;��H;�H;��H;j�H;F�H;?�H;d�H;��H;�H;��H;'�H;��H;��H;~�H;b�H;~�H;��H;��H;%�H;��H;�H;��H;g�H;?�H;F�H;h�H;��H;�H;��H;}�H;}�H;z�H;��H;�H;� I;�I;�I;�	I;�I;�I;�I;�I;�I;�I;I;V I;N"I;�#I;�$I;�%I;      �I;tI;�I;�I;�I;�I;0I;I;�I;3I;�I;�
I;VI;�I;�I;� I;7�H;��H;��H;��H;��H; �H;��H;/�H;��H;��H;��H;��H;�H;L�H;��H;U�H;��H;��H;S�H;G�H;P�H;G�H;S�H;��H;��H;Y�H;��H;N�H;�H;��H;��H;��H;��H;.�H;��H; �H;��H;��H;��H;��H;6�H;� I;�I;�I;VI;�
I;�I;4I;�I;I;0I;�I;�I;�I;�I;lI;      �I;�I;I;II;2I;�I;I;(I;I;�I;�
I;?I;�I;jI;I;��H;��H;��H;��H;��H;��H;N�H;��H;��H;Y�H;H�H;P�H;��H;��H;�H;��H;"�H;��H;��H;F�H;.�H;+�H;/�H;F�H;~�H;��H;%�H;��H;�H;��H;��H;N�H;G�H;Z�H;��H;��H;N�H;��H;��H;��H;��H;��H;��H;I;hI;�I;AI;�
I;�I;I;'I;I;�I;'I;HI;I;�I;      jI;II;�I;�I;�I;eI;�I;�I;�I;�I;�	I;ZI;�I;�I;� I;K�H;'�H;�H;�H;b�H;��H;)�H;��H;C�H;9�H;K�H;N�H;k�H;��H;	�H;��H;�H;��H;f�H;N�H;-�H;�H;-�H;N�H;f�H;��H;�H;��H;�H;��H;k�H;M�H;M�H;9�H;A�H;��H;)�H;��H;b�H;�H;�H;&�H;K�H;� I;�I;�I;ZI;�	I;�I;�I;�I;�I;jI;�I;�I;�I;AI;      �I;�I;I;HI;2I;�I;I;(I;I;�I;�
I;AI;�I;hI;I;��H;��H;��H;��H;��H;��H;N�H;��H;��H;Z�H;H�H;P�H;��H;��H;�H;��H;"�H;��H;��H;F�H;.�H;+�H;/�H;F�H;~�H;��H;%�H;��H;�H;��H;��H;N�H;G�H;Y�H;��H;��H;N�H;��H;��H;��H;��H;��H;��H;I;hI;�I;AI;�
I;�I;I;'I;I;�I;'I;II;I;�I;      �I;tI;�I;�I;�I;�I;0I;I;�I;3I;�I;�
I;WI;�I;�I;� I;6�H;��H;��H;��H;��H; �H;��H;/�H;��H;��H;��H;��H;�H;L�H;��H;V�H;��H;��H;S�H;G�H;P�H;G�H;S�H;��H;��H;Y�H;��H;N�H;�H;��H;��H;��H;��H;-�H;��H; �H;��H;��H;��H;��H;6�H;� I;�I;�I;WI;�
I;�I;4I;�I;I;0I;�I;�I;�I;�I;lI;      �%I;�%I;�$I;�#I;V"I;S I;I;�I;�I;�I;�I;�I;�I;�	I;�I;�I;� I;�H;��H;z�H;��H;}�H;��H;�H;��H;j�H;F�H;?�H;d�H;��H;�H;��H;'�H;��H;��H;~�H;b�H;~�H;��H;��H;%�H;��H;�H;��H;g�H;?�H;F�H;j�H;��H;�H;��H;}�H;}�H;z�H;��H;�H;� I;�I;�I;�	I;�I;�I;�I;�I;�I;�I;I;W I;K"I;�#I;�$I;�%I;      J2I;2I;1I;�/I;�-I;R+I;�(I;_%I;"I;]I;�I;�I;	I;2I;�I;I;�I;�I;��H;�H;��H;Z�H;L�H;��H;��H;V�H;%�H;�H;��H;A�H;��H;��H;q�H;+�H;��H;��H;��H;��H;��H;+�H;p�H;��H;��H;B�H;��H;�H;"�H;S�H;��H;��H;J�H;Z�H;��H;�H;��H;�I;�I;I;�I;3I;	I;�I;�I;_I;"I;^%I;�(I;S+I;�-I;�/I;1I;2I;      �CI;�CI;�BI;�@I;'>I;
;I;h7I;L3I;�.I;)*I;h%I;� I;�I;(I;�I;QI;A
I;jI;�I;�H;��H;��H;u�H;m�H;a�H;��H;4�H; �H;��H;��H;�H;��H;��H;��H;T�H;!�H;�H;!�H;T�H;��H;��H;��H;�H;��H;��H; �H;3�H;��H;^�H;m�H;t�H;��H;��H;}�H;�I;kI;@
I;OI;�I;(I;�I;� I;h%I;)*I;�.I;L3I;h7I;;I;%>I;�@I;�BI;�CI;      \I;�[I;ZI;�WI;^TI;.PI;aKI;FI;r@I;g:I;84I;�-I;�'I;�!I;"I;�I;{I;�I;1I;5I;� I;B�H;D�H;��H;^�H;t�H;��H;*�H;��H;��H;��H;�H;��H;�H;��H;��H;��H;��H;��H;�H;��H;�H;��H;��H;��H;)�H;��H;q�H;[�H;��H;A�H;B�H;� I;5I;1I;�I;zI;�I;"I;�!I;�'I;�-I;54I;j:I;r@I; FI;aKI;.PI;[TI;�WI;ZI;�[I;      X|I;�{I;�yI;�vI;HrI;�lI;dfI;Z_I;�WI;�OI;�GI;�?I;�7I;�/I; (I;-!I;�I;�I;*I;'
I;�I;{I;��H;��H;��H;��H;t�H;��H;�H;��H;��H;��H;<�H;��H;L�H;�H;�H;�H;L�H;��H;<�H;��H;��H;��H;�H;��H;r�H;��H;��H;��H;��H;zI;�I;$
I;)I;�I;�I;/!I;"(I;�/I;�7I;�?I;�GI;�OI;�WI;^_I;ffI;�lI;IrI;�vI;�yI;�{I;      ��I;0�I;��I;ȘI;1�I;�I;��I;u�I;�vI;�kI;*aI;nVI;LI;�AI;78I;/I;�&I;�I;�I;�I;�I;�I;cI;��H;�H;�H;��H;��H;��H;�H;��H;��H;��H;e�H;�H;��H;��H;��H;�H;e�H;��H;��H;��H;�H;��H;��H;��H;
�H;�H;��H;`I;�I;�I;�I;�I;�I;�&I;/I;78I;�AI;LI;nVI;*aI;�kI;�vI;w�I;��I;�I;/�I;ØI;��I;0�I;      ��I;C�I;%�I;u�I;�I;�I;f�I;e�I;��I;=�I;��I;VtI;pfI;YI;�LI;�@I;�5I;�+I;�"I;�I;�I;}I;�I;I;��H;D�H;)�H;��H;��H;��H;'�H;��H;�H;=�H;��H;��H;g�H;��H;��H;?�H;�H;��H;&�H;��H;��H;��H;)�H;D�H;��H;I;�I;{I;�I;�I;�"I;�+I;�5I;�@I;�LI;YI;pfI;UtI;��I;>�I;��I;g�I;f�I;�I;��I;s�I;#�I;K�I;      j�H;��H;\�H;.I;�%I;�HI;�hI;K�I;�I;��I;'�I;�I;1�I;�vI;]fI;�VI;�HI;E<I;�0I;p&I;PI;zI;�I;�I;I;0�H;H�H;*�H;��H;v�H;��H;5�H;"�H;G�H;��H;Q�H;Q�H;P�H;��H;G�H;"�H;4�H;��H;r�H;��H;)�H;E�H;/�H;{I;�I;�I;zI;JI;n&I;�0I;F<I;�HI;�VI;]fI;�vI;1�I;�I;*�I;��I;�I;M�I;�hI;�HI;�%I;,I;Y�H;��H;      �fF;(zF;.�F;�G;`sG;��G;ZH;��H;�I;�WI;��I;�I;НI;�I;�I;BsI;�`I;yPI;�AI;�4I;I)I;>I;�I;aI;�I;�I;-�H;B�H;
�H;��H;r�H;��H;V�H;k�H;��H;N�H;Q�H;M�H;��H;k�H;S�H;��H;o�H;��H;
�H;B�H;,�H;�I;�I;]I;�I;>I;D)I;�4I;�AI;zPI;�`I;BsI;�I;�I;НI;�I;��I;�WI;�I;��H;ZH;�G;dsG;�G;-�F;zF;      �@@;�p@;��@;��A;��B;pD;�EE;egF;�dG;73H;��H;79I;syI;�I;�I;ۑI;�~I;�iI;�VI;TFI;�7I;=+I;� I;dI;�I;�I;�I;��H;�H; �H;a�H;`�H;��H;��H;��H;^�H;;�H;]�H;��H;��H;��H;`�H;_�H;��H;�H;��H;I;�I;�I;cI;~ I;;+I;�7I;RFI;�VI;�iI;�~I;ّI;�I;�I;uyI;69I;��H;73H;�dG;ggF;�EE;pD;��B;��A;��@;�p@;      �2;�%3;�U4;�16;֍8;U7;;��=;�@;C;�E;T�F;��G;�H;�<I;�I;țI;V�I;u�I;�pI;�[I;xII;�9I;`,I;� I;`I;cI;�I;I;��H;��H;��H;i�H;|�H;�H;*�H;��H;A�H;��H;-�H;�H;|�H;i�H;��H;��H;��H;I;�I;aI;^I;� I;],I;�9I;vII;�[I;�pI;v�I;T�I;ɛI;�I;�<I;�H;��G;S�F;~E;C;�@;��=;S7;;�8;�16;�U4;z%3;      ��;8�;�;:�;�#;�);	�.;�W4;i|9;~�=;n�A;�D;��F;�H;��H;�_I;�I;��I;��I;�uI;�^I;&KI;g:I;b,I;} I;�I;�I;�I;cI;��H;C�H;r�H;I�H;��H;��H;��H;��H;��H;��H;��H;I�H;r�H;C�H;��H;bI;�I;�I;�I;| I;],I;f:I;&KI;�^I;�uI;��I;��I;�I;�_I;��H;�H;ߟF;�D;o�A;|�=;i|9;�W4;�.;�);�#;:�;w;(�;      	��:���:��:�
�:�+�:��;�;�;��&;��/;}=7;�D=;��A;�E;�7G;��H;�8I;-�I;G�I;�I;>xI;�_I;%KI;�9I;;+I;@I;zI;}I;�I;~I;B�H;��H;Y�H;{�H;�H;N�H;(�H;L�H;�H;{�H;Y�H;��H;@�H;xI;�I;{I;vI;@I;7+I;�9I;"KI;�_I;9xI;�I;F�I;-�I;�8I;��H;�7G;�E;��A;�D=;}=7;��/;��&;�;�;��;,�:�
�:��:���:      P�x9��9h��9
:��^:� �:Wʼ:Q�:��;�h;�#;�</;�;8;��>;�oC;�fF;|(H;�I;�I;�I;�I;?xI;�^I;}II;�7I;M)I;LI;�I;�I;�I;� I;��H;��H;v�H;��H;��H;��H;��H;��H;x�H;��H;��H;� I;�I;�I;�I;JI;L)I;�7I;wII;�^I;>xI;�I;�I;�I;�I;z(H;�fF;�oC;��>;�;8;�</;�#;�h;��;Q�:Yʼ:�:��^: 
:X��9���9      ׯ����������`ct��D�`$�8��&:���:���:�Z;�C;r�&;�'3;X<;��A;!�E;��G;�I;�|I;�I;�I;�uI;�[I;NFI;�4I;p&I;�I;�I;"
I;3I;x�H;�H;v�H;��H;��H;_�H;��H;��H;v�H;�H;y�H;3I; 
I;�I;�I;j&I;�4I;MFI;�[I;�uI;�I;�I;�|I;I;��G;"�E;��A;X<;�'3;r�&;�C;�Z;���:���:��&:`$�8�D�Hct��𳺺�����      �M����D���jg��`7}�=�D�]���w��������9��:��:J	;S�;/�.;2�9;)�@;0^E;��G;�I;�I;I�I;��I;�pI;�VI;�AI;�0I;�"I;�I;,I;.I;�I;��H;��H;��H;��H;�H;��H;��H;��H;��H;�I;.I;)I;�I;�"I;�0I;�AI;�VI;�pI;��I;G�I;�I;�I;��G;0^E;)�@;2�9;0�.;Q�;J	;��:��:���9����w��[��9�D�\7}�jg��B�����      ��?��<<���1��h!��z��B�N���n��P�-��ﳺH|���&:֏�:���:��;Z�+;�8;z�@;0^E;��G;�I;-�I;��I;u�I;�iI;|PI;H<I;�+I;�I;�I;�I;jI;�I;�H;��H;��H;�H;��H;��H;�H;�I;kI;�I;�I;�I;�+I;E<I;}PI;�iI;q�I;��I;-�I;�I;��G;/^E;{�@;�8;Z�+;��;���:֏�:�&:H|���ﳺO�-��n��N���B黬z��h!���1��<<�      _��L���I��v�������^��75��z�t�̻�눻kR�Hct���x9���:�m�:i;��*;�8;+�@;%�E;|(H;�8I;�I;W�I;�~I;�`I;�HI;�5I;�&I;�I;wI;<
I;�I;� I;0�H;��H;#�H;��H;2�H;� I;�I;:
I;wI;�I;�&I;�5I;�HI;�`I;�~I;R�I;��I;�8I;z(H;%�E;+�@;�8;��*;i;�m�:���:��x9Hct�kR��눻t�̻�z��75��^����v����I��N��      '��`��
�
���Y��FC���t����|���?���	���ЗV�����@�8�:C�:i;_�+;5�9;��A;�fF;��H;�_I;̛I;ؑI;DsI;�VI;�@I;/I;-!I;�I;KI;I;�I;� I;��H;G�H;��H;� I;�I;I;KI;�I;-!I;/I;�@I;�VI;FsI;ّI;țI;�_I;��H;�fF;��A;5�9;_�+;i;C�:8�:@�����ЗV�����	���?���|��t��EC��Y��
����
�a�      ��t��p�-�d� �Q�{�9�]*����`�ҼwI���o���'��ڻ,6}�����5�0�:�m�:��;,�.;]<;�oC;�7G;��H;�I;�I;�I;_fI;�LI;:8I;(I;I;�I;�I;�I;�I;	I;� I;	I;�I;�I;�I;�I;I;(I;58I;�LI;]fI;�I;�I;�I;��H;�7G;�oC;`<;+�.;��;�m�:0�:�5����,6}��ڻ��'�	�o�wI��_�Ҽ���]*�|�9� �Q�-�d��p�      ��Ž6���̷�S���z����}��Q�T�'����$C��&\��#<<�|>�hn����� ����:���:P�;�'3;��>;�E;�H;�<I;�I;�I;�vI;YI;�AI;�/I;�!I;!I;/I;�	I;�I;aI;�I;aI;�I;�	I;-I;"I;�!I;�/I;�AI;YI;�vI;�I;�I;�<I;�H;�E;��>;�'3;P�;���:���: ����hn��|>�#<<�&\��$C�����T�'��Q���}��z��S��̷�6���      d.��3�ɤ�W����ψŽ85�����XG�1��^kּB����xC�{>�+6}����� �x9܏�:L	;v�&;�;8;��A;�F;�H;vyI;ԝI;5�I;qfI;LI;�7I;�'I;�I;	I;�I;QI;�I;�I;�I;QI;�I;I;�I;�'I;�7I; LI;pfI;1�I;םI;yyI;�H;��F;��A;�;8;v�&;L	;ޏ�:��x9����+6}�{>��xC�B���^kּ1��XG����85��ψŽ��W��ɤ��3�      Jx��s���d�O�N�a�3�}I����I����z����\�A*��ݼB���#<<��ڻЗV�Dct��&:��:�C;�</;�D=;�D;��G;59I;�I;�I;TtI;mVI;�?I;�-I;� I;�I;�I;�
I;8I;SI;8I;�
I;�I;�I;� I;�-I;�?I;kVI;TtI;�I;�I;79I;��G;�D;�D=;�</;�C;��:$�&:Hct�їV��ڻ#<<�B����ݼA*���\��z��I������}I�a�3�O�N���d��s�      .l¾(��V������������d���7�y��9Sؽ[���d�A*�_kּ&\����'���kR�P|����:�Z;�#;z=7;r�A;T�F;��H;��I;(�I;�I;-aI;�GI;34I;b%I;�I;�I;�I;�
I;�	I;�
I;�I;�I;�I;e%I;34I;�GI;*aI;�I;'�I;��I;��H;Q�F;n�A;z=7;�#;�Z;��:H|��lR�����'�&\��_kּA*��d�[��9Sؽy����7��d���������V���(��      �V������������Ͼ�d���ǆ�F�N��3��c�[����\�0��$C���o���	��눻�ﳺ���9���:�h;��/;��=;�E;93H;�WI;��I;9�I; lI;�OI;c:I;(*I;_I;�I;1I;�I;�I;�I;1I;�I;]I;(*I;d:I;�OI;�kI;9�I;��I;�WI;=3H;~E;~�=;��/;�h;���:���9�ﳺ�눻��	��o�$C��1����\�[���cི3�F�N��ǆ��d����Ͼ���������      �,b�ƽ\��>M���5�=��3r��'l¾Ꝓ�$&W��3�9Sؽ�z��XG����wI����?�t�̻Q�-�������:��;��&;g|9;
C;�dG;�I;}�I;��I;�vI;�WI;l@I;�.I;"I;�I;�I;I;�I;I;�I;�I;�!I;�.I;l@I;�WI;�vI;��I;z�I;�I;�dG;C;d|9;��&;��;���:���O�-�v�̻��?�wI�����XG��z��9Sؽ�3�$&W�Ꝓ�'l¾3r��=����5��>M�ƽ\�      ���&��\���N䂿Ľ\���1�����J˾Ꝓ�F�N�y��I������T�'�_�Ҽ��|��z��n���w����&:Q�:�;�W4;�@;hgF;��H;M�I;`�I;u�I;W_I;FI;H3I;^%I;�I; I; I;�I;!I;�I;�I;^%I;H3I;FI;W_I;r�I;`�I;K�I;��H;kgF;�@;�W4;�;Q�:��&:�w���n���z���|�_�ҼT�'����I���y��F�N�Ꝓ��J˾�����1�Ľ\�N䂿\���&��      !}߿�$ڿ0�ʿ����
����Ps�RX:����'l¾�ǆ���7����85���Q�����t���75�N��b���$�8Mʼ:��;�.;��=;�EE;ZH;�hI;f�I;��I;bfI;\KI;e7I;�(I;I;/I; I;�I; I;/I;I;�(I;e7I;]KI;bfI;��I;f�I;�hI;ZH;�EE;��=; �.;��;Sʼ:�$�8b��L���75��t������Q�85�������7��ǆ�'l¾���RX:��Ps�
�������0�ʿ�$ڿ      {�����p������ſ&���Ps���1�3r���d���d�}I�ψŽ��}�]*�EC���^��B�@�D��D�� �:��;�);Q7;;mD;��G;�HI;�I;�I;�lI;1PI;
;I;V+I;[ I;�I;�I;kI;�I;�I;[ I;S+I;;I;1PI;�lI;�I;�I;�HI;��G;oD;L7;;�);��; �:�D�@�D��B��^�FC��]*���}�ψŽ}I��d��d��3r����1��Ps�&����ſ��꿄p����      ��7��3�آ%�{��<����ſ
���Ľ\�=����Ͼ����a�3��轻z��{�9�Y�ἔ���z�_7}�hct���^:�+�:�#;ڍ8;��B;bsG;�%I;�I;2�I;?rI;STI;$>I;�-I;Q"I;�I;$I;�I;$I;�I;O"I;�-I;%>I;STI;>rI;/�I;�I;�%I;`sG;��B;֍8;��#;�+�:��^:hct�_7}��z����Y��{�9��z����a�3�������Ͼ=��Ľ\�
�����ſ�<��{�آ%��3�      /�_��+Y��lG�f.�{���꿲���O䂿��5���󾏰��O�N�W��S���Q����v����h!�kg����$
:�
�:A�;�16;��A;�G;.I;y�I;ƘI;�vI;�WI;�@I;�/I;�#I;�I;HI;�I;HI;�I;�#I;�/I;�@I;�WI;�vI;ØI;y�I;.I;�G;��A;�16;D�;�
�:0
:��kg���h!�v������ �Q�S��W��O�N���������5�O䂿�������{�f.��lG��+Y�      Ҭ��%}�?tf��lG�آ%��p�0�ʿ\����>M����V�����d�ɤ�̷�-�d��
�I����1�H��������9���:p;�U4;��@;0�F;^�H; �I;��I;�yI;�YI;�BI;1I;�$I;�I;I;�I;I;�I;�$I;1I;�BI;�YI;�yI;��I; �I;^�H;0�F;��@;�U4;s;���: ��9���H�����1��I���
�-�d�̷�ɤ���d�V�������>M�\���0�ʿ�p�آ%��lG�?tf�%}�      T���E���%}��+Y��3�����$ڿ&��ƽ\����(���s��3�6����p�a�N���<<������ؘ�9���:'�;w%3;�p@;zF;��H;=�I;6�I;�{I;�[I;�CI;�1I;�%I;cI;�I;DI;�I;fI;�%I;�1I;�CI;�[I;�{I;3�I;=�I;��H;zF;�p@;s%3;,�;���:ؘ�9������<<�N��a��p�6����3��s�(�����ƽ\�&���$ڿ����3��+Y�%}�E���      �Aq���i���U�H:�@�����>���w���}A�e5�� ���^Z�����A���]�����d��?",��5���Ѻ���9>��:z�;|Y4;��@;�VF;��H;�GI;�bI;LOI;\:I;*I;_I;�I;
I;�I;�I;�I;
I;�I;]I;*I;\:I;KOI;�bI;�GI;��H;�VF;��@;zY4;}�;>��:���9�Ѻ�5��>",��d������]��A������^Z�� ��e5�}A�w���>�������@�H:���U���i�      ��i���b�\�O�.5�3i�������������q<����f��b
V�HE	�!���IY�h9�>�����(��R��l�Ⱥ��:���:<�;b�4;��@;�hF;ؗH;QII;�bI;�NI;�9I;�)I;'I;�I;�I;�I;�I;�I;�I;�I;%I;�)I;�9I;�NI;�bI;QII;ؗH;�hF;��@;^�4;B�;���:��:p�Ⱥ�R����(�?���h9��IY�!��HE	�b
V�f������q<������������3i�.5�\�O���b�      ��U�\�O�J-?�/�'���O�῵欿b�{�ga/���뾞���I����d���ZN�Z5������0H�H ��҈��$�":��:��;��5;�`A;��F;u�H;WMI;7bI;�MI;�8I; )I;I;$I;I;EI;GI;EI;}I;$I;~I;!)I;�8I;�MI;5bI;WMI;u�H;��F;�`A;��5;��;��:$�":ֈ��H ��0H�����Z5���ZN�d������I�������ga/�b�{��欿O����/�'�J-?�\�O�      H:�.5�/�'��������lȿ���n$_���Y�Ҿݕ���6�����*���`=�8�漨)��=G�6������Q:5�:/0";2�7;�&B;,�F;��H;,SI;�`I;�KI;^7I;�'I;|I;XI;�I;�I;�
I;�I;�I;XI;yI;�'I;^7I;�KI;�`I;,SI;��H;+�F;�&B;-�7;00";3�:��Q: ��6��<G��)��8���`=��*������6�ݕ��Y�Ҿ��n$_����lȿ�������/�'�.5�      @�3i�������K�ѿl������q<��:��a����q����Wн罅���'�Qb̼�zl��.���X�(��F�:��; �&;�9;jC;�MG;�H;yYI;�^I;�HI;$5I;&I;"I;HI;�I;�
I;�	I;�
I;�I;HI;!I;&I;#5I;�HI;�^I;yYI;�H;�MG;fC;�9;#�&;��;F�:0���X��.���zl�Qb̼��'�罅��Wн����q��a���:��q<���l���K�ѿ������3i�      �������O��lȿl���������O���|]׾|����I�����A��>�d�l�y֮��QH��jλ�$��#�ӱ�:�N;�+;<;?4D; �G;�I;�^I;�[I;#EI;c2I;�#I;�I;�I;�I;�	I;�I;�	I;�I;�I;�I;�#I;c2I; EI;�[I;�^I;�I;��G;<4D;<;�+;�N;ױ�: $��$��jλ RH�y֮�l�=�d��A������I�|���|]׾����O�����l���lȿO�Ῥ��      >��������欿�������O��x����� ���l���"��ܽ���`=����q���k"�R���ۺ��9�?�:�L;Ϲ0;�>;�ME;�#H;&I;bI;GWI;�@I;4/I;�!I;{I;CI;LI;�I;�I;�I;LI;BI;{I;�!I;4/I;�@I;CWI;bI;&I;�#H;�ME;�>;͹0;�L;�?�:�9�ۺR���k"�q������`=����ܽ��"��l�� ����뾂x���O�������欿����      w�������b�{�n$_��q<������~��	w���6�����!���h����޷��x d�b.��_^e�H[���Z:υ�:�, ;��5;�A;WF;�H;!AI;�bI;�QI;,<I;�+I;�I;LI;xI;�	I;*I;nI;*I;�	I;xI;JI;�I;�+I;,<I;�QI;�bI;AI;�H;WF;�A;��5;�, ;υ�:��Z:H[�^^e�b.��x d�޷������h�!�������6�	w��~��������q<�n$_�b�{�����      }A��q<�ga/����:�|]׾� ��	w��>�EE	�����ڽ����3�Z�꼓���",��W��%����P�	��:�M
;�f);��:;`@C;7@G;��H;�TI;
`I;jKI;!7I;�'I;�I;�I;}I;I;�I;�I;�I;I;}I;�I;�I;�'I;!7I;gKI;
`I;�TI;��H;4@G;]@C;��:;�f);�M
;��:��P�#���W��",�����Z�꼘�3�ڽ������EE	�>�	w��� ��|]׾�:���ga/��q<�      e5�������Y�Ҿ�a��|����l��6�EE	���Ƚk���aG����`֮��W�{��0�k�����d,:��:8�;Փ1;��>;wE;h�G;cI;c_I;�ZI;zDI;�1I;r#I;�I;8I;D
I;KI;I;^I;I;KI;D
I;7I;�I;q#I;�1I;wDI;�ZI;b_I;cI;f�G;uE;��>;ԓ1;8�;��:�d,:���2�k�{���W�`֮�����aG�k����ȽEE	��6��l�|����a��Y�Ҿ������      � ��f�����ݕ����q��I���"���������k���ZN�Y�¼C�y��$��Q��M� � |W�B�:c0;e�&;#x8;� B;ǛF;�H;�@I;4bI;�RI;\=I;Q,I;I;&I;�I;I;wI;[I;�I;[I;wI;I;�I;(I;I;Q,I;X=I;�RI;2bI;�@I;�H;F;� B;"x8;d�&;b0;B�: pW�N� ��Q���$�C�y�¼Y��ZN�k������������"��I���q�ݕ�����f��      �^Z�b
V��I��6�������ܽ!��ڽ���aG�Y��ȼ|)��q�(�L��G5������Z:��:TS;J'1;�=;�D;l�G;1�H;YI;Z^I;�II;76I;�&I;�I;�I;�
I;�I;�I;� I;��H;� I;�I;�I;�
I;�I;�I;�&I;66I;�II;W^I;YI;.�H;j�G;�D;�=;J'1;RS;��:��Z:���G5�L��p�(�|)���ȼY��aG�ڽ��!���ܽ������6��I�b
V�      ���HE	��������Wн�A�����h���3����¼|)��$x/���һ7�X��"����9���:�>;yf);�`9;�&B;��F;�}H;7I;�aI;�UI;�@I;/I;<!I;�I;dI;"I;�I;� I;��H;<�H;��H;� I;�I;"I;fI;�I;<!I;/I;�@I;�UI;�aI;7I;�}H;�F;�&B;�`9;wf);�>;���:��9�"��9�X���һ$x/�|)��¼�����3��h��󑽢A���Wн��콻��HE	�      �A��!��d���*��罅�=�d��`=����Z��`֮�B�y�p�(���һb]e�t���0�f9'��:q�;�1";`�4;�m?;E;��G;��H;�WI;�^I;JKI;�7I;4(I;�I;gI;�
I;bI;^I;��H;�H;}�H;�H;��H;\I;bI;�
I;gI;�I;3(I;�7I;IKI;�^I;�WI;��H;��G;E;�m?;`�4;�1";s�;%��:0�f9r���b]e���һp�(�C�y�`֮�Z�꼗���`=�=�d�罅��*��d��!��      �]��IY��ZN��`=���'�l����߷�������W��$�L��:�X�|����9���:���:��;�0;!�<;��C;cG;>�H;@I;maI;UI;~@I;P/I;�!I;�I;QI;�I;�I;"�H;��H;L�H;��H;L�H;��H;#�H;�I;�I;QI;�I;�!I;P/I;}@I;UI;laI;@I;9�H;cG;��C;"�<;�0;��;���:���:�9z���:�X�L���$��W�����߷�����l���'��`=��ZN��IY�      ���h9�X5��8��Qb̼y֮�p��x d� ",�|���Q��G5�#���f9���:	�:N�;
�-;��:;"LB;|VF;XKH; I;]I;f\I;�HI;G6I;`'I;]I;�I;[
I;�I;< I;�H;��H;��H;+�H;��H;��H;�H;; I;�I;[
I;�I;YI;`'I;D6I;�HI;d\I;]I;I;YKH;zVF;"LB;��:;�-;M�;	�:���:0�f9#��G5��Q��|�� ",�x d�p��x֮�Qb̼8��X5��h9�      �d��=��������)���zl��QH��k"�b.���W��0�k�N� ������9#��:���:K�;�-;�9;�aA;��E;h�G;��H;FSI;W`I;+PI;�<I;�,I;�I;tI;NI;�I;�I;��H;��H;�H;��H;��H;��H;�H;��H;��H;�I;�I;NI;qI;�I;�,I;�<I;+PI;R`I;ASI;��H;g�G;��E;�aA;
�9;�-;J�;���:%��:��9���N� �0�k��W��b.���k"��QH��zl��)������?���      @",���(�/H�<G��.���jλR��b^e�&����� xW�x�Z:���:o�;��;�-;�9;�A;dE;e�G;��H;�GI;9aI;�UI;�BI;�1I;-$I;I;-I;�I;4I;��H;��H;�H;I�H;U�H;(�H;U�H;I�H;�H;��H;��H;4I;�I;*I;I;)$I;�1I;�BI;�UI;6aI;�GI;��H;g�G;dE;�A;�9;�-;��;p�;���:|�Z: xW����#��c^e�R���jλ�.��<G�/H���(�      �5���R��D ��
6���X��$��ۺH[���P��d,:B�:��:�>;�1";�0;��:;�aA;dE;6�G;��H;	>I;n`I;�YI;1GI;"6I;�'I;0I;�I;;I;�I; I;C�H;a�H;6�H;��H;��H;��H;��H;��H;6�H;_�H;E�H; I;�I;9I;�I;-I;�'I;$6I;/GI;�YI;p`I;>I;��H;7�G;dE;�aA;��:;�0;�1";�>;��:B�:�d,:��P�H[��ۺ�$��X�
6��D ���R��      �ѺJ�Ⱥ̈�� ��8��@$����9��Z:��:��:`0;NS;sf);Y�4;�<;LB;��E;a�G;��H;�:I;�_I;�[I;dJI;F9I;�*I; I;6I;@I;�I;PI;*�H;��H;P�H;m�H;8�H;q�H;(�H;t�H;8�H;m�H;P�H;��H;+�H;MI;�I;@I;4I;I;�*I;B9I;cJI;�[I;�_I;�:I;��H;d�G;��E;LB;�<;Z�4;sf);NS;`0;��:��:��Z:���9$��� ��ʈ��^�Ⱥ      ���9<�:4�":��Q:6�:۱�:�?�:ǅ�:�M
;5�;d�&;E'1;�`9;�m?;��C;xVF;h�G;��H;>I;�_I;T\I;�KI;W;I;-I;!I;3I;�I;'I;�I;�H;u�H;��H;w�H;��H;��H;�H;��H;�H;��H;��H;v�H;��H;u�H;�H;�I;'I;�I;2I;!I;-I;V;I;�KI;Q\I;�_I;	>I;��H;g�G;zVF;��C;�m?;�`9;G'1;a�&;4�;�M
;˅�:�?�:ᱩ:8�:��Q:<�":��:      N��:���:�:!�:��;�N;�L;�, ;�f);ӓ1;&x8;�=;�&B;E;cG;VKH;��H;�GI;n`I;�[I;�KI;�;I;..I;q"I;vI;WI;\	I;�I;��H;-�H;�H;��H;��H;\�H;�H;��H;��H;��H;�H;\�H;��H;��H;�H;)�H;��H;�I;X	I;WI;yI;n"I;,.I;�;I;�KI;�[I;n`I;�GI;��H;UKH;eG;E;�&B;�=;#x8;ԓ1;�f);�, ;�L;�N;��;!�:�:���:      }�;@�;��;(0";�&;�+;й0;��5;��:;��>;� B;�D;�F;��G;=�H;I;BSI;7aI;�YI;dJI;V;I;0.I;�"I;BI;I;=
I;nI;��H;��H;��H;��H;��H;:�H;�H;1�H;��H;��H;��H;3�H;�H;9�H;��H;��H;��H;��H;��H;lI;@
I;I;?I;�"I;0.I;U;I;gJI;�YI;9aI;ASI;I;=�H;��G;�F;�D;� B;��>;��:;��5;ҹ0;�+;"�&;(0";��;4�;      �Y4;u�4;�5;2�7;�9;<;�>;�A;`@C;vE;țF;l�G;�}H;��H;@I;]I;V`I;�UI;0GI;C9I;-I;p"I;?I;eI;�
I;�I;- I;)�H;��H;'�H;��H;5�H;��H;��H;�H;��H;��H;��H;�H;��H;��H;7�H;��H;%�H;��H;)�H;, I;�I;�
I;aI;@I;q"I;-I;C9I;1GI;�UI;U`I;]I;@I;��H;�}H;l�G;śF;uE;^@C;�A;�>;<;��9;1�7;�5;g�4;      ��@;��@;�`A;�&B;jC;?4D;�ME;WF;6@G;e�G;�H;1�H;7I;�WI;maI;f\I;0PI;�BI;(6I;�*I;!I;zI;I;�
I;.I;^ I;s�H;&�H;b�H; �H;@�H;��H;��H;��H;!�H;��H;��H;��H;!�H;��H;��H;��H;A�H; �H;`�H;&�H;p�H;^ I;1I;�
I;I;|I;!I;�*I;(6I;�BI;.PI;d\I;naI;�WI;7I;1�H;�H;b�G;4@G;WF;�ME;?4D;lC;�&B;�`A;��@;      �VF;�hF;�F;,�F;�MG;��G;�#H;�H;��H;_I;�@I;YI;�aI;�^I;UI;�HI;�<I;�1I;�'I;�I;0I;VI;<
I;�I;W I;��H;W�H;��H;-�H;:�H;��H;��H;�H;��H;D�H;��H;��H;��H;G�H;��H;|�H;��H;��H;9�H;-�H;��H;U�H;��H;Z I;�I;<
I;VI;,I;�I;�'I;�1I;�<I;�HI;UI;�^I;�aI;YI;�@I;\I;��H;�H;�#H;��G;�MG;+�F;�F;�hF;      ��H;חH;s�H;��H;�H;�I;&I;AI;�TI;e_I;4bI;Z^I;�UI;JKI;~@I;G6I;�,I;)$I;.I;8I;�I;[	I;lI;0 I;l�H;Z�H;��H;P�H;j�H;��H;j�H;M�H;z�H;��H;y�H;"�H;�H;#�H;w�H;��H;w�H;M�H;j�H;��H;j�H;S�H;��H;X�H;o�H;. I;lI;\	I;�I;8I;.I;*$I;�,I;F6I;~@I;JKI;�UI;Z^I;4bI;b_I;�TI;AI;&I;�I;"�H;��H;r�H;ؗH;      �GI;OII;]MI;%SI;vYI;�^I;bI;�bI;`I;�ZI;�RI;�II;�@I;�7I;P/I;^'I;�I;I;�I;BI;&I;�I;��H;,�H;!�H;��H;Q�H;F�H;��H;j�H;A�H;I�H;��H;�H;��H;�H;u�H;�H;��H;�H;��H;J�H;C�H;g�H;��H;G�H;Q�H;��H;#�H;-�H;��H;�I;%I;BI;�I;I;�I;^'I;R/I;�7I;�@I;�II;�RI;�ZI;`I;�bI;bI;�^I;�YI;&SI;]MI;\II;      cI;�bI;/bI;�`I;�^I;�[I;GWI;�QI;jKI;zDI;[=I;:6I;/I;3(I;�!I;ZI;tI;)I;:I;�I;�I;��H;��H;��H;\�H;0�H;g�H;��H;]�H;@�H;6�H;y�H;��H;j�H;�H;��H;��H;��H;�H;j�H;��H;z�H;6�H;?�H;^�H;��H;j�H;.�H;_�H;��H;��H;��H;�I;�I;=I;,I;sI;YI;�!I;4(I;/I;96I;Z=I;wDI;jKI;�QI;GWI;�[I;�^I;�`I;2bI;�bI;      VOI;�NI;�MI;�KI;�HI;'EI;�@I;.<I;(7I;�1I;Z,I;�&I;?!I;�I;�I;�I;QI;�I;�I;QI;�H;*�H;��H;)�H;�H;7�H;��H;g�H;?�H;?�H;h�H;��H;6�H;��H;��H;b�H;]�H;b�H;��H;��H;3�H;��H;h�H;=�H;=�H;k�H;��H;7�H;�H;(�H;��H;*�H;�H;PI;�I;�I;QI;�I;�I;�I;?!I;�&I;X,I;�1I;(7I;3<I;�@I;'EI;�HI;�KI;�MI;�NI;      _:I;	:I;�8I;h7I;.5I;`2I;;/I;�+I;�'I;x#I;I;�I;�I;nI;RI;_
I;�I;3I; I;.�H;{�H;�H;��H;��H;=�H;��H;g�H;D�H;5�H;k�H;��H;/�H;��H;O�H;�H;��H;��H;��H;�H;Q�H;��H;0�H;��H;i�H;6�H;D�H;h�H;��H;?�H;��H;��H;�H;x�H;.�H; I;3I;�I;_
I;TI;mI;�I;�I;I;x#I;�'I;�+I;;/I;`2I;.5I;j7I;�8I;	:I;      %*I;�)I;')I;�'I;&I;�#I;�!I;�I;�I;�I;+I;�I;gI;I;�I;�I;�I;��H;I�H;��H;��H;��H;��H;:�H;��H;��H;K�H;J�H;w�H;��H;,�H;��H;/�H;��H;��H;��H;w�H;��H;��H;��H;,�H;��H;/�H;��H;z�H;J�H;K�H;��H;��H;:�H;��H;��H;��H;��H;I�H;��H;�I;�I;�I;I;iI;�I;*I;�I;�I;�I;�!I;�#I;&I;�'I;$)I;�)I;      `I;7I;�I;�I;,I;~I;yI;PI;�I;8I;�I;�
I;%I;fI;�I;> I;��H;��H;b�H;S�H;{�H;��H;:�H;��H;��H;~�H;x�H;��H;��H;9�H;��H;2�H;��H;��H;M�H;D�H;Q�H;D�H;M�H;��H;��H;3�H;��H;:�H;��H;��H;w�H;~�H;��H;��H;9�H;��H;{�H;U�H;b�H;��H;��H;> I;�I;hI;#I;�
I;�I;:I;�I;QI;{I;�I;%I;�I;�I;0I;      �I;�I;I;`I;OI;�I;CI;I;�I;F
I;#I;�I;�I;aI;&�H;�H;��H;�H;:�H;s�H;��H;]�H;�H;��H;��H;��H;��H;�H;h�H;��H;N�H;��H;��H;\�H;!�H;	�H;��H;	�H;#�H;^�H;��H;��H;N�H;��H;k�H;�H;��H;��H;��H;��H;�H;]�H;��H;s�H;:�H;�H;��H;�H;%�H;aI;�I;�I;"I;D
I;�I;I;EI;�I;EI;`I;I;�I;      I;�I;�I;�I;�I;�I;PI;�	I;%I;NI;�I;�I;� I;��H;��H;��H;�H;E�H;��H;>�H;��H;��H;1�H;
�H;�H;B�H;s�H;��H;�H;��H;�H;��H;L�H;$�H;�H;��H;��H;��H;�H;$�H;I�H;��H;�H;��H;�H;��H;s�H;B�H;�H;�H;1�H;��H;��H;>�H;��H;H�H;�H;��H;��H;��H;� I;�I;~I;OI;%I;�	I;PI;�I;�I;�I;�I;�I;      �I;�I;LI;�I;�
I;�	I;�I;3I;�I;I;bI;� I;��H;�H;O�H;��H;��H;O�H;��H;x�H;�H;��H;��H;��H;��H;��H; �H;�H;��H;b�H;��H;��H;C�H;�H;��H;��H;��H;��H;��H;	�H;B�H;��H;��H;c�H;��H;�H; �H;��H;��H;��H;��H;��H;�H;x�H;��H;Q�H;��H;��H;O�H;�H;��H;� I;`I;I;�I;2I;�I;�	I;�
I;�I;JI;�I;      �I;�I;SI;�
I;�	I;�I;�I;rI;�I;]I;�I;��H;@�H;��H;��H;1�H;��H; �H;��H;,�H;��H;��H;��H;��H;��H;��H;�H;{�H;��H;`�H;��H;}�H;P�H;��H;��H;��H;��H;��H;��H;��H;N�H;~�H;��H;b�H;��H;{�H;�H;��H;��H;��H;��H;��H;��H;,�H;��H;!�H;��H;1�H;��H;��H;@�H;��H;�I;`I;�I;qI;�I;�I;�	I;�
I;RI;�I;      �I;�I;LI;�I;�
I;�	I;�I;3I;�I;I;bI;� I;��H;�H;O�H;��H;��H;O�H;��H;x�H; �H;��H;��H;��H;��H;��H; �H;�H;��H;b�H;��H;��H;B�H;�H;��H;��H;��H;��H;��H;	�H;B�H;��H;��H;c�H;��H;�H; �H;��H;��H;��H;��H;��H;�H;x�H;��H;Q�H;��H;��H;P�H;�H;��H;� I;bI;I;�I;2I;�I;�	I;�
I;�I;HI;�I;      I;�I;�I;�I;�I;�I;PI;�	I;%I;NI;~I;�I;� I;��H;��H;��H;�H;G�H;��H;>�H;��H;��H;1�H;	�H;�H;B�H;s�H;��H;�H;��H;�H;��H;L�H;$�H;�H;��H;��H;��H;�H;$�H;I�H;��H;�H;��H;�H;��H;s�H;B�H;�H;�H;1�H;��H;��H;>�H;��H;H�H;�H;��H;��H;��H;� I;�I;~I;OI;%I;�	I;PI;�I;�I;�I;�I;�I;      �I;�I;I;`I;NI;�I;CI;I;�I;D
I;#I;�I;�I;aI;&�H;�H;��H;�H;:�H;s�H;��H;]�H;�H;��H;��H;��H;��H;�H;h�H;��H;N�H;��H;��H;^�H;#�H;	�H;��H;	�H;!�H;\�H;��H;��H;N�H;��H;k�H;�H;��H;��H;��H;��H;�H;]�H;��H;s�H;:�H;�H;��H;�H;%�H;aI;�I;�I;#I;F
I;�I;�I;CI;�I;BI;`I;I;�I;      cI;7I;�I;�I;*I;~I;{I;PI;�I;8I;�I;�
I;#I;hI;�I;> I;��H;��H;b�H;S�H;}�H;��H;:�H;��H;��H;�H;z�H;��H;��H;9�H;��H;2�H;��H;��H;M�H;D�H;Q�H;D�H;M�H;��H;��H;5�H;��H;:�H;��H;��H;w�H;|�H;��H;��H;9�H;��H;{�H;U�H;b�H;��H;��H;> I;�I;fI;#I;�
I;�I;:I;�I;MI;yI;I;%I;�I;�I;5I;      %*I;�)I;')I;�'I;&I;�#I;�!I;�I;�I;�I;+I;�I;iI;I;�I;�I;�I;��H;I�H;��H;��H;��H;��H;:�H;��H;��H;K�H;J�H;w�H;��H;/�H;��H;.�H;��H;��H;��H;w�H;��H;��H;��H;,�H;��H;,�H;��H;z�H;J�H;K�H;��H;��H;:�H;��H;��H;��H;��H;I�H;��H;�I;�I;�I;I;iI;�I;+I;�I;�I;�I;�!I;�#I;&I;�'I;&)I;�)I;      _:I;	:I;�8I;j7I;15I;`2I;;/I;�+I;�'I;v#I;I;�I;�I;nI;TI;`
I;�I;2I; I;.�H;|�H;�H;��H;��H;?�H;��H;h�H;D�H;5�H;k�H;��H;/�H;��H;Q�H;�H;��H;��H;��H;�H;O�H;��H;0�H;��H;h�H;6�H;D�H;g�H;��H;=�H;��H;��H;�H;x�H;.�H; I;3I;�I;_
I;RI;nI;�I;�I;I;y#I;�'I;�+I;;/I;`2I;-5I;h7I;�8I;	:I;      OOI;�NI;�MI;�KI;�HI;!EI;�@I;0<I;)7I;�1I;X,I;�&I;@!I;�I;�I;�I;SI;�I;�I;SI;�H;*�H;��H;(�H;�H;9�H;��H;k�H;?�H;@�H;h�H;��H;4�H;��H;��H;b�H;]�H;b�H;��H;��H;4�H;��H;h�H;=�H;?�H;g�H;��H;6�H;�H;(�H;��H;*�H;�H;QI;�I;�I;PI;�I;�I;�I;@!I;�&I;Z,I;�1I;*7I;3<I;�@I;$EI;�HI;�KI;�MI;�NI;      	cI;�bI;5bI;�`I;�^I;�[I;JWI;�QI;iKI;wDI;[=I;:6I;/I;3(I;�!I;YI;tI;*I;=I;�I;�I;��H;��H;��H;_�H;0�H;i�H;��H;^�H;@�H;6�H;w�H;��H;j�H;�H;��H;��H;��H;�H;j�H;��H;z�H;6�H;?�H;]�H;��H;i�H;.�H;\�H;��H;��H;��H;�I;�I;:I;*I;sI;\I;�!I;3(I;/I;:6I;[=I;yDI;lKI;�QI;KWI;�[I;�^I;�`I;5bI;�bI;      �GI;RII;]MI;&SI;yYI;�^I;bI;�bI;`I;�ZI;�RI;�II;�@I;�7I;R/I;^'I;�I;I;�I;CI;*I;�I;��H;-�H;#�H;��H;Q�H;G�H;��H;k�H;C�H;I�H;��H;�H;��H;�H;u�H;�H;��H;�H;��H;J�H;A�H;g�H;��H;F�H;Q�H;��H;!�H;,�H;��H;�I;#I;BI;�I;I;�I;`'I;P/I;�7I;�@I;�II;�RI;�ZI;`I;�bI;bI;�^I;�YI;%SI;]MI;\II;      ��H;ؗH;r�H;��H;�H;�I;&I;AI;�TI;c_I;4bI;Z^I;�UI;JKI;~@I;G6I;�,I;)$I;.I;9I;�I;\	I;nI;1 I;o�H;Z�H;��H;S�H;k�H;��H;j�H;M�H;x�H;��H;w�H;#�H;�H;"�H;y�H;��H;x�H;N�H;j�H;��H;i�H;P�H;��H;Z�H;l�H;- I;kI;[	I;�I;8I;.I;*$I;�,I;F6I;~@I;JKI;�UI;Z^I;5bI;c_I;�TI;AI;&I;�I;�H;��H;n�H;ϗH;      �VF;�hF;�F;+�F;�MG;��G;�#H;�H;��H;]I;�@I;YI;�aI;�^I;UI;�HI;�<I;�1I;�'I;�I;0I;VI;<
I;�I;Z I;��H;W�H;��H;.�H;:�H;��H;��H;~�H;��H;D�H;��H;��H;��H;F�H;��H;|�H;��H;��H;7�H;,�H;��H;U�H;��H;W I;�I;<
I;VI;,I;�I;�'I;�1I;�<I;�HI;UI;�^I;�aI;YI;�@I;]I;��H;�H;�#H;��G;�MG;.�F;�F;�hF;      ��@;��@;�`A;�&B;lC;?4D;�ME;WF;4@G;d�G;�H;1�H;7I;�WI;naI;f\I;/PI;�BI;(6I;�*I;!I;|I;I;�
I;1I;^ I;r�H;&�H;c�H;"�H;A�H;��H;��H;��H; �H;��H;��H;��H;!�H;��H;��H;��H;@�H;�H;_�H;&�H;p�H;^ I;.I;�
I;I;zI;!I;�*I;(6I;�BI;.PI;f\I;naI;�WI;7I;1�H;�H;d�G;4@G;WF;�ME;?4D;jC;�&B;�`A;��@;      �Y4;q�4;�5;.�7;�9;<;�>;�A;a@C;wE;ǛF;l�G;�}H;��H;@I;]I;V`I;�UI;1GI;C9I;-I;q"I;BI;cI;�
I;�I;- I;)�H;��H;(�H;��H;6�H;��H;��H;�H;��H;��H;��H;�H;��H;��H;6�H;��H;$�H;��H;)�H;, I;�I;�
I;bI;=I;p"I;-I;C9I;0GI;�UI;U`I;]I;@I;��H;�}H;l�G;ǛF;uE;a@C;�A;�>;<;��9;.�7;
�5;e�4;      z�;N�;��;&0";�&;�+;Թ0;��5;��:;��>;� B;�D;�F;��G;=�H;I;BSI;6aI;�YI;eJI;Y;I;0.I;�"I;BI;I;?
I;oI;��H;��H;��H;��H;��H;:�H;�H;3�H;��H;��H;��H;1�H;�H;9�H;��H;��H;��H;��H;��H;kI;?
I;I;=I;�"I;0.I;R;I;eJI;�YI;9aI;BSI;I;>�H;��G;�F;�D;� B;��>;��:;��5;Թ0;�+;�&;(0";��;<�;      N��:���:�:!�:��;�N;�L;�, ;�f);ԓ1;%x8;�=;�&B;E;cG;VKH;��H;�GI;n`I;�[I;�KI;�;I;/.I;r"I;yI;VI;\	I;�I;��H;-�H;�H;��H;��H;\�H;�H;��H;��H;��H;�H;\�H;��H;��H;�H;)�H;��H;�I;X	I;WI;vI;n"I;,.I;�;I;�KI;�[I;n`I;�GI;��H;VKH;eG;E;�&B;�=;%x8;ӓ1;�f);�, ;�L;�N;��;!�:�:���:      ���9�:H�":��Q:8�:ͱ�:�?�:υ�:�M
;5�;c�&;G'1;�`9;�m?;��C;zVF;h�G;��H;	>I;�_I;S\I;�KI;W;I;-I;!I;3I;�I;'I;�I;�H;u�H;��H;w�H;��H;��H;�H;��H;�H;��H;��H;w�H;��H;u�H;�H;�I;'I;�I;3I;!I;-I;V;I;�KI;Q\I;�_I;>I;��H;g�G;xVF;��C;�m?;�`9;G'1;c�&;4�;�M
;υ�:�?�:߱�:B�:��Q:H�":�:      �ѺJ�ȺĈ��"��$��@$��9��Z:��:��:`0;NS;sf);Z�4;�<;LB;��E;c�G;��H;�:I;�_I;�[I;eJI;F9I;�*I;I;6I;@I;�I;PI;+�H;��H;R�H;m�H;8�H;u�H;(�H;r�H;8�H;m�H;O�H;��H;*�H;MI;�I;@I;4I; I;�*I;B9I;aJI;�[I;�_I;�:I;��H;c�G;��E;LB;�<;Y�4;sf);NS;_0;��:��:��Z:�9 $���"��Ȉ��d�Ⱥ      �5���R��D ��
6���X��$��ۺH[� �P��d,:B�:��:�>;�1";�0;��:;�aA;dE;7�G;��H;	>I;p`I;�YI;3GI;$6I;�'I;0I;�I;;I;�I; I;C�H;a�H;6�H;��H;��H;��H;��H;��H;6�H;_�H;E�H; I;�I;9I;�I;-I;�'I;"6I;-GI;�YI;n`I;>I;��H;6�G;dE;�aA;��:;�0;�1";�>;��:B�:�d,:��P�H[��ۺ�$��X�
6��D ���R��      @",���(�/H�<G��.���jλR��b^e�%����� xW���Z:���:o�;��;�-;�9;�A;dE;e�G;��H;�GI;9aI;�UI;�BI;�1I;-$I;I;,I;�I;4I;��H;��H;�H;I�H;U�H;(�H;U�H;K�H;�H;��H;��H;4I;�I;*I;I;*$I;�1I;�BI;�UI;6aI;�GI;��H;g�G;dE;�A;�9;�-;��;o�;���:|�Z: xW����%��b^e�R���jλ�.��<G�/H���(�      �d��=��������)���zl��QH��k"�b.���W��0�k�M� ������9%��:���:J�;�-;	�9;�aA;��E;h�G;��H;FSI;V`I;+PI;�<I;�,I;�I;tI;NI;�I;�I;��H;��H;�H;��H;��H;��H;�H;��H;��H;�I;�I;NI;qI;�I;�,I;�<I;+PI;R`I;ASI;��H;g�G;��E;�aA;
�9;�-;K�;���:#��:��9���N� �2�k��W��a.���k"��QH��zl��)������?���      ���h9�X5��8��Qb̼y֮�p��x d� ",�|���Q��G5�#���f9���:	�:N�;
�-;��:;"LB;{VF;YKH;I;]I;d\I;�HI;G6I;`'I;]I;�I;[
I;�I;< I;�H;��H;��H;+�H;��H;��H;�H;; I;�I;[
I;�I;YI;`'I;D6I;�HI;f\I;]I;I;XKH;zVF;"LB;��:;�-;M�;	�:���:�f9#��G5��Q��|�� ",�x d�p��x֮�Qb̼8��X5��h9�      �]��IY��ZN��`=���'�l����߷�������W��$�L��:�X�z����9���:���:��;�0;!�<;��C;cG;>�H;@I;laI;UI;~@I;P/I;�!I;�I;QI;�I;�I;#�H;��H;L�H;��H;L�H;��H;#�H;�I;�I;QI;�I;�!I;P/I;}@I;UI;maI;@I;9�H;cG;��C;"�<;�0;��;���:���:�9|���:�X�L���$��W�����߷�����l���'��`=��ZN��IY�      �A��!��d���*��罅�=�d��`=����Z��`֮�C�y�q�(���һd]e�r���0�f9'��:q�;�1";_�4;�m?;E;��G;��H;�WI;�^I;JKI;�7I;4(I;�I;gI;�
I;cI;^I;��H;�H;}�H;�H;��H;\I;aI;�
I;gI;�I;3(I;�7I;IKI;�^I;�WI;��H;��G;E;�m?;_�4;�1";t�;%��:0�f9t���d]e���һp�(�C�y�`֮�Z�꼗���`=�=�d�罅��*��d��!��      ���HE	��������Wн�A�����h���3����¼|)��$x/���һ9�X��"����9���:�>;wf);�`9;�&B;��F;�}H;7I;�aI;�UI;�@I;/I;<!I;�I;dI;"I;�I;� I;��H;<�H;��H;� I;�I; I;dI;�I;<!I;/I;�@I;�UI;�aI;7I;�}H;�F;�&B;�`9;wf);�>;���:��9�"��7�X���һ$x/�|)��¼�����3��h��󑽢A���Wн��콻��HE	�      �^Z�b
V��I��6�������ܽ!��ڽ���aG�Y��ȼ|)��q�(�L��G5������Z:��:RS;G'1;�=;�D;k�G;.�H;YI;Z^I;�II;76I;�&I;�I;�I;�
I;�I;�I;� I;��H;� I;�I;�I;�
I;�I;�I;�&I;66I;�II;W^I;YI;1�H;j�G;�D;�=;J'1;TS;��:��Z:���G5�L��q�(�|)���ȼY��aG�ڽ��!���ܽ������6��I�b
V�      � ��f�����ݕ����q��I���"���������k���ZN�Y�¼D�y��$��Q��M� � xW�B�:c0;c�&;"x8;� B;ǛF;�H;�@I;4bI;�RI;[=I;Q,I;I;&I;�I;I;wI;[I;�I;[I;wI;I;�I;'I;I;Q,I;Z=I;�RI;2bI;�@I;�H;ěF;� B;#x8;d�&;b0;B�: pW�N� ��Q���$�D�y�¼Y��ZN�k������������"��I���q�ݕ�����f��      e5�������Y�Ҿ�a��|����l��6�EE	���Ƚk���aG����`֮��W�{��0�k�����d,:��:6�;ԓ1;��>;wE;f�G;cI;c_I;�ZI;zDI;�1I;q#I;�I;8I;D
I;KI;I;^I;I;KI;D
I;7I;�I;r#I;�1I;wDI;�ZI;b_I;cI;h�G;vE;��>;Փ1;8�;��:�d,:���2�k�|���W�`֮�����aG�k����ȽEE	��6��l�|����a��Y�Ҿ������      }A��q<�ga/����:�}]׾� ��	w��>�EE	�����ڽ����3�Z�꼓���",��W��%����P�	��:�M
;�f);��:;`@C;4@G;��H;�TI;
`I;jKI;7I;�'I;�I;�I;}I;I;�I;�I;�I;I;}I;�I;�I;�'I;!7I;gKI;
`I;�TI;��H;7@G;]@C;��:;�f);�M
;��:��P�#���W��",�����Z�꼘�3�ڽ������EE	�>�	w��� ��|]׾�:���ga/��q<�      w�������b�{�n$_��q<������~��	w���6�����!���h����޷��x d�a.��_^e�H[���Z:˅�:�, ;��5;�A;WF;�H;AI;�bI;�QI;,<I;�+I;�I;LI;zI;�	I;*I;nI;,I;�	I;zI;JI;�I;�+I;,<I;�QI;�bI;AI;�H;WF;�A;��5;�, ;Ӆ�:��Z:H[�^^e�b.��x d�޷������h�!�������6�	w��~��������q<�n$_�b�{�����      >��������欿�������O��x����� ���l���"��ܽ���`=����q���k"�R���ۺ���9�?�:�L;Ϲ0;�>;�ME;�#H;&I;bI;EWI;�@I;4/I;!I;|I;CI;LI;�I;�I;�I;LI;CI;yI;�!I;4/I;�@I;GWI;bI;&I;�#H;�ME;�>;͹0;�L;�?�:�9�ۺR���k"�q������`=����ܽ��"��l�� ����뾂x���O�������欿����      �������O��lȿl���������O���|]׾|����I�����A��>�d�l�y֮��QH��jλ�$� $�ͱ�:�N;�+;<;<4D; �G;�I;�^I;�[I;#EI;c2I;�#I;�I;�I;�I;�	I;�I;�	I;�I;�I;I;�#I;c2I; EI;�[I;�^I;�I;��G;?4D;<;�+;�N;ױ�:$��$��jλ RH�y֮�l�>�d��A������I�|���|]׾����O�����l���lȿO�Ῥ��      @�3i�������K�ѿl������q<��:��a����q����Wн罅���'�Qb̼�zl��.���X�0��B�:��; �&;�9;fC;�MG;�H;yYI;�^I;�HI;#5I;&I;"I;HI;�I;�
I;�	I;�
I;�I;HI;!I;&I;$5I;�HI;�^I;yYI;�H;�MG;jC;�9;#�&;��;J�:0���X��.���zl�Qb̼��'�罅��Wн����q��a���:��q<���l���K�ѿ������3i�      H:�.5�/�'��������lȿ���n$_���Y�Ҿݕ���6�����*���`=�8�漨)��<G�6������Q:3�:-0";1�7;�&B;,�F;��H;,SI;�`I;�KI;^7I;�'I;zI;XI;�I;�I;�
I;�I;�I;XI;zI;�'I;^7I;�KI;�`I;,SI;��H;,�F;�&B;.�7;20";5�:��Q: ��6��<G��)��8���`=��*������6�ݕ��Y�Ҿ��n$_����lȿ�������/�'�.5�      ��U�\�O�J-?�/�'���N�῵欿b�{�ga/���뾞���I����d���ZN�Z5������0H�H ��ֈ�� �":��:��;��5;�`A;��F;u�H;WMI;6bI;�MI;�8I;!)I;I;$I;I;EI;GI;EI;I;$I;~I; )I;�8I;�MI;5bI;WMI;u�H;�F;�`A;��5;��;��:$�":ֈ��I ��0H�����Z5���ZN�d������I�������ga/�b�{��欿N����/�'�J-?�\�O�      ��i���b�\�O�.5�3i�������������q<����f��b
V�HE	�!���IY�h9�>�����(��R��l�Ⱥ��:���:<�;b�4;��@;�hF;ؗH;QII;�bI;�NI;�9I;�)I;'I;�I;�I;�I;�I;�I;�I;�I;%I;�)I;�9I;�NI;�bI;QII;חH;�hF;��@;`�4;B�;���:��:p�Ⱥ�R����(�?���h9��IY�!��HE	�b
V�f������q<������������3i�.5�\�O���b�      �>���8���*�O������˿p��G�b�E\�6m־^��S�:��J�)��F�B�:��}������/������t�>:�t�:lp ;�J6;%EA;�IF;�NH;!�H;"I;�I;.I;�I;�I;I;� I;��H;H�H;��H;� I;I;�I;�I;.I;�I;"I;!�H;�NH;�IF;%EA;�J6;op ;�t�:x�>:����/�����~���:��F�B�)���J�S�:�^��6m־E\�G�b�p���˿����O���*���8�      ��8��4��g&�7��>����<ƿ򲗿�>]�î�R�Ѿ�p���*7����&W��MR?��|�l8�������:����G:� �:!;/�6;:lA;�YF;�TH;��H;8"I;�I;
I;�I;dI;I;� I;��H;0�H;��H;� I;I;cI;�I;
I;�I;5"I;��H;�TH;�YF;:lA;,�6;!;� �:�G:>��������l8���|�MR?�&W�����*7��p��R�Ѿî��>]�򲗿�<ƿ>���7���g&��4�      ��*��g&��#�v�W[�rL�������M�s5��>ľ����,��D�꒐��5�/�ݼ���q
���x��sk�d�b:�l�:&#;�7;��A;�F;�dH;�I;w"I;I;�I;]I;I;�I;> I;��H;��H;��H;< I;�I;I;]I;�I;I;t"I;�I;�dH;�F;��A;�7;(#;�l�:d�b:�sk���x��q
���/�ݼ�5�꒐��DὫ�,����>ľs5���M����rL��W[�v��#��g&�      O�7��v����˿B1��9�y�Ŏ6��z �����3�l�+��ͽ$�����&���˼6�k������X�Ԙ �Ƶ�:k�;2&;�9;��B;/�F;�}H;
I;�"I;LI;�I;�I;�I;fI;��H;C�H;��H;C�H;��H;fI;�I;�I;�I;KI;�"I;
I;�}H;/�F;��B;�9;4&;k�;ȵ�:�� ���X����6�k���˼��&�$����ͽ+�3�l������z �Ŏ6�9�y�B1���˿���v�7��      ����>���W[忷˿�T���}�R�®��E۾ԗ����M���	������j��3�d����O�$�׻}�/�������:� 
;/*;z;;kC;�'G;�H;I;$"I;I;�I;�
I;�I;�I;d�H;��H;�H;��H;c�H;�I;�I;�
I;�I;I;""I;I;�H;�'G;kC;w;;2*;� 
;���:��|�/�$�׻��O�d���3���j������	���M�ԗ���E۾®�}�R���T���˿W[�>���      �˿�<ƿrL��B1����>]���)�%��ֳ���{���,�s��(��Q`I��J���,���3/��+��� ��169
5�:	�;!p.;@.=;�aD;�G;��H;I;^!I;yI;lI;�	I;�I;	I;��H;1�H;��H;1�H;��H;	I;�I;�	I;kI;vI;Y!I;I;��H;	�G;�aD;<.=;p.;	�;5�:p169� ��+���3/��,���J��Q`I�(��s�齥�,���{�ֳ�%����)��>]��B1��rL���<ƿ      p��򲗿���9�y�}�R���)�ov��>ľ^���I�Yl����������&�ѮҼ�}�%B�����������!:G+�:[z;�3;{j?;�\E;�G;��H;�I;�I;�I;�I;�I;�I;: I;��H;��H;��H;��H;��H;: I;�I;�I;�I;�I;�I;�I;��H;�G;�\E;wj?;�3;Zz;G+�:��!:��������%B��}�ѮҼ��&��������Yl��I�^���>ľov���)�}�R�9�y����򲗿      G�b��>]���M�Ŏ6�®�%���>ľ$q��{�Z�+�S9ݽ!W����L����F����G��׻�;�xm�Ɋ:�i;=P$;��7;��A;/JF;RCH;	�H;� I;�I;�I;6I;KI;�I;7�H;�H;��H;/�H;��H;�H;7�H;�I;LI;6I;�I;�I;� I;�H;PCH;.JF;��A;��7;;P$;�i;Ɋ:�m��;��׻��G�F�������L�!W��S9ݽ+�{�Z�$q���>ľ%��®�Ŏ6���M��>]�      E\�î�s5��z ��E۾ֳ�^��{�Z�M?#����A����j�$��Aϼ����������~lۺ0;�9�4�:w�;��,;��;;U�C;�G;m�H;�I;�!I;�I;]I;GI;�I;^I;<�H;%�H;��H;@�H;��H;#�H;<�H;^I;�I;EI;\I;�I;�!I;�I;l�H;�G;T�C;��;;~�,;x�;�4�:0;�9zlۺ����������Aϼ$����j��A�����M?#�{�Z�^��ֳ��E۾�z �s5�î�      6m־R�Ѿ�>ľ����ԗ����{��I�+�����V���{�>�/�"���,��4=�.�һ4�@�h� ���k:M�:,b;��3;Rj?;�2E;�G;��H;PI;� I;�I;�I;?	I;I;  I;�H;�H;��H;v�H;��H;�H;�H;��H;I;?	I;�I;�I;� I;NI;��H;�G;�2E;Pj?;��3;,b;K�:��k:d� �6�@�.�һ4=��,��"��>�/��{��V�����+��I���{�ԗ�������>ľR�Ѿ      ^���p����3�l���M���,�Yl�S9ݽ�A���{���5��J��;���T[�?������O���Q�9�:��;H*;B�9;|kB;��F;�NH;��H;; I;�I;�I;;I;-I;]I;�H;��H;��H;��H;��H;��H;��H;��H;~�H;`I;*I;;I;�I;�I;9 I;��H;�NH;�F;ykB;B�9;F*;��;�:�Q�9�O������?��T[�;���J����5��{��A��S9ݽYl���,���M�3�l����p��      S�:��*7���,�+���	�s�齃���!W����j�>�/��J���I����k�a��-��2��`���4Ɋ:�o�:5;}r3;@�>;K�D;��G;i�H;*I;J!I;�I;�I;�
I;I;~ I;��H;��H;��H;��H;��H;��H;��H;��H;��H;� I;I;�
I;�I;�I;H!I;(I;g�H;��G;H�D;?�>;}r3;4;�o�::Ɋ:p���2���-��a���k��I���J��>�/���j�!W������s�齃�	�+���,��*7�      �J�����D��ͽ���(�������L�$��#��;����k����TI����/��/��>:���:�B;��,;��:;O�B;�xF;�<H;�H;'I;�I;I;bI;�I;�I;��H;��H;W�H;��H;��H;��H;��H;��H;W�H;��H;��H;�I;�I;_I;I;�I;&I;�H;�<H;�xF;M�B;��:;��,;�B;���:�>:�/���/�TI�������k�;��"��$����L����(������ͽ�D����      )��%W��钐�$�����j�P`I���&����Aϼ�,���T[�a�TI��1;��mk�L:f5�:�;*&;��6;�!@;V2E;��G;��H;I;!I;nI;/I;I;WI;� I;��H;%�H;��H;��H;��H;h�H;��H;��H;��H;%�H;��H;� I;XI;I;.I;mI;!I;I;��H;�G;V2E;�!@;��6;*&;�;d5�:L:�mk�0;�TI��a��T[��,��Aϼ�����&�P`I���j�$���钐�%W��      F�B�MR?��5���&��3��J��ѮҼF�����5=�?��-����/��mk����9�׳:��;U!;z3;�=;��C;@�F;4dH;�H;�I;0I;�I;CI;�I;�I;d�H;�H;��H;��H;b�H;��H;Z�H;��H;c�H;��H;��H;"�H;d�H;�I;�I;CI;�I;0I;�I;�H;/dH;?�F;��C;�=;z3;X!;��;�׳:���9�mk���/��-��?�5=����F��ѮҼ�J���3���&��5�MR?�      :���|�.�ݼ��˼d���,����}���G����.�һ����2���/�H:�׳:&�;�b;ӣ0;�<;ˮB;�IF;�H;H�H;�I;� I;;I;XI;{
I;�I;A I;O�H;s�H;,�H;G�H;B�H;��H;\�H;��H;B�H;F�H;*�H;t�H;O�H;A I;�I;{
I;UI;9I;� I;�I;C�H;�H;�IF;ɮB;�<;գ0;�b;'�;�׳:L:�/�2������.�һ�����G���}��,��d����˼.�ݼ�|�      ~���k8����6�k���O��3/�$B��׻����4�@��O��p����>:d5�:��;�b;��/;M;;]�A;��E;�G;�H;�
I;� I;I;I; I;�I;�I;��H;]�H;��H;��H;�H;6�H;��H;T�H;��H;6�H; �H;��H;��H;]�H;��H;�I;�I;�I;I;I;� I;�
I;�H;�G;��E;^�A;P;;��/;�b;��;d5�:�>:`����O��4�@������׻$B��3/���O�6�k���l8��      ������q
����&�׻�+�������;�~lۺt� ��Q�90Ɋ:���:�;U!;ѣ0;N;;ߓA;�pE;��G;�H;�H;�I;YI;xI;DI;�I;�I;#�H;d�H;��H;%�H;B�H;�H; �H;��H;^�H;��H; �H;�H;A�H;'�H;��H;c�H;�H;�I;�I;DI;xI;UI;�I;�H;�H;��G;�pE;�A;M;;ѣ0;U!;�;���:0Ɋ:�Q�9p� �xlۺ�;������+��#�׻����q
���      /�������x���X���/�� ������m�@;�9x�k:�:�o�:�B;*&;z3;�<;]�A;�pE;�tG;}H;L�H;KI;�I;eI;I;�
I;I;s I;r�H;F�H;��H;��H;��H;��H;	�H;��H;��H;��H;	�H;��H;��H;��H;��H;C�H;n�H;s I;I;�
I;I;aI;�I;KI;J�H;}H;�tG;�pE;\�A;�<;~3;*&;�B;�o�:�:x�k:H;�9�m침���ۺ ��/���X���x����      ��������sk�ؘ � ��P169��!: Ɋ:�4�:I�:��;1;��,;�6;�=;®B;��E;��G;}H;��H;�I;5 I;�I;|I;�I;KI;�I;j�H;�H;^�H;�H;3�H;��H;��H;�H;��H;��H;��H;�H;��H;��H;4�H;�H;]�H;�H;j�H;�I;JI;�I;xI;�I;5 I;�I;��H;}H;��G;��E;ĮB;�=;�6;��,;1;��;I�:�4�: Ɋ:��!:p169���ؘ ��sk�0���      ��>:X�G:p�b:���:���:5�:G+�:�i;u�;*b;F*;yr3;��:;�!@;��C;�IF;�G;�H;K�H;�I;? I;eI;]I;�I;6I;�I;C�H;��H;��H;��H;m�H;��H;��H;��H;6�H;��H;��H;��H;6�H;��H;��H;��H;m�H;��H;��H;��H;@�H;�I;6I;�I;\I;eI;< I;�I;L�H;��H;�G;�IF;��C;�!@;��:;zr3;D*;(b;w�;�i;G+�:5�:���:���:|�b:�G:      �t�:�:�l�:a�;� 
;�;_z;BP$;��,;��3;E�9;@�>;M�B;V2E;@�F;�H;�H;�H;KI;5 I;dI;�I;[I;�I;I;��H;E�H;p�H;��H;��H;�H;��H;��H;��H;Y�H;�H;��H;�H;Y�H;��H;��H;��H;�H;��H;��H;r�H;D�H;��H;I;�I;ZI;�I;bI;8 I;KI;	�H;�H;�H;A�F;V2E;M�B;@�>;D�9;��3;��,;AP$;az;�;� 
;a�;�l�:	�:      np ;	!;$#;*&;%*;p.;�3;�7;��;;Pj?;|kB;K�D;�xF;��G;1dH;C�H;�
I;�I;�I;�I;]I;\I;I;{I;W�H;��H;��H;K�H;�H;7�H;��H;��H;��H;�H;w�H;=�H;(�H;=�H;w�H;�H;��H;��H;��H;5�H;�H;K�H;��H;��H;Y�H;xI;I;^I;YI;�I;�I;�I;�
I;A�H;3dH;��G;�xF;K�D;{kB;Nj?;��;;�7;�3;!p.;/*;*&;(#;�!;      �J6;A�6;�7;�9;z;;<.=;�j?;��A;V�C;�2E;��F;��G;�<H;��H;�H;�I;� I;YI;dI;zI;�I;�I;yI;o�H;��H;��H;��H;Q�H;_�H;��H;��H;��H;��H;J�H;��H;��H;l�H;��H;��H;J�H;��H;��H;��H;��H;]�H;Q�H;��H;��H;��H;m�H;xI;�I;�I;{I;dI;ZI;� I;�I;�H;��H;�<H;��G;�F;�2E;V�C;��A;�j?;=.=;�;;�9;�7;2�6;      -EA;ElA;��A;��B;kC;�aD;�\E;+JF;�G;�G;�NH;i�H;�H;I;�I;� I;%I;xI;I;�I;9I;I;Z�H;��H;�H;��H;Z�H;m�H;��H;��H;��H;��H;��H;��H;�H;��H;��H;��H;�H;��H;��H;��H;��H;��H;��H;n�H;W�H;��H;�H;��H;\�H;I;7I;�I;I;|I;"I;� I;�I;I;�H;k�H;�NH;��G;�G;-JF;�\E;�aD;kC;��B;��A;ElA;      �IF;�YF;��F;-�F;�'G; �G;�G;ICH;g�H;��H;��H;(I;!I;!I;-I;8I;I;@I;�
I;HI;~I;��H;��H;��H;��H;��H;��H;��H;��H;��H;��H;��H;X�H;��H;u�H;W�H;H�H;W�H;v�H;��H;V�H;��H;��H;��H;��H;��H;��H;��H;��H;��H;��H;��H;zI;HI;�
I;BI;I;5I;-I;!I;#I;(I;��H;��H;g�H;ICH;�G; �G;�'G;+�F;��F;�YF;      OH;�TH;�dH;�}H;�H;��H;��H;�H;�I;QI;: I;L!I;�I;nI;�I;WI;�I;�I;I;�I;A�H;E�H;��H;��H;V�H;��H; �H;��H;��H;��H;��H;�H;��H;-�H;��H;��H;��H;��H;��H;,�H;��H;�H;��H;��H;��H;��H;��H;��H;W�H;��H;��H;H�H;A�H;�I;I;�I;�I;WI;�I;nI;�I;L!I;9 I;NI;�I;�H;��H;��H;�H;�}H;�dH;�TH;      �H;��H;�I;�	I;I;I;�I;!I;�!I;� I;�I;�I;I;0I;CI;z
I;�I;�I;p I;l�H;��H;p�H;K�H;T�H;j�H;��H;��H;��H;��H;��H;�H;q�H;�H;��H;q�H;A�H;9�H;A�H;q�H;��H;
�H;q�H;�H;��H;��H;��H;��H;��H;k�H;T�H;K�H;r�H;��H;m�H;r I;�I;�I;z
I;CI;0I;I;�I;�I;� I;�!I;!I;�I;I;I; 
I;�I;��H;      0"I;<"I;p"I;�"I;!"I;Y!I;�I;�I;�I;�I;�I;�I;`I;I;�I;�I;�I;�H;o�H;�H;��H;��H;�H;c�H;��H;��H;��H;��H;��H;�H;e�H;��H;��H;2�H;��H;��H;��H;��H;��H;2�H;�H;��H;e�H;
�H;��H;��H;��H;��H;��H;c�H;�H;��H;��H;�H;p�H;"�H;�I;�I;�I;I;_I;�I;�I;�I;�I;�I;�I;Y!I;("I;�"I;t"I;3"I;      �I;�I;$I;LI;I;|I;�I;�I;fI;�I;BI;�
I;�I;_I;�I;C I;��H;^�H;B�H;`�H;��H;��H;3�H;��H;��H;��H;��H;��H;
�H;W�H;��H;{�H;�H;��H;��H;��H;p�H;��H;��H;��H;�H;~�H;��H;V�H;�H;��H;��H;��H;��H;��H;2�H;��H;��H;`�H;B�H;a�H;��H;B I;�I;^I;�I;�
I;@I;�I;gI;�I;�I;|I;I;LI;"I;�I;      3I;I;�I;�I;�I;iI;�I;=I;NI;C	I;3I; I;�I;� I;i�H;V�H;c�H;��H;��H;�H;r�H;�H;��H;��H;��H;��H;��H;�H;d�H;��H;_�H;��H;��H;v�H;D�H;'�H;�H;'�H;D�H;v�H;��H;�H;_�H;��H;e�H;�H;��H;��H;��H;��H;��H;�H;o�H;�H;��H;��H;c�H;V�H;i�H;� I;�I; I;2I;D	I;OI;=I;�I;kI;�I;�I;�I;I;      �I;�I;dI;�I;�
I;�	I;�I;PI;�I;I;cI;� I;��H;��H;%�H;{�H;��H;'�H;��H;;�H;��H;��H;��H;��H;��H;��H;�H;r�H;��H;|�H;��H;��H;[�H;4�H;��H;��H;��H;��H;��H;4�H;X�H;��H;��H;~�H;��H;r�H;�H;��H;��H;��H;��H;��H;��H;;�H;��H;(�H;��H;{�H;%�H;��H;��H;� I;cI;I;�I;PI;�I;�	I;�
I;�I;bI;�I;      �I;vI;I;�I;�I;�I;�I;�I;cI;  I;��H;�H;��H;(�H;��H;0�H;��H;>�H;��H;��H;��H;��H;��H;��H;��H;W�H;��H;�H;��H;�H;��H;\�H;�H;��H;��H;��H;��H;��H;��H;��H;�H;_�H;��H;�H;��H;�H;��H;V�H;��H;��H;��H;��H;��H;��H;��H;?�H;��H;0�H;��H;)�H;��H;�H;��H; I;cI;�I;�I;�I;�I;�I;I;qI;      ,I;I;�I;mI;�I;I;< I;>�H;?�H;�H;��H;��H;Z�H;��H;��H;N�H;&�H;�H;��H;��H;��H;��H;�H;N�H;|�H;��H;)�H;��H;2�H;��H;s�H;2�H;��H;��H;��H;��H;r�H;��H;��H;��H;��H;8�H;t�H;��H;5�H;��H;)�H;��H;}�H;N�H;�H;��H;��H;��H;��H;�H;%�H;N�H;��H;��H;X�H;��H;��H;�H;A�H;>�H;< I;I;�I;nI;�I;I;      � I;� I;H I;��H;�H;��H;�H;�H;,�H;	�H;��H;��H;��H;��H;h�H;I�H;=�H;�H;�H;�H;=�H;Y�H;v�H;��H;�H;q�H;��H;q�H;��H;��H;B�H;��H;��H;��H;l�H;b�H;d�H;b�H;l�H;��H;��H;�H;C�H;��H;��H;q�H;��H;q�H;�H;��H;v�H;Y�H;:�H;�H;�H;�H;;�H;I�H;f�H;��H;��H;��H;��H;	�H;,�H;�H;�H;��H;u�H;��H;H I;� I;      ��H;��H;��H;D�H;��H;*�H;��H;��H;��H;��H;��H;��H;��H;��H;��H;��H;��H;~�H;��H;��H;��H;�H;=�H;��H;��H;R�H;��H;C�H;��H;��H;'�H;��H;��H;��H;b�H;H�H;H�H;H�H;b�H;��H;��H;��H;'�H;��H;��H;C�H;��H;P�H;��H;��H;=�H;�H;��H;��H;��H;�H;��H;��H;��H;��H;��H;��H;��H;��H;��H;��H;��H;.�H;��H;D�H;��H;��H;      D�H;:�H;�H;��H;/�H;}�H;��H;6�H;F�H;v�H;��H;��H;��H;o�H;^�H;a�H;Y�H;U�H;��H;��H;��H;��H;'�H;p�H;��H;D�H;��H;=�H;��H;t�H;�H;��H;��H;w�H;d�H;I�H;E�H;I�H;d�H;w�H;��H;��H;�H;v�H;��H;=�H;��H;E�H;��H;n�H;'�H;��H;��H;��H;��H;W�H;X�H;a�H;^�H;p�H;��H;��H;��H;x�H;H�H;4�H;��H;��H;$�H;��H;�H;2�H;      ��H;��H;��H;D�H;��H;*�H;��H;��H;��H;��H;��H;��H;��H;��H;��H;��H;��H;~�H;��H;��H;��H;�H;<�H;��H;��H;R�H;��H;C�H;��H;��H;'�H;��H;��H;��H;b�H;H�H;H�H;H�H;b�H;��H;��H;��H;'�H;��H;��H;C�H;��H;P�H;��H;��H;=�H;�H;��H;��H;��H;�H;��H;��H;��H;��H;��H;��H;��H;��H;��H;��H;��H;.�H;��H;D�H;��H;��H;      � I;� I;F I;��H;}�H;��H;�H;�H;,�H;�H;��H;��H;��H;��H;f�H;I�H;=�H;�H;�H;�H;>�H;Y�H;v�H;��H;�H;q�H;��H;q�H;��H;��H;C�H; �H;��H;��H;l�H;b�H;d�H;b�H;l�H;��H;��H;�H;C�H;��H;��H;q�H;��H;q�H;�H;��H;v�H;Y�H;:�H;�H;�H;�H;;�H;I�H;f�H;��H;��H;��H;��H;	�H;,�H;�H;�H;��H;u�H;��H;F I;� I;      -I;I;�I;nI;�I;I;< I;>�H;@�H;�H;��H;��H;X�H;��H;��H;N�H;&�H;�H;��H;��H;��H;��H;�H;P�H;}�H;��H;)�H;��H;0�H;��H;t�H;5�H;��H;��H;��H;��H;r�H;��H;��H;��H;��H;6�H;s�H;��H;5�H;��H;)�H;��H;|�H;M�H;�H;��H;��H;��H;��H;�H;%�H;N�H;��H;��H;Z�H;��H;��H;�H;A�H;@�H;< I;I;�I;mI;�I;I;      �I;vI;I;�I;�I;�I;�I;�I;cI;  I;��H;�H;��H;(�H;��H;0�H;��H;>�H;��H;��H;��H;��H;��H;��H;��H;W�H;��H;�H;��H;�H;��H;^�H;�H;��H;��H;��H;��H;��H;��H;��H;�H;a�H;��H;�H;��H;�H;��H;W�H;��H;��H;��H;��H;��H;��H;��H;>�H;��H;0�H;��H;(�H;��H;�H;��H; I;eI;�I;�I;�I;�I;�I;I;tI;      �I;�I;dI;�I;�
I;�	I;�I;SI;�I;I;cI;� I;��H;��H;%�H;{�H;��H;'�H;��H;=�H;��H;��H;��H;��H;��H;��H;�H;r�H;��H;|�H;��H;��H;Z�H;4�H;��H;��H;��H;��H;��H;4�H;X�H;��H;��H;~�H;��H;r�H;�H;��H;��H;��H;��H;��H;��H;;�H;��H;(�H;��H;{�H;#�H;��H;��H;� I;cI;I;�I;PI;�I;�	I;�
I;�I;dI;�I;      3I;I;�I;�I;�I;iI;�I;=I;OI;C	I;3I;I;�I;� I;i�H;W�H;c�H;��H;��H;�H;r�H;�H;��H;��H;��H;��H;��H;�H;c�H;��H;_�H;��H;��H;v�H;D�H;'�H;�H;'�H;D�H;v�H;��H;��H;_�H;��H;e�H;�H;��H;��H;��H;��H;��H;�H;o�H;�H;��H;��H;b�H;V�H;i�H;� I;�I;!I;2I;D	I;NI;?I;�I;kI;�I;�I;�I;I;      �I;�I;$I;KI;I;wI;�I;�I;gI;�I;@I;�
I;�I;_I;�I;B I;��H;`�H;B�H;a�H;��H;��H;3�H;��H;��H;��H;��H;��H;
�H;W�H;��H;{�H;�H;��H;��H;��H;p�H;��H;��H;��H;�H;|�H;��H;V�H;�H;��H;��H;��H;��H;��H;2�H;��H;��H;`�H;B�H;`�H;��H;E I;�I;^I;�I;�
I;BI;�I;iI;�I;�I;zI;I;KI;$I;�I;      )"I;9"I;w"I;�"I;&"I;W!I;�I;�I;�I;�I;�I;�I;`I;I;�I;�I;�I;�H;p�H;�H;��H;��H;�H;c�H;��H;��H;��H;��H;��H;�H;e�H;��H;��H;2�H;��H;��H;��H;��H;��H;2�H;��H;��H;e�H;
�H;��H;��H;��H;��H;��H;c�H;�H;��H;��H;�H;o�H;!�H;�I;�I;�I;I;_I;�I;�I;�I;�I;�I;�I;X!I;%"I;�"I;y"I;8"I;      �H;��H;�I; 
I;I;I;�I;!I;�!I;� I;�I;�I;I;2I;AI;z
I;�I;�I;r I;m�H;��H;r�H;K�H;T�H;k�H;��H;��H;��H;��H;��H;�H;q�H;
�H;��H;p�H;C�H;9�H;A�H;q�H;��H;�H;r�H;�H;��H;��H;��H;��H;��H;j�H;T�H;J�H;p�H;��H;l�H;p I;�I;�I;{
I;CI;/I;I;�I;�I;� I;�!I;!I;�I; I;I;�	I;�I;��H;      OH;�TH;�dH;�}H;�H;��H;��H;�H;�I;PI;9 I;L!I;�I;nI;�I;XI;�I;�I;I;�I;F�H;H�H;��H;��H;W�H;��H;�H;��H;��H;��H;��H;�H;��H;,�H;��H;��H;��H;��H;��H;,�H;��H;�H;��H;��H;��H;��H;��H;��H;V�H;��H;��H;E�H;@�H;�I;I;�I;�I;UI;�I;nI;�I;L!I;; I;PI;�I;	�H;��H;��H;�H;�}H;�dH;�TH;      �IF;�YF; �F;-�F;�'G;�G;�G;LCH;f�H;��H;��H;'I;$I;!I;,I;6I;I;AI;�
I;HI;~I;��H;��H;��H;��H;��H;��H;��H;��H;��H;��H;��H;W�H;��H;t�H;W�H;H�H;W�H;v�H;��H;V�H;��H;��H;��H;��H;��H;��H;��H;��H;��H;��H;��H;zI;HI;�
I;AI;I;8I;-I;!I;!I;(I;��H;��H;g�H;KCH;�G;�G;�'G;.�F; �F;�YF;      -EA;ElA;��A;��B;kC;�aD;�\E;-JF;�G; �G;�NH;k�H;�H;I;�I;� I;#I;zI;I;�I;9I;I;]�H;��H;�H;��H;Z�H;n�H;��H;��H;��H;��H;��H;��H;�H;��H;��H;��H;�H;��H;��H;��H;��H;��H;��H;m�H;X�H;��H;�H;��H;Y�H;I;7I;�I;I;{I;"I;� I;�I;I;�H;k�H;�NH; �G;�G;-JF;�\E;�aD;kC;��B;��A;ClA;      �J6;=�6;��7;�9;v;;@.=;}j?;��A;X�C;�2E;��F;��G;�<H;��H;�H;�I;� I;WI;dI;{I;�I;�I;yI;o�H;��H;��H;��H;Q�H;`�H;��H;��H;��H;��H;I�H;��H;��H;l�H;��H;��H;J�H;��H;��H;��H;��H;\�H;Q�H;��H;��H;��H;n�H;xI;�I;�I;zI;dI;ZI;� I;�I;�H;��H;�<H;��G;�F;�2E;Y�C;��A;}j?;A.=;�;;�9;��7;2�6;      kp ;!;4#;(&;%*;%p.;�3;�7;��;;Pj?;{kB;K�D;�xF;��G;3dH;C�H;�
I;�I;�I;�I;]I;^I;I;{I;Y�H;��H;��H;K�H;
�H;9�H;��H;��H;��H;�H;w�H;=�H;(�H;=�H;w�H;�H;��H;��H;��H;5�H;�H;K�H;��H;��H;W�H;xI;I;\I;YI;�I;�I;�I;�
I;C�H;3dH;��G;�xF;K�D;|kB;Mj?;��;;��7;�3;%p.;)*;(&;*#;!;      �t�:�:�l�:a�;� 
;�;az;AP$;��,;��3;E�9;@�>;M�B;V2E;@�F;�H;�H;�H;KI;7 I;eI;�I;\I;�I;I;��H;H�H;r�H;��H;��H;�H;��H;��H;��H;X�H;�H;��H;�H;Y�H;��H;��H;��H;�H;��H;��H;p�H;B�H;��H;I;�I;XI;�I;bI;7 I;KI;	�H;�H;�H;A�F;V2E;M�B;B�>;D�9;��3;��,;BP$;_z;�;� 
;a�;�l�:�:      t�>:@�G:��b:���:���:5�:I+�:�i;u�;*b;F*;zr3;��:;�!@;��C;�IF;�G;�H;L�H;�I;> I;eI;]I;�I;6I;I;C�H;��H;��H;��H;m�H;��H;��H;��H;6�H;��H;��H;��H;6�H;��H;��H;��H;m�H;��H;��H;��H;A�H;�I;6I;�I;\I;eI;< I;�I;K�H;��H;�G;�IF;��C;�!@;��:;yr3;D*;(b;w�;�i;K+�:5�:���:���:��b:�G:      ��������sk��� ���� 169��!:Ɋ:�4�:K�:��;1;��,;�6;�=;ĮB;��E;��G;}H;��H;�I;5 I;�I;|I;�I;JI;�I;j�H;�H;`�H;�H;3�H;��H;��H;�H;��H;��H;��H;�H;��H;��H;4�H;�H;\�H;�H;j�H;�I;JI;�I;xI;�I;5 I;�I;��H;}H;��G;��E;®B;�=;�6;��,;.;��;E�:�4�:
Ɋ:��!:p169����� ��sk�4���      /�������x���X���/�� ������m�@;�9x�k:�:�o�:�B;*&;|3;�<;]�A;�pE;�tG;}H;L�H;KI;�I;eI;I;�
I;I;s I;p�H;F�H;��H;��H;��H;��H;	�H;��H;��H;��H;	�H;��H;��H;��H;��H;C�H;n�H;s I;I;�
I;I;aI;�I;KI;H�H;}H;�tG;�pE;\�A;�<;|3;*&;�B;�o�:�:x�k:H;�9�m침���ܺ �}�/���X���x����      ������q
����&�׻�+�������;�zlۺp� ��Q�90Ɋ:���:�;U!;ѣ0;M;;��A;�pE;��G;�H;�H;�I;YI;xI;BI;�I;�I;"�H;d�H;��H;%�H;B�H;�H; �H;��H;^�H;��H;!�H;�H;A�H;'�H;��H;c�H;!�H;�I;�I;DI;xI;UI;�I;�H;�H;��G;�pE;��A;M;;ѣ0;W!;�;���:0Ɋ:�Q�9t� �xlۺ�;������+��#�׻����q
���      ~���k8����6�k���O��3/�$B��׻����4�@��O��`����>:d5�:��;�b;��/;M;;^�A;��E;�G;�H;�
I;� I;I;I;�I;�I;�I;��H;]�H;��H;��H; �H;6�H;��H;T�H;��H;6�H; �H;��H;��H;]�H;��H;�I;�I;�I;I;I;� I;�
I;�H;߿G;��E;]�A;P;;��/;�b;��;d5�:�>:p����O��7�@������׻$B��3/���O�6�k���l8��      :���|�.�ݼ��˼d���,����}���G����.�һ����2���/�H:�׳:'�;�b;ӣ0;�<;ɮB;�IF;�H;G�H;�I;� I;8I;XI;{
I;�I;? I;O�H;s�H;,�H;F�H;B�H;��H;\�H;��H;B�H;G�H;*�H;t�H;O�H;B I;�I;{
I;UI;<I;� I;�I;C�H;�H;�IF;ɮB;�<;գ0;�b;&�;�׳:@:�/�2������/�һ�����G���}��,��d����˼.�ݼ�|�      F�B�MR?��5���&��3��J��ѮҼF�����5=�?��-����/��mk����9�׳:��;U!;z3;�=;��C;?�F;4dH;�H;�I;/I;�I;CI;�I;�I;d�H;�H;��H;��H;c�H;��H;Z�H;��H;b�H;��H;��H;"�H;d�H;�I;�I;CI;�I;1I;�I;�H;/dH;@�F;��C;�=;z3;X!;��;�׳:���9�mk���/��-��?�6=����F��ѮҼ�J���3���&��5�MR?�      )��%W��钐�$�����j�P`I���&����Aϼ�,���T[�a�TI��1;��mk�L:f5�:�;*&;��6;�!@;V2E;��G;��H;I;!I;nI;.I;I;WI;� I;��H;%�H;��H;��H;��H;h�H;��H;��H;��H;"�H;��H;� I;XI;I;/I;mI;!I;I;��H;�G;V2E;�!@;��6;*&;�;d5�:L:�mk�1;�TI��a��T[��,��Aϼ�����&�P`I���j�$���钐�%W��      �J�����D��ͽ���(�������L�$��"��;����k����TI����/��/��>:���:�B;��,;��:;M�B;�xF;�<H;�H;$I;�I;I;`I;�I;�I;��H;��H;W�H;��H;��H;��H;��H;��H;W�H;��H;��H;�I;�I;_I;I;�I;)I;�H;�<H;�xF;O�B;��:;��,;�B;���:�>:�/���/�TI�������k�;��"��$����L����(������ͽ�D����      S�:��*7���,�+���	�s�齃���!W����j�>�/��J���I����k�a��-��2��`���6Ɋ:�o�:4;zr3;?�>;K�D;��G;g�H;(I;J!I;�I;�I;�
I;I;~ I;��H;��H;��H;��H;��H;��H;��H;��H;��H;~ I;I;�
I;�I;�I;H!I;(I;i�H;��G;H�D;@�>;}r3;4;�o�::Ɋ:p���4���-��a���k��I���J��>�/���j�!W������s�齃�	�+���,��*7�      ^���p����3�l���M���,�Yl�S9ݽ�A���{���5��J��;���T[�?������O���Q�9�:��;C*;B�9;|kB;��F;�NH;��H;; I;�I;�I;;I;*I;]I;�H;��H;��H;��H;��H;��H;��H;��H;~�H;_I;-I;;I;�I;�I;: I;��H;�NH;�F;ykB;B�9;F*;��;�:�Q�9�O������?��T[�;���J����5��{��A��S9ݽYl���,���M�3�l����p��      6m־R�Ѿ�>ľ����ԗ����{��I�+�����V���{�>�/�"���,��4=�.�һ4�@�h� ���k:M�:*b;��3;Qj?;�2E;�G;��H;PI;� I;�I;�I;?	I;I;��H;�H;�H;��H;v�H;��H;�H;�H;��H;I;?	I;�I;�I;� I;NI;��H;�G;�2E;Qj?;��3;,b;K�:��k:d� �6�@�.�һ4=��,��"��>�/��{��V�����+��I���{�ԗ�������>ľR�Ѿ      E\�î�s5��z ��E۾ֳ�^��{�Z�M?#����A����j�$��Aϼ����������~lۺ0;�9�4�:u�;~�,;��;;U�C;�G;l�H;�I;�!I;�I;\I;EI;�I;_I;<�H;#�H;��H;@�H;��H;%�H;<�H;\I;�I;GI;\I;�I;�!I;�I;l�H;�G;T�C;��;;��,;x�;�4�:0;�9zlۺ����������Aϼ$����j��A�����M?#�{�Z�^��ֳ��E۾�z �s5�î�      G�b��>]���M�Ŏ6�®�%���>ľ$q��{�Z�+�S9ݽ!W����L����F����G��׻�;��m�Ɋ:�i;;P$;��7;��A;.JF;PCH;	�H;� I;�I;�I;6I;KI;�I;9�H;�H;��H;/�H;��H;�H;9�H;�I;KI;6I;�I;�I;� I;�H;OCH;/JF;��A;��7;=P$;�i;
Ɋ:�m��;��׻��G�F�������L�!W��S9ݽ+�{�Z�$q���>ľ%��®�Ŏ6���M��>]�      p��򲗿���9�y�}�R���)�ov��>ľ^���I�Yl����������&�ѮҼ�}�%B�����������!:A+�:Zz;�3;{j?;�\E;�G;��H;�I;�I;�I;�I;�I;�I;; I;��H;��H;��H;��H;��H;: I;�I;�I;�I;�I;�I;�I;��H;�G;�\E;xj?;�3;[z;I+�:��!:��������%B��}�ѮҼ��&��������Yl��I�^���>ľov���)�}�R�9�y����򲗿      �˿�<ƿrL��B1����>]���)�%��ֳ���{���,�s��(��Q`I��J���,���3/��+��� �p1695�:	�;p.;@.=;�aD;
�G;��H;I;\!I;yI;kI;�	I;�I;	I;��H;1�H;��H;2�H;��H;	I;�I;�	I;lI;vI;Y!I;I;��H;
�G;�aD;<.=;!p.;	�;5�:p169� ��+���3/��,���J��Q`I�(��s�齥�,���{�ֳ�%����)��>]��B1��rL���<ƿ      ����>���W[忷˿�T���}�R�®��E۾ԗ����M���	������j��3�d����O�$�׻|�/������:� 
;/*;z;;kC;�'G;�H;I;%"I;I;�I;�
I;�I;�I;d�H;��H;�H;��H;c�H;�I;�I;�
I;�I;I;""I;I;�H;�'G;kC;w;;2*;� 
;���:��}�/�#�׻��O�d���3���j������	���M�ԗ���E۾®�}�R���T���˿W[�>���      O�7��v����˿B1��9�y�Ŏ6��z �����3�l�+��ͽ$�����&���˼6�k������X�ؘ �µ�:k�;2&;�9;��B;/�F;�}H;
I;�"I;NI;�I;�I;�I;fI;��H;C�H;��H;C�H;��H;fI;�I;�I;�I;KI;�"I;
I;�}H;/�F;��B;�9;4&;k�;ȵ�:ؘ ���X����6�k���˼��&�$����ͽ+�3�l������z �Ŏ6�9�y�B1���˿���v�7��      ��*��g&��#�v�W[�rL�������M�s5��>ľ����,��D�꒐��5�/�ݼ���q
���x��sk�`�b:�l�:(#;�7;��A;�F;�dH;�I;w"I;I;�I;]I;I;�I;> I;��H;��H;��H;> I;�I;I;]I;�I;I;t"I;�I;�dH;�F;��A;�7;(#;�l�:d�b:�sk���x��q
���/�ݼ�5�꒐��DὫ�,����>ľs5���M����rL��W[�v��#��g&�      ��8��4��g&�7��>����<ƿ򲗿�>]�î�R�Ѿ�p���*7����&W��MR?��|�l8�������:����G:� �:!;/�6;:lA;�YF;�TH;��H;8"I;�I;
I;�I;dI;I;� I;��H;0�H;��H;� I;I;cI;�I;
I;�I;5"I;��H;�TH;�YF;:lA;-�6;!;� �:�G:>��������l8���|�MR?�&W�����*7��p��R�Ѿî��>]�򲗿�<ƿ>���7���g&��4�      ��!$������꿰�ſ�ޞ�'3s��2�?����� j���{HͽƸ����'�@<ͼi�n�V���Q^��,.����:�W;�S%;|o8;��A;vDF;�H;��H;�H;	�H;a�H;X�H;`�H;��H;�H;��H;F�H;��H;�H;��H;^�H;Y�H;a�H;�H;�H;��H;�H;uDF;��A;{o8;�S%;�W;���:�,.�Q^�T���j�n�@<ͼ��'�Ƹ��{Hͽ�� j���?����2�'3s��ޞ���ſ������!$�      !$�������忉�����!cm�W�-�����Rh��Xde�#-�تɽ�v��(�$�~�ɼpmj�)����X���(Ɔ:�x;^�%;J�8;�B;�RF;H;E�H;k�H;�H;��H;\�H;R�H;��H;��H;��H;A�H;��H;��H;��H;P�H;]�H;��H;�H;i�H;E�H;H;�RF;�B;G�8;d�%;�x;(Ɔ:���X�(���qmj�~�ɼ(�$��v��تɽ#-�Xde�Rh������W�-�!cm��������忞����      ��������� �ԿNw�����<�\�"����m��\0X�����;����w����������]��黣F����0ʒ:�;U�';׏9;9pB;�zF;�!H;��H;O�H;2�H;��H;b�H;W�H;��H;��H;��H;,�H;��H;��H;��H;V�H;b�H;��H;/�H;L�H;��H;�!H;�zF;9pB;ԏ9;X�';�;,ʒ:��깣F��黤�]����������w��;�����\0X�m�����"�<�\����Nw�� �Կ��𿞏�      ����� �Կp���ޞ�bF�i�C�.E�$�;�I���D���"��g�c�|��֯���J��ѻ��)�p{K�d��:9�
;
N*;��:;�C;$�F;�8H;m�H;��H;��H;��H;[�H;W�H;��H;��H;��H;�H;��H;��H;��H;V�H;[�H;��H;��H;��H;m�H;�8H;#�F;�C;��:;N*;9�
;d��:�{K���)��ѻ��J��֯�|�g�c�"�����D��I��$�;.E�i�C�bF��ޞ�p�� �Կ��      ��ſ���Nw���ޞ�����@�W�7�%�����jɰ��|x�h{+�ӱ����J��  �˶��P�1�����*��$
9<�:΅;.�-;��<;��C;�G;�TH;e�H;�H;�H;��H;q�H;O�H;��H;��H;��H;�H;��H;��H;��H;N�H;r�H;��H;�H;�H;e�H;�TH;�G;��C;��<;1�-;̅;<�:�$
9�*����Q�1�ʶ���  ��J���ӱ�h{+��|x�jɰ�����6�%�@�W������ޞ�Nw�����      �ޞ�������bF�A�W�X�-����AKɾ�G����O����ƽǸ��τ-���ۼㄼ,4�ǐ��ζ�(^:C��:�;Ɩ1;d>;��D;�\G;[sH;��H;��H;z�H;<�H;��H;E�H;��H;��H;��H;��H;��H;��H;��H;E�H;��H;<�H;w�H;~�H;��H;YsH;�\G;��D;d>;Ŗ1;�;E��:$^:�ζ�ǐ�,4�ㄼ��ۼ΄-�Ǹ��ƽ�����O��G��AKɾ���X�-�A�W�bF�������      (3s�!cm�<�\�j�C�7�%�����TҾl�� j��C(����_P����[�{������Y�$��;X���<��k:���:� ;�5;_R@;}uE;�G;I�H;_�H;��H;�H;_�H;��H;A�H;��H;��H;u�H;��H;u�H;��H;��H;A�H;��H;_�H;�H;��H;_�H;G�H;�G;{uE;\R@;�5;� ;���:�k:��<�8X�$����Y����{���[�_P����콬C(� j�l���TҾ���7�%�j�C�<�\�!cm�      �2�W�-�"�.E�����AKɾl����s�9�5���w㻽�v��	z0��;��+���*����6�@5S��M�:{�	;��(;7�9;�/B;�DF;lH;�H;��H;��H;��H;��H;��H;-�H;O�H;\�H;Y�H;v�H;W�H;\�H;N�H;*�H;��H;��H;��H;��H;��H;�H;kH;�DF;�/B;7�9;��(;|�	;�M�:@5S�6�����*��+���;�	z0��v��w㻽��9�5���s�l��AKɾ����.E�"�W�-�      ?����������$�;jɰ��G�� j�9�5��	�ЪɽZ����J�r���沼��]�����	x�����n:��:�v;��/;�-=;��C;^�F;7IH;��H;=�H;��H;8�H;��H;��H;�H;#�H;)�H;2�H;A�H;2�H;)�H;"�H;�H;��H;��H;7�H;��H;;�H;��H;7IH;[�F;��C;�-=;��/;�v;	��:�n:����	x������]��沼r���J�Z���Ъɽ�	�:�5� j��G��jɰ�$�;��徹���      ��Rh��m���I���|x���O��C(���Ъɽ����SDX�H��%<ͼㄼ�X!��s���W��rK����:�y;0�#;!I6;OR@;�PE;��G;��H;��H;G�H;�H;��H;��H;��H;��H;�H;��H;��H;��H;��H;��H;�H;��H;��H;��H;��H;�H;G�H;��H;��H;��G;�PE;NR@;!I6;.�#;�y;���:�rK��W��s���X!�ㄼ%<ͼH��SDX�����Ъɽ���C(���O��|x��I��m��Rh��       j�Xde�\0X��D�h{+�������x㻽Z���SDX������ۼȾ��}�;�2>ۻ�X���y��?":��:��;��-;��;;�B;�zF;�H;��H;��H;;�H; �H;�H;�H;��H;��H;��H;��H;��H;��H;��H;��H;��H;��H;��H;�H;�H;��H;;�H;��H;��H;�H;�zF;�B;��;;�-;��;��:�?":��y��X�2>ۻ}�;�Ⱦ����ۼ���SDX�Z���x㻽��콄��h{+��D�\0X�Xde�      ��#-������Ա�ƽ_P���v���J�H����ۼ
��[�J�����p+��*rѺ�+
9+N�:�;� $;%�5;�?;��D;z\G;fH;�H;��H;��H;��H;6�H;�H;q�H;��H;{�H;t�H;��H;Y�H;��H;u�H;{�H;��H;t�H;�H;8�H;��H;��H;��H;�H;fH;v\G;��D;�?;%�5;� $;�;1N�:`+
9,rѺp+������[�J�
����ۼH���J��v��_P��ƽԱ轅����#-�      {Hͽتɽ�;��"����Ǹ����[�	z0�r��%<ͼȾ��[�J����j��M*���Z��:�b�:r�;�/;�L<;'C;GmF;��G;!�H;$�H;*�H;)�H;^�H;o�H;�H;D�H;Q�H;<�H;6�H;$�H;�H;$�H;6�H;:�H;N�H;F�H;�H;o�H;]�H;(�H;&�H;#�H;�H;��G;CmF;'C;�L<;
�/;r�;�b�:V��:p�M*��j����[�J�Ⱦ��%<ͼr��	z0���[�Ǹ����"���;��تɽ      Ƹ���v����w�g�c��J�΄-�{��;缃沼ㄼ|�;������j��x5��깼?Q:���:�i;N*;��8;��@;�PE;�uG;WiH;��H;��H;.�H;@�H;��H;��H;�H;�H;��H;��H;��H;��H;��H;��H;��H;��H;��H;�H;�H;��H;��H;@�H;*�H;��H;��H;TiH;�uG;�PE;��@;��8;N*;�i;���:�?Q:ؾ�w5��j������|�;�ㄼ�沼�;�{�΄-��J�g�c���w��v��      ��'�(�$����|��  ���ۼ����+����]��X!�3>ۻp+��N*��깐�>:*��:2�;S�%;	�5;��>;�(D;*�F;�!H;N�H;p�H;�H;��H;��H;	�H;��H;��H;��H;��H;��H;��H;o�H;��H;o�H;��H;��H;��H;��H;��H;��H;�H;��H;��H;�H;n�H;J�H;�!H;*�F;�(D;��>;�5;V�%;0�;*��:��>:��N*�p+��4>ۻ�X!���]��+�������ۼ�  �|����(�$�      @<ͼ~�ɼ�����֯�˶��ㄼ��Y��*�����s���X�,rѺ���?Q:0��:��
;n�#;��3;�c=;"$C;DDF; �G;/�H;�H;/�H;W�H;�H;w�H;D�H;��H;��H;��H;X�H;s�H;-�H;�H;*�H;�H;-�H;s�H;W�H;��H;��H;��H;?�H;w�H;�H;W�H;.�H; �H;+�H; �G;?DF;"$C;�c=;��3;n�#;��
;0��:�?Q:��,rѺ�X��s������*���Y�ㄼ˶���֯�����~�ɼ      j�n�omj���]���J�R�1�,4�"������	x��W���y�`+
9T��:���:4�;i�#;t�2;�<;�pB;G�E;ύG;�eH;�H;U�H;��H;�H;��H;��H;\�H;j�H;Z�H;1�H;�H;��H;��H;��H;��H;��H;��H;��H;�H;2�H;Z�H;i�H;Z�H;��H;��H;�H;��H;Q�H;�H;�eH;̍G;H�E;�pB;�<;x�2;k�#;4�;���:V��:�+
9��y��W��	x����!��+4�R�1���J���]�qmj�      X���)������ѻ���ǐ�<X�	6���� sK��?":+N�:�b�:�i;T�%;�3;�<;b0B;��E;�\G;�HH;d�H;��H;~�H;�H;Y�H;^�H;��H;9�H;<�H;�H;��H;��H;��H;u�H;s�H;P�H;s�H;u�H;��H;��H;��H;�H;;�H;6�H;��H;[�H;Z�H;�H;z�H;��H;d�H;�HH;�\G;E;e0B;�<;~�3;T�%;�i;�b�:+N�:�?":�rK����
6�<X�
ǐ�����ѻ��.���      Q^��X��F���)��*��ζ���<�@6S��n:~��:��:�;n�;	N*;�5;�c=;�pB;��E;�JG;s8H;��H;��H;3�H;M�H;��H;�H;��H;�H;�H;��H;��H;��H;y�H;&�H;�H;�H;��H;�H;�H;%�H;w�H;��H;��H;��H;�H;�H;��H;�H;��H;H�H;0�H;��H;��H;v8H;�JG;ÇE;�pB;�c=;�5;	N*;n�;�;��:~��:�n:@6S���<��ζ��*���)��F��X�      �,.�̪���김{K�`$
9 ^:��k:�M�:��:�y;��;� $;�/;��8;��>;$C;D�E;�\G;p8H;�H;(�H;B�H;��H;X�H;��H;v�H;��H;��H;��H;��H;^�H;5�H;�H;��H;��H;��H;��H;��H;��H;��H;�H;7�H;^�H;��H;��H;��H;��H;v�H;��H;R�H;��H;D�H;%�H;�H;r8H;�\G;G�E;$C;��>;��8;�/;� $;��;�y;��:�M�:��k:$^: %
9�{K������      ���:HƆ:2ʒ:T��:,�:I��:���:x�	;�v;0�#;�-;!�5;�L<;��@;�(D;?DF;΍G;�HH;��H;'�H;��H;n�H;��H;��H;C�H;��H;��H;��H;��H;F�H;)�H;��H;��H;��H;U�H;G�H;G�H;G�H;V�H;��H;��H;��H;)�H;C�H;��H;��H;��H;��H;C�H;�H;��H;n�H;��H;(�H;��H;�HH;΍G;?DF;�(D;��@;�L<;#�5;�-;.�#;�v;x�	;���:Q��:,�:X��:6ʒ:&Ɔ:      �W;�x;&�;/�
;̅;�;"� ;��(;��/; I6;��;;�?;%C;�PE;-�F;�G;�eH;d�H;��H;D�H;n�H;��H;S�H;�H;��H;��H;��H;��H;�H;��H;��H;m�H;B�H;0�H;��H;��H;��H;��H;��H;0�H;A�H;m�H;��H;��H;�H;��H;��H;��H;��H;�H;S�H;��H;m�H;E�H;��H;e�H;�eH;�G;.�F;�PE;(C;�?;��;;!I6;��/;��(;"� ;�;��;.�
;'�;�x;      �S%;`�%;T�';N*;&�-;Ɩ1;�5;4�9;�-=;LR@;�B;��D;DmF;�uG;�!H;+�H;�H;��H;3�H;��H;��H;U�H;)�H;��H;��H;��H;`�H;�H;��H;��H;K�H;�H;��H;��H;��H;��H;|�H;��H;��H;��H;��H;�H;L�H;��H;��H;�H;[�H;��H;��H;��H;)�H;V�H;��H;��H;3�H;��H;�H;*�H;�!H;�uG;DmF;��D;�B;LR@;�-=;4�9;�5;Ȗ1;0�-;N*;W�';S�%;      �o8;X�8;ۏ9;��:;��<;d>;fR@;�/B;��C;�PE;�zF;y\G;��G;WiH;M�H; �H;Q�H;~�H;J�H;U�H;}�H;�H;��H;��H;��H;r�H;�H;��H;��H;:�H;��H;��H;��H;X�H;R�H;F�H;"�H;F�H;T�H;V�H;��H;��H;��H;7�H;��H;��H;�H;r�H;��H;��H;��H;�H;{�H;V�H;L�H;�H;Q�H;�H;N�H;WiH;��G;y\G;�zF;�PE;��C;�/B;fR@;d>;��<;��:;ޏ9;J�8;      ��A;�B;$pB;�C;��C;��D;|uE;�DF;\�F;��G;�H;fH;�H;��H;q�H;1�H;��H;�H;��H;��H;E�H;��H;��H;��H;Q�H;��H;��H;��H;0�H;��H;��H;n�H;<�H;�H;��H;��H;��H;��H;��H;�H;:�H;p�H;��H;��H;/�H;��H;��H;��H;S�H;��H;��H;��H;E�H;��H;��H;#�H;��H;/�H;q�H;��H;�H; fH;�H;��G;[�F;�DF;|uE;��D;��C;�C;'pB;�B;      �DF;�RF;�zF;!�F;�G;�\G;�G;dH;6IH;��H;��H;
�H;�H;��H;�H;T�H;�H;V�H;��H;s�H;��H;��H;��H;p�H;��H;��H;��H;)�H;��H;��H;J�H;�H;��H;��H;��H;��H;��H;��H;��H;��H;��H;�H;J�H;��H;��H;)�H;��H;��H;��H;o�H;��H;��H;��H;u�H;��H;V�H;�H;T�H;�H;��H;�H;
�H;��H;��H;6IH;dH;�G;�\G;�G;!�F;�zF;�RF;      H;H;�!H;�8H;�TH;^sH;M�H;�H;��H;��H;��H;��H;&�H;-�H;��H;�H;��H;Z�H;��H;��H;��H;��H;]�H;�H;��H;��H;�H;��H;z�H;H�H;�H;��H;��H;w�H;^�H;9�H;M�H;;�H;^�H;w�H;��H;��H;�H;G�H;x�H;��H;�H;��H;��H;�H;[�H;��H;��H;��H;��H;]�H;��H;�H;��H;-�H;&�H;��H;��H;��H;��H;�H;P�H;[sH;�TH;�8H;�!H;!H;      ��H;H�H;��H;h�H;e�H;��H;c�H;��H;?�H;L�H;@�H;��H;(�H;B�H;��H;v�H;��H;��H;�H;��H;��H;��H;�H;��H;��H;*�H;��H;��H;9�H;��H;��H;z�H;T�H;!�H;�H;�H;�H;�H;�H;#�H;S�H;{�H;��H;��H;7�H;��H;��H;*�H;��H;��H;�H;��H;��H;��H;�H;��H;��H;v�H;��H;A�H;)�H;��H;>�H;K�H;A�H;��H;d�H;��H;p�H;h�H;��H;T�H;      �H;n�H;H�H;��H;�H;��H;��H; �H;��H;	�H; �H;��H;]�H;��H;�H;D�H;\�H;5�H;�H;��H;��H;�H;��H;��H;)�H;��H;u�H;9�H;��H;��H;l�H;5�H; �H;��H;��H;��H;��H;��H;��H;��H;��H;8�H;m�H;��H;��H;9�H;w�H;��H;,�H;��H;��H;�H;��H;��H;�H;8�H;\�H;C�H;�H;��H;]�H;��H;��H;�H; �H;��H;��H;�H;�H;��H;L�H;f�H;      �H;$�H;<�H;��H;�H;~�H;�H;��H;A�H;��H;�H;B�H;t�H;��H;��H;��H;l�H;6�H;��H;��H;E�H;��H;��H;:�H;��H;��H;F�H;��H;��H;c�H;2�H;��H;��H;��H;��H;��H;w�H;��H;��H;��H;��H;��H;4�H;c�H;��H;��H;C�H;��H;��H;;�H;��H;��H;C�H;��H;��H;8�H;l�H;��H;��H;��H;t�H;B�H;�H;��H;B�H;��H;�H;�H;�H;��H;8�H;#�H;      e�H;��H;��H;��H;�H;<�H;i�H;��H;��H;��H;	�H;�H;�H;�H;��H;��H;^�H;�H;��H;d�H;.�H;��H;I�H;��H;��H;K�H;��H;��H;j�H;5�H;��H;��H;��H;y�H;V�H;`�H;^�H;`�H;W�H;z�H;��H;��H;��H;5�H;m�H;��H;��H;J�H;��H;��H;I�H;��H;,�H;d�H;��H;�H;_�H;��H;��H;�H;�H;�H;	�H;��H;��H;��H;i�H;=�H;	�H;��H;��H;��H;      c�H;m�H;g�H;c�H;w�H;��H;��H;��H;��H;��H;��H;z�H;G�H;�H;��H;��H;9�H;��H;��H;>�H;��H;o�H;�H;��H;k�H;�H;��H;}�H;5�H;��H;��H;��H;z�H;F�H;1�H;0�H;3�H;0�H;1�H;F�H;y�H;��H;��H;��H;6�H;}�H;��H;	�H;m�H;��H;�H;q�H;��H;>�H;��H;��H;8�H;��H;��H;�H;H�H;z�H;��H;��H;��H;��H;��H;��H;u�H;c�H;g�H;i�H;      d�H;e�H;`�H;a�H;Z�H;B�H;B�H;4�H;
�H;��H;��H;��H;T�H;�H;��H;\�H;�H;��H;|�H;�H;��H;D�H;��H;��H;6�H;��H;��H;W�H;�H;��H;��H;|�H;4�H;)�H;)�H;�H;��H;�H;)�H;)�H;1�H;��H;��H;��H;�H;X�H;��H;��H;7�H;��H;��H;D�H;��H;�H;|�H;��H;�H;\�H;��H;�H;R�H;��H;��H;��H;
�H;4�H;B�H;G�H;U�H;a�H;`�H;^�H;      ��H;��H;��H;��H;��H;��H;��H;W�H;(�H;	�H;��H;��H;?�H;��H;��H;x�H;��H;��H;)�H;��H;��H;3�H;��H;]�H;�H;��H;t�H;!�H;��H;��H;w�H;H�H;%�H;�H;�H;��H;��H;��H;�H;�H;#�H;J�H;y�H;��H;��H;!�H;t�H;��H;�H;\�H;��H;3�H;��H;��H;)�H;��H;��H;x�H;��H;��H;?�H;��H;��H;�H;)�H;W�H;��H;��H;��H;��H;��H;��H;      �H;�H;��H;��H;��H;��H;��H;h�H;3�H;��H;��H;��H;?�H;��H;��H;5�H;��H;r�H;�H;��H;]�H;��H;��H;X�H;��H;��H;[�H;�H;��H;��H;T�H;5�H;'�H;�H;��H;��H;��H;��H;��H;�H;&�H;8�H;V�H;��H;��H;�H;Z�H;��H;��H;V�H;��H;��H;Z�H;��H;�H;s�H;��H;5�H;��H;��H;=�H;��H;��H;��H;3�H;g�H;��H;��H;��H;��H;��H;
�H;      ��H;��H;��H;��H;��H;��H;|�H;d�H;>�H;��H;��H;��H;+�H;��H;s�H;�H;��H;o�H;�H;��H;N�H;��H;��H;M�H;��H;��H;9�H;�H;��H;��H;`�H;4�H;�H;��H;��H;��H;��H;��H;��H;��H;�H;8�H;`�H;��H;��H;�H;8�H;��H;��H;J�H;��H;��H;L�H;��H;�H;p�H;��H;�H;t�H;��H;)�H;��H;��H;��H;>�H;c�H;|�H;��H;��H;��H;��H;��H;      F�H;L�H;<�H;�H;�H;��H;��H;�H;H�H;��H;��H;b�H;�H;��H;��H;1�H;��H;I�H;��H;��H;I�H;��H;z�H;'�H;��H;��H;L�H;�H;��H;}�H;a�H;:�H;��H;��H;��H;��H;��H;��H;��H;��H;��H;;�H;a�H;}�H;��H;�H;J�H;��H;��H;$�H;{�H;��H;I�H;��H;��H;J�H;��H;1�H;��H;��H;�H;c�H;��H;��H;K�H;}�H;��H;��H;�H;�H;;�H;C�H;      ��H;��H;��H;��H;��H;��H;|�H;d�H;>�H;��H;��H;��H;)�H;��H;t�H;�H;��H;o�H;�H;��H;O�H;��H;��H;K�H;��H;��H;9�H;�H;��H;��H;`�H;5�H;�H;��H;��H;��H;��H;��H;��H;��H;�H;7�H;`�H;��H;��H;�H;8�H;��H;��H;J�H;��H;��H;L�H;��H;�H;p�H;��H;�H;s�H;��H;+�H;��H;��H;��H;>�H;c�H;|�H;��H;��H;��H;��H;��H;      �H;�H;��H;��H;��H;��H;��H;h�H;3�H;��H;��H;��H;=�H;��H;��H;5�H;��H;r�H;�H;��H;^�H;��H;��H;X�H;��H;��H;[�H;�H;��H;��H;V�H;5�H;'�H;�H;��H;��H;��H;��H;��H;�H;&�H;:�H;T�H;��H;��H;�H;Z�H;��H;��H;U�H;��H;��H;Z�H;��H;�H;s�H;��H;5�H;��H;��H;?�H;��H;��H;��H;3�H;g�H;��H;��H;��H;��H;��H;�H;      ��H;��H;��H;��H;��H;��H;��H;W�H;(�H;�H;��H;��H;?�H;��H;��H;x�H;��H;��H;)�H;��H;��H;3�H;��H;]�H;�H;��H;t�H;!�H;��H;��H;y�H;H�H;%�H;�H;�H;��H;��H;��H;�H;�H;#�H;J�H;w�H;��H;��H;!�H;v�H;��H;�H;[�H;��H;3�H;��H;��H;)�H;��H;��H;x�H;��H;��H;?�H;��H;��H;	�H;)�H;W�H;��H;��H;��H;��H;��H;��H;      g�H;d�H;a�H;d�H;Z�H;D�H;D�H;3�H;
�H;��H;��H;��H;R�H;�H;��H;\�H;�H;��H;|�H;�H;��H;D�H;��H;��H;7�H;��H;��H;X�H;�H;��H;��H;}�H;3�H;'�H;)�H;�H;��H;�H;)�H;'�H;1�H;��H;��H;��H;�H;W�H;��H;��H;6�H;��H;��H;D�H;��H;�H;|�H;��H;�H;\�H;��H;��H;R�H;��H;��H;��H;�H;2�H;D�H;E�H;R�H;d�H;]�H;c�H;      c�H;m�H;i�H;b�H;w�H;��H;��H;��H;��H;��H;��H;z�H;G�H;�H;��H;��H;8�H;��H;��H;?�H;��H;q�H;�H;��H;m�H;�H;��H;}�H;4�H;��H;��H;��H;z�H;F�H;1�H;0�H;3�H;0�H;1�H;F�H;w�H;��H;��H;��H;6�H;}�H;��H;	�H;k�H;��H;�H;o�H;��H;>�H;��H;��H;8�H;��H;��H;�H;G�H;z�H;��H;��H;��H;��H;��H;��H;u�H;b�H;g�H;i�H;      e�H;��H;��H;��H;�H;;�H;i�H;��H;��H;��H;	�H;�H;�H;�H;��H;��H;^�H;�H;��H;d�H;0�H;��H;K�H;��H;��H;K�H;��H;��H;l�H;6�H;��H;��H;��H;z�H;W�H;`�H;^�H;`�H;V�H;y�H;��H;��H;��H;4�H;l�H;��H;��H;J�H;��H;��H;G�H;��H;,�H;d�H;��H;�H;^�H;��H;��H;�H;�H;�H;�H;��H;��H;��H;i�H;=�H;	�H;��H;��H;��H;      �H;$�H;;�H;��H;�H;z�H;!�H;��H;B�H;��H;�H;B�H;t�H;��H;��H;��H;m�H;6�H;��H;��H;H�H;��H;��H;;�H;��H;��H;F�H;��H;��H;e�H;4�H;��H;��H;��H;��H;��H;w�H;��H;��H;��H;��H;��H;2�H;b�H;��H;��H;C�H;��H;��H;:�H;��H;��H;C�H;��H;��H;8�H;j�H;��H;��H;��H;t�H;B�H;�H;��H;C�H;��H;�H;|�H;�H;��H;;�H;#�H;      �H;k�H;O�H;��H;�H;{�H;��H;��H;��H;�H; �H;��H;]�H;��H;�H;C�H;^�H;6�H;�H;��H;��H;�H;��H;��H;,�H;��H;u�H;9�H;��H;��H;m�H;5�H; �H;��H;��H;��H;��H;��H;��H;��H;��H;6�H;l�H;��H;��H;9�H;w�H;��H;)�H;��H;��H;�H;��H;��H;�H;6�H;\�H;F�H;�H;��H;]�H;��H; �H;�H; �H;�H;��H;�H;�H;��H;P�H;j�H;      ��H;I�H;��H;h�H;f�H;��H;d�H;��H;?�H;K�H;@�H;��H;)�H;A�H;��H;v�H;��H;��H;�H;��H;��H;��H;�H;��H;��H;*�H;��H;��H;9�H;��H;��H;{�H;T�H;!�H;�H;�H;�H;�H;�H;!�H;S�H;{�H;��H;��H;9�H;��H;��H;*�H;��H;��H;�H;��H;��H;��H;�H;��H;��H;w�H;��H;@�H;(�H;��H;>�H;L�H;B�H;��H;c�H;��H;q�H;h�H;��H;Q�H;       H;H;�!H;�8H;�TH;YsH;N�H;�H;��H;��H;��H;��H;&�H;-�H;��H;�H;��H;[�H;��H;��H;��H;��H;]�H;�H;��H;��H;�H;��H;x�H;H�H;�H;��H;��H;w�H;^�H;;�H;M�H;8�H;^�H;v�H;��H;��H;�H;G�H;x�H;��H;�H;��H;��H;�H;[�H;��H;��H;��H;��H;[�H;��H;�H;��H;-�H;&�H;��H;��H;��H;��H;�H;L�H;XsH;�TH;�8H;�!H;H;      �DF;�RF;�zF;#�F;�G;�\G;�G;fH;4IH;��H;��H;�H; �H;��H;�H;V�H;�H;U�H;��H;u�H;��H;��H;��H;p�H;��H;��H;��H;)�H;��H;��H;J�H;�H;��H;��H;��H;��H;��H;��H;��H;��H;��H;�H;J�H;��H;��H;)�H;��H;��H;��H;o�H;��H;��H;��H;s�H;��H;W�H;�H;T�H;�H;��H;�H;
�H;��H;��H;4IH;eH;�G;�\G;�G;#�F;�zF;�RF;      ��A;�B;%pB;�C;��C;��D;|uE;�DF;[�F;��G;�H; fH;�H;��H;q�H;1�H;��H; �H;��H;��H;H�H;��H;��H;��H;S�H;��H;��H;��H;/�H;��H;��H;n�H;:�H;�H;��H;��H;��H;��H;��H;�H;:�H;q�H;��H;��H;-�H;��H;��H;��H;Q�H;��H;��H;��H;C�H;��H;��H;!�H;��H;1�H;q�H;��H;�H;fH;�H;��G;\�F;�DF;|uE;��D;��C;�C;'pB;�B;      �o8;U�8;�9;��:;��<;d>;bR@;�/B;��C;�PE;�zF;y\G;��G;WiH;N�H;�H;Q�H;}�H;L�H;V�H;�H;�H;��H;��H;��H;p�H;�H;��H;��H;:�H;��H;��H;��H;U�H;Q�H;G�H;"�H;F�H;T�H;X�H;��H;��H;��H;7�H;��H;��H;�H;r�H;��H;��H;��H;�H;{�H;U�H;J�H;�H;P�H; �H;M�H;WiH;��G;y\G;�zF;�PE;��C;�/B;`R@;d>;��<;��:;�9;I�8;      �S%;o�%;c�';N*;'�-;̖1;#�5;4�9;�-=;LR@;�B;��D;CmF;�uG;�!H;+�H;�H;��H;3�H;��H;��H;V�H;*�H;��H;��H;��H;`�H;�H;��H;��H;L�H;�H;��H;��H;��H;��H;|�H;��H;��H;��H;��H;�H;K�H;��H;��H;�H;]�H;��H;��H;��H;'�H;U�H;��H;��H;3�H;��H;�H;+�H;�!H;�uG;CmF;��D;�B;JR@;�-=;5�9;#�5;̖1;,�-;N*;[�';]�%;      �W;�x;$�;.�
;΅;�;"� ;��(;��/;!I6;��;;�?;(C;�PE;-�F; �G;�eH;d�H;��H;D�H;n�H;��H;U�H;�H;��H;��H;��H;��H;�H;��H;��H;m�H;B�H;0�H;��H;��H;��H;��H;��H;0�H;A�H;m�H;��H;��H;�H;��H;��H;��H;��H;�H;P�H;��H;m�H;E�H;��H;e�H;�eH;�G;.�F;�PE;%C;�?;��;; I6;��/;��(;"� ;�;�;/�
;&�;�x;      ���:<Ɔ::ʒ:X��:,�:=��:���:{�	;�v;.�#;�-;#�5;�L<;��@;�(D;?DF;ύG;�HH;��H;(�H;��H;n�H;��H;��H;C�H;��H;��H;��H;��H;F�H;)�H;��H;��H;��H;V�H;G�H;G�H;G�H;U�H;��H;��H;��H;)�H;C�H;��H;��H;��H;��H;C�H;}�H;��H;n�H;��H;(�H;��H;�HH;̍G;?DF;�(D;��@;�L<;!�5;�-;-�#;�v;{�	;���:I��:4�:V��:>ʒ:$Ɔ:      �,.�Ȫ�p�깠{K��$
9^:�k:�M�:	��:�y;��;� $;�/;��8;��>;$C;E�E;�\G;r8H;�H;(�H;D�H;��H;X�H;��H;v�H;��H;��H;��H;��H;^�H;5�H;�H;��H;��H;��H;��H;��H;��H;��H;�H;7�H;^�H;��H;��H;��H;��H;v�H;��H;R�H;��H;B�H;%�H;�H;p8H;�\G;E�E;$C;��>;��8;�/;� $;��;�y;	��:�M�:�k:(^: %
9�{K�������      Q^��X��F���)��*��ζ���<� 6S��n:~��:��:�;n�;	N*;�5;�c=;�pB;E;�JG;t8H;��H;��H;3�H;L�H;��H; �H;��H;�H;�H;��H;��H;��H;y�H;%�H;�H;�H;��H;�H;�H;&�H;w�H;��H;��H;��H;�H;�H;��H;�H;��H;H�H;.�H;��H;��H;v8H;�JG;E;�pB;�c=;�5;	N*;n�;�;��:~��:�n: 6S���<��ζ��*���)��F��X�      W���*������ѻ���ǐ�;X�	6�����rK��?":/N�:�b�:�i;T�%;~�3;�<;c0B;E;�\G;�HH;d�H;��H;~�H;�H;W�H;^�H;��H;9�H;<�H;�H;��H;��H;��H;u�H;s�H;P�H;s�H;u�H;��H;��H;��H;�H;;�H;6�H;��H;[�H;Z�H;�H;x�H;��H;d�H;�HH;�\G;��E;c0B;�<;�3;T�%;�i;�b�:+N�:�?": sK����	6�;X�
ǐ�����ѻ��.���      j�n�omj���]���J�R�1�,4� ������	x��W���y�`+
9V��:���:4�;k�#;x�2;�<;�pB;H�E;΍G;�eH;�H;U�H;��H;�H;��H;��H;[�H;j�H;Z�H;2�H;�H;��H;��H;��H;��H;��H;��H;��H;�H;2�H;Z�H;i�H;Z�H;��H;��H;�H;��H;Q�H;�H;�eH;΍G;J�E;�pB;�<;t�2;i�#;4�;���:T��:`+
9��y��W��	x����"��+4�Q�1���J���]�rmj�      @<ͼ}�ɼ�����֯�˶��ㄼ��Y��*�����s���X�,rѺ���?Q:0��:��
;o�#;��3;�c=;"$C;ADF; �G;.�H;�H;.�H;V�H;�H;w�H;C�H;��H;��H;��H;X�H;s�H;-�H;�H;*�H;�H;-�H;s�H;W�H;��H;��H;��H;@�H;w�H;�H;X�H;/�H; �H;+�H; �G;ADF;"$C;�c=;��3;l�#;��
;0��:�?Q:��,rѺ�X��s������*���Y�ㄼ˶���֯�����~�ɼ      ��'�(�$����|��  ���ۼ����+����]��X!�4>ۻp+��N*��깐�>:*��:2�;S�%;�5;��>;�(D;*�F;�!H;N�H;n�H;�H;��H;��H;�H;��H;��H;��H;��H;��H;��H;o�H;��H;o�H;��H;��H;��H;��H;��H;��H;�H;��H;��H;�H;p�H;J�H;�!H;*�F;�(D;��>;	�5;V�%;0�;*��:��>:��N*�p+��3>ۻ�X!���]��+�������ۼ�  �|����(�$�      Ƹ���v����w�g�c��J�΄-�{��;缃沼ㄼ|�;������j��x5�ؾ깼?Q:���:�i;N*;��8;��@;�PE;�uG;WiH;��H;��H;-�H;@�H;��H;��H;�H;�H;��H;��H;��H;��H;��H;��H;��H;��H;��H;�H;�H;��H;��H;@�H;-�H;��H;��H;TiH;�uG;�PE;��@;��8;N*;�i;���:�?Q:��x5��j������}�;�ㄼ�沼�;�{�΄-��J�g�c���w��v��      {Hͽتɽ�;��"����Ǹ����[�	z0�r��%<ͼȾ��[�J����j��M*���V��:�b�:r�;
�/;�L<;'C;GmF;��G;�H;"�H;*�H;(�H;]�H;o�H;�H;D�H;N�H;:�H;6�H;$�H;�H;$�H;6�H;<�H;O�H;D�H;�H;o�H;[�H;)�H;'�H;$�H;!�H;��G;CmF;'C;�L<;
�/;r�;�b�:V��:��K*��j����[�J�Ⱦ��%<ͼr��	z0���[�Ǹ����"���;��تɽ      ��#-������Ա�ƽ_P���v���J�H����ۼ
��[�J�����p+��,rѺ�+
9/N�:�;� $;#�5;�?;��D;y\G;fH;�H;��H;��H;��H;8�H;�H;q�H;��H;|�H;u�H;��H;Y�H;��H;t�H;{�H;��H;r�H;�H;8�H;��H;��H;��H;
�H;fH;w\G;��D;�?;%�5;� $;�;1N�:`+
9,rѺp+������[�J�
����ۼH���J��v��_P��ƽԱ轅����#-�       j�Xde�\0X��D�h{+�������x㻽Z���SDX������ۼȾ��}�;�2>ۻ�X���y��?":��:��;�-;��;;�B;�zF;�H;��H;��H;;�H;��H;�H;�H;��H;��H;��H;��H;��H;��H;��H;��H;��H;��H;��H;�H;�H;��H;;�H;��H;��H;�H;�zF;�B;��;;�-;��;��:�?":��y��X�2>ۻ~�;�Ⱦ����ۼ���SDX�Z���x㻽��콄��h{+��D�\0X�Xde�      ��Rh��m���I���|x���O��C(���Ъɽ����SDX�H��%<ͼㄼ�X!��s���W��rK����:�y;-�#;!I6;OR@;�PE;��G;��H;��H;G�H;�H;��H;��H;��H;��H;�H;��H;��H;��H;��H;��H;�H;��H;��H;��H;��H;�H;G�H;��H;��H;��G;�PE;NR@;!I6;0�#;�y;���:�rK��W��s���X!�ㄼ%<ͼH��SDX�����Ъɽ���C(���O��|x��I��m��Rh��      ?����������$�;jɰ��G�� j�9�5��	�ЪɽZ����J�r���沼��]�����	x�����n:��:�v;��/;�-=;��C;[�F;7IH;��H;;�H;��H;7�H;��H;��H;�H;"�H;)�H;2�H;A�H;2�H;)�H;#�H; �H;��H;��H;7�H;��H;=�H;��H;7IH;^�F;��C;�-=;��/;�v;	��:�n:����	x������]��沼r���J�Z���Ъɽ�	�9�5� j��G��jɰ�$�;��徹���      �2�W�-�"�.E�����AKɾl����s�9�5���w㻽�v��	z0��;��+���*����6�@5S��M�:z�	;��(;7�9;�/B;�DF;kH;�H;��H;��H;��H;��H;��H;,�H;O�H;]�H;W�H;v�H;\�H;\�H;P�H;,�H;��H;��H;��H;��H;��H;�H;iH;�DF;�/B;7�9;��(;|�	;�M�:@5S�6�����*��+���;�	z0��v��w㻽��9�5���s�l��AKɾ����.E�"�W�-�      (3s�!cm�<�\�j�C�7�%�����TҾl�� j��C(����_P����[�{������Y�#��9X���<��k:���:� ;�5;_R@;{uE;�G;I�H;_�H;��H;�H;_�H;��H;B�H;��H;��H;u�H;��H;u�H;��H;��H;@�H;��H;_�H;�H;��H;_�H;G�H;�G;}uE;]R@;�5;� ;���:�k:��<�8X�$����Y����{���[�_P����콬C(� j�l���TҾ���7�%�j�C�<�\�!cm�      �ޞ�������bF�@�W�X�-����AKɾ�G����O����ƽǸ��΄-���ۼㄼ+4�ǐ��ζ�$^:;��:�;Ė1;d>;��D;�\G;[sH;��H;��H;z�H;<�H;��H;G�H;��H;��H;��H;��H;��H;��H;��H;D�H;��H;<�H;w�H;~�H;��H;YsH;�\G;��D;d>;Ɩ1;�;E��:$^:�ζ�ǐ�,4�ㄼ��ۼτ-�Ǹ��ƽ�����O��G��AKɾ���X�-�A�W�bF�������      ��ſ���Nw���ޞ�����@�W�7�%�����jɰ��|x�h{+�ӱ����J��  �ʶ��P�1�����*��$
98�:̅;.�-;��<;��C;�G;�TH;e�H;�H;�H;��H;q�H;O�H;��H;��H;��H;�H;��H;��H;��H;N�H;r�H;��H;�H;�H;e�H;�TH;�G;��C;��<;1�-;΅;@�:p$
9�*����Q�1�˶���  ��J���ӱ�h{+��|x�jɰ�����7�%�@�W������ޞ�Nw�����      ����� �Կp���ޞ�bF�i�C�.E�$�;�I���D���"��g�c�|��֯���J��ѻ��)�p{K�^��:9�
;
N*;��:;�C;#�F;�8H;m�H;��H;��H;��H;[�H;W�H;��H;��H;��H;�H;��H;��H;��H;V�H;Y�H;��H;��H;��H;m�H;�8H;#�F;�C;��:;N*;9�
;f��:�{K���)��ѻ��J��֯�|�g�c�"�����D��I��$�;.E�i�C�bF��ޞ�p�� �Կ��      ��������� �ԿNw�����<�\�"����m��\0X�����;����w����������]��黣F����*ʒ:�;U�';׏9;9pB;�zF;�!H;��H;O�H;2�H;��H;b�H;W�H;��H;��H;��H;,�H;��H;��H;��H;V�H;b�H;��H;/�H;L�H;��H;�!H;�zF;9pB;ԏ9;X�';�;0ʒ:��깣F��黤�]����������w��;�����\0X�m�����"�<�\����Nw�� �Կ��𿞏�      !$�������忉�����!cm�W�-�����Rh��Xde�#-�تɽ�v��(�$�~�ɼpmj�)����X���(Ɔ:�x;^�%;J�8;�B;�RF;H;E�H;k�H;�H;��H;\�H;R�H;��H;��H;��H;A�H;��H;��H;��H;P�H;]�H;��H;�H;i�H;E�H;H;�RF;�B;G�8;d�%;�x;(Ɔ:���X�(���qmj�~�ɼ(�$��v��تɽ#-�Xde�Rh������W�-�!cm��������忞����      gܿ5�ֿ�aǿ?^��1���\o���7����iþ�(���-=��` �A���_�1]�-p���I�D�ѻ_�)�@�R���:Y�
;�*;6�:;�B;VIF;A�G;�lH;E�H;��H;z�H;��H;��H;��H;��H;C�H;��H;C�H;��H;��H;��H;��H;z�H;��H;B�H;�lH;C�G;VIF;�B;3�:;�*;Y�
;��:`�R�_�)�C�ѻ�I�-p��1]��_�A���` ��-=��(���iþ����7�\o�1���?^���aǿ5�ֿ      5�ֿEpѿ�¿������bXi�ҕ3��
�XD��Gl��B�9��.���R��#\� �cx��)�E��ͻ��$����	��:g�;��*;O�:;,�B;7UF;��G;fnH;�H;�H;��H;��H;��H;��H;��H;X�H;��H;X�H;��H;��H;��H;��H;��H;�H;ݡH;fnH;��G;6UF;,�B;J�:;��*;g�;��: ����$��ͻ*�E�cx�� �#\��R���.��B�9�Gl��XD���
�ҕ3�bXi��������¿Fpѿ      �aǿ�¿����������"Y��f'�����:o���.}��k/����&ڟ�$<Q�-#�ע��(;� ����� "7�1�:�;�,;��;;�C;VwF;5�G;�rH;l�H;ѸH;O�H;4�H;0�H;��H;��H;��H;�H;��H;��H;��H;.�H;5�H;O�H;θH;i�H;�rH;5�G;UwF;�C;��;;�,;�;1�: #7�������(;�ע�-#�$<Q�&ڟ�����k/��.}�:o�������f'��"Y�����������¿      ?^������l���\o���@�+�&�޾����;ce�2����ڽ����g@������R���O*�:G��ƛ���G^9f��:/;�d.;�<;אC;K�F;��G;�yH;ץH;H�H;^�H;��H;��H;�H;,�H;��H;O�H;��H;,�H;�H;��H;��H;^�H;G�H;ԥH;�yH;��G;K�F;ԐC;�<;�d.;/;h��:�G^9ƛ��8G���O*��R������g@�������ڽ1��;ce�����&�޾+���@�\o�l�������      1����������\o��!J�M�#��\��XD������|PH�����b�� C��� +���ټ%����ݿ��Ĭ��p�:g��:s�;�Y1;*>;�0D;��F;�H;��H;�H;<�H;��H;��H;C�H;��H;��H;��H;��H;��H;��H;��H;B�H;��H;��H;:�H;�H;��H;�H;��F;�0D;&>;�Y1;s�;i��:h�:Ƭ��ܿ����%����ټ� +� C���b�����|PH�����XD���\��M�#��!J�\o��������      \o�bXi��"Y���@�M�#��
��о�A���i���(����xr���_��5��ɺ�l�`��<��D�d���\�P�X:�P�:a;�4;�?;��D;�8G;�0H;֋H;��H;��H;B�H;��H;��H;5�H;��H;H�H;��H;H�H;��H;5�H;��H;��H;B�H;��H;��H;֋H;�0H;�8G;��D;ۧ?;�4;a;�P�:L�X:��\�B�d��<��l�`��ɺ��5��_�xr�������(��i��A���о�
�M�#���@��"Y�bXi�      ��7�ҕ3��f'�+��\���о�����.}��-=�}
���Ľ\��,:�����������7�GĻ��$��M��A��:�{;�D&;8,8;AJA;7�E;�G;�LH;"�H;��H;e�H;�H;B�H;��H;��H;Z�H;��H;R�H;��H;Z�H;��H;��H;C�H;�H;c�H;��H;"�H;�LH;�G;3�E;=JA;5,8;�D&;�{;9��:�M����$�GĻ��7���������,:�\����Ľ}
��-=��.}������о�\��+��f'�ҕ3�      ���
�����&�޾XD���A���.}�*�D�jt���ڽ�!��\����Z�ļ�
v�6�������IɺhT�9=��:C(;�-;Ƌ;;��B;�IF;��G;NfH;ٝH;-�H;`�H;�H;��H;��H;��H;��H;,�H;��H;,�H;��H;��H;��H;��H;�H;^�H;*�H;؝H;MfH;��G;�IF;��B;Ƌ;;�-;E(;;��:hT�9�Iɺ����6���
v�Z�ļ���\��!����ڽjt�*�D��.}��A��XD��&�޾�����
�      �iþXD��:o�����������i��-=�jt����R��jys�z +����w񗼌(;��ѻ�s@�4�!��4j:.Q�:�;�D3;u�>;EFD;��F;�	H;n|H;ϥH;��H;h�H;/�H;0�H;��H;X�H;n�H;��H;"�H;��H;n�H;W�H;��H;1�H;.�H;g�H;��H;ϥH;j|H;�	H;��F;BFD;t�>;�D3;�;,Q�:�4j:0�!��s@��ѻ�(;�w����z +�jys��R����jt��-=��i���������:o��XD��      �(��Gl���.}�;ce�|PH���(�}
���ڽ�R���{�D�6�� �+p��Z�`�Ũ��,���HҺ�N^9:�;�~(;c�8;JA;7|E;OjG;�=H;y�H;�H;b�H;��H;d�H;��H;��H;�H;��H;-�H;��H;-�H;��H;�H;��H;��H;d�H;��H;\�H;�H;x�H;�=H;LjG;5|E;JA;c�8;�~(;�;: O^9�HҺ�,��Ũ�Z�`�*p��� �C�6��{��R����ڽ}
���(�|PH�;ce��.}�Gl��      �-=�B�9��k/�2��������Ľ�!��jys�D�6�$#��ɺ��vz����/^��@�$�P}���r:f��:�;�Y1;2I=;ixC;]wF;_�G;AfH;��H;��H;��H;��H;��H;�H;�H;��H;��H;��H;��H;��H;��H;��H;�H;�H;��H;��H;��H;��H;~�H;?fH;Z�G;XwF;fxC;2I=;�Y1;�;f��:��r:P}�@�$�/^������vz��ɺ�$#�C�6�jys��!����Ľ����2���k/�B�9�      �` ��.�������ڽ�b��xr��\��\�z +�� ��ɺ�=��O*�4ͻ�5R��ƅ���:���:��;�);*u8;��@;�*E;�8G;�$H;��H;z�H;2�H;d�H;��H;��H;��H;:�H;��H;-�H;�H;\�H;�H;-�H;��H;:�H;��H;��H;��H;c�H;0�H;v�H;��H;}$H;�8G;�*E;��@;*u8;�);��;���:��:�ƅ��5R�4ͻ�O*�=��ɺ�� �z +�\�\��xr���b����ڽ��.��      A���R��&ڟ�����!C���_�,:�������+p���vz��O*��4ֻ�k�ګ����09��:61;�� ;�D3;{�=;�C;"lF;��G;]H;ؗH;��H;>�H;}�H;��H;��H;�H;6�H;G�H;��H;��H;��H;��H;��H;G�H;6�H;�H;��H;��H;|�H;>�H;��H;חH;�\H;��G;lF;�C;{�=;�D3;�� ;81;��:��09ګ���k��4ֻ�O*��vz�*p����輥��,:��_�!C������&ڟ��R��      �_�#\�#<Q�g@�� +��5�����Z�ļv�Z�`����4ͻ�k��Hɺ Z6���:<Q�:W�;e.;��:;V�A;d|E;�NG;'H;>�H;	�H;��H;��H;j�H;��H;��H;o�H;5�H;�H;L�H;��H;=�H;��H;L�H;�H;5�H;r�H;��H;��H;g�H;��H;��H;�H;<�H;|'H;�NG;c|E;V�A;��:;e.;[�;:Q�:��: Y6��Hɺ�k�3ͻ���Y�`�v�[�ļ�����5�� +�g@�#<Q�#\�      1]� �-#�������ټ�ɺ������
v��(;�ƨ�0^���5R�ޫ�� \6� ��:C��:.�;U�*;,8;�!@;��D;��F;6�G;fH;ęH;ͰH;޿H;��H;"�H;�H;_�H;��H;
�H;��H;��H;d�H;��H;d�H;��H;��H;
�H;��H;_�H; �H;�H;��H;ݿH;ͰH;H;fH;.�G;��F;��D;�!@;,8;X�*;,�;?��: ��: \6�ޫ���5R�0^��ƨ��(;��
v������ɺ���ټ����-#� �      -p��cx��
ע��R��&��m�`���7�7���ѻ�,��?�$��ƅ���09��:G��:�;(;�Z6;��>;�C;,IF;�G;)EH;��H;��H;�H;O�H;j�H;T�H;7�H;�H;��H;��H;M�H;(�H;��H;��H;��H;(�H;L�H;��H;��H;�H;7�H;N�H;h�H;M�H;�H;�H;��H;#EH;�G;)IF;�C;��>;�Z6;(;�;G��:��:��09�ƅ�?�$��,���ѻ7����7�l�`�&���R��
ע�cx��      �I�(�E��(;��O*����<��GĻ�����s@��HҺ@}�:��:8Q�:.�;(;B�5;�>;rC;q�E;�cG;z$H;8|H;x�H;^�H;��H;��H;y�H;�H;^�H;��H;��H;��H;��H;~�H;	�H;0�H;	�H;~�H;��H;��H;��H;��H;\�H;�H;y�H;��H;��H;]�H;s�H;2|H;z$H;�cG;t�E;rC;>;C�5;(;.�;:Q�:��:��:X}��HҺ�s@�����GĻ�<�����O*��(;�*�E�      H�ѻ�ͻ���9G��࿐�Q�d���$��Iɺ<�!��N^9��r:���:61;U�;V�*;�Z6;�>;n�B;��E;9G;�	H;?nH;W�H;��H;�H;��H;��H;�H;��H;A�H;��H;��H;=�H;9�H;��H;B�H;e�H;A�H;��H;9�H;<�H;��H;��H;@�H;��H;�H;��H;��H;�H;��H;S�H;?nH;�	H; 9G;��E;n�B; >;�Z6;V�*;W�;61;���:��r:�N^90�!��Iɺ��$�L�d�ݿ��8G������ͻ      X�)���$���ƛ��Ԭ����\��M��HT�9�4j:釶:f��:��;�� ;e.;,8;��>;oC;��E;�)G;��G;RdH;��H;֫H;��H;��H;x�H;�H;�H;��H;��H;��H;��H;��H;��H;=�H;r�H;��H;r�H;=�H;��H;��H;��H;��H;��H;��H;�H;�H;x�H;��H;��H;ҫH;��H;NdH;��G;�)G;êE;oC;��>;,8;e.;�� ;��;b��::�4j:HT�9�M����\�Ȭ��ě������$�      @�R� �� "7��G^9\�:@�X:5��:/��:&Q�:�;�;�);�D3;��:;�!@;�C;p�E;9G;��G;�`H;��H;Y�H;[�H;��H;��H;v�H;��H;��H;��H;�H;��H;I�H;)�H;��H;j�H;��H;��H;��H;k�H;��H;(�H;J�H;��H;�H;��H;��H;��H;u�H;��H;��H;X�H;Y�H;��H;�`H;��G;9G;p�E;�C;�!@;��:;�D3;�);�;�;&Q�:/��:5��:L�X:��:�G^9 "7����      ��:'��:3�:T��:S��:�P�:�{;@(;�;�~(;�Y1;&u8;x�=;T�A;��D;(IF;�cG;�	H;QdH;��H;��H;�H;q�H;4�H;�H;��H;��H;��H;e�H;&�H;��H;��H;��H;&�H;��H;��H;��H;��H;��H;&�H;��H;��H;��H;#�H;b�H;��H;��H;��H;�H;0�H;r�H;�H;��H;��H;RdH;�	H;�cG;)IF;��D;V�A;z�=;'u8;�Y1;�~(;�;@(;�{;Q�:U��:X��:3�:��:      ]�
;��;)�;$;r�;a;�D&;�-;�D3;d�8;8I=;��@;�C;d|E;��F;�G;z$H;?nH;��H;[�H;�H;��H;z�H;_�H;��H;��H;$�H;��H;��H;I�H;_�H;5�H;��H;]�H;��H;��H;��H;��H;��H;]�H;��H;6�H;a�H;E�H;��H;��H;!�H;��H;��H;[�H;x�H;��H;�H;\�H;��H;@nH;z$H;�G;��F;d|E;�C;��@;6I=;f�8;�D3;�-;�D&;a;��;$;*�;|�;      �*;��*;�,;�d.;�Y1;�4;8,8;ċ;;u�>;JA;ixC;�*E;lF;�NG;4�G;%EH;5|H;W�H;իH;]�H;r�H;{�H;�H;:�H;7�H;��H;M�H;+�H;��H;�H;��H;��H;"�H;y�H;��H;��H;��H;��H;��H;y�H;"�H;��H;��H;�H;��H;+�H;J�H;��H;9�H;9�H;�H;|�H;n�H;`�H;֫H;W�H;3|H;%EH;4�G;�NG;lF;�*E;gxC;JA;u�>;ċ;;9,8;�4;�Y1;�d.;�,;��*;      H�:;X�:;��;;�<;)>;ݧ?;GJA;��B;EFD;5|E;\wF;�8G;��G;'H;fH;��H;w�H;��H;��H;��H;/�H;\�H;9�H;$�H;Z�H;��H;��H;r�H;��H;��H;V�H;��H;\�H;��H;��H;��H;�H;��H;��H;��H;Y�H;��H;V�H;��H;��H;t�H;��H;��H;[�H;!�H;9�H;_�H;/�H;��H;��H;��H;u�H;��H;fH;�'H;��G;�8G;ZwF;5|E;FFD;��B;EJA;ݧ?;1>;�<;��;;L�:;      ��B;6�B;�C;ؐC;�0D;��D;5�E;�IF;��F;LjG;\�G;�$H; ]H;@�H;řH;��H;b�H;�H;��H;��H;�H;��H;=�H;_�H;��H;��H;:�H;��H;i�H;6�H;��H;�H;m�H;��H;��H;��H;��H;��H;��H;��H;m�H;�H;��H;5�H;f�H;��H;:�H;��H;��H;^�H;<�H;��H;�H;��H;��H;�H;a�H;��H;řH;?�H; ]H;�$H;\�G;IjG;��F;�IF;6�E;��D;�0D;ڐC;�C;7�B;      aIF;DUF;JwF;E�F;��F;�8G;�G;��G;�	H;�=H;?fH;��H;՗H;�H;ʰH;�H;��H;��H;t�H;t�H;|�H;��H;��H;��H;��H;7�H;g�H;J�H;��H;��H;�H;`�H;t�H;��H;��H;��H;��H;��H;��H;��H;r�H;a�H;�H;��H;��H;J�H;d�H;:�H;��H;��H;��H;��H;x�H;u�H;u�H;��H;��H;�H;˰H;�H;՗H;��H;?fH;�=H;�	H;��G;�G;�8G;��F;H�F;LwF;7UF;      N�G;��G;5�G;��G;�H;�0H;�LH;NfH;n|H;y�H;~�H;{�H;��H;��H;ݿH;O�H;��H;��H;�H;��H;��H;"�H;L�H;��H;4�H;i�H;<�H;��H;��H;��H;!�H;m�H;��H;��H;��H;��H;��H;��H;��H;��H;��H;n�H;!�H;��H;��H;��H;;�H;h�H;:�H;��H;J�H;$�H;��H;��H;�H;��H;��H;M�H;ݿH;��H;��H;{�H;~�H;w�H;p|H;MfH;�LH;�0H;�H;��G;6�G;��G;      �lH;hnH;�rH;�yH;��H;؋H;(�H;��H;ӥH;�H;��H;7�H;>�H;��H;��H;j�H;x�H;�H;�H;��H;��H;��H;)�H;u�H;|�H;L�H;��H;r�H;��H;*�H;G�H;v�H;��H;��H;��H;��H;��H;��H;��H;��H;��H;x�H;H�H;&�H;��H;r�H;��H;L�H;~�H;v�H;+�H;��H;��H;��H;�H;�H;x�H;j�H;��H;��H;<�H;6�H;��H;�H;ԥH;�H;(�H;֋H;��H;�yH;�rH;snH;      Z�H;�H;g�H;ۥH;�H;��H;��H;/�H;��H;c�H;��H;h�H;}�H;h�H;!�H;R�H;�H;��H;��H;��H;c�H;��H;��H;��H;b�H;�H;��H;��H;
�H;N�H;j�H;��H;��H;��H;��H;��H;��H;��H;��H;��H;��H;��H;k�H;N�H;
�H;��H;��H;��H;e�H;��H;��H;��H;b�H;��H;��H;��H;�H;T�H;!�H;h�H;}�H;e�H;��H;`�H;��H;.�H;°H;��H;�H;ۥH;j�H;ܡH;      ��H;��H;ڸH;J�H;J�H;��H;l�H;e�H;r�H;��H;��H;��H;��H;��H;�H;:�H;_�H;;�H;��H;�H;#�H;E�H;�H;��H;,�H;��H;��H;(�H;N�H;a�H;��H;�H;��H;��H;��H;��H;��H;��H;��H;��H;��H;��H;��H;a�H;L�H;(�H;��H;��H;.�H;��H;�H;F�H;%�H;�H;��H;=�H;^�H;:�H;�H;��H;��H;��H;��H;��H;t�H;h�H;j�H;��H;H�H;K�H;׸H;�H;      �H;��H;\�H;g�H;��H;A�H; �H;�H;6�H;j�H;��H;��H;��H;��H;c�H;�H;��H;��H;��H;��H;��H;_�H;��H;[�H;��H;�H;�H;I�H;j�H;��H;��H;��H;{�H;}�H;��H;��H;m�H;��H;��H;}�H;x�H;��H;��H;��H;m�H;I�H;�H;�H;��H;Y�H;��H;a�H;��H;��H;��H;��H;��H;�H;c�H;��H;��H;��H;��H;j�H;8�H;�H; �H;D�H;��H;i�H;]�H;��H;      ��H;��H;<�H;��H;��H;��H;D�H;��H;5�H;��H;#�H;��H;�H;x�H;��H;��H;��H;��H;��H;S�H;��H;9�H;��H;��H;�H;`�H;m�H;y�H;��H;��H;��H;��H;|�H;v�H;��H;n�H;d�H;n�H;��H;v�H;y�H;��H;��H;��H;��H;y�H;m�H;^�H;�H;��H;��H;:�H;��H;S�H;��H;��H;��H;��H;��H;y�H;�H;��H;#�H;��H;7�H;��H;D�H;��H;��H;��H;=�H;��H;      ��H;��H;8�H;��H;N�H;��H;��H;��H;��H;��H;�H;E�H;<�H;:�H;�H;��H;��H;9�H;��H;.�H;��H;��H;#�H;`�H;h�H;u�H;��H;��H;��H;��H;{�H;�H;��H;�H;]�H;]�H;��H;]�H;]�H;�H;}�H;��H;{�H;��H;��H;��H;��H;t�H;j�H;`�H;"�H;��H;��H;/�H;��H;<�H;��H;��H;�H;:�H;;�H;C�H;�H;��H;��H;��H;��H;�H;G�H;��H;8�H;��H;      ��H;��H;��H;�H;��H;/�H;��H;��H;]�H;�H;��H;��H;K�H;�H;��H;U�H;��H;:�H;��H;��H;,�H;`�H;y�H;��H;��H;��H;��H;��H;��H;��H;|�H;x�H;{�H;h�H;Y�H;^�H;c�H;^�H;Y�H;h�H;y�H;{�H;|�H;��H;��H;��H;��H;��H;��H;��H;y�H;`�H;,�H;��H;��H;<�H;��H;U�H;��H;�H;K�H;��H;��H;�H;`�H;��H;��H;3�H;��H;�H;��H;��H;      ��H;��H;��H;4�H;��H;��H;c�H;��H;w�H;�H;��H;;�H;��H;S�H;��H;2�H;��H;��H;>�H;t�H;��H;��H;��H;��H;��H;��H;��H;��H;��H;��H;��H;��H;\�H;Y�H;d�H;Y�H;=�H;Y�H;d�H;Z�H;Y�H;��H;��H;��H;��H;��H;��H;��H;��H;��H;��H;��H;��H;t�H;>�H;��H;��H;2�H;��H;S�H;��H;;�H;��H;�H;w�H;��H;c�H;��H;��H;5�H;��H;��H;      =�H;c�H;��H;��H;��H;C�H;��H;7�H;��H;.�H;��H;*�H;��H;��H;k�H;��H;�H;=�H;u�H;��H;��H;��H;��H;��H;��H;��H;��H;��H;��H;��H;��H;r�H;\�H;c�H;Z�H;V�H;E�H;V�H;Z�H;`�H;Z�H;u�H;��H;��H;��H;��H;��H;��H;��H;��H;��H;��H;��H;��H;u�H;>�H;�H;��H;j�H;��H;��H;*�H;��H;1�H;��H;6�H;��H;G�H;��H;��H;��H;[�H;      ��H;�H;�H;R�H;��H;��H;W�H;��H;)�H;��H;��H;i�H;��H;D�H;��H;��H;7�H;^�H;��H;��H;��H;��H;��H;�H;��H;��H;��H;��H;��H;��H;o�H;k�H;��H;e�H;=�H;G�H;@�H;G�H;=�H;e�H;��H;m�H;o�H;��H;��H;��H;��H;��H;��H;�H;��H;��H;��H;��H;��H;`�H;6�H;��H;��H;D�H;��H;i�H;��H;��H;*�H;��H;W�H;��H;��H;R�H;�H;�H;      =�H;c�H;��H;��H;��H;C�H;��H;7�H;��H;.�H;��H;*�H;��H;��H;j�H;��H;�H;=�H;u�H;��H;��H;��H;��H;��H;��H;��H;��H;��H;��H;��H;��H;r�H;\�H;c�H;Z�H;V�H;E�H;V�H;Z�H;`�H;Z�H;u�H;��H;��H;��H;��H;��H;��H;��H;��H;��H;��H;��H;��H;u�H;>�H;�H;��H;k�H;��H;��H;*�H;��H;0�H;��H;6�H;��H;G�H;��H;��H;��H;Z�H;      ��H;��H;��H;5�H;��H;��H;b�H;��H;w�H;�H;��H;;�H;��H;S�H;��H;2�H;��H;��H;>�H;t�H;��H;��H;��H;��H;��H;��H;��H;��H;��H;��H;��H;��H;\�H;Z�H;d�H;Y�H;=�H;Y�H;d�H;Y�H;Y�H;��H;��H;��H;��H;��H;��H;��H;��H;��H;��H;��H;��H;t�H;>�H;��H;��H;2�H;��H;S�H;��H;;�H;��H;�H;w�H;��H;c�H;��H;��H;5�H;��H;��H;      ��H;��H;��H;�H;��H;/�H;��H;��H;]�H;�H;��H;��H;K�H;
�H;��H;U�H;��H;:�H;��H;��H;/�H;`�H;y�H;��H;��H;��H;��H;��H;��H;��H;|�H;x�H;{�H;h�H;Y�H;^�H;c�H;^�H;Y�H;h�H;y�H;{�H;|�H;��H;��H;��H;��H;��H;��H;��H;y�H;`�H;,�H;��H;��H;<�H;��H;U�H;��H;�H;K�H;��H;��H;�H;^�H;��H;��H;3�H;��H;�H;��H;��H;      ��H;��H;:�H;��H;N�H;��H;��H;��H;��H;��H;�H;C�H;;�H;:�H;�H;��H;��H;9�H;��H;.�H;��H;��H;#�H;`�H;j�H;u�H;��H;��H;��H;��H;{�H;�H;�H;}�H;]�H;]�H;��H;\�H;]�H;}�H;}�H;��H;{�H;��H;��H;��H;��H;t�H;h�H;^�H;"�H;��H;��H;/�H;��H;;�H;��H;��H;�H;:�H;;�H;E�H;�H;��H;��H;��H;��H;�H;F�H;��H;5�H;��H;      ��H;��H;=�H;��H;��H;��H;I�H;��H;5�H;��H;#�H;��H;�H;x�H;��H;��H;��H;��H;��H;S�H;��H;:�H;��H;��H;�H;`�H;m�H;y�H;��H;��H;��H;��H;y�H;v�H;��H;n�H;d�H;n�H;��H;v�H;y�H;��H;��H;��H;��H;y�H;m�H;^�H;�H;��H;��H;9�H;��H;S�H;��H;��H;��H;��H;��H;x�H;�H;��H;"�H;��H;7�H;��H;G�H;��H;��H;��H;=�H;��H;      �H;��H;\�H;i�H;��H;A�H; �H;�H;8�H;h�H;��H;��H;��H;��H;c�H;�H;��H;��H;��H;��H;��H;a�H;��H;\�H;��H;�H;�H;I�H;j�H;��H;��H;��H;y�H;}�H;��H;��H;m�H;��H;��H;}�H;x�H;��H;��H;��H;k�H;I�H;�H;�H;��H;Y�H;��H;_�H;��H;��H;��H;��H;��H;�H;c�H;��H;��H;��H;��H;k�H;8�H;�H; �H;D�H;��H;g�H;\�H;��H;      ��H;��H;ڸH;J�H;H�H;��H;m�H;h�H;r�H;��H;��H;��H;��H;��H;�H;:�H;_�H;;�H;��H;�H;(�H;F�H;�H;��H;.�H;��H;��H;(�H;L�H;c�H;��H;�H;��H;��H;��H;��H;��H;��H;��H;��H;��H;��H;��H;`�H;N�H;(�H;��H;��H;,�H;��H;�H;E�H;#�H;�H;��H;=�H;^�H;;�H;�H;��H;��H;��H;��H;��H;u�H;i�H;m�H;��H;F�H;J�H;ظH;�H;      S�H;�H;m�H;ڥH;�H;��H;İH;/�H;��H;`�H;��H;g�H;}�H;h�H;!�H;T�H;�H;��H;��H;��H;h�H;��H;��H;��H;e�H;�H;��H;��H;	�H;O�H;k�H;��H;��H;��H;��H;��H;��H;��H;��H;��H;��H;��H;j�H;L�H;
�H;��H;��H;��H;b�H;��H;��H;��H;b�H;��H;��H;��H;�H;T�H;!�H;h�H;}�H;h�H;��H;b�H;��H;/�H;İH;��H;�H;֥H;q�H;ߡH;      �lH;inH;�rH;�yH;��H;֋H;(�H;�H;ӥH;�H;��H;6�H;<�H;��H;��H;j�H;y�H;�H;�H;��H;��H;��H;+�H;v�H;~�H;J�H;��H;r�H;��H;*�H;H�H;x�H;��H;��H;��H;��H;��H;��H;��H;��H;��H;x�H;G�H;(�H;��H;r�H;��H;L�H;|�H;u�H;(�H;��H;��H;��H;�H;�H;v�H;k�H;��H;��H;>�H;6�H;��H;�H;ԥH;�H;(�H;ՋH;��H;�yH;�rH;qnH;      H�G;��G;6�G;��G;�H;�0H;�LH;NfH;n|H;x�H;~�H;{�H;��H;��H;ݿH;N�H;��H;��H;�H;��H;��H;$�H;L�H;��H;:�H;h�H;<�H;��H;��H;��H;!�H;n�H;��H;��H;��H;��H;��H;��H;��H;��H;��H;n�H;!�H;��H;��H;��H;;�H;i�H;4�H;��H;J�H;"�H;��H;��H;�H;��H;��H;N�H;ݿH;��H;��H;{�H;��H;x�H;p|H;NfH;�LH;�0H;�H;��G;4�G;��G;      gIF;AUF;UwF;I�F;��F;�8G;�G;��G;�	H;�=H;?fH;��H;՗H;�H;ʰH;�H;��H;��H;u�H;u�H;}�H;��H;��H;��H;��H;9�H;g�H;J�H;��H;��H;�H;`�H;t�H;��H;��H;��H;��H;��H;��H;��H;q�H;a�H;�H;��H;��H;J�H;e�H;9�H;��H;��H;��H;��H;y�H;t�H;t�H;��H;��H;�H;ʰH;�H;ԗH;��H;?fH;�=H;�	H;��G;�G;�8G;��F;G�F;UwF;3UF;      ��B;6�B;�C;ڐC;�0D;��D;6�E;�IF;��F;KjG;]�G;�$H; ]H;?�H;řH;��H;b�H;�H;��H;��H;�H;��H;=�H;_�H;��H;��H;;�H;��H;i�H;6�H;��H;�H;m�H;��H;��H;��H;��H;��H;��H;��H;k�H;�H;��H;5�H;f�H;��H;9�H;��H;��H;_�H;<�H;��H;�H;��H;��H;�H;`�H;��H;řH;?�H; ]H;�$H;\�G;KjG;��F;�IF;5�E;��D;�0D;ؐC;�C;6�B;      K�:;W�:;��;;�<;&>;�?;BJA;��B;GFD;7|E;\wF;�8G;��G;�'H;fH;��H;w�H;��H;��H;��H;2�H;_�H;:�H;$�H;[�H;��H;��H;t�H;��H;��H;V�H;��H;Z�H;��H;��H;��H;�H;��H;��H;��H;Z�H;��H;V�H;��H;��H;r�H;��H;��H;Z�H;"�H;7�H;\�H;-�H;��H;��H;��H;u�H;��H;fH;~'H;��G;�8G;ZwF;3|E;FFD;��B;AJA;�?;4>;�<;��;;I�:;      �*;��*;�,;�d.;�Y1;�4;=,8;ċ;;u�>;JA;gxC;�*E;lF;�NG;4�G;&EH;5|H;U�H;֫H;^�H;t�H;|�H;�H;<�H;9�H;��H;M�H;+�H;��H;�H;��H;��H;"�H;y�H;��H;��H;��H;��H;��H;y�H;!�H;��H;��H;�H;��H;+�H;J�H;��H;7�H;7�H; �H;{�H;n�H;^�H;իH;Y�H;5|H;%EH;5�G;�NG;lF;�*E;gxC;JA;u�>;Ƌ;;=,8;�4;�Y1;�d.;�,;��*;      ]�
;��;'�;$;t�;a;�D&;�-;�D3;f�8;8I=;��@;�C;d|E;��F;�G;x$H;?nH;��H;[�H;�H;��H;z�H;_�H;��H;��H;$�H;��H;��H;I�H;a�H;6�H;��H;]�H;��H;��H;��H;��H;��H;]�H;��H;5�H;_�H;E�H;��H;��H;!�H;��H;��H;\�H;w�H;��H;�H;\�H;��H;@nH;x$H;�G;��F;d|E;�C;��@;6I=;d�8;�D3;�-;�D&;a;��;$;)�;{�;      ��:��:;�:X��:U��:�P�:�{;C(;�;�~(;�Y1;'u8;x�=;V�A;��D;)IF;�cG;�	H;RdH;��H;��H;�H;t�H;4�H;�H;��H;��H;��H;c�H;&�H;��H;��H;��H;%�H;��H;��H;��H;��H;��H;&�H;��H;��H;��H;#�H;b�H;��H;��H;��H;�H;0�H;p�H;�H;��H;��H;QdH;�	H;�cG;(IF;��D;T�A;z�=;&u8;�Y1;�~(;�;C(;�{;�P�:]��:T��:?�:��:      P�R� �� 7�pG^9t�:<�X:;��:1��:,Q�:�;�;�);�D3;��:;�!@;�C;p�E;9G;��G;�`H;��H;Y�H;[�H;��H;��H;u�H;��H;��H;��H;�H;��H;I�H;)�H;��H;k�H;��H;��H;��H;j�H;��H;(�H;J�H;��H;�H;��H;��H;��H;v�H;��H;��H;X�H;Y�H;��H;�`H;��G;9G;p�E;�C;�!@;��:;�D3;�);�;�;*Q�:7��:9��:L�X:��:pG^9 7����      X�)���$���ě��Ь����\��M��HT�9�4j::f��:��;�� ;e.;,8;��>;oC;��E;�)G;��G;QdH;��H;֫H;��H;��H;w�H;�H;�H;��H;��H;��H;��H;��H;��H;=�H;r�H;��H;r�H;=�H;��H;��H;��H;��H;��H;��H;�H;	�H;x�H;��H;��H;ҫH;��H;OdH;��G;�)G;êE;nC;��>;,8;e.;�� ;��;f��:釶:�4j:PT�9�M����\�Ƭ��ƛ������$�      G�ѻ�ͻ���9G��࿐�Q�d���$��Iɺ<�!��N^9��r:���:61;U�;V�*;�Z6; >;m�B;��E;9G;�	H;?nH;W�H;��H;�H;��H;��H;�H;��H;A�H;��H;��H;=�H;9�H;��H;B�H;e�H;B�H;��H;9�H;<�H;��H;��H;@�H;��H;�H;��H;��H;�H;��H;U�H;?nH;�	H; 9G;��E;n�B;�>;�Z6;V�*;U�;61;���:��r:�N^90�!��Iɺ��$�N�d�ܿ��:G������ͻ      �I�(�E��(;��O*����<��GĻ�����s@��HҺ@}�:��::Q�:.�;(;C�5; >;qC;r�E;�cG;z$H;8|H;w�H;]�H;��H;��H;y�H;�H;^�H;��H;��H;��H;��H;~�H;
�H;0�H;	�H;~�H;��H;��H;��H;��H;\�H;�H;y�H;��H;��H;^�H;t�H;2|H;z$H;�cG;t�E;rC;>;C�5;(;.�;8Q�:��:��:P}��HҺ�s@�����GĻ�<�����O*��(;�+�E�      -p��cx��
ע��R��&��m�`���7�6���ѻ�,��?�$��ƅ���09��:G��:�;(;�Z6;��>;�C;+IF;�G;&EH;��H;�H;�H;O�H;h�H;R�H;7�H;�H;��H;��H;L�H;(�H;��H;��H;��H;(�H;M�H;��H;��H;�H;7�H;O�H;j�H;M�H;�H;��H;��H;#EH;�G;)IF;�C;��>;�Z6;(;�;G��:��:��09�ƅ�?�$��,���ѻ6����7�l�`�&���R��
ע�cx��      1]� �-#�������ټ�ɺ������
v��(;�ƨ�0^���5R�ޫ�� \6�"��:?��:.�;S�*;,8;�!@;��D;��F;5�G;fH;��H;ʰH;޿H;��H;"�H;�H;_�H;��H;
�H;��H;��H;d�H;��H;d�H;��H;��H;
�H;��H;_�H; �H;�H;��H;ݿH;ΰH;ęH;fH;1�G;��F;��D;�!@;,8;X�*;,�;C��: ��: \6�ޫ���5R�0^��ƨ��(;��
v������ɺ���ټ����-#� �      �_�"\�#<Q�g@�� +��5�����Z�ļv�Y�`����4ͻ�k��Hɺ Y6���:<Q�:Z�;e.;��:;T�A;c|E;�NG;'H;<�H;�H;��H;��H;g�H;��H;��H;o�H;6�H;�H;L�H;��H;=�H;��H;L�H;�H;3�H;q�H;��H;��H;h�H;��H;��H;
�H;>�H;|'H;�NG;d|E;W�A;��:;e.;Z�;:Q�:��: Z6��Hɺ�k�4ͻ���Y�`�v�[�ļ�����5�� +�g@�#<Q�#\�      A���R��&ڟ�����!C���_�,:�������*p���vz��O*��4ֻ�k�ګ����09��:61;�� ;�D3;z�=;�C;!lF;��G;�\H;חH;��H;>�H;}�H;��H;��H;�H;6�H;G�H;��H;��H;��H;��H;��H;G�H;5�H;�H;��H;��H;{�H;>�H;��H;ڗH;]H;��G;lF;�C;{�=;�D3;�� ;81;��:��09ث���k��4ֻ�O*��vz�+p����輥��,:��_�!C������&ڟ��R��      �` ��.�������ڽ�b��xr��\��\�z +�� ��ɺ�=��O*�4ͻ�5R��ƅ���:���:��;�);&u8;��@;�*E;�8G;}$H;��H;y�H;0�H;d�H;��H;��H;��H;;�H;��H;-�H; �H;\�H; �H;-�H;��H;8�H;��H;��H;��H;c�H;2�H;y�H;��H;�$H;�8G;�*E;��@;*u8;�);��;���:��:�ƅ��5R�4ͻ�O*�=��ɺ�� �z +�\�\��xr���b����ڽ��.��      �-=�B�9��k/�2��������Ľ�!��jys�C�6�$#��ɺ��vz����.^��@�$�@}���r:f��:�;�Y1;2I=;ixC;\wF;Z�G;@fH;��H;��H;��H;��H;��H;�H;�H;��H;��H;��H;��H;��H;��H;��H;�H;�H;��H;��H;��H;��H;~�H;AfH;_�G;YwF;fxC;2I=;�Y1;�;f��:��r:X}�A�$�/^������vz��ɺ�$#�C�6�jys��!����Ľ����2���k/�B�9�      �(��Gl���.}�;ce�|PH���(�}
���ڽ�R���{�D�6�� �*p��Z�`�Ũ��,���HҺ�N^9:�;�~(;c�8;JA;7|E;LjG;�=H;y�H;�H;_�H;��H;d�H;��H;��H;�H;��H;-�H;��H;-�H;��H;�H;��H;��H;d�H;��H;]�H;�H;x�H;�=H;OjG;5|E;JA;c�8;�~(;�;: O^9�HҺ�,��Ũ�Z�`�+p��� �D�6��{��R����ڽ}
���(�|PH�;ce��.}�Gl��      �iþXD��:o�����������i��-=�jt����R��jys�z +����w񗼌(;��ѻ�s@�4�!��4j:.Q�:�;�D3;u�>;EFD;��F;�	H;m|H;ϥH;��H;g�H;.�H;0�H;��H;W�H;n�H;��H;"�H;��H;n�H;X�H;��H;0�H;/�H;g�H;��H;ϥH;l|H;�	H;��F;CFD;t�>;�D3;�;,Q�:�4j:0�!��s@��ѻ�(;�w����z +�jys��R����jt��-=��i���������:o��XD��      ���
�����&�޾XD���A���.}�*�D�jt���ڽ�!��\����Z�ļ�
v�6�������IɺhT�9=��:B(;�-;Ƌ;;��B;�IF;��G;NfH;؝H;-�H;^�H;�H;��H;��H;��H;��H;,�H;��H;-�H;��H;��H;��H;��H;�H;`�H;*�H;ٝH;MfH;��G;�IF;��B;Ƌ;;�-;E(;;��:hT�9�Iɺ����6���
v�Z�ļ���\��!����ڽjt�*�D��.}��A��XD��&�޾�����
�      ��7�ҕ3��f'�+��\���о�����.}��-=�}
���Ľ\��,:�����������7�GĻ��$��M��;��:�{;�D&;8,8;AJA;3�E;�G;�LH;"�H;��H;e�H;�H;B�H;��H;��H;Z�H;��H;R�H;��H;Z�H;��H;��H;B�H;�H;c�H;��H;"�H;�LH;�G;7�E;>JA;6,8;�D&;�{;;��:�M����$�GĻ��7���������,:�\����Ľ}
��-=��.}������о�\��+��f'�ҕ3�      \o�bXi��"Y���@�M�#��
��о�A���i���(����xr���_��5��ɺ�l�`��<��C�d���\�L�X:�P�:a;�4;�?;��D;�8G;�0H;֋H;��H;��H;B�H;��H;�H;5�H;��H;H�H;��H;J�H;��H;5�H;��H;��H;B�H;��H;��H;֋H;�0H;�8G;��D;ݧ?;�4;a;�P�:L�X:��\�B�d��<��l�`��ɺ��5��_�xr�������(��i��A���о�
�M�#���@��"Y�bXi�      1����������\o��!J�M�#��\��XD������|PH�����b�� C��� +���ټ%����ݿ��Ƭ��h�:a��:s�;�Y1;*>;�0D;��F;�H;��H;�H;<�H;��H;��H;C�H;��H;��H;��H;��H;��H;��H;��H;B�H;��H;��H;:�H;�H;��H;�H;��F;�0D;'>;�Y1;s�;i��:h�:Ĭ��ܿ����%����ټ� +� C���b�����|PH�����XD���\��M�#��!J�\o��������      ?^������l���\o���@�+�&�޾����;ce�1����ڽ����g@������R���O*�9G��ƛ���G^9b��:/;�d.;�<;ԐC;K�F;��G;�yH;֥H;J�H;^�H;��H;��H;�H;,�H;��H;O�H;��H;,�H;�H;��H;��H;^�H;G�H;ԥH;�yH;��G;K�F;אC;�<;�d.;/;h��:�G^9ƛ��8G���O*��R������g@�������ڽ2��;ce�����&�޾+���@�\o�l�������      �aǿ�¿����������"Y��f'�����:o���.}��k/����&ڟ�$<Q�-#�ע��(;������ #7�+�:�;�,;��;;�C;VwF;5�G;�rH;l�H;ѸH;O�H;4�H;0�H;��H;��H;��H;�H;��H;��H;��H;.�H;5�H;O�H;θH;i�H;�rH;5�G;UwF;�C;��;;�,;�;1�: #7�������(;�ע�-#�$<Q�&ڟ�����k/��.}�:o�������f'��"Y�����������¿      5�ֿEpѿ�¿������bXi�ҕ3��
�XD��Gl��B�9��.���R��#\� �bx��)�E��ͻ��$���	��:g�;��*;O�:;,�B;7UF;��G;fnH;�H;�H;��H;��H;��H;��H;��H;X�H;��H;X�H;��H;��H;��H;��H;��H;�H;ݡH;fnH;��G;6UF;,�B;L�:;��*;g�;��: ����$��ͻ*�E�cx�� �#\��R���.��B�9�Gl��XD���
�ҕ3�bXi��������¿Epѿ      �?��~h��?v��� ��:�X��O/�1y�C�;Ⱆ��+X����ѽ����an;�]�������B(�К���� �e9D�:;�Y.;j�<;�WC;9[F;�G;;0H;�jH;d�H;��H;ǵH;_�H;��H;��H;��H;��H;��H;��H;��H;]�H;ɵH;��H;b�H;~jH;;0H;�G;7[F;�WC;g�<;�Y.;;F�: �e9��Κ���B(�����]��an;������ѽ���+X�Ⱆ�C�;1y��O/�:�X�� ��?v��~h��      ~h��1���c�����y�YvS�rM+��v�9ɾ�����T�"]�\ν����z\8�����x���%�D���6��@�9�-�:��;��.;3�<;oC;�dF;�G;�1H;0kH;֌H;�H;�H;��H;�H;��H;�H;��H;�H;��H;�H;��H;�H;�H;ьH;-kH;�1H;�G;�dF;oC;/�<;��.;��;�-�:0�96��D����%��x�����z\8�����\ν"]��T�����9ɾ�v�rM+�YvS���y�c���1���      ?v��c���X ��c�h�8E�Y��l���~㼾���nH�Ո�{�ý�Ȅ��s/��o��#�����J���кH�9�g�:m;m0;9]=;�C;2�F;��G;W6H;lmH;V�H;ߥH;ǶH;6�H;|�H;�H;?�H;�H;?�H;	�H;|�H;4�H;ǶH;ߥH;Q�H;imH;W6H;��G;1�F;�C;5]=;p0;m;�g�:0�9�кJ������#���o��s/��Ȅ�{�ýՈ��nH���~㼾l���Y��8E�c�h�X ��c���      � ����y�c�h��N��O/����D�߾B���*|��6�r}�䳽lSt�>�!�qrμ@F{��_��X������8 :X��:[;�2;�O>;�D;~�F;��G;S=H;�pH;��H;��H;�H;�H;�H;��H;��H;��H;��H;��H;�H;�H;�H;��H;��H;�pH;S=H;��G;{�F;�D;�O>;�2;[;^��:0 :�����X���_�@F{�qrμ=�!�lSt�䳽r}��6��*|�B��D�߾����O/��N�c�h���y�      :�X�YvS�8E��O/��S�JW����������NS\��� ���<����Y�{��Ѓ����]�w����b��Y�0�Y:��:�`;|�4;�?;v�D;�F;1�G;@FH;�uH;�H;ʩH;ǹH;M�H;�H;]�H;S�H;3�H;S�H;[�H;�H;L�H;ɹH;ʩH;�H;�uH;@FH;1�G;�F;u�D;�?;~�4;�`;��:(�Y:�Y�
�b�x�����]�Ѓ��{���Y�<����当� �NS\���������JW���S��O/�8E�YvS�      �O/�rM+�Y�����JW��9ɾC���Mw�� :�k��y�ý�L��^n;�`���sv���E<��˻��-����y�:�^;�%;7;��@;Q5E;�"G;2�G;tPH;D{H;�H;��H;��H;��H;2�H;K�H; �H;��H; �H;K�H;0�H;��H;��H;��H;�H;@{H;tPH;0�G;�"G;O5E;��@;7;�%;�^;�y�:����-��˻�E<�sv��_���^n;��L��y�ýk��� :��Mw�C��9ɾJW�����Y��rM+�      1y��v�l���E�߾����C��@����nH���F὞u����d�0O�jrμI"��������l�뺐t89�;�:��;�+;�|:;�7B;'�E;IbG;�H;)[H;��H;Z�H;֯H;3�H;��H;��H;C�H;�H;��H;�H;C�H;��H;��H;5�H;֯H;X�H;��H;)[H;�H;GbG;#�E;�7B;�|:;�+;��;�;�:�t89h��������I"��jrμ0O���d��u��F����nH�@���C������E�߾l����v�      C�;9ɾ~㼾B�������Mw��nH�����Z�䳽̕��s\8�p#������
^N�B���b��Hx��5:U��:R�;�0;]]=;j�C;�[F; �G;*H;fH;��H;T�H;{�H;��H;T�H;�H;i�H;�H;��H;�H;i�H;�H;R�H;��H;y�H;T�H;��H;fH;*H;�G;�[F;f�C;[]=;�0;S�;Q��:�5:�Hx��b�A��
^N�����p#��s\8�̕��䳽�Z񽲯��nH��Mw�����B��~㼾9ɾ      Ⱆ��������*|�NS\�� :����Z�n$�������K�v���Oļ����������&�����/�:�^;��#;�G6;x�?;&�D;��F;��G;4@H;�pH;�H;��H;L�H;��H;e�H;��H;��H;�H;��H;�H;��H;��H;d�H;��H;L�H;��H;�H;�pH;1@H;��G;��F;"�D;v�?;�G6;��#;�^;�/�:���&������������Oļv���K�����n$���Z���� :�OS\��*|�������      �+X��T��nH��6��� �k��F�䳽�����mR����ټ�����E<��?ݻd\�~����!:e�:��;P�,;��:;�7B;ǲE;�LG;rH;�SH;�{H;��H;�H;N�H;x�H;��H;H�H;�H;+�H;��H;+�H;�H;F�H;��H;{�H;L�H;�H;��H;�{H;�SH;pH;�LG;ĲE;�7B;��:;P�,;��;e�:�!:����d\��?ݻ�E<�����ټ����mR�����䳽F�k���� ��6��nH��T�      ��"]�Ո�r}���z�ý�u��̕���K�����o�iv���&R���H^��<�� �=�F��:�B;t";��4;��>;}D;ÁF;1�G;*H;�dH;��H;L�H;��H;d�H;f�H;��H;�H;Z�H;G�H;�H;E�H;Z�H;�H;��H;i�H;c�H;��H;I�H;��H;�dH;*H;.�G;��F;xD;��>;��4;r";�B;L��: �=�<��H^�����&R�iv���o�����K�̕���u��z�ý��r}�Ո�"]�      �ѽ\ν{�ý䳽<����L����d�s\8�w��ټiv����Y��_������� [�H�Y:���:xm;�r-;9�:;��A;koE;�"G;��G;�GH;�sH; �H;ǦH;�H;c�H;Q�H;��H;��H;��H;`�H;$�H;`�H;��H;��H;��H;S�H;a�H;�H;ĦH; �H;�sH;�GH;��G;�"G;goE;��A;9�:;�r-;xm;���:@�Y:$[��������_���Y�iv��ټv��s\8���d��L��<���䳽{�ý\ν      ���������Ȅ�lSt��Y�^n;�1O�q#���Oļ�����&R��_������N3�L�Y��4:^�:��;@&;H6;�X?;�D;exF;�G;m!H;�^H;��H;(�H;	�H;w�H;=�H;4�H;�H;I�H;�H;��H;F�H;��H;�H;G�H;�H;6�H;=�H;w�H;�H;(�H;��H;�^H;i!H;�G;axF;�D;�X?;
H6;@&;��;Z�:�4:P�Y��N3������_��&R������Oļq#��1O�^n;��Y�lSt��Ȅ�����      an;�z\8��s/�=�!�{��_���jrμ��������E<��������N3��Gx���9@�:_;{ ;\2;��<;#�B;߲E;h5G;<�G;kFH;�qH;؎H;��H;�H;��H;��H;��H;3�H;��H;Q�H;��H;@�H;��H;Q�H;��H;3�H;��H;��H;��H;�H;~�H;֎H;�qH;iFH;9�G;d5G;߲E;#�B;��<;\2;} ;_;D�:��9�Gx��N3��������E<��������jrμ_���|��=�!��s/�z\8�      ]������o�qrμу��sv��I"��^N�����?ݻH^�� ��T�Y���9<�:(��:�;z�.;�|:;%?A;��D;_�F;�G;*H;SaH;N�H;��H;�H;q�H;R�H;p�H;��H;.�H;O�H;��H;��H;�H;��H;��H;O�H;.�H;��H;n�H;O�H;m�H;�H;��H;N�H;PaH;*H;�G;_�F;��D;&?A;�|:;{�.;�;(��:<�:��9T�Y� ��H^���?ݻ���^N�I"��sv��у��qrμ�o����      �����x���#��?F{���]��E<����C�뻚���d\�:��$[��4:>�:.��:�[;��,;�8;O!@;1D;�[F;T{G;+H;zPH;MvH;�H;v�H;2�H;c�H;��H;��H;�H;�H;��H;��H;��H;��H;��H;��H;��H;�H;�H;��H;��H;^�H;2�H;s�H;�H;KvH;tPH;&H;T{G;�[F;1D;O!@;�8;��,;�[;0��:@�:�4:$[�:��d\�����D�뻟���E<���]�?F{��#���x��      �B(��%�����_�z����˻����b�&����� �=�H�Y:Z�:_;�;��,;;`8;��?;��C;�F; GG;�G;'@H;]kH;7�H;<�H;(�H;��H;��H;��H;��H;N�H;��H;�H;��H;��H;��H;��H;��H;�H;��H;P�H;��H;��H;��H;��H;#�H;<�H;5�H;YkH; @H;�G;GG;�F;��C;��?;=`8;��,;�;_;Z�:H�Y: �=�|���&��b�����˻x����_�����%�      Қ��F���J���X���b���-�r�뺘Hx�����!:H��:���:��;z ;z�.;�8;��?;(�C;�E;l#G;�G;2H;"bH;~�H;��H;��H;�H;�H;��H;M�H;k�H;m�H;!�H;L�H;��H;n�H;��H;n�H;��H;J�H; �H;m�H;k�H;K�H;��H;�H;޷H;��H;��H;z�H;bH;2H;�G;m#G;�E;)�C;��?;�8;z�.;} ;��;���:L��:�!:����Hx�p����-�
�b��X��J��J���      
��<���к����4�Y����t89�5:�/�:e�:�B;xm;@&;\2;�|:;L!@;��C;�E;�G;�G;�(H;0[H;�zH;r�H;�H;׳H;��H;��H;��H;��H;��H;.�H;��H;b�H;�H;2�H;��H;2�H;��H;b�H;��H;/�H;��H;��H;��H;��H;��H;׳H;�H;n�H;�zH;0[H;�(H;�G;�G;�E;�C;L!@;�|:;\2;@&;zm;�B;e�:�/�:�5:�t89����Y������к<��       �e9��98�9( :�Y:�y�:�;�:I��:�^;��;p";�r-;H6;��<;"?A; 1D;�F;i#G;�G;%H;�WH;�vH;��H;w�H;}�H;��H;D�H;��H;��H;o�H;
�H;��H;��H;]�H;B�H;��H;-�H;��H;A�H;_�H;��H;��H;
�H;l�H;��H;��H;A�H;��H;|�H;s�H;��H;�vH;�WH;%H;�G;j#G;�F; 1D;$?A;��<;H6;�r-;p";��;�^;I��:�;�:�y�:D�Y:( :@�9h�9      P�:�-�:�g�:H��:��:�^;��;O�;��#;R�,;��4;5�:;�X?; �B;��D;�[F; GG;�G;�(H;�WH;�uH;ÌH;K�H;2�H;Y�H;0�H;��H;$�H;�H;��H;��H;�H;��H;%�H;�H;��H;��H;��H;�H;%�H;��H;�H;��H;��H;�H;$�H;��H;0�H;Y�H;.�H;I�H;ÌH;�uH;�WH;�(H; �G;GG;�[F;��D; �B;�X?;5�:;��4;P�,;��#;N�;��;�^;��:N��:�g�:�-�:      ;��;m;[;�`;�%;�+;�0;�G6;��:;��>;��A;�D;ݲE;_�F;S{G;}�G;2H;1[H;�vH;H;��H;��H;�H;��H;��H;��H;��H;��H;�H;t�H;o�H;��H;��H;��H;��H;�H;��H;��H;��H;��H;o�H;u�H;�H;��H;��H;��H;��H;��H;��H;��H;��H;��H;�vH;1[H;2H;}�G;Q{G;`�F;�E;�D;��A;��>;��:;�G6;�0;�+;�%;�`;[;m;��;      �Y.;��.;l0;�2;v�4;7;�|:;[]=;y�?;�7B;}D;koE;bxF;h5G;�G;'H;$@H; bH;�zH;��H;I�H;��H;��H;�H;��H;��H;�H;-�H;V�H;��H;��H;��H;��H;}�H;$�H;W�H;~�H;U�H;$�H;}�H;��H;��H;��H;��H;T�H;.�H;��H;��H;��H;�H;��H;��H;G�H;��H;�zH;#bH;$@H;&H;�G;h5G;bxF;moE;{D;�7B;y�?;[]=;�|:;ā7;��4;�2;m0;��.;      z�<;<�<;=]=;�O>;
�?;��@;�7B;f�C;#�D;ŲE;��F;�"G;�G;:�G;*H;wPH;ZkH;��H;q�H;t�H;,�H;�H;�H;m�H;j�H;p�H;��H;��H;Y�H;s�H;2�H;G�H;B�H;�H;x�H;��H;��H;��H;{�H;�H;A�H;H�H;2�H;p�H;V�H;��H;��H;r�H;m�H;l�H;�H;�H;+�H;v�H;q�H;��H;ZkH;wPH;*H;:�G;�G;�"G;��F;ŲE;%�D;f�C;�7B;��@;�?;�O>;@]=;0�<;      �WC;oC;��C;�D;v�D;Q5E;&�E;�[F;��F;�LG;0�G;��G;k!H;mFH;SaH;NvH;;�H;��H;�H;��H;\�H;��H;��H;q�H;.�H;A�H;{�H;��H;"�H;��H;�H;��H;��H;m�H;��H;�H;	�H;�H;��H;m�H;��H;��H;�H;��H;�H;��H;x�H;A�H;1�H;q�H;��H;��H;[�H;��H;�H;��H;8�H;NvH;TaH;kFH;i!H;��G;0�G;�LG;��F;�[F;&�E;S5E;x�D;�D;�C;oC;      D[F;�dF;$�F;z�F;�F;�"G;GbG;�G;��G;rH;
*H;�GH;�^H;�qH;J�H;�H;:�H;��H;ӳH;��H;-�H;��H;��H;o�H;:�H;c�H;��H;��H;��H;��H;��H;��H;\�H;��H;�H;K�H;K�H;K�H;�H;��H;[�H;��H;��H;��H;��H;��H;��H;d�H;<�H;o�H;��H;��H;)�H;��H;ԳH;��H;9�H;�H;J�H;�qH;�^H;�GH;
*H;rH;��G;�G;GbG;�"G;$�F;{�F;(�F;�dF;      �G;�G;��G;��G;4�G;4�G;�H;*H;2@H;�SH;�dH;�sH;��H;֎H;��H;v�H;(�H;ݷH;��H;G�H;��H;��H;��H;��H;t�H;��H;��H;z�H;��H;��H;��H;2�H;��H;�H;<�H;n�H;��H;n�H;:�H;�H;��H;4�H;��H;��H;��H;z�H;��H;��H;v�H;��H;��H;��H;��H;G�H;��H;�H;(�H;t�H;��H;֎H;��H;�sH;�dH;�SH;5@H;*H;�H;2�G;:�G;��G;��G;
�G;      30H;�1H;^6H;P=H;@FH;vPH;-[H;$fH;qH;�{H;��H;&�H;(�H;��H;�H;4�H;��H;�H;��H;��H;"�H;��H;.�H;��H;��H;��H;x�H;��H;��H;��H;8�H;��H;��H;H�H;{�H;��H;�H;��H;{�H;G�H;��H;��H;9�H;��H;��H;��H;x�H;��H;��H;��H;.�H;��H;!�H;��H;��H;�H;��H;4�H;�H;��H;&�H;&�H;��H;�{H;qH;$fH;-[H;vPH;KFH;N=H;`6H;�1H;      �jH;1kH;hmH;�pH;�uH;@{H;��H;��H; �H;H;K�H;ʦH;�H;�H;o�H;b�H;��H;��H;��H;��H;�H;��H;S�H;\�H;�H;��H;��H;��H;��H;&�H;��H;��H;.�H;k�H;��H;��H;��H;��H;��H;k�H;+�H;��H;��H;&�H;��H;��H;��H;��H;�H;\�H;S�H;��H;�H;��H;��H;��H;��H;b�H;o�H;�H;�H;ȦH;I�H;��H;#�H;��H;��H;C{H;�uH;�pH;imH;(kH;      o�H;یH;_�H;��H;�H;��H;b�H;[�H;��H;#�H;��H;,�H;}�H;��H;T�H;��H;��H;H�H;��H;r�H;��H;�H;��H;s�H;��H;��H;��H;��H;$�H;��H;��H;5�H;j�H;��H;��H;��H;��H;��H;��H;��H;g�H;6�H;��H;��H;$�H;��H;��H;��H;��H;s�H;��H;�H;��H;r�H;��H;J�H;��H;��H;T�H;��H;}�H;,�H;��H;#�H;��H;^�H;b�H;�H;��H;��H;\�H;،H;      ��H;�H;�H;��H;٩H;��H;�H;��H;U�H;S�H;k�H;n�H;D�H;��H;r�H;��H;��H;k�H;��H;�H;��H;u�H;��H;6�H;�H;��H;��H;9�H;��H;��H;/�H;b�H;��H;��H;��H;��H;��H;��H;��H;��H;��H;c�H;/�H;��H;��H;;�H;��H;��H;�H;6�H;��H;v�H;��H;�H;��H;k�H;��H;��H;t�H;��H;D�H;m�H;j�H;S�H;U�H;��H;�H;��H;שH;��H;�H;�H;      ԵH;"�H;ζH;�H;˹H;��H;6�H;��H;��H;{�H;o�H;Z�H;9�H;��H;��H;�H;W�H;n�H;4�H;��H;�H;s�H;��H;K�H;��H;��H;1�H;��H;��H;6�H;]�H;{�H;��H;��H;��H;��H;��H;��H;��H;��H;��H;|�H;_�H;7�H;��H;��H;1�H;��H;��H;K�H;��H;s�H;�H;��H;4�H;o�H;W�H;�H;��H;��H;9�H;[�H;o�H;{�H;��H;��H;6�H;��H;ʹH;�H;϶H;�H;      d�H;��H;>�H;�H;W�H;��H;��H;\�H;l�H;��H;��H;��H;�H;:�H;4�H;�H;��H;�H;��H;��H;��H;��H;��H;I�H;��H;^�H;��H;��H;0�H;p�H;��H;��H;��H;��H;��H;��H;��H;��H;��H;��H;��H;��H;��H;q�H;2�H;��H;��H;\�H;��H;H�H;��H;��H;��H;��H;��H; �H;��H;�H;2�H;;�H;�H;��H;��H;��H;l�H;[�H;��H;��H;P�H;�H;>�H;��H;      ��H;�H;x�H;�H;�H;,�H;��H;�H;��H;J�H;�H;��H;J�H;��H;V�H;��H;�H;L�H;f�H;f�H;,�H;��H;z�H;�H;f�H;��H;�H;G�H;j�H;��H;��H;��H;��H;��H;��H;��H;��H;��H;��H;��H;��H;��H;��H;��H;m�H;G�H;�H;��H;h�H;�H;z�H;��H;*�H;f�H;f�H;M�H;�H;��H;T�H;��H;L�H;��H;�H;J�H;��H;�H;��H;0�H;�H;�H;x�H;�H;      ��H;��H;�H;��H;x�H;D�H;L�H;t�H;��H;�H;_�H;��H;�H;X�H;��H;��H;��H;��H;��H;K�H;�H;��H;#�H;~�H;��H;	�H;:�H;|�H;��H;��H;��H;��H;��H;��H;��H;��H;��H;��H;��H;��H;��H;��H;��H;��H;��H;|�H;7�H;	�H;��H;}�H;#�H;��H;�H;K�H;��H;��H;��H;��H;��H;X�H;�H;��H;^�H;�H;��H;t�H;L�H;H�H;m�H;��H;�H;��H;      ��H;�H;F�H;��H;a�H;�H;�H;�H;�H;+�H;N�H;k�H;��H;��H;��H;��H;��H;j�H;4�H;��H;��H;��H;W�H;��H;�H;J�H;n�H;��H;��H;��H;��H;��H;��H;��H;��H;��H;��H;��H;��H;��H;��H;��H;��H;��H;��H;��H;m�H;H�H;�H;��H;W�H;��H;��H;��H;4�H;k�H;��H;��H;��H;��H;��H;k�H;L�H;.�H;�H;�H;�H;�H;U�H;��H;F�H;�H;      ��H;��H;+�H;��H;D�H;��H;��H;��H;��H;��H;�H;.�H;K�H;I�H;�H;�H;��H;��H;��H;4�H;��H;�H;~�H;��H;�H;J�H;��H;��H;��H;��H;��H;��H;��H;��H;��H;��H;��H;��H;��H;��H;��H;��H;��H;��H;��H;��H;��H;K�H;�H;��H;~�H;�H;��H;4�H;��H;��H;��H;�H;�H;I�H;K�H;.�H;�H;��H;��H;��H;��H;��H;7�H;��H;*�H;��H;      ��H;�H;F�H;��H;b�H;�H;�H;�H;�H;+�H;N�H;k�H;��H;��H;��H;��H;��H;j�H;4�H;��H;��H;��H;W�H;��H;�H;J�H;n�H;��H;��H;��H;��H;��H;��H;��H;��H;��H;��H;��H;��H;��H;��H;��H;��H;��H;��H;��H;m�H;J�H;�H;��H;W�H;��H;��H;��H;4�H;k�H;��H;��H;��H;��H;��H;k�H;N�H;,�H;�H;�H;�H;�H;U�H;��H;C�H;�H;      ��H;��H;�H;��H;x�H;D�H;L�H;w�H;��H;�H;^�H;��H;�H;X�H;��H;��H;��H;��H;��H;K�H;
�H;��H;#�H;~�H;��H;	�H;9�H;|�H;��H;��H;��H;��H;��H;��H;��H;��H;��H;��H;��H;��H;��H;��H;��H;��H;��H;|�H;7�H;	�H;��H;{�H;#�H;��H;�H;K�H;��H;��H;��H;��H;��H;X�H;�H;��H;^�H;�H;��H;s�H;L�H;H�H;n�H;��H;�H;��H;       �H;�H;x�H;�H;�H;,�H;��H;�H;��H;J�H;�H;��H;L�H;��H;T�H;��H;�H;L�H;f�H;f�H;/�H;��H;z�H;�H;h�H;��H;�H;G�H;j�H;��H;��H;��H;��H;��H;��H;��H;��H;��H;��H;��H;��H;��H;��H;��H;m�H;G�H;�H;��H;f�H;�H;z�H;��H;*�H;f�H;f�H;M�H;�H;��H;T�H;��H;J�H;��H;�H;J�H;��H;�H;��H;0�H;�H;�H;v�H;�H;      f�H;��H;>�H; �H;U�H;��H;��H;[�H;l�H;��H;��H;��H;�H;;�H;2�H;�H;��H;�H;��H;��H;�H;��H;��H;H�H;��H;^�H;��H;��H;0�H;p�H;��H;��H;��H;��H;��H;��H;��H;��H;��H;��H;��H;��H;��H;q�H;2�H;��H;��H;\�H;��H;F�H;��H;��H;��H;��H;��H;�H;��H;�H;4�H;:�H;	�H;��H;��H;��H;l�H;X�H;��H;��H;N�H; �H;;�H;��H;      ԵH;"�H;ѶH;�H;͹H;��H;:�H;��H;��H;z�H;m�H;Z�H;9�H;��H;��H;�H;W�H;n�H;4�H;��H;�H;s�H;��H;K�H;��H;��H;1�H;��H;��H;6�H;_�H;{�H;��H;��H;��H;��H;��H;��H;��H;��H;��H;|�H;]�H;7�H;��H;��H;1�H;��H;��H;K�H;��H;s�H;�H;��H;4�H;o�H;W�H;�H;��H;��H;9�H;[�H;m�H;{�H;��H;��H;:�H;��H;ʹH;�H;϶H;�H;      ��H;�H;�H;��H;٩H;��H;�H;��H;U�H;R�H;k�H;m�H;D�H;��H;t�H;��H;��H;j�H;��H;�H;��H;v�H;��H;7�H;�H;��H;��H;;�H;��H;��H;/�H;b�H;��H;��H;��H;��H;��H;��H;��H;��H;��H;c�H;/�H;��H;��H;9�H;��H;��H;�H;6�H;��H;u�H;��H;�H;��H;k�H;��H;��H;r�H;��H;D�H;n�H;j�H;U�H;U�H;��H;�H;��H;שH;��H;�H;�H;      h�H;یH;_�H;��H;��H;�H;e�H;^�H;��H;"�H;��H;,�H;}�H;��H;T�H;��H;��H;H�H;��H;s�H;��H;�H;��H;s�H;��H;��H;��H;��H;$�H;��H;��H;5�H;i�H;��H;��H;��H;��H;��H;��H;��H;i�H;6�H;��H;��H;$�H;��H;��H;��H;��H;s�H;��H;�H;��H;r�H;��H;J�H;��H;��H;T�H;��H;}�H;,�H;��H;"�H;��H;^�H;d�H;�H;��H;��H;]�H;ڌH;      �jH;-kH;omH;�pH;�uH;={H;��H;��H; �H;��H;K�H;ʦH;	�H;�H;o�H;b�H;��H;��H;��H;��H;�H;��H;T�H;\�H;�H;��H;��H;��H;��H;'�H;��H;��H;,�H;k�H;��H;��H;��H;��H;��H;k�H;,�H;��H;��H;$�H;��H;��H;��H;��H;�H;\�H;Q�H;��H;�H;��H;��H;��H;��H;c�H;n�H;�H;�H;ʦH;K�H;��H;"�H;��H;��H;?{H;�uH;�pH;pmH;-kH;      30H;�1H;^6H;N=H;AFH;vPH;-[H;&fH;qH;�{H;��H;&�H;&�H;��H;�H;4�H;��H;�H;��H;��H;'�H;��H;/�H;��H;��H;��H;x�H;��H;��H;��H;9�H;��H;��H;F�H;z�H;��H;�H;��H;{�H;H�H;��H;��H;8�H;��H;��H;��H;x�H;��H;��H;��H;-�H;��H; �H;��H;��H;�H;��H;5�H;�H;��H;(�H;&�H;��H;�{H;qH;&fH;-[H;sPH;LFH;P=H;`6H;�1H;      �G;
�G;��G;��G;3�G;0�G;�H;*H;2@H;�SH;�dH;�sH;��H;֎H;��H;v�H;)�H;ݷH;��H;G�H;��H;��H; �H;��H;v�H;��H;��H;z�H;��H;��H;��H;4�H;��H;�H;:�H;n�H;��H;m�H;<�H;�H;��H;4�H;��H;��H;��H;z�H;��H;��H;t�H;��H;��H;��H;��H;G�H;��H;޷H;&�H;t�H;��H;֎H;��H;�sH;�dH;�SH;4@H;*H;�H;0�G;4�G;��G;��G;�G;      J[F;�dF;1�F;~�F; �F;�"G;GbG;�G;��G;sH;
*H;�GH;�^H;�qH;H�H;�H;:�H;��H;ԳH;��H;.�H;��H;��H;p�H;<�H;c�H;��H;��H;��H;��H;��H;��H;\�H;��H;�H;K�H;K�H;K�H;�H;��H;Z�H;��H;��H;��H;��H;��H;��H;d�H;:�H;n�H;��H;��H;)�H;��H;ӳH;��H;9�H;�H;J�H;�qH;�^H;�GH;
*H;pH;��G;�G;IbG;�"G;$�F;{�F;1�F;�dF;      �WC;oC; �C;�D;x�D;Q5E;&�E;�[F;��F;�LG;1�G;��G;i!H;kFH;TaH;OvH;:�H;��H;�H;��H;]�H;��H;��H;r�H;1�H;?�H;{�H;��H;"�H;��H;�H;��H;��H;m�H;��H;�H;	�H;�H;��H;l�H;��H;��H;�H;��H;�H;��H;x�H;A�H;.�H;q�H;��H;��H;[�H;��H;�H;��H;8�H;NvH;SaH;kFH;k!H;��G;0�G;�LG;��F;�[F;&�E;Q5E;v�D;�D; �C;oC;      }�<;:�<;E]=;�O>;�?;��@;�7B;i�C;%�D;ȲE;��F;�"G;�G;:�G;*H;wPH;[kH;~�H;q�H;v�H;/�H;�H;�H;m�H;m�H;p�H;��H;��H;Y�H;s�H;2�H;G�H;B�H;�H;x�H;��H;��H;��H;z�H;�H;A�H;H�H;2�H;p�H;V�H;��H;��H;p�H;j�H;m�H;�H;�H;)�H;t�H;q�H;��H;YkH;wPH;*H;:�G;�G;�"G;��F;ŲE;&�D;i�C;�7B;��@;�?;�O>;E]=;/�<;      �Y.; �.;~0;�2;v�4;ȁ7;�|:;[]=;y�?;�7B;{D;moE;axF;h5G;�G;'H;$@H; bH;�zH;��H;L�H;��H;��H;�H;��H;��H;�H;.�H;V�H;��H;��H;��H;��H;}�H;$�H;W�H;~�H;U�H;$�H;}�H;��H;��H;��H;��H;S�H;-�H;��H;��H;��H;�H;��H;��H;E�H;��H;�zH;"bH;&@H;'H;�G;h5G;axF;moE;{D;�7B;y�?;[]=;�|:;ȁ7;|�4;�2;s0;��.;      ;��;m;[;�`;�%;�+;�0;�G6;��:;��>;��A;�D;�E;_�F;S{G;}�G;2H;1[H;�vH;ÌH;��H;��H;�H;��H;��H;��H;��H;��H; �H;u�H;o�H;��H;��H;��H;��H;�H;��H;��H;��H;��H;o�H;t�H;�H;��H;��H;��H;��H;��H; �H;��H;��H;��H;�vH;1[H;2H;|�G;S{G;`�F;ݲE;�D;��A;��>;��:;�G6;�0;�+;�%;�`;[;m;��;      D�:�-�:�g�:N��:��:�^;��;P�;��#;R�,;��4;5�:;�X?; �B;��D;�[F; GG;�G;�(H;�WH;�uH;ÌH;K�H;2�H;Y�H;.�H;��H;$�H;�H;��H;��H;�H;��H;#�H;�H;��H;��H;��H;�H;%�H;��H;�H;��H;��H;�H;$�H;��H;0�H;Y�H;.�H;I�H;ÌH;�uH;�WH;�(H;�G;GG;�[F;��D; �B;�X?;5�:;��4;N�,;��#;P�;��;�^;��:J��:�g�:�-�:      �e9��9`�9$ :4�Y:�y�:�;�:M��:�^;��;p";�r-;	H6;��<;$?A; 1D;�F;i#G;�G;%H;�WH;�vH;��H;w�H;|�H;��H;D�H;��H;��H;o�H;
�H;��H;��H;_�H;A�H;��H;-�H;��H;B�H;]�H;��H;��H;
�H;l�H;��H;��H;A�H;��H;}�H;s�H;��H;�vH;�WH;%H;�G;j#G;�F;1D;"?A;��<;H6;�r-;o";��;�^;O��:�;�:�y�:P�Y:$ :H�9X�9      
��<���к����0�Y����t89�5:�/�:e�:�B;xm;@&;\2;�|:;L!@;�C;�E;�G;�G;�(H;0[H;�zH;r�H;�H;ֳH;��H;��H;��H;��H;��H;.�H;��H;b�H;��H;2�H;��H;2�H;�H;b�H;��H;/�H;��H;��H;��H;��H;��H;ٳH;�H;n�H;�zH;0[H;�(H;�G;�G;�E;�C;L!@;�|:;\2;@&;xm;�B;e�:�/�:�5:�t89����Y������к<��      Қ��F���J���X���b���-�n�뺘Hx�����!:H��:���:��;z ;z�.;�8;��?;(�C;�E;l#G;�G;2H;"bH;}�H;��H;��H;�H;�H;��H;M�H;k�H;k�H;!�H;J�H;��H;n�H;��H;n�H;��H;L�H; �H;n�H;k�H;K�H;��H;�H;޷H;��H;��H;|�H;bH;2H;�G;m#G;�E;)�C;��?;�8;z�.;z ;��;���:H��:�!:����Hx�n����-�
�b��X��J��J���      �B(��%�����_�x����˻����b�&�|��� �=�H�Y:Z�:_;�;��,;=`8;��?;��C;�F; GG;�G;'@H;]kH;5�H;:�H;(�H;��H;��H;��H;��H;P�H;��H;�H;��H;��H;��H;��H;��H;�H;��H;P�H;��H;��H;��H;��H;#�H;<�H;7�H;YkH;"@H;�G;GG;�F;��C;��?;;`8;��,;�;_;Z�:H�Y: �=�����&��b�����˻x����_�����%�      �����x���#��?F{���]��E<����C�뻚���d\�:�� [��4:>�:0��:�[;��,;�8;O!@;1D;�[F;T{G;(H;xPH;KvH;�H;v�H;2�H;b�H;��H;��H;�H;�H;��H;��H;��H;��H;��H;��H;��H;�H;�H;��H;��H;^�H;2�H;s�H;�H;MvH;vPH;&H;T{G;�[F;1D;O!@;�8;��,;�[;.��:>�:�4:$[�:��d\�����C�뻟���E<���]�?F{��#���x��      ]������o�qrμу��tv��I"��^N�����?ݻH^�� ��T�Y���9<�:(��:�;x�.;�|:;%?A;��D;_�F;�G;*H;PaH;M�H;��H;�H;q�H;Q�H;n�H;��H;/�H;O�H;��H;��H;�H;��H;��H;P�H;.�H;��H;p�H;Q�H;n�H;�H;��H;N�H;SaH;*H;�G;_�F;��D;&?A;�|:;{�.;�;(��:<�:��9T�Y� ��H^���?ݻ���^N�I"��sv��у��qrμ�o����      an;�z\8��s/�=�!�{��_���jrμ��������E<��������N3��Gx���9D�:_;{ ;\2;��<; �B;߲E;h5G;<�G;iFH;�qH;؎H;~�H;�H;��H;��H;��H;4�H;��H;Q�H;��H;@�H;��H;Q�H;��H;2�H;��H;��H;��H;�H;��H;֎H;�qH;kFH;9�G;d5G;߲E;#�B;��<;\2;~ ;_;@�:��9�Gx��N3��������E<��������jrμ_���{��=�!��s/�z\8�      ���������Ȅ�lSt��Y�^n;�1O�q#���Oļ�����&R��_������N3�L�Y��4:^�:��;@&;H6;�X?;�D;exF;�G;i!H;�^H;��H;(�H;�H;w�H;=�H;4�H;�H;G�H;�H;��H;F�H;��H;�H;I�H;�H;4�H;=�H;w�H;�H;(�H;��H;�^H;m!H;�G;axF;�D;�X?;H6;@&;��;Z�:�4:L�Y��N3������_��&R������Oļq#��1O�^n;��Y�lSt��Ȅ�����      �ѽ\ν{�ý䳽<����L����d�s\8�w��ټiv����Y��_�������$[�H�Y:���:xm;�r-;6�:;��A;joE;�"G;��G;�GH;�sH; �H;ŦH;�H;a�H;P�H;��H;��H;��H;a�H;$�H;a�H;��H;��H;��H;S�H;c�H;�H;ŦH; �H;�sH;�GH;��G;�"G;goE;��A;9�:;�r-;xm;���:@�Y:([��������_���Y�iv��ټv��s\8���d��L��<���䳽{�ý\ν      ��"]�Ո�r}���z�ý�u��̕���K�����o�iv���&R���H^��<�� �=�H��:�B;t";��4;��>;{D;��F;.�G;*H;�dH;��H;L�H;��H;c�H;f�H;��H;�H;Z�H;E�H;�H;G�H;Z�H;�H;��H;i�H;d�H;��H;I�H;��H;�dH;*H;1�G;��F;zD;��>;��4;s";�B;L��: �=�>��H^�����&R�iv���o�����K�̕���u��z�ý��r}�Ո�"]�      �+X��T��nH��6��� �k��F�䳽�����mR����ټ�����E<��?ݻd\�|���|!:e�:��;N�,;��:;�7B;ǲE;�LG;rH;�SH;�{H;��H;�H;L�H;z�H;��H;F�H;�H;+�H;��H;+�H;�H;H�H;��H;x�H;N�H;�H;��H;�{H;�SH;rH;�LG;ĲE;�7B;��:;P�,;��;e�:�!:����d\��?ݻ�E<�����ټ����mR�����䳽F�k���� ��6��nH��T�      Ⱆ��������*|�NS\�� :����Z�n$�������K�v���Oļ����������&�����/�:�^;��#;�G6;x�?;&�D;��F;��G;2@H;�pH;�H;��H;L�H;��H;e�H;��H;��H;�H;��H;�H;��H;��H;d�H;��H;L�H;��H;�H;�pH;1@H;��G;��F;"�D;v�?;�G6;��#;�^;�/�:���&������������Oļv���K�����n$���Z���� :�OS\��*|�������      C�;9ɾ~㼾B�������Mw��nH�����Z�䳽̕��s\8�p#������
^N�B���b��Hx��5:U��:P�;�0;[]=;i�C;�[F;�G;*H;fH;��H;T�H;y�H;��H;T�H;	�H;j�H;�H;��H;
�H;i�H;	�H;R�H;��H;{�H;T�H;��H;fH;*H;�G;�[F;f�C;]]=;�0;S�;Q��:�5:�Hx��b�B��
^N�����p#��s\8�̕��䳽�Z񽲯��nH��Mw�����B��~㼾9ɾ      1y��v�l���E�߾����C��@����nH���FὟu����d�0O�jrμI"��������j�뺐t89�;�:�;�+;�|:;�7B;#�E;GbG;�H;)[H;��H;Z�H;֯H;2�H;��H;��H;C�H;�H;��H;�H;C�H;��H;~�H;3�H;֯H;X�H;��H;)[H;�H;GbG;'�E;�7B;�|:;�+;��;�;�:�t89h��������I"��jrμ0O���d��u��F����nH�@���C������E�߾l����v�      �O/�rM+�Y�����JW��9ɾC���Mw�� :�k��y�ý�L��^n;�_���sv���E<��˻��-����y�:�^;�%;��7;��@;O5E;�"G;1�G;tPH;C{H;�H;��H;��H;��H;0�H;K�H; �H;��H;!�H;K�H;2�H;��H;��H;��H;�H;@{H;tPH;1�G;�"G;Q5E;��@;7;�%;�^;�y�:����-��˻�E<�sv��`���^n;��L��y�ýk��� :��Mw�C��9ɾJW�����Y��rM+�      :�X�YvS�8E��O/��S�JW����������NS\��� ���<����Y�{��Ѓ����]�w����b��Y�(�Y:��:�`;|�4;�?;u�D;�F;0�G;@FH;�uH;�H;ʩH;ƹH;M�H;�H;\�H;S�H;3�H;S�H;\�H;�H;L�H;ɹH;ʩH;�H;�uH;@FH;3�G;�F;v�D;	�?;~�4;�`;��:(�Y:�Y�
�b�x�����]�Ѓ��{���Y�<����当� �NS\���������JW���S��O/�8E�YvS�      � ����y�c�h��N��O/����D�߾B���*|��6�r}�䳽lSt�>�!�qrμ@F{��_��X������4 :V��:[;�2;�O>;�D;}�F;��G;S=H;�pH;��H;��H;�H;�H;�H;��H;��H;��H;��H;��H;�H;�H;�H;��H;��H;�pH;S=H;��G;}�F;�D;�O>;�2;[;^��:4 :�����X���_�@F{�qrμ>�!�lSt�䳽r}��6��*|�B��D�߾����O/��N�c�h���y�      ?v��c���X ��c�h�8E�Y��l���~㼾���nH�Ո�{�ý�Ȅ��s/��o��#�����J���к0�9�g�:m;m0;9]=;�C;2�F;��G;W6H;lmH;U�H;ߥH;ǶH;6�H;|�H;�H;>�H;�H;?�H;�H;|�H;4�H;ǶH;ߥH;R�H;imH;W6H;��G;1�F;�C;5]=;p0;m;�g�:8�9�кJ������#���o��s/��Ȅ�{�ýՈ��nH���~㼾l���Y��8E�c�h�X ��c���      ~h��1���c�����y�YvS�rM+��v�9ɾ�����T�"]�\ν����z\8�����x���%�D���6��8�9�-�:��;��.;3�<;oC;�dF;�G;�1H;0kH;֌H;�H;�H;��H;�H;��H;�H;��H;�H;��H;�H;��H;�H;�H;ӌH;-kH;�1H;�G;�dF;oC;0�<;��.;��;�-�:0�96��D����%��x�����z\8�����\ν"]��T�����9ɾ�v�rM+�YvS���y�c���1���      HEb�c]��N���7����u� ���˾��,�j��!,�s���N��Gm�-��:,˼��x�X���1��ڥ��(�:��:�;[�1;J,>;��C;�wF;	�G;� H;?H;iH;g�H;��H;P�H;0�H;��H;A�H;��H;B�H;��H;0�H;O�H;��H;g�H;iH;	?H;� H;	�G;�wF;��C;G,>;_�1;�;��: �:ڥ���1��X����x�:,˼-��Gm�N��s����!,�,�j�����˾u� ������7��N�c]�      c]�g�W��TI�v3� E�������Ǿx����f�:)�(��v;���Fi��k���Ǽ�[t�J�	�$Ȅ��W����:(��:��;qJ2;gZ>;]	D;�F;W�G;+H;�?H;�iH;��H;��H;��H;M�H;��H;l�H;��H;l�H;��H;M�H;��H;��H;��H;�iH;�?H;-H;W�G;�F;]	D;cZ>;vJ2;��;(��:��:�W��$Ȅ�J�	��[t���Ǽ�k��Fi�v;��(��:)��f�x�����Ǿ���� E�v3��TI�g�W�      �N��TI���;�1�'�l��쾂���z󐾶Z��K ��s�C����&^���"����g����¨u�� ���3<:=��:;}g3;
�>;�BD;˖F;��G;�H;_BH;�kH;j�H;��H;@�H;�H;��H;��H;[�H;��H;��H;�H;?�H;��H;j�H;�kH;ZBH;�H;��G;ʖF;�BD;�>;�g3;;?��:�3<:� ����u������g��"����&^�C����s潧K ��Z�z󐾂�����l�1�'���;��TI�      ��7�v3�1�'����u� ��{Ծ"���I���|�F�����ӽ���a�L�Lv��뮼PT����PV�0�=�(*i:���:�z ;�$5;ï?;!�D;�F;
�G;�H;�FH;�nH;��H;��H;��H;��H;J�H;i�H;�H;i�H;J�H;��H;��H;��H;��H;�nH;�FH;�H;
�G;�F; �D;��?;�$5;�z ;���: *i:4�=��PV���PT��뮼Lv�a�L�����ӽ���|�F�I���"����{Ծu� ����1�'�v3�      ��� E�l�u� �X�ݾm���X͓��f��>/�����'���섽R�6��t�w��\�:�Tʻk.�Xڷ��t�:�;��$;�Y7;o�@;
E;3�F;M�G;�H;PLH;�rH;ƏH;ߤH;5�H;0�H;D�H;]�H;��H;\�H;C�H;0�H;4�H;�H;ƏH;�rH;MLH;�H;N�G;2�F;
E;k�@;�Y7;��$;�;�t�:Xڷ�k.�Tʻ\�:�w���t�R�6��섽�'������>/��f�X͓�m���Y�ݾu� �l� E�      u� ��������{Ծm���x���]�x��SC��^��޽B���{�e�*��E�Ѽ&G������R�������8)��:�Y;j�);�9;�A;҄E;�G;2�G;|!H;SSH;�wH;��H;��H;R�H;��H;��H;��H;��H;��H;��H;��H;R�H;��H;��H;�wH;OSH;|!H;1�G;�G;фE;�A;�9;j�);�Y;'��:��8����R�����&G��E�Ѽ)��{�e�B����޽�^��SC�]�x�x���m����{Ծ�쾤���      ��˾��Ǿ����"���X͓�]�x���J��K �p��� ������?����뮼*�[�����2|�nW����:��:�';�/;~g<;�C;�F;�NG;��G;A-H;�[H;�}H;ٗH;ڪH;͸H;��H;�H;��H;�H;��H;�H;��H;͸H;ܪH;ٗH;�}H;[H;A-H;��G;�NG;�F;�C;|g<;�/;�';��:��:hW���2|����*�[��뮼���?���� ��p����K ���J�]�x�X͓�"���������Ǿ      ��x���z�I����f��SC��K �qn���Ž����Z��k� }ռ-X��`y-�$���V.�����P�:�+�:��;84;O�>;D;�wF;G�G;��G;�9H;kdH;��H;��H;r�H;��H;��H;��H;d�H;��H;d�H;��H;��H;�H;t�H;��H;��H;hdH;�9H;��G;G�G;�wF;D;O�>;84;��;�+�:�P�:���W.�$���_y-�-X�� }ռ�k��Z�����Žqn���K ��SC��f�I���z�x���      ,�j��f��Z�|�F��>/��^�p����ŽH ���Fi��Q+�}t�pT��n�W�����1���Ⱥ Y�9�P�:�Y;��(;"�8;A;�E;�F;�G;�H;GH;�mH;��H;ԡH;Q�H;~�H;��H;��H;�H;�H;�H;��H;��H;~�H;R�H;ѡH;��H;�mH;GH;�H;�G;�F;�E;A;"�8;��(;�Y;�P�:Y�9�Ⱥ�1�����n�W�oT��}t�Q+��Fi�H ���Žp����^��>/�|�F��Z��f�      �!,�:)��K ��������޽ ������Fi��0����鷼��x�����.��<�(�x��t+i:Ý�:Z�;��0;e�<;�C;��E;&=G;�G;%H;vTH;�wH;��H;(�H;_�H;��H;P�H;��H;��H;��H;��H;��H;P�H;��H;`�H;(�H;��H;�wH;vTH;%H;�G;"=G;��E;�C;e�<;��0;X�;Ý�:x+i:x��=�(��.�������x�鷼����0��Fi���� ���޽�������K �:)�      s���(��s��ӽ�'��B�������Z��Q+�����"��G����0���׻��b�W���Y�9
��:H`;�*';Z7;$$@;@�D;�F;,�G;��G;K8H;bH;�H;j�H;��H;��H;��H;��H;��H;`�H;L�H;`�H;��H;��H;��H;��H;��H;j�H;�H;bH;I8H;��G;)�G;�F;=�D;$$@;Z7;�*';H`;��:�Y�9W����b���׻��0�G���"������Q+��Z����B����'���ӽ�s�(��      N��v;��C�������섽{�e��?��k�~t�鷼G���e7�����Ǆ�B0� �t�bu�:>,�:�;�1;n�<;{�B;@�E;G;
�G;tH;�JH;qoH;�H;��H;'�H;��H;��H;0�H;��H; �H;��H;�H;��H;/�H;��H;��H;'�H;��H;�H;ooH;�JH;sH;�G;G;=�E;{�B;n�<;�1;�;D,�:`u�: �t�D0��Ǆ���껂e7�G��鷼}t��k��?�{�e��섽���C���v;��      Hm��Fi��&^�a�L�R�6�*���� }ռpT����x���0�������� ���׷�ho`:��:7�;E�*;V�8;)�@;Q�D;�F;~G;��G;�1H;�[H;�|H;ҕH;�H;��H;��H;��H;��H;��H;��H;��H;��H;��H;��H;��H;��H;��H;�H;ЕH;�|H;�[H;�1H;��G;~G;{�F;Q�D;)�@;T�8;E�*;:�;��:lo`:�׷����������껿�0���x�oT��!}ռ��*��R�6�a�L��&^��Fi�      -���k��Kv��t�E�Ѽ�뮼-X��n�W������׻�Ǆ����@��t5<:���:�Y;�t%;%5;�Z>;aC;��E;L*G;}�G;*H;HH;�lH;�H;�H;֯H;�H;��H;��H;�H;��H;��H;@�H;��H;��H;�H;��H;��H;�H;ԯH;�H;�H;~lH;HH;(H;y�G;G*G;��E;aC;�Z>;%5;�t%;�Y;���:|5<:0������Ǆ���׻���m�W�-X���뮼D�Ѽ�t�Kv���k�      :,˼��Ǽ�"���뮼w��&G��*�[�ay-�����.����b�D0��׷�p5<:*M�:];��!;�J2;�g<;h0B;DCE;C�F;e�G;�G;�4H;�\H;|H;��H;��H;m�H;��H;R�H;��H;a�H;b�H;�H;��H;�H;d�H;b�H;��H;U�H;��H;i�H;��H;��H;|H;�\H;�4H;�G;]�G;C�F;CCE;j0B;�g<; K2;��!;];*M�:t5<:�׷�D0㺸�b��.�����ay-�*�[�%G��w���뮼�"����Ǽ      ��x��[t���g�PT�^�:�������&����1��<�(�
W����t�ho`:���:];){ ;��0;v;;=A;/�D;�wF;�cG;j�G;�!H;�MH;�oH;��H;��H;ٯH;��H;x�H;��H;m�H;��H;�H;��H;7�H;��H;�H;�H;k�H;��H;w�H;��H;үH;��H;��H;�oH;�MH;�!H;f�G;�cG;�wF;/�D;=A;y;;��0;({ ;];���:ho`:��t�W��;�(��1��'���������]�:�PT���g��[t�      X��H�	������ Tʻ�R���2|�X.��Ⱥx���Y�9bu�:��:�Y;��!;��0;�:;˵@;"CD;�2F;�8G;��G;�H;@H;:dH;؀H;��H;Z�H;\�H;_�H;��H;�H;��H;�H;��H;�H;��H;�H;��H;�H;��H;�H;��H;]�H;W�H;W�H;��H;ڀH;:dH;{@H;�H;��G;�8G;�2F;"CD;ε@;�:;��0;��!;�Y;��:du�:�Y�9p���ȺY.��2|��R��Tʻ�����J�	�      �1��%Ȅ���u��PV�r.����rW������X�9p+i:��:>,�:7�;�t%;�J2;t;;ɵ@;�D;%F;@G;��G;�H;�5H;�ZH;IxH;T�H;=�H;)�H;(�H;k�H;��H;-�H;B�H;;�H;P�H;k�H;��H;k�H;P�H;:�H;A�H;.�H;�H;j�H;$�H;)�H;:�H;T�H;HxH;�ZH;�5H;�H;��G;@G;%F;�D;ɵ@;t;;�J2;�t%;7�;>,�:��:x+i:Y�9���pW�����j.��PV���u�*Ȅ�      ʥ���W��� ��8�=��ڷ���8�:�P�:�P�:���:F`;�;C�*;%5;�g<;=A;CD;%F;�G;��G;|�G;�-H;/SH;mqH;��H;ҝH;��H;(�H;M�H;�H;�H;��H;f�H;��H;��H;��H;��H;��H;��H;��H;d�H;��H;�H;�H;I�H;(�H;��H;ԝH;��H;iqH;*SH;�-H;y�G;��G;�G;'F;CD;=A;�g<;%5;C�*;�;H`;���:�P�:�P�:�:@�8Xڷ�4�=�� ���W��      $�:ܡ:�3<:$*i:�t�:!��:��:�+�:�Y;\�;�*';�1;P�8;�Z>;g0B;)�D;�2F;=G;��G;1�G;�)H;�NH;�lH;_�H;z�H;��H;��H;B�H;��H;�H;J�H;;�H;C�H;k�H;��H;��H;��H;��H;��H;k�H;B�H;=�H;L�H;�H;��H;@�H;��H;��H;x�H;[�H;�lH;�NH;�)H;2�G;��G;=G;�2F;*�D;g0B;�Z>;P�8;�1;�*';Z�;�Y;�+�:��:'��:�t�:$*i:�3<:��:      ��:@��:I��:���:�;�Y;�';��;��(;��0;Z7;j�<;(�@;aC;CCE;�wF;�8G;��G;}�G;�)H;�LH;jH;H�H;p�H;��H;�H;ϾH;v�H;:�H;��H;&�H;g�H;��H;��H;��H;��H;��H;��H;��H;��H;��H;h�H;&�H;��H;6�H;v�H;ξH;�H;��H;k�H;H�H;jH;�LH;�)H;}�G;��G;�8G;�wF;BCE;aC;(�@;j�<;�Y7;��0;��(;��;�';�Y;�;���:C��:��:      �;��;*;�z ;��$;s�);�/;?4;$�8;e�<;*$@;}�B;Q�D;��E;D�F;�cG;��G;�H;�-H;�NH;jH;^�H;ɔH;äH;�H;ԼH;��H;��H;]�H;�H;��H;B�H;^�H;��H;��H;~�H;��H;~�H;��H;��H;\�H;B�H;��H;��H;Y�H;��H;��H;ּH;�H;��H;ŔH;\�H;jH;�NH;�-H;�H;��G;�cG;E�F;��E;R�D;~�B;)$@;g�<;&�8;<4;�/;s�);��$;�z ;*;��;      c�1;sJ2;}g3;�$5;�Y7;�9;�g<;O�>;A;�C;?�D;@�E;~�F;J*G;c�G;i�G;�H;�5H;/SH;�lH;H�H;ʔH;?�H;�H;��H;}�H;u�H;G�H;�H;��H;��H;��H;��H;��H;��H;>�H;��H;>�H;��H;��H;��H;��H;��H;��H;�H;G�H;r�H;��H;��H;�H;<�H;ɔH;F�H;�lH;/SH;�5H;�H;g�G;a�G;L*G;~�F;@�E;@�D;�C;A;N�>;�g<;
�9;�Y7;�$5;�g3;dJ2;      \,>;pZ>;�>;��?;n�@;�A;�C;D;�E;��E;�F;G;~G;z�G;	�G;�!H;{@H;�ZH;jqH;^�H;k�H;¤H;�H;0�H;��H;��H;`�H;*�H;�H;�H;~�H;L�H;��H;��H;v�H;��H;
�H;��H;x�H;��H;��H;O�H;|�H;�H;�H;*�H;]�H;��H;��H;/�H;�H;¤H;i�H;_�H;lqH;�ZH;{@H;�!H;	�G;z�G;~G;G;�F;��E;�E;D;�C;�A;u�@;��?;�>;dZ>;      ��C;d	D;|BD;$�D;
E;ԄE;�F;�wF;�F;$=G;(�G;
�G;��G;+H;�4H;�MH;?dH;JxH;��H;��H;��H;�H;��H;��H;_�H;�H;��H;��H;��H;��H;��H;��H;��H;o�H;�H;r�H;|�H;r�H;�H;n�H;��H;��H;��H;��H;��H;��H;��H;�H;_�H;��H;��H;�H;��H;��H;�H;MxH;<dH;�MH;�4H;-H;��G;
�G;(�G;"=G;�F;�wF;�F;ՄE;
E;$�D;|BD;e	D;      �wF;�F;��F;�F;2�F;�G;�NG;C�G;}�G;�G;��G;vH;�1H;HH;�\H;�oH;׀H;Q�H;НH;��H;�H;ѼH;z�H;��H;
�H;��H;Q�H;L�H;��H;��H;G�H;��H;e�H;)�H;��H;��H;��H;��H;��H;)�H;c�H;��H;I�H;��H;��H;L�H;O�H;��H;�H;��H;|�H;ӼH;޳H;��H;НH;S�H;׀H;�oH;�\H;HH;�1H;vH;��G;�G;�G;C�G;�NG;�G;9�F;�F;��F;�F;      �G;Z�G;��G;�G;P�G;6�G;��G;��G;�H;%H;L8H;�JH;�[H;�lH;|H;��H;��H;:�H;��H;��H;ѾH;��H;t�H;b�H;��H;T�H;6�H;��H;{�H;(�H;g�H;B�H;�H;��H;�H;8�H;F�H;8�H;�H;��H;�H;A�H;i�H;(�H;{�H;��H;3�H;S�H;��H;a�H;t�H;��H;ξH;��H;��H;=�H;��H;��H;|H;�lH;�[H;�JH;L8H;%H;�H;��G;��G;5�G;W�G;�G;��G;[�G;      � H;.H;�H;�H;�H;|!H;G-H;�9H;GH;zTH;bH;uoH;�|H;	�H;��H;��H;W�H;'�H;'�H;D�H;u�H;��H;I�H;-�H;��H;N�H;��H;��H;�H;9�H;9�H;�H;��H;�H;L�H;��H;��H;��H;L�H;�H;��H;�H;9�H;7�H;	�H;��H;��H;N�H;��H;-�H;G�H;��H;t�H;D�H;'�H;'�H;U�H;��H;��H;�H;�|H;uoH;bH;yTH;GH;�9H;G-H;z!H;�H;�H;�H;9H;      "?H;�?H;\BH;�FH;OLH;RSH;�[H;ldH;�mH;�wH;�H;�H;ҕH;�H;��H;ׯH;]�H;$�H;L�H;��H;9�H;\�H;�H;�H;��H;��H;y�H;�H;U�H;&�H;��H;��H;�H;j�H;��H;��H;��H;��H;��H;j�H;�H;��H;��H;%�H;V�H;�H;y�H;��H;��H;�H;�H;]�H;7�H;��H;L�H;%�H;\�H;ׯH;��H;�H;ҕH;�H;�H;�wH;�mH;kdH;�[H;SSH;VLH;�FH;\BH;�?H;      iH;�iH;�kH;�nH;�rH;xH;�}H;��H;��H;�H;r�H;ΡH;�H;ۯH;n�H;��H;b�H;g�H;�H;"�H;��H; �H;��H;�H;��H;��H;'�H;9�H;%�H;�H;��H;�H;X�H;��H;��H;��H;��H;��H;��H;��H;T�H;�H;��H; �H;#�H;7�H;$�H;��H;��H;�H;��H; �H;��H;#�H;�H;h�H;`�H;��H;n�H;گH;�H;͡H;r�H;�H;��H;��H;�}H;xH;�rH;�nH;�kH;�iH;      k�H;�H;u�H;��H;ԏH;��H;�H;ǜH;ۡH;/�H;��H;0�H;��H;�H;��H;�H;��H;��H;�H;Q�H;,�H;��H;��H;��H;��H;L�H;f�H;:�H;��H;��H;�H;f�H;��H;��H;�H;�H;�H;�H;�H;��H;��H;h�H;�H;��H;��H;:�H;f�H;I�H;��H;��H;��H;��H;*�H;Q�H;�H;�H;��H;~�H;��H;�H;��H;/�H;��H;/�H;ۡH;ƜH;�H;��H;ҏH;��H;w�H;�H;      ��H;�H;��H;��H;�H;��H;ݪH;{�H;U�H;`�H;��H;��H;��H;��H;Y�H;��H;�H;.�H;��H;C�H;m�H;G�H;��H;Q�H;��H;��H;B�H;�H;��H;�H;b�H;��H;��H;�H;�H;:�H;V�H;:�H;�H;�H;��H;��H;c�H;�H;��H;�H;A�H;��H;��H;Q�H;��H;F�H;m�H;D�H;��H;0�H;	�H;��H;X�H;��H;��H;��H;��H;`�H;V�H;z�H;ߪH;��H;�H;��H; �H; �H;      W�H;��H;J�H;��H;?�H;R�H;ѸH;��H;��H;��H;��H;��H;��H;��H;��H;q�H;��H;>�H;i�H;I�H;��H;^�H;��H;��H;��H;h�H;�H;��H;�H;^�H;��H;��H;�H;/�H;T�H;H�H;<�H;H�H;T�H;/�H;�H;��H;��H;^�H;�H;��H;�H;e�H;��H;��H;��H;]�H;��H;L�H;i�H;?�H;��H;q�H;��H;��H;��H;��H;��H;��H;��H;��H;ѸH;V�H;8�H;��H;L�H;��H;      A�H;[�H;�H;��H;:�H;��H;��H;��H;��H;Q�H;��H;5�H;��H;�H;f�H;��H;��H;;�H;��H;u�H;��H;��H;��H;��H;h�H;*�H;��H;�H;i�H;��H;��H;�H;(�H;<�H;f�H;t�H;R�H;t�H;f�H;<�H;'�H;	�H;��H;��H;l�H;�H;��H;'�H;j�H;��H;��H;��H;��H;u�H;��H;=�H;��H;��H;f�H;�H;��H;5�H;��H;Q�H;��H;��H;��H;��H;0�H;��H;�H;S�H;      ��H;�H;��H;Q�H;_�H;��H;�H;��H;��H;��H;��H;��H;��H;��H;i�H;�H;��H;M�H;��H;��H;��H;��H;��H;|�H;�H;��H; �H;L�H;��H;��H;�H;�H;Q�H;i�H;K�H;i�H;��H;i�H;K�H;i�H;N�H; �H;�H;��H;��H;L�H;��H;��H;�H;{�H;��H;��H;��H;��H;��H;N�H;��H;�H;h�H;��H;��H;��H;��H;��H;��H;��H;�H;��H;T�H;S�H;��H;
�H;      ;�H;u�H;��H;l�H;m�H;��H;��H;p�H;�H;��H;g�H;(�H;��H;��H;$�H;��H;�H;g�H;��H;��H;��H;�H;>�H;��H;n�H;��H;8�H;��H;��H;��H;�H;?�H;G�H;w�H;i�H;`�H;p�H;`�H;i�H;t�H;F�H;A�H;�H;��H;��H;��H;6�H;��H;o�H;��H;>�H;�H;��H;��H;��H;i�H;�H;��H;$�H;��H;��H;(�H;e�H;��H;�H;m�H;��H;��H;`�H;l�H;��H;k�H;      ��H;��H;j�H;�H;��H;��H;�H;��H;�H;��H;Q�H;��H;��H;I�H;��H;>�H;��H;��H;��H;��H;��H;��H;��H;�H;v�H;��H;F�H;��H;��H;�H; �H;]�H;<�H;V�H;��H;q�H;\�H;q�H;��H;V�H;9�H;_�H; �H;�H;��H;��H;D�H;��H;v�H;�H;��H;��H;��H;��H;��H;��H;��H;>�H;��H;I�H;��H;��H;Q�H;��H;�H;��H;�H;��H;��H;�H;j�H;��H;      ;�H;u�H;��H;m�H;n�H;��H;��H;p�H;�H;��H;g�H;(�H;��H;��H;$�H;��H;�H;g�H;��H;��H;��H;�H;>�H;��H;o�H;��H;8�H;��H;��H;��H;�H;?�H;G�H;w�H;i�H;`�H;p�H;`�H;i�H;t�H;F�H;A�H;�H;��H;��H;��H;6�H;��H;n�H;��H;>�H;�H;��H;��H;��H;i�H;�H;��H;$�H;��H;��H;(�H;g�H;��H;�H;m�H;��H;��H;b�H;l�H;��H;k�H;      ��H;�H;��H;S�H;_�H;��H;�H;��H;��H;��H;��H;��H;��H;��H;h�H;�H;��H;M�H;��H;��H;��H;��H;��H;|�H;�H;��H; �H;L�H;��H;��H;�H;�H;Q�H;i�H;K�H;i�H;��H;i�H;K�H;i�H;N�H;!�H;�H;��H;��H;L�H;��H;��H;�H;y�H;��H;��H;��H;��H;��H;N�H;��H;�H;h�H;��H;��H;��H;��H;��H;��H;��H;�H;��H;T�H;Q�H;��H;
�H;      B�H;[�H;�H;��H;:�H;��H;��H;��H;��H;Q�H;��H;5�H;��H;�H;f�H;��H;��H;;�H;��H;t�H;��H;��H;��H;��H;j�H;)�H;��H;�H;i�H;��H;��H;�H;(�H;<�H;f�H;t�H;R�H;r�H;f�H;<�H;'�H;	�H;��H;��H;l�H;�H;��H;*�H;h�H;��H;��H;��H;��H;u�H;��H;=�H;��H;��H;f�H;�H;��H;5�H;��H;Q�H;��H;��H;��H;��H;/�H;��H;�H;S�H;      Z�H;��H;L�H;��H;>�H;T�H;ѸH;��H;��H;��H;��H;��H;��H;��H;��H;q�H;��H;>�H;i�H;J�H;��H;]�H;��H;��H;��H;g�H;�H;��H;�H;^�H;��H;��H;�H;.�H;T�H;H�H;<�H;H�H;T�H;.�H;�H;��H;��H;_�H;�H;��H;�H;g�H;��H;��H;��H;^�H;��H;J�H;i�H;>�H;��H;q�H;��H;��H;��H;��H;��H;��H;��H;��H;ѸH;X�H;5�H;��H;I�H;��H;      ��H;�H; �H;��H;�H;��H;�H;|�H;V�H;`�H;��H;��H;��H;��H;X�H;��H;�H;.�H;��H;F�H;q�H;F�H;��H;Q�H;��H;��H;A�H;�H;��H;�H;c�H;��H;��H;�H;�H;:�H;V�H;:�H;�H;�H;��H;��H;b�H;�H;��H;�H;A�H;��H;��H;Q�H;��H;G�H;k�H;C�H;��H;0�H;	�H;��H;X�H;��H;��H;��H;��H;b�H;X�H;z�H;�H;��H;�H;��H; �H;��H;      k�H;�H;u�H;��H;ԏH;��H;�H;ǜH;ۡH;-�H;��H;/�H;��H;�H;��H;�H;��H;~�H;�H;Q�H;.�H;��H;��H;��H;��H;J�H;f�H;:�H;��H;��H;�H;f�H;��H;��H;�H;�H;�H;�H;�H;��H;��H;h�H;�H;��H;��H;:�H;f�H;J�H;��H;��H;��H;��H;)�H;Q�H;�H;��H;��H;�H;��H;�H;��H;0�H;��H;0�H;ۡH;ǜH;�H;��H;ҏH;��H;u�H;�H;      iH;�iH;�kH;�nH;�rH;�wH;�}H;��H;��H;�H;r�H;ΡH;�H;ۯH;n�H;��H;b�H;g�H;�H;#�H;��H; �H;��H;�H;��H;��H;&�H;7�H;%�H;�H;��H;�H;U�H;��H;��H;��H;��H;��H;��H;��H;U�H;�H;��H; �H;%�H;9�H;$�H;��H;��H;�H;��H; �H;��H;"�H;�H;h�H;`�H;��H;n�H;گH;�H;ΡH;r�H;�H;��H;��H;�}H;xH;�rH;�nH;�kH;�iH;      ?H;�?H;cBH;�FH;VLH;OSH;�[H;ndH;�mH;�wH;�H;�H;ҕH;�H;��H;ׯH;]�H;$�H;L�H;��H;=�H;]�H;�H;�H;��H;��H;y�H;�H;V�H;&�H;��H;��H;�H;j�H;��H;��H;��H;��H;��H;j�H;�H;��H;��H;%�H;U�H;�H;{�H;��H;��H;�H;�H;\�H;6�H;��H;L�H;%�H;\�H;ٯH;��H;�H;ҕH;�H;�H;�wH;�mH;ldH;�[H;RSH;QLH;�FH;dBH;�?H;      � H;/H;�H;�H;�H;z!H;G-H;�9H;GH;yTH;bH;uoH;�|H;	�H;��H;��H;W�H;%�H;'�H;D�H;y�H;��H;I�H;-�H;��H;N�H;��H;��H;�H;:�H;9�H;�H;��H;�H;J�H;��H;��H;��H;L�H;�H;��H;�H;9�H;6�H;	�H;��H;��H;O�H;��H;-�H;G�H;��H;r�H;D�H;'�H;'�H;U�H;��H;��H;�H;�|H;uoH;bH;zTH;GH;�9H;G-H;y!H;�H;�H;�H;9H;      �G;[�G;��G;�G;P�G;4�G;��G;��G;�H;%H;L8H;�JH;�[H;�lH;|H;��H;��H;;�H;��H;��H;ӾH;��H;u�H;a�H;��H;S�H;6�H;��H;|�H;*�H;i�H;A�H;�H;��H;�H;8�H;F�H;6�H;�H;��H;�H;D�H;g�H;'�H;y�H;��H;4�H;T�H;��H;a�H;r�H;��H;ξH;��H;��H;;�H;��H;��H;|H;�lH;�[H;�JH;N8H;%H;�H;��G;��G;1�G;Q�G;�G;��G;S�G;      �wF;�F;ɖF;�F;4�F;�G;�NG;F�G;|�G;�G;��G;tH;�1H;HH;�\H;�oH;׀H;Q�H;НH;��H;�H;ӼH;}�H;��H;�H;��H;Q�H;L�H;��H;��H;I�H;��H;d�H;)�H;��H;��H;��H;��H;��H;)�H;c�H;��H;G�H;��H;��H;L�H;P�H;��H;
�H;��H;z�H;ѼH;޳H;��H;НH;Q�H;րH;�oH;�\H;HH;�1H;vH;��G;�G;}�G;E�G;�NG;�G;9�F;�F;ɖF;�F;      ��C;d	D;zBD;$�D;
E;ԄE;�F;�wF;�F;$=G;)�G;
�G;��G;-H;�4H;�MH;>dH;JxH;�H;��H;��H;�H;��H;��H;_�H;�H;��H;��H;��H;��H;��H;��H;��H;n�H;�H;s�H;|�H;r�H;�H;n�H;��H;��H;��H;��H;��H;��H;��H;�H;_�H;��H;��H;�H;��H;��H;��H;MxH;<dH;�MH;�4H;*H;��G;
�G;(�G;"=G;�F;�wF;�F;ԄE;
E;$�D;|BD;d	D;      _,>;nZ>;�>;��?;j�@;�A;�C;D;�E;��E;�F;G;~G;z�G;	�G;�!H;|@H;�ZH;lqH;_�H;m�H;¤H;�H;2�H;��H;��H;`�H;*�H;�H;�H;|�H;M�H;��H;��H;u�H;��H;
�H;��H;x�H;��H;��H;M�H;~�H;�H;�H;*�H;^�H;��H;��H;0�H;�H;¤H;i�H;^�H;jqH;�ZH;y@H;�!H;	�G;z�G;~G;G;�F;��E;�E;D;�C;�A;y�@;��?;�>;cZ>;      \�1;�J2;�g3;�$5;�Y7;�9;�g<;O�>;A;�C;@�D;A�E;}�F;L*G;c�G;i�G;�H;�5H;/SH;�lH;K�H;ɔH;?�H;�H;��H;~�H;v�H;G�H;�H;��H;��H;��H;��H;��H;��H;>�H;��H;>�H;��H;��H;��H;��H;��H;��H;�H;G�H;r�H;~�H;��H;�H;<�H;ʔH;D�H;�lH;/SH;�5H;�H;i�G;d�G;J*G;}�F;@�E;?�D;�C;A;N�>;�g<;�9;�Y7;�$5;�g3;qJ2;      �;��;*;�z ;��$;q�);�/;?4;$�8;g�<;*$@;~�B;R�D;��E;D�F;�cG;��G;�H;�-H;�NH;jH;\�H;ǔH;äH;�H;ԼH;��H;��H;\�H;�H;��H;B�H;]�H;��H;��H;~�H;��H;~�H;��H;��H;]�H;C�H;��H;��H;Y�H;��H;��H;ּH;�H;¤H;ŔH;^�H;jH;�NH;�-H;�H;��G;�cG;E�F;��E;Q�D;~�B;)$@;e�<;&�8;=4;�/;s�);��$;�z ;*;��;      ��:4��:Q��:���:�;�Y;�';��;��(;��0;Z7;j�<;(�@;aC;CCE;�wF;�8G;��G;}�G;�)H;�LH;jH;J�H;n�H;��H;�H;ϾH;v�H;9�H;��H;&�H;g�H;��H;��H;��H;��H;��H;��H;��H;��H;��H;j�H;&�H;��H;6�H;v�H;ξH;�H;��H;k�H;G�H;jH;�LH;�)H;}�G;��G;�8G;�wF;CCE;aC;(�@;j�<;Z7;��0;��(;��;�';�Y;�;���:K��:��:       �:�:�3<:*i:�t�:��:��:�+�:�Y;\�;�*';�1;P�8;�Z>;g0B;*�D;�2F;<G;��G;1�G;�)H;�NH;�lH;_�H;x�H;��H;��H;@�H;��H;�H;L�H;<�H;C�H;k�H;��H;��H;��H;��H;��H;k�H;B�H;<�H;J�H;�H;��H;B�H;��H;��H;z�H;\�H;�lH;�NH;�)H;2�G;��G;?G;�2F;)�D;g0B;�Z>;P�8;�1;�*';Z�;�Y;�+�:��:'��:�t�:*i:�3<:��:      ʥ���W��� ��4�=��ڷ���8�:�P�:�P�:���:H`;�;C�*;%5;�g<;=A; CD;%F;�G;��G;|�G;�-H;/SH;lqH;��H;ҝH;��H;(�H;L�H;�H;�H;��H;f�H;��H;��H;��H;��H;��H;��H;��H;d�H;��H;�H;�H;J�H;(�H;��H;ԝH;��H;iqH;*SH;�-H;z�G;��G;�G;'F;CD;=A;�g<;%5;C�*;�;F`;���:�P�:�P�:�:`�8Xڷ�8�=�� ���W��      �1��%Ȅ���u��PV�p.����pW������X�9x+i:��:>,�:7�;�t%;�J2;t;;ɵ@;�D;%F;@G;��G;�H;�5H;�ZH;HxH;S�H;=�H;)�H;'�H;k�H;�H;-�H;B�H;:�H;P�H;k�H;��H;k�H;P�H;;�H;A�H;.�H;��H;j�H;$�H;)�H;:�H;V�H;IxH;�ZH;�5H;�H;��G;AG;%F;�D;ɵ@;t;;�J2;�t%;7�;>,�:��:p+i:Y�9���nW�����k.��PV���u�*Ȅ�      Y��H�	������Tʻ�R���2|�X.��Ⱥp���Y�9du�:��:�Y;��!;��0;�:;ɵ@;"CD;�2F;�8G;��G;�H;@H;:dH;׀H;��H;W�H;Z�H;_�H;��H;�H;��H;�H;��H;�H;��H;�H;��H;��H;��H;�H;��H;]�H;Y�H;Z�H;��H;ڀH;:dH;{@H;�H;��G;�8G;�2F;"CD;ε@;�:;��0;��!;�Y;��:bu�:�Y�9|���ȺY.��2|��R��Tʻ�����K�	�      ��x��[t���g�PT�]�:�������&����1��:�(�W����t�ho`:���:];({ ;��0;w;;=A;/�D;�wF;�cG;i�G;�!H;�MH;�oH;��H;��H;֯H;��H;w�H;��H;m�H;�H;�H;��H;7�H;��H;�H;��H;k�H;��H;x�H;��H;ԯH;��H;��H;�oH;�MH;�!H;f�G;�cG;�wF;/�D;=A;w;;��0;){ ;];���:ho`: �t�
W��>�(��1��&���������^�:�PT���g��[t�      :,˼��Ǽ�"���뮼w��&G��+�[�ay-�����.����b�D0��׷�t5<:*M�:];��!;�J2;�g<;h0B;CCE;C�F;c�G;
�G;�4H;�\H;|H;��H;��H;j�H;��H;Q�H;��H;b�H;d�H;�H;��H;�H;b�H;b�H;��H;U�H;��H;k�H;��H;��H;|H;�\H;�4H;�G;`�G;C�F;CCE;j0B;�g<; K2;��!;];*M�:l5<:�׷�D0㺹�b��.�����ay-�+�[�&G��w���뮼�"����Ǽ      -���k��Kv��t�E�Ѽ�뮼-X��n�W������׻�Ǆ����@��|5<:���:�Y;�t%;%5;�Z>;aC;��E;L*G;{�G;(H;HH;�lH;�H;�H;֯H;�H;��H;��H;�H;��H;��H;@�H;��H;��H;�H;��H;��H;�H;֯H;�H;�H;�lH;HH;*H;y�G;G*G;��E;aC;�Z>;%5;�t%;�Y;���:t5<:H������Ǆ���׻���m�W�-X���뮼D�Ѽ�t�Kv���k�      Hm��Fi��&^�a�L�R�6�*���� }ռpT����x���0������������׷�ho`:��:9�;E�*;T�8;(�@;Q�D;�F;~G;��G;�1H;�[H;�|H;ѕH;�H;��H;��H;��H;��H;��H;��H;��H;��H;��H;��H;��H;��H;��H;�H;ЕH;�|H;�[H;�1H;��G;~G;{�F;Q�D;)�@;T�8;E�*;:�;��:ho`:�׷� ��������껿�0���x�pT�� }ռ��)��R�6�a�L��&^��Fi�      N��v;��C�������섽{�e��?��k�~t�鷼G���e7�����Ǆ�B0� �t�du�:>,�:�;�1;j�<;{�B;@�E;G;�G;sH;�JH;ooH;�H;��H;'�H;��H;��H;0�H;��H; �H;��H;!�H;��H;0�H;��H;��H;'�H;��H;�H;qoH;�JH;sH;
�G;G;=�E;{�B;n�<;�1;�;D,�:`u�:@�t�B0��Ǆ���껃e7�G��鷼~t��k��?�{�e��섽���C���v;��      s���(��s��ӽ�'��B�������Z��Q+�����"��G����0���׻��b�W���Y�9��:H`;�*';�Y7;$$@;@�D;�F;)�G;��G;K8H;bH;�H;j�H;��H;��H;��H;��H;��H;`�H;L�H;`�H;��H;��H;��H;��H;��H;j�H;�H;bH;K8H;��G;,�G;�F;=�D;$$@;Z7;�*';H`;��:�Y�9
W����b���׻��0�G���"������Q+��Z����B����'���ӽ�s�(��      �!,�:)��K ��������޽ ������Fi��0����鷼��x�����.��=�(�x��p+i:Ý�:Z�;��0;e�<;�C;��E;"=G;�G;%H;vTH;�wH;��H;(�H;]�H;��H;P�H;��H;��H;��H;��H;��H;P�H;��H;_�H;(�H;��H;�wH;vTH;%H;�G;&=G;��E;�C;e�<;��0;X�;Ý�:x+i:|��=�(��.�������x�鷼����0��Fi���� ���޽�������K �:)�      ,�j��f��Z�|�F��>/��^�p����ŽH ���Fi��Q+�}t�oT��n�W�����1���Ⱥ Y�9�P�:�Y;��(;"�8;A;�E;�F;}�G;�H;GH;�mH;��H;ѡH;O�H;�H;��H;��H;�H;�H;�H;��H;��H;|�H;Q�H;ԡH;��H;�mH;GH;�H;}�G;�F;�E;A;"�8;��(;�Y;�P�:Y�9�Ⱥ�1�����n�W�pT��}t�Q+��Fi�H ���Žp����^��>/�|�F��Z��f�      ��x���z�I����f��SC��K �qn���Ž����Z��k� }ռ-X��_y-�$���V.�����P�:�+�:��;84;O�>;D;�wF;G�G;��G;�9H;kdH;��H;��H;r�H;��H;��H;��H;d�H;��H;f�H;��H;��H;�H;r�H;��H;��H;hdH;�9H;��G;F�G;�wF;D;P�>;84;��;�+�:�P�:���X.�$���`y-�-X�� }ռ�k��Z�����Žqn���K ��SC��f�I���z�x���      ��˾��Ǿ����"���X͓�]�x���J��K �p��� ������?����뮼*�[�����2|�jW����:��:�';�/;~g<;�C;�F;�NG;��G;A-H;�[H;�}H;ٗH;ڪH;θH;��H;�H;��H;�H;��H;�H;��H;̸H;ڪH;ٗH;�}H;�[H;A-H;��G;�NG;�F;�C;|g<;�/;�';��:��:hW���2|����*�[��뮼���?���� ��p����K ���J�]�x�X͓�"���������Ǿ      u� ��������{Ծm���x���]�x��SC��^��޽B���{�e�*��E�Ѽ&G������R�������8'��:�Y;j�);�9;�A;фE;�G;2�G;|!H;SSH;�wH;��H;��H;T�H;��H;��H;��H;��H;��H;��H;��H;Q�H;��H;��H;�wH;OSH;|!H;1�G;�G;҄E;�A;�9;j�);�Y;'��:��8����R�����&G��E�Ѽ*��{�e�B����޽�^��SC�]�x�x���m����{Ծ�쾤���      ��� E�l�u� �X�ݾm���X͓��f��>/�����'���섽R�6��t�w��\�:�Tʻk.�Xڷ��t�:�;��$;�Y7;o�@;
E;3�F;M�G;�H;PLH;�rH;ƏH;ߤH;5�H;0�H;D�H;\�H;��H;]�H;C�H;0�H;4�H;�H;ƏH;�rH;OLH;�H;N�G;2�F;
E;m�@;�Y7;��$;�;�t�:Xڷ�k.�Tʻ\�:�w���t�R�6��섽�'������>/��f�X͓�m���X�ݾu� �l� E�      ��7�v3�1�'����u� ��{Ծ"���I���|�F�����ӽ���a�L�Lv��뮼PT����PV�4�=�(*i:���:�z ;�$5;ï?; �D;�F;
�G;�H;�FH;�nH;��H;��H;��H;��H;J�H;i�H;�H;i�H;J�H;��H;��H;��H;��H;�nH;�FH;�H;
�G;�F;!�D;��?;�$5;�z ;���: *i:0�=��PV���PT��뮼Lv�a�L�����ӽ���|�F�I���"����{Ծu� ����1�'�v3�      �N��TI���;�1�'�l��쾂���z󐾶Z��K ��s�C����&^���"����g����¨u�� ���3<:;��:;}g3;
�>;�BD;˖F;��G;�H;]BH;�kH;j�H;�H;@�H;�H;��H;��H;[�H;��H;��H;�H;?�H;��H;j�H;�kH;\BH;�H;��G;ʖF;�BD;�>;�g3;;?��:�3<:� ����u������g��"����&^�C����s潧K ��Z�z󐾂�����l�1�'���;��TI�      c]�g�W��TI�v3� E�������Ǿx����f�:)�(��v;���Fi��k���Ǽ�[t�J�	�$Ȅ��W����:(��:��;qJ2;gZ>;]	D;�F;W�G;-H;�?H;�iH;��H;��H;��H;M�H;��H;l�H;��H;l�H;��H;M�H;��H;��H;��H;�iH;�?H;+H;U�G;�F;]	D;cZ>;vJ2;��;(��:��:�W��$Ȅ�J�	��[t���Ǽ�k��Fi�v;��(��:)��f�x�����Ǿ���� E�v3��TI�g�W�      3�$��� ����%��B��*�þ�*��4Dx���=�����Pν	���''K��c�"��r�V����	E^�P�S�8x[:���:)e;m�4;V`?;�mD;��F;evG;L�G;�H;�OH;�sH;��H;��H;��H;/�H;��H;\�H;��H;/�H;��H;��H;��H;�sH;�OH;�H;L�G;evG;��F;�mD;R`?;p�4;)e;���:4x[:P�S�E^����r�V�"���c�''K�	����Pν�����=�4Dx��*��*�þB��%������� �      �� ����T��P��2������0��8�s�ڀ:�i9� �ʽ4Z���G��8�.���5S�����/X�,�D�$Cd:�B�:! ;4�4;ڈ?;D;_�F;(yG;��G;� H;TPH;StH;K�H;�H;�H;m�H;��H;o�H;��H;n�H;�H;�H;N�H;StH;QPH;� H;��G;(yG;]�F;D;ֈ?;:�4;! ;�B�:Cd:,�D��/X���껰5S�.���8��G�4Z�� �ʽi9�ڀ:�8�s��0�����2��P��T�����      ���T��:�
������Yؾ"���॒���f���0�][�R8��Ґ����>�����MȤ��6H�]�ܻ�qF�p����}:��:~";m�5;�?;��D;�F;$�G;��G;{#H;�RH;�uH;��H;��H;��H;�H;)�H;��H;)�H;�H;��H;��H;��H;�uH;�RH;x#H;��G;$�G;�F;��D;�?;p�5;~";��:��}:p���qF�^�ܻ�6H�MȤ�������>�Ґ��R8��][���0���f�॒�"����Yؾ����:�
�T��      %��P������AI�*�þ�R��=���wS��Q"��s������}��0��켋�����6�B�ƻ.}*�`���3�:�x;v%;m7;�@;�D;�F;��G;��G;>(H;VH;�xH;��H;~�H;ڲH;�H;��H;��H;��H;�H;ܲH;}�H;��H;�xH;VH;:(H;��G;��G;�F;�D;�@;m7;v%;�x;/�:`���,}*�B�ƻ��6��������0���}�����s��Q"�wS�=����R��*�þAIᾦ���P��      B��2�很Yؾ*�þĪ�~쏾�k�ڀ:���~�ؽ�����c�`y���Ҽ ���D� �b��� 8(7��:��
;�(;�_9;ΘA;�\E;��F;ޝG;��G;�.H;�ZH;&|H;.�H;��H;��H;M�H;�H;��H;�H;L�H;��H;��H;/�H;&|H;�ZH;�.H;��G;��G;��F;�\E;ɘA;�_9;�(;��
;��: 8(7��b�C� � �����Ҽ`y��c�����~�ؽ��ڀ:��k�~쏾Ī�*�þ�Yؾ2��      *�þ���"����R��~쏾8�s��H�����������ѐ����D��c�����@�f�S,�����P���9(��:�;Dj-;��;;��B;�E;�G;��G;��G;�6H;�`H;��H;��H;�H;��H;�H;��H;�H;��H;�H;��H;�H;��H;��H;�`H;�6H;��G;��G;�G;�E;��B;��;;Dj-;�;$��:�9�P�����S,�@�f������c���D�ѐ�������������H�8�s�~쏾�R��"������      �*���0��॒�=����k��H��#%�\[��Pν
t��d�f�6/%���伈���v�=��?ػzFL�l�D�΍R:R�:L�;W2;��=;ݚC;�0F;�GG;��G;[H;"@H;�gH;��H;n�H;�H;иH;��H;+�H;��H;+�H;��H;иH;�H;o�H;��H;�gH;@H;ZH;��G;�GG;�0F;ؚC;��=;W2;M�;L�:΍R:d�D�zFL��?ػv�=��������6/%�d�f�
t���Pν\[��#%��H��k�=���॒��0��      4Dx�8�s���f�wS�ڀ:����\[��7ս�榽��}���;��8�W�����r����6G�����ʬ�_��:9�;�}$;�6;9�?;�D;�F;�pG;��G;"H;dJH;noH;y�H;��H;7�H;u�H;��H;��H;d�H;��H;��H;u�H;5�H;��H;y�H;noH;`JH;"H;��G;�pG;�F;�D;9�?;�6;�}$;8�;_��:�ʬ����6G�������r�X����8���;���}��榽�7ս\[����ڀ:�wS���f�8�s�      ��=�ڀ:���0��Q"��������Pν�榽B����G�4����Ҽ ��KE:�:�ܻ�D^������i:~��:�;X|,;֡:;��A;jiE;��F;Z�G;��G;�(H;tUH;�wH;��H;c�H;ͳH;0�H;�H;��H;Q�H;��H;�H;/�H;̳H;e�H;��H;�wH;pUH;�(H;��G;Z�G;��F;eiE;��A;֡:;Z|,;�;~��:�i:�����D^�:�ܻKE:� ����Ҽ4����G�B���榽�Pν�������Q"���0�ڀ:�      ���j9�][��s�~�ؽ���
t����}� �G������2c��X�V�E,��*�����@����:V��:� ;��3;�0>; �C;F;9G;n�G;�H;*8H;�`H;:�H;*�H;7�H;��H;'�H;��H;�H;P�H;�H;��H;&�H;��H;:�H;*�H;:�H;�`H;)8H;�H;n�G;9G;F;��C;�0>;��3; ;V��:��:P������*��E,�X�V�2c���������G���}�
t������ؽ�s�][�j9�      �Pν �ʽR8���������ѐ��e�f���;�4�����EȤ�6�f�)��Jߵ�Jo5���D���-:y��:�>;�+;�_9;�A;��D;P�F;�vG;�G;SH;�GH;�lH;��H;ўH;2�H;g�H;1�H;��H;?�H;c�H;?�H;��H;0�H;d�H;4�H;ўH;��H;�lH;�GH;QH;�G;�vG;K�F;��D;�A;�_9;�+;�>;��:��-:��D�Io5�Iߵ�)��6�f�EȤ����4����;�e�f�ѐ���������R8�� �ʽ      	���4Z��Ґ����}��c���D�6/%��8���Ҽ2c��6�f�����ƻr/X�8���H��9C�:W�;�";��3;e>;rYC;��E;	G;&�G;��G;�,H;>WH;OxH;đH;o�H;&�H;K�H;)�H;o�H;}�H;n�H;}�H;p�H;)�H;K�H;'�H;m�H;ÑH;MxH;>WH;�,H;��G;$�G;G;��E;rYC;e>;��3;�";Z�;A�:P��98���r/X��ƻ���5�f�2c����Ҽ�8�6/%���D��c���}�Ґ��5Z��      ('K��G���>��0�`y��c����X��� ��Y�V�(���ƻ�od�`�º �(7�4�:���:¡;Q.;	�:;<zA;`�D;�F;�nG;x�G;,H;�@H;_fH;��H;g�H;�H;�H;#�H;)�H;��H;��H;x�H;��H;��H;(�H;#�H;�H;�H;f�H;��H;_fH;�@H;,H;u�G;}nG;��F;`�D;<zA;�:;Q.;ġ;���:�4�: �(7`�º�od��ƻ(��X�V� ��X�����优c�ay��0���>��G�      �c��8���������Ҽ����������r�JE:�E,�Hߵ�r/X�`�º@Ĭ���}:?�:;g�);Nm7;E�?;��C;8F;�)G;H�G;��G;@*H;�SH;�tH;��H;��H;.�H;�H;��H;�H;M�H;��H;��H;��H;M�H;�H;��H;�H;.�H;��H;��H;�tH;�SH;@*H;��G;E�G;�)G;8F;��C;C�?;Nm7;j�);;=�:��}: Ĭ�`�ºq/X�Hߵ�D,�JE:���r�����������Ҽ�켻����8�      "��.��NȤ����� ���A�f�w�=����;�ܻ�*��Jo5�:��� �(7��}:�n�:I�;�>&;��4;�=;��B;�E;E�F;ʁG;,�G;kH;�AH;�eH;z�H;�H;��H;�H;��H;]�H;��H;��H;��H;��H;��H;��H;��H;\�H;��H;�H;��H;�H;z�H;�eH;�AH;hH;&�G;āG;E�F;�E;��B;�=;��4;�>&;K�;�n�:��}: �(7:���Jo5��*��:�ܻ���w�=�@�f� �������MȤ�.��      q�V��5S��6H���6�E� �T,��?ػ8G���D^������D�H��9�4�:;�:L�;%;��3;A�<;�B;�E;1�F;�XG;<�G;� H;�0H;�WH;�vH;-�H;��H;��H;νH;�H;��H;��H;��H;��H;w�H;��H;��H;��H;��H;�H;ͽH;��H;��H;,�H;�vH;�WH;�0H;z H;8�G;�XG;.�F;�E;�B;B�<;��3;%;L�;?�:�4�:H��9��D�����D^�9G���?ػS,�E� ���6��6H��5S�      ��ﻧ��_�ܻD�ƻd󩻲��wFL��������@����-:C�:���:;�>&;��3;~9<;:�A;�D;yZF;T5G;3�G;�G;�!H;nJH;nkH;߅H;��H;��H;ظH;&�H;��H;��H;�H;��H;��H;/�H;��H;��H;�H;��H; �H;&�H;ָH;��H;��H;ۅH;okH;mJH;�!H;�G;3�G;S5G;yZF;�D;<�A;~9<;��3;�>&;;���:C�:��-:0���������wFL����c�D�ƻ_�ܻ���      E^��/X��qF�,}*�$���P��t�D� ˬ��i:��:}��:W�;¡;f�);��4;>�<;9�A;L�D;�9F;G;��G;|�G;vH;U?H;�aH;P}H;��H;��H;ֳH;�H; �H;��H;��H;W�H;��H;^�H;��H;^�H;��H;V�H;��H;��H;��H;�H;ӳH;��H;��H;Q}H;�aH;P?H;sH;|�G;��G;G;�9F;N�D;7�A;>�<;��4;g�);¡;X�;��:��:�i:@ˬ�p�D��P����,}*��qF�0X�      <�S�@�D�P��p��� 3(7�9ލR:Y��:���:V��:�>;�";Q.;Pm7;�=;�B;�D;�9F;RG;U�G;��G;�H;�6H;�YH;vH;\�H;,�H;;�H;>�H;��H;^�H;��H;U�H;s�H;��H;��H;2�H;��H;��H;s�H;T�H;��H;]�H;��H;;�H;:�H;'�H;^�H;vH;�YH;�6H;�H;��G;V�G;RG;�9F;
�D;�B;�=;Nm7;Q.;�";�>;V��:���:W��:ލR:H�9 9(7h���P��<�D�      8x[:\Cd:��}:1�:��:��:H�:5�;�;� ;�+;��3;�:;>�?;��B;�E;uZF;G;Q�G;��G;zH;�1H;TH;�pH;�H;��H;#�H;��H;��H;��H;:�H;�H;��H;]�H;1�H;Q�H;��H;Q�H;1�H;\�H;��H;�H;:�H;��H;��H;��H;!�H;��H;�H;�pH;TH;�1H;wH;��G;R�G;G;wZF;�E;��B;>�?;�:;��3;�+;� ;�;5�;H�:$��:��:/�:��}:<Cd:      ��:�B�:��:�x;��
;�;M�;�}$;U|,;��3;�_9;b>;9zA;��C;�E;/�F;S5G;��G;��G;{H;�/H;-QH;?mH;��H;ٗH;ЧH;��H;7�H;��H;T�H;��H;��H;��H; �H;��H;��H;��H;��H;��H;�H;��H;��H;��H;Q�H;��H;9�H;��H;ЧH;ٗH;��H;<mH;.QH;�/H;}H;��G;��G;Q5G;1�F;�E;��C;:zA;b>;�_9;��3;Z|,;�}$;N�;�;��
;�x;��:�B�:      1e;; ;�";n%;�(;Kj-;a2;��6;١:;�0>;�A;rYC;^�D;8F;F�F;�XG;0�G;~�G;�H;�1H;+QH;lH;��H;��H;s�H;j�H;�H;��H;��H;K�H;��H;�H;��H;��H;��H;��H;��H;��H;��H;��H;��H;�H;��H;G�H;��H;��H;�H;m�H;t�H;��H;��H;lH;+QH;�1H;�H;�G;2�G;�XG;G�F;8F;`�D;rYC;�A;�0>;ܡ:;�6;`2;Mj-;#�(;n%;�";4 ;      u�4;6�4;m�5;m7;�_9;��;;��=;9�?;��A;��C;��D;��E;��F;�)G;ȁG;9�G;�G;wH;�6H;TH;?mH;��H;�H;E�H;��H;��H;d�H;o�H;�H;��H;T�H;)�H;p�H;��H;��H;��H;��H;��H;��H;��H;n�H;)�H;T�H;��H;�H;o�H;a�H;��H;��H;E�H;�H;��H;;mH;TH;�6H;yH;�G;8�G;ȁG;�)G;��F;��E;��D;��C;��A;8�?;��=;��;;�_9;m7;p�5;(�4;      j`?;�?;�?;�@;͘A;��B;�C;�D;hiE;F;L�F;	G;}nG;F�G;(�G;} H;�!H;U?H;�YH;�pH;��H;��H;E�H;��H;˺H;g�H;��H;C�H;��H;��H;��H;��H;��H;�H;��H;r�H;��H;q�H;��H;	�H;��H;��H;��H;��H;��H;C�H;��H;g�H;κH;��H;C�H;��H;��H;�pH;�YH;V?H;�!H;} H;)�G;F�G;}nG;	G;L�F;F;hiE;�D;�C;��B;ԘA;�@;�?;ڈ?;      �mD;D;{�D;�D;�\E;�E;�0F;��F;��F;9G;�vG;&�G;u�G;��G;kH;�0H;rJH;�aH;$vH; �H;ݗH;w�H;��H;ӺH;)�H;�H;��H;O�H;%�H;6�H;��H;{�H;��H;�H;��H;"�H;e�H;!�H;��H;�H;��H;}�H;��H;6�H;#�H;O�H;��H;�H;*�H;ҺH;��H;x�H;ۗH;"�H;%vH;�aH;qJH;�0H;kH;��G;u�G;&�G;�vG;9G;��F;��F;�0F;�E;�\E;�D;y�D;D;      ��F;k�F;ܮF;�F;��F;�G;�GG;�pG;X�G;n�G;�G;��G;+H;?*H;�AH;�WH;kkH;M}H;Z�H;��H;̧H;i�H;��H;e�H;��H;t�H;��H;��H;��H;P�H;L�H;��H;��H;��H;t�H;��H;�H;��H;u�H;��H;��H;��H;N�H;P�H;��H;��H;��H;u�H;�H;d�H;��H;j�H;ɧH;��H;Z�H;N}H;kkH;�WH;�AH;?*H;+H;��G;�G;m�G;Z�G;�pG;�GG;�G;��F;�F;ܮF;`�F;      svG;-yG;#�G;��G;�G;��G;�G;��G;��G;�H;PH;�,H;�@H;�SH;�eH;�vH;߅H;��H;*�H;%�H;��H;�H;d�H;��H;��H; �H;��H;��H;�H;�H;��H;��H;��H;��H;�H;a�H;a�H;a�H;�H;�H;��H;��H;��H;�H;�H;��H;��H;��H;��H;��H;b�H;�H;��H;&�H;,�H;��H;߅H;�vH;�eH;�SH;�@H;�,H;PH;�H;��G;��G;�G;��G;�G;��G;$�G;+yG;      B�G;��G;��G;��G;��G;��G;`H;(H;�(H;-8H;�GH;DWH;`fH;�tH;z�H;,�H;��H;��H;9�H;��H;7�H;��H;q�H;F�H;J�H;��H;��H;��H;��H;��H;��H;��H;��H;�H;��H;��H;��H;��H;��H;�H;��H;��H;��H;��H;��H;��H;��H;��H;L�H;H�H;o�H;��H;6�H;��H;9�H;��H;��H;-�H;{�H;�tH;_fH;DWH;�GH;-8H;�(H;(H;`H;��G;��G;��G;��G;��G;      �H;� H;y#H;A(H;�.H;�6H;%@H;dJH;tUH;�`H;�lH;QxH;��H;��H;�H;��H;��H;ӳH;>�H;��H;��H;��H;�H;��H;�H;��H;�H;��H;p�H;��H;��H;��H;,�H;��H;��H;�H;.�H;�H;��H;��H;)�H;��H;��H;��H;o�H; �H;�H;��H; �H;��H;�H;��H;��H;��H;>�H;ӳH;��H;��H;�H;��H;��H;QxH;�lH;�`H;wUH;dJH;%@H;�6H;�.H;A(H;y#H;� H;      �OH;[PH;�RH;VH;�ZH;�`H;�gH;uoH;�wH;B�H;��H;БH;k�H;��H;��H;��H;ڸH;�H;��H;��H;T�H;H�H;��H;��H;-�H;N�H;�H;��H;��H;��H;��H;)�H;��H;�H;;�H;^�H;s�H;^�H;;�H;�H;��H;)�H;��H;��H;��H;��H;�H;L�H;/�H;��H;��H;H�H;T�H;��H;��H;�H;ظH;��H;��H;��H;k�H;БH;��H;B�H;�wH;voH;�gH;�`H;�ZH;VH;�RH;XPH;      �sH;etH;�uH;�xH;5|H;��H;ɅH;��H;��H;-�H;՞H;x�H;�H;3�H;�H;սH;,�H;��H;`�H;A�H;��H;��H;T�H;��H;��H;O�H;��H;��H;��H;��H;�H;��H;�H;N�H;��H;��H;��H;��H;��H;N�H;�H;��H;�H;��H;��H;��H;��H;N�H;��H;��H;P�H;��H;��H;B�H;a�H;��H;*�H;ԽH;�H;2�H;�H;w�H;՞H;.�H;��H;��H;ʅH;��H;3|H;�xH;�uH;etH;      �H;W�H;��H;��H;5�H;��H;p�H;��H;f�H;7�H;7�H;-�H;�H;�H;��H;�H;�H;��H;��H;�H;��H;"�H;*�H;��H;x�H;��H;��H;��H;��H;*�H;��H;�H;J�H;��H;��H;��H;��H;��H;��H;��H;G�H;�H;��H;,�H;��H;��H;��H;��H;{�H;��H;'�H;"�H;��H;�H;��H;��H;�H;�H;��H;�H;�H;.�H;7�H;7�H;h�H;��H;p�H;��H;2�H;��H;��H;S�H;      ��H;�H;�H;��H;��H;�H;�H;?�H;ҳH;��H;g�H;S�H;(�H;��H;`�H;��H;��H;��H;V�H;��H;��H;��H;q�H;��H;��H;��H;��H;��H;0�H;��H;�H;N�H;��H;��H;��H;��H;	�H;��H;��H;��H;��H;P�H;�H;��H;1�H;��H;��H;��H;��H;��H;p�H;��H;��H;��H;X�H;��H;��H;��H;_�H;��H;(�H;R�H;g�H;��H;ҳH;<�H;�H;�H;��H;��H;�H;	�H;      ʰH;�H;��H;߲H;��H;��H;ָH;}�H;5�H;(�H;7�H;/�H;+�H;�H;��H;��H;�H;W�H;v�H;e�H;'�H;��H;��H;�H;�H;��H;|�H;�H;��H;�H;L�H;��H;��H;��H;��H;�H;�H;�H;��H;��H;��H;��H;J�H;�H;��H;�H;|�H;��H;�H;�H;��H;��H;&�H;e�H;w�H;Y�H;�H;��H;��H;�H;+�H;/�H;5�H;(�H;6�H;|�H;ָH;��H;��H;�H;��H;�H;      .�H;��H;�H;��H;f�H;ݾH;��H;��H; �H;��H;�H;z�H;��H;T�H;��H;��H;��H;��H;��H;9�H;��H;��H;��H;�H;��H;r�H;�H;��H;��H;=�H;��H;��H;��H;��H;�H;�H;�H;�H;�H;��H;��H;��H;��H;=�H;��H;��H;�H;t�H;��H;��H;��H;��H;��H;9�H;��H;��H;��H;��H;��H;T�H;��H;z�H;��H;��H; �H;��H;��H;�H;[�H;��H;�H;z�H;      ��H;��H;1�H;�H;+�H;��H;4�H;�H;�H;�H;F�H;��H;��H;��H;��H;��H;��H;Z�H;��H;[�H;��H;��H;��H;w�H;�H;��H;`�H;��H;�H;_�H;��H;��H;��H;�H;�H;/�H;'�H;/�H;�H;�H;��H;��H;��H;a�H;�H;��H;^�H;��H;�H;u�H;��H;��H;��H;[�H;��H;\�H;��H;��H;��H;��H;��H;��H;F�H;�H;�H;�H;4�H;��H;�H;�H;3�H;��H;      _�H;v�H;��H;��H;��H;�H;��H;i�H;X�H;P�H;j�H;w�H;|�H;��H;��H;~�H;7�H;��H;4�H;��H;��H;��H;��H;��H;a�H;�H;`�H;��H;/�H;z�H;��H;��H;�H;�H;�H;(�H;0�H;(�H;�H;�H;�H;��H;��H;z�H;2�H;��H;^�H;�H;a�H;��H;��H;��H;��H;��H;4�H;��H;6�H;~�H;��H;��H;|�H;w�H;j�H;S�H;Y�H;g�H;��H;�H;��H;��H;��H;l�H;      ��H;��H;1�H;�H;+�H;��H;4�H;�H;�H;�H;F�H;��H;��H;��H;��H;��H;��H;Z�H;��H;[�H;��H;��H;��H;w�H;�H;��H;`�H;��H;�H;_�H;��H;��H;��H;�H;�H;/�H;'�H;/�H;�H;�H;��H;��H;��H;a�H;�H;��H;^�H;��H;�H;w�H;��H;��H;��H;[�H;��H;\�H;��H;��H;��H;��H;��H;��H;G�H;�H;�H;�H;5�H;��H;�H;�H;0�H;��H;      ,�H;��H;�H;��H;f�H;ݾH;��H;��H;�H;��H;��H;z�H;��H;T�H;��H;��H;��H;��H;��H;9�H;��H;��H;��H;�H;��H;t�H;�H;��H;��H;=�H;��H;��H;��H;��H;�H;�H;�H;�H;�H;��H;��H;��H;��H;?�H;��H;��H;�H;t�H;��H;��H;��H;��H;��H;9�H;��H;��H;��H;��H;��H;T�H;��H;z�H;��H;��H; �H;��H;��H;�H;[�H;��H;�H;x�H;      ̰H;�H;��H;�H;��H;��H;ָH;}�H;5�H;(�H;7�H;/�H;+�H;�H;��H;��H;�H;W�H;w�H;d�H;*�H;��H;��H;�H;�H;��H;|�H;�H;��H;�H;J�H;��H;��H;��H;��H;�H;�H;�H;��H;��H;��H;��H;L�H;�H;��H;�H;|�H;��H;�H;�H;��H;��H;&�H;e�H;v�H;Z�H;�H;��H;��H;�H;+�H;/�H;7�H;(�H;6�H;|�H;ָH;��H;��H;߲H;��H;�H;      ��H;�H;�H;��H;��H;�H;�H;>�H;ҳH;��H;g�H;R�H;&�H;��H;_�H;��H;��H;��H;X�H;��H;��H;��H;q�H;��H;��H;��H;��H;��H;0�H;��H;�H;N�H;��H;��H;��H;��H;	�H;��H;��H;��H;��H;Q�H;�H;��H;1�H;��H;��H;��H;��H;��H;p�H;��H;��H;��H;V�H;��H;��H;��H;`�H;��H;&�H;S�H;g�H;��H;ҳH;;�H;�H;�H;�H;��H;�H;�H;      �H;W�H;��H;��H;5�H;��H;s�H;��H;f�H;9�H;7�H;-�H;�H;�H;��H;�H;�H;��H;��H;�H;��H;"�H;*�H;��H;{�H;��H;��H;��H;��H;*�H;��H;�H;I�H;��H;��H;��H;��H;��H;��H;��H;G�H;�H;��H;,�H;��H;��H;��H;��H;x�H;��H;)�H;"�H;��H;�H;��H;��H;�H;�H;��H;�H;�H;.�H;7�H;9�H;h�H;��H;s�H;��H;1�H;��H;��H;S�H;      �sH;etH;�uH;�xH;5|H;��H;ʅH;��H;��H;-�H;՞H;w�H;�H;3�H;�H;սH;*�H;��H;a�H;B�H;��H;��H;T�H;��H;��H;O�H;��H;��H;��H;��H;�H;��H;�H;N�H;��H;��H;��H;��H;��H;N�H;�H;��H;�H;��H;��H;��H;��H;N�H;��H;��H;Q�H;��H;��H;A�H;`�H;��H;*�H;սH;�H;3�H;�H;x�H;ӞH;.�H;��H;��H;ɅH;��H;3|H;�xH;�uH;dtH;      �OH;ZPH;�RH;VH;�ZH;�`H;�gH;xoH;�wH;A�H;��H;БH;k�H;��H;��H;��H;ڸH;�H;��H;��H;X�H;H�H;��H;��H;/�H;M�H;�H;��H;��H;��H;��H;)�H;��H;�H;;�H;^�H;s�H;^�H;;�H;�H;��H;*�H;��H;��H;��H;��H;�H;M�H;-�H;��H;��H;H�H;R�H;��H;��H;�H;ظH;��H;��H;��H;k�H;БH;��H;A�H;�wH;xoH;�gH;�`H;�ZH;VH;�RH;ZPH;      �H;� H;�#H;?(H;�.H;�6H;)@H;fJH;tUH;�`H;�lH;SxH;��H;��H;�H;��H;��H;ҳH;>�H;��H;��H;��H;�H;��H; �H;��H;�H; �H;o�H;��H;��H;��H;*�H;��H;��H;�H;.�H;�H;��H;��H;*�H;��H;��H;��H;o�H;��H;�H;��H;�H;��H;�H;��H;��H;��H;>�H;ԳH;��H;��H;�H;��H;��H;QxH;�lH;�`H;vUH;dJH;'@H;�6H;�.H;<(H;�#H;� H;      B�G;��G;��G;��G;��G;��G;`H;)H;�(H;-8H;�GH;DWH;_fH;�tH;{�H;-�H;��H;��H;9�H;��H;;�H;��H;q�H;F�H;L�H;��H;��H;��H; �H;��H;��H;��H;��H;�H;��H;��H;��H;��H;��H;�H;��H;��H;��H;��H;��H;��H;��H;��H;J�H;H�H;o�H;��H;6�H;��H;9�H;��H;��H;-�H;z�H;�tH;`fH;DWH;�GH;-8H;�(H;(H;`H;��G;��G;��G;��G;��G;      nvG;.yG;%�G;��G;��G;��G;�G;��G;��G;�H;PH;�,H;�@H;�SH;�eH;�vH;߅H;��H;,�H;&�H;��H;�H;d�H;��H;��H; �H;��H;��H;�H;�H;��H;��H;��H;�H;�H;a�H;a�H;`�H;�H;�H;��H;��H;��H;�H;�H;��H;��H; �H;��H;��H;b�H;�H;��H;%�H;*�H;��H;ޅH;�vH;�eH;�SH;�@H;�,H;QH;�H;��G;��G;�G;��G;�G;��G;$�G;&yG;      ��F;g�F;�F;	�F;��F;�G;�GG;�pG;X�G;n�G;�G;��G;+H;?*H;�AH;�WH;mkH;M}H;Z�H;��H;ϧH;j�H;��H;d�H;�H;t�H;��H;��H;��H;Q�H;N�H;��H;��H;��H;r�H;��H;�H;��H;u�H;��H;��H;��H;L�H;M�H;��H;��H;��H;u�H;��H;d�H;��H;i�H;ȧH;��H;Z�H;N}H;jkH;�WH;�AH;?*H;+H;��G;�G;m�G;X�G;�pG;�GG;�G;��F;�F;�F;]�F;      �mD;D;y�D;�D;�\E;�E;�0F;�F;��F;9G;�vG;&�G;u�G;��G;kH;�0H;qJH;�aH;%vH;"�H;ޗH;x�H; �H;ӺH;*�H;�H;��H;O�H;&�H;7�H;��H;|�H;��H;�H;��H;"�H;e�H;!�H;��H;�H;��H;}�H;��H;4�H;"�H;O�H;��H;�H;)�H;ҺH;��H;w�H;ۗH;"�H;$vH;�aH;pJH;�0H;kH;��G;u�G;&�G;�vG;9G;��F;��F;�0F;�E;�\E;�D;y�D;D;      p`?;�?;�?;�@;ɘA;��B;ޚC;�D;jiE;F;N�F;	G;~nG;F�G;)�G;} H;�!H;S?H;�YH;�pH;��H;��H;F�H;��H;κH;e�H;��H;C�H;��H;��H;��H;��H;��H;�H;��H;r�H;��H;q�H;��H;�H;��H;��H;��H;��H;��H;C�H;��H;g�H;˺H;��H;B�H;��H;��H;�pH;�YH;V?H;�!H;} H;(�G;F�G;}nG;	G;K�F;F;jiE;�D;ޚC;��B;ؘA;�@;�?;׈?;      n�4;A�4;��5;
m7;�_9;��;;��=;9�?;��A;��C;��D;��E;��F;�)G;ȁG;9�G;�G;uH;�6H;TH;@mH;��H;�H;F�H;��H;��H;d�H;o�H;�H;��H;T�H;)�H;q�H;��H;��H;��H;��H;��H;��H;��H;n�H;)�H;T�H;��H;�H;o�H;b�H;��H;��H;C�H;�H;��H;;mH;TH;�6H;yH;�G;9�G;ʁG;�)G;��F;��E;��D;��C;��A;8�?;��=;��;;�_9;
m7;t�5;3�4;      1e;: ;�";n%;�(;Kj-;`2;��6;١:;�0>;�A;rYC;`�D;9F;F�F;�XG;0�G;~�G;�H;�1H;.QH;lH;��H;��H;t�H;k�H;�H;��H;��H;K�H;��H;�H;��H;��H;��H;��H;��H;��H;��H;��H;��H;�H;��H;G�H;��H;��H;�H;k�H;s�H;��H;��H;lH;+QH;�1H;�H;�G;/�G;�XG;G�F;7F;^�D;tYC;�A;�0>;ܡ:;��6;a2;Kj-;!�(;n%;�";6 ;      ���:�B�:��:�x;��
;�;Q�;�}$;W|,;��3;�_9;b>;:zA;��C;�E;1�F;S5G;��G;��G;{H;�/H;.QH;=mH;��H;ٗH;ϧH;��H;9�H;��H;T�H;��H;��H;��H;�H;��H;��H;��H;��H;��H; �H;��H;��H;��H;Q�H;��H;7�H;��H;ЧH;ٗH;��H;=mH;-QH;�/H;}H;��G;��G;Q5G;/�F;�E;��C;9zA;b>;�_9;��3;W|,;�}$;Q�;�;��
;�x;��:�B�:      4x[:dCd:��}:+�:��:��:L�:7�;�;� ;�+;��3;�:;>�?;��B;�E;wZF;G;R�G;��G;{H;�1H;TH;�pH;�H;��H;#�H;��H;��H;��H;:�H;�H;��H;\�H;1�H;R�H;��H;R�H;1�H;]�H;��H;�H;:�H;��H;��H;��H;!�H;��H;�H;�pH;TH;�1H;xH;��G;Q�G;G;uZF;�E;��B;>�?;�:;��3;�+;� ;�;7�;L�:$��:��:+�:��}:8Cd:      <�S�@�D�P��h��� 4(7�9ލR:[��:���:V��:�>;�";Q.;Nm7;�=;�B;�D;�9F;RG;U�G;��G;�H;�6H;�YH;vH;[�H;*�H;:�H;>�H;��H;]�H;��H;U�H;s�H;��H;��H;2�H;��H;��H;s�H;T�H;��H;^�H;��H;;�H;;�H;)�H;^�H;vH;�YH;�6H;�H;��G;V�G;RG;�9F;
�D;�B;�=;Nm7;Q.;�";�>;V��:���:Y��:ލR:H�9 9(7p���P��<�D�      E^��/X��qF�,}*�%���P��p�D� ˬ��i:��:}��:X�;¡;f�);��4;>�<;9�A;L�D;�9F;G;��G;|�G;vH;U?H;�aH;N}H;��H;��H;ԳH;�H;��H;��H;��H;V�H;��H;^�H;��H;^�H;��H;W�H;��H;��H; �H;�H;ӳH;��H;��H;Q}H;�aH;P?H;sH;|�G;��G;G;�9F;N�D;7�A;>�<;��4;f�);¡;W�;}��:��:�i:@ˬ�p�D��P����,}*��qF�0X�      ��ﻨ��_�ܻE�ƻd󩻳��wFL�������� ����-:C�:���:;�>&;��3;�9<;9�A;�D;yZF;S5G;3�G;�G;�!H;mJH;nkH;߅H;��H;��H;ظH;&�H;��H;��H;�H;��H;��H;/�H;��H;��H;�H;��H; �H;&�H;׸H;��H;��H;ۅH;okH;nJH;�!H;�G;3�G;S5G;{ZF;�D;<�A;~9<;��3;�>&;;���:C�:��-:P���������wFL����c�D�ƻ_�ܻ���      r�V��5S��6H���6�D� �T,��?ػ8G���D^�����D�P��9�4�:;�:L�;%;��3;A�<;�B;�E;/�F;�XG;;�G;~ H;�0H;�WH;�vH;,�H;��H;��H;ͽH;�H;��H;��H;��H;��H;w�H;��H;��H;��H;��H;�H;νH;��H;��H;-�H;�vH;�WH;�0H;| H;8�G;�XG;/�F;�E;�B;B�<;��3;%;N�;;�:�4�:H��9��D�����D^�8G���?ػS,�E� ���6��6H��5S�      "��.��NȤ����� ���A�f�w�=����<�ܻ�*��Jo5�8��� �(7��}:�n�:K�;�>&;��4;�=;��B;�E;E�F;ʁG;,�G;hH;�AH;�eH;z�H;�H;��H;�H;��H;_�H;��H;��H;��H;��H;��H;��H;��H;]�H;��H;�H;��H;�H;z�H;�eH;�AH;kH;(�G;ƁG;E�F;�E;��B;�=;��4;�>&;I�;�n�:��}: �(7:���Jo5��*��;�ܻ���w�=�@�f� �������NȤ�.��      �c��8���������Ҽ����������r�JE:�D,�Hߵ�r/X�^�º@Ĭ���}:=�:;i�);Nm7;B�?;��C;8F;�)G;H�G;��G;?*H;�SH;�tH;��H;��H;.�H;�H;��H;�H;M�H;��H;��H;��H;M�H;�H;��H;�H;.�H;��H;��H;�tH;�SH;@*H;��G;E�G;�)G;8F;��C;B�?;Nm7;j�);;?�:��}:`Ĭ�`�ºr/X�Iߵ�E,�JE:���r�����������Ҽ�켻����8�      ('K��G���>��0�`y��c����X��� ��X�V�(���ƻ�od�`�º �(7�4�:���:¡;Q.;�:;:zA;`�D;��F;�nG;u�G;+H;�@H;_fH;��H;f�H;�H;�H;#�H;(�H;��H;��H;x�H;��H;��H;)�H;"�H;�H;�H;g�H;��H;_fH;�@H;/H;x�G;{nG;��F;`�D;<zA;�:;Q.;ġ;���:�4�: �(7`�º�od��ƻ(��X�V� ��X�����优c�`y��0���>��G�      	���4Z��Ґ����}��c���D�6/%��8���Ҽ2c��5�f�����ƻr/X�6���P��9C�:X�;�";��3;b>;rYC;��E;G;$�G;��G;�,H;>WH;OxH;đH;m�H;%�H;L�H;*�H;p�H;�H;n�H;�H;o�H;)�H;I�H;'�H;o�H;đH;MxH;>WH;�,H;��G;&�G;G;��E;rYC;f>;��3;�";Z�;A�:@��96���r/X��ƻ���6�f�2c����Ҽ�8�6/%���D��c���}�Ґ��5Z��      �Pν �ʽR8���������ѐ��e�f���;�4�����EȤ�6�f�(��Jߵ�Io5���D���-:}��:�>;�+;�_9;�A;��D;P�F;�vG;�G;SH;�GH;�lH;��H;ўH;2�H;e�H;0�H;��H;?�H;c�H;?�H;��H;1�H;e�H;3�H;ўH;��H;�lH;�GH;QH;�G;�vG;K�F;��D;�A;�_9;�+;�>;��:��-:��D�Jo5�Jߵ�)��6�f�EȤ����4����;�e�f�ѐ���������R8�� �ʽ      ���j9�][��s�~�ؽ���
t����}� �G������2c��X�V�E,��*�����@����:V��:� ;��3;�0>;��C;F;9G;n�G;�H;)8H;�`H;:�H;*�H;7�H;��H;&�H;��H;�H;P�H;�H;��H;'�H;��H;9�H;*�H;:�H;�`H;*8H;�H;n�G;9G;F; �C;�0>;��3; ;V��:��:`������*��E,�X�V�2c������� �G���}�
t������ؽ�s�][�j9�      ��=�ڀ:���0��Q"��������Pν�榽B����G�4����Ҽ ��KE:�:�ܻ�D^������i:~��:�;W|,;֡:;��A;jiE;��F;Z�G;��G;�(H;sUH;�wH;��H;c�H;ϳH;/�H;�H;��H;Q�H;��H;�H;0�H;̳H;c�H;��H;�wH;qUH;�(H;��G;Z�G;��F;eiE;��A;֡:;Z|,;�;~��:�i:�����D^�:�ܻKE:� ����Ҽ4����G�B���榽�Pν�������Q"���0�ڀ:�      4Dx�8�s���f�wS�ڀ:����\[��7ս�榽��}���;��8�X�����r����6G�����ʬ�_��:9�;�}$;�6;9�?;�D;�F;�pG;��G;"H;cJH;noH;y�H;��H;7�H;v�H;��H;��H;d�H;��H;��H;v�H;5�H;��H;y�H;noH;bJH;"H;��G;�pG;�F;�D;9�?;�6;�}$;8�;_��:�ʬ����6G�������r�X����8���;���}��榽�7ս\[����ڀ:�wS���f�8�s�      �*���0��॒�=����k��H��#%�\[��Pν
t��d�f�6/%���伈���v�=��?ػzFL�h�D�΍R:N�:J�;W2;��=;ݚC;�0F;�GG;��G;ZH;"@H;�gH;��H;n�H;�H;ѸH;��H;+�H;��H;+�H;��H;иH;�H;n�H;��H;�gH; @H;[H;��G;�GG;�0F;ښC;��=;W2;M�;L�:΍R:`�D�|FL��?ػv�=��������6/%�d�f�
t���Pν\[��#%��H��k�=���॒��0��      *�þ���"����R��~쏾8�s��H�����������ѐ����D��c�����@�f�S,�����P���9$��:�;Dj-;��;;��B;�E;�G;��G;��G;�6H;�`H;��H;��H;�H;��H;�H;��H;�H;��H;�H;��H;�H;��H;��H;�`H;�6H;��G;��G;�G;�E;��B;��;;Dj-;�;&��:�9�P�����S,�@�f������c���D�ѐ�������������H�8�s�~쏾�R��"������      B��2�很Yؾ*�þĪ�~쏾�k�ڀ:���~�ؽ�����c�`y���Ҽ ���C� �b��� 8(7��:��
;�(;�_9;ΘA;�\E;��F;ޝG;��G;�.H;�ZH;&|H;.�H;��H;��H;M�H;�H;��H;�H;L�H;��H;��H;/�H;&|H;�ZH;�.H;��G;��G;��F;�\E;˘A;�_9;�(;��
;��: 8(7��c�D� � �����Ҽ`y��c�����~�ؽ��ڀ:��k�~쏾Ī�*�þ�Yؾ2��      %��P������AI�*�þ�R��=���wS��Q"��s������}��0��켋�����6�B�ƻ,}*�`���1�:�x;v%;m7;�@;�D;�F;��G;��G;<(H;VH;�xH;��H;~�H;ܲH;�H;��H;��H;��H;�H;ڲH;}�H;��H;�xH;VH;;(H;��G;��G;�F;�D;�@;m7;v%;�x;/�:`���,}*�C�ƻ��6��������0���}�����s��Q"�wS�=����R��*�þAIᾦ���P��      ���T��:�
������Yؾ"���॒���f���0�][�R8��Ґ����>�����MȤ��6H�]�ܻ�qF�p����}:��:~";m�5;�?;��D;�F;$�G;��G;{#H;�RH;�uH;��H;��H;��H;�H;)�H;��H;)�H;�H;��H;��H;��H;�uH;�RH;x#H;��G;$�G;�F;��D;�?;p�5;~";��:��}:p���qF�^�ܻ�6H�MȤ�������>�Ґ��R8��][���0���f�॒�"����Yؾ����:�
�T��      �� ����T��P��2������0��8�s�ڀ:�i9� �ʽ4Z���G��8�.���5S�����/X�,�D�$Cd:�B�:! ;4�4;ڈ?;D;_�F;(yG;��G;� H;TPH;StH;K�H;�H;�H;m�H;��H;o�H;��H;n�H;�H;�H;N�H;StH;QPH;� H;��G;'yG;]�F;D;׈?;:�4;! ;�B�: Cd:,�D��/X���껰5S�.���8��G�4Z�� �ʽi9�ڀ:�8�s��0�����2��P��T�����      IF�Yh����YVھ:�������~���S��#��o��<S��r₽6�6�u���my��YFB��Eֻ�A?���	��Y�:���:~�";�46;k@;��D;۩F;�nG; �G;CH;>@H;!gH;��H;f�H;ƩH;�H;�H;��H;�H;�H;ƩH;d�H;��H;!gH;<@H;@H; �G;�nG;۩F;��D;g@;�46;~�";���:�Y�:��	��A?��EֻYFB�my��u���6�6�r₽<S���o���#��S��~������:��YVھ��Yh��      Yh���b���쾪*־�v��*���*��*�O�X� �s��r���؀�K�3���Cݜ�?�>�Q�ѻۡ9�P���po�:E% ;�M#;�6;\A@;"�D;կF;/qG;|�G;YH;	AH;�gH;�H;ŚH;�H;Q�H;.�H;�H;.�H;Q�H;�H;ĚH;��H;�gH;AH;VH;|�G;/qG;կF;"�D;VA@;��6;�M#;F% ;lo�:P���ڡ9�R�ѻ?�>�Cݜ���J�3��؀��r��s�X� �*�O�*��*����v���*־���b��      ���쾶�޾25ʾO;���:��,�v��E�b'����u����u���+��W��A����4���Ļ9)��i���W�:j�; %;"l7;5�@;$�D;�F;	xG;��G;{H;jCH;ciH;R�H;ɛH;ܪH;��H;˺H;��H;˺H;��H;ܪH;țH;R�H;ciH;eCH;xH;��G;xG;�F;$�D;1�@;%l7; %;i�;�W�:�i��9)���Ļ��4��A���W缇�+���u�u�����b'��E�,�v��:��O;��25ʾ��޾��      YVھ�*־25ʾu��������M���9b��5�����ս����Xc�	��Жռ�I��W�$�jT���Z�`Z��`�:
�;��';X�8;0RA;�9E;��F;��G;!�G;�H;3GH;JlH;��H;q�H;�H;�H;˻H;��H;˻H;�H;�H;p�H;��H;JlH;2GH;�H;!�G;��G;��F;�9E;+RA;\�8;��';�;\�:`Z���Z�jT��X�$��I��Жռ	���Xc������ս���5��9b��M������u���25ʾ�*־      :���v��O;������UP��H�r�}�H�X� ���8@��ԓ����K�d� ־���s�t���񕻒ܺ06u9c&�:0�;J�+;��:;�"B;��E;�F;��G;�G;tH;bLH;5pH;�H;��H;ۭH;t�H;�H;��H;�H;r�H;ܭH;��H;�H;4pH;^LH;sH;�G;��G;�F;��E;�"B;��:;J�+;1�;]&�: 6u9�ܺ��t����s� ־�d���K�ԓ��8@����X� �}�H�H�r�UP������O;���v��      ����+����:���M��H�r�*�O�#,�Z�
��gٽsĥ���u�|1�o���.Ϥ���P�[�.o�Zp���:���:Q;[�/;s�<;!C;P�E;�!G;Y�G;7�G;�%H;�RH;uH;7�H;~�H;�H;@�H;��H;>�H;��H;@�H;�H;|�H;:�H;uH;�RH;�%H;7�G;W�G;�!G;O�E;C;s�<;[�/;Q;���:�:Vp���.o�[򻮎P�.Ϥ�o���|1���u�tĥ��gٽZ�
�#,�*�O�H�r��M���:��*���      �~��*��,�v��9b�}�H�#,�OZ����:S��z^����N������μ�I���%+����̝.� ���
k~:���:Cm;��3;R�>;[�C;vPF;�FG;x�G;#�G;�/H;0ZH;�zH;��H;��H;��H;]�H;b�H;�H;a�H;]�H;��H;��H;��H;�zH;/ZH;�/H;#�G;v�G;�FG;tPF;U�C;R�>;��3;Dm;���:
k~:���Ν.�����%+��I����μ�����N�z^��:S�����OZ�#,�}�H��9b�,�v�*��      �S�*�O��E��5�X� �Z�
���罨9��*l���Xc���(��������[�����ݎ�#ܺP<9V��:[�	;]d';� 8;u�@;��D;�F;YjG;��G;�H;�:H;qbH;�H;F�H;i�H;~�H;��H;q�H;�H;q�H;��H;~�H;h�H;F�H;�H;pbH;�:H;�H;��G;YjG;�F;��D;u�@;� 8;_d';Y�	;V��:`<9&ܺ�ݎ������[��������(��Xc�*l���9�����Z�
�X� ��5��E�*�O�      �#�X� �b'������gٽ:S��*l��T�j�G�3��i��վ�}���
(���ĻYA?�L�B�N�@:�[�:6Q;"�.;�;;�tB;A�E;��F;i�G;*�G;H;�FH;WkH;H;_�H;G�H;��H;J�H;��H;2�H;��H;I�H;��H;G�H;_�H;H;VkH;�FH;H;'�G;i�G;��F;>�E;�tB;�;;$�.;5Q;�[�:V�@:L�B�XA?���Ļ
(�}����վ��i�F�3�S�j�*l��:S���gٽ����b'�X� �      �o��s��置�ս9@��tĥ�{^���Xc�G�3���	�Ό˼�]��UFB��Z򻬜��QӺ ��8��:��;�M#;�=5;>?;��C;�@F;A:G;,�G;Q�G;k'H;�RH;�tH;�H;��H;c�H;�H;��H;
�H;~�H;
�H;��H;�H;b�H;��H;�H;�tH;�RH;k'H;P�G;+�G;>:G;�@F;��C;>?;�=5;�M#;��;��:���8QӺ�����Z�UFB��]��Ό˼��	�G�3��Xc�{^��tĥ�9@����ս���s�      <S���r��v�����ԓ����u���N���(��i�Ό˼�A����P�hs��2|�����\:`�:��;�n-;	�:;�A;�,E;��F;goG;.�G;�H;8H;}_H;@~H;)�H;>�H;��H;L�H;��H;w�H;��H;v�H;��H;K�H;��H;A�H;)�H;=~H;{_H;8H;�H;.�G;doG;��F;�,E;�A;�:;�n-;��;d�:\:����1|��hs���P��A��͌˼�i���(���N���u�ԓ�����v���r��      r₽�؀���u��Xc���K�|1�������վ��]����P����>T����9���o�H4�9�&�:w�	;~%;z�5;��>;ջC;�F;�!G;ۚG;�G;{H;�HH;lH;هH;��H;έH;�H;��H;��H;��H;�H;��H;��H;��H;�H;ѭH;��H;هH;lH;�HH;yH;�G;՚G;�!G;�F;ԻC;��>;w�5;~%;z�	;�&�:H4�9��o���9�>T�������P��]���վ�����|1���K��Xc���u��؀�      6�6�J�3���+�	��d�o�����μ���}���UFB�hs�?T���D��{���;u9�q�:���:�Y;u0;�;;B;":E;�F;5hG;�G;D�G;�0H;�XH;ixH;[�H;��H;>�H;5�H;�H;P�H;g�H;u�H;g�H;O�H;�H;5�H;@�H;��H;[�H;gxH;�XH;�0H;F�G;�G;0hG;�F;":E;B;�;;u0;�Y;���:�q�:�;u9�{���D�?T��hs�UFB�}��������μo���e�	����+�K�3�      u�����W�Жռ�վ�.Ϥ��I����[�	(��Z����9��{���<9~X�:�X�:^Q;],;��8;�A@;7BD;�@F;�,G;��G;��G;�H;EH;]hH;p�H;��H;��H;��H;_�H;\�H;�H;��H;��H;��H;�H;Z�H;_�H;��H;��H;��H;n�H;ZhH;	EH;�H;��G;��G;�,G;�@F;7BD;�A@;��8;`,;^Q;�X�:�X�:�<9�{����9���Z�(���[��I��-Ϥ� ־�Жռ�W���      my��Dݜ��A���I����s���P��%+������Ļ����2|���o��;u9~X�: ,�:u;);�6;��>;�PC;��E;)�F;�xG;e�G;�H;�1H;SXH;>wH;�H;R�H;@�H;��H;U�H;~�H;��H;#�H;��H;#�H;��H;}�H;T�H;��H;@�H;P�H;�H;=wH;QXH;�1H;�H;a�G;�xG;)�F;��E;�PC;��>;��6;);t; ,�:~X�:�;u9��o�2|�������Ļ����%+���P���s��I���A��Eݜ�      YFB�@�>���4�X�$�u��[�����ݎ�ZA?�SӺ����@4�9�q�:�X�:t;��';�=5;��=;0�B;PGE;|�F;�UG;Z�G;�G;�H;�HH;OjH;5�H;��H;��H;p�H;��H;�H;}�H;I�H;Z�H;�H;Z�H;I�H;{�H;�H;��H;p�H;��H;��H;5�H;KjH; IH;�H;�G;V�G;�UG;x�F;PGE;0�B;��=;�=5;��';w;�X�:�q�:H4�9����PӺXA?��ݎ����[�u��X�$���4�A�>�      �EֻM�ѻ��ĻlT���񕻱.o�ɝ.�$ܺP�B� ��8\:�&�:���:\Q;);�=5;;=;L#B;��D;vF;#7G;��G;��G;�H;�:H;O^H;�zH;7�H;��H;�H;G�H;�H;��H;X�H;��H;g�H;��H;e�H;��H;X�H;��H;�H;G�H;��H;��H;6�H;�zH;Q^H;�:H;�H;��G;��G; 7G;vF;��D;O#B;;=;�=5;);^Q;���:�&�:\: ��8H�B�&ܺȝ.��.o���lT����ĻS�ѻ      �A?�ܡ9�9)��Z��ܺvp��(��� <9F�@:��:d�:x�	;�Y;\,;�6;��=;J#B;�D;�XF;"G;��G;V�G;�H;0/H;�SH;�qH;�H;��H;��H;��H;��H;�H;��H;	�H;��H;W�H;��H;U�H;��H;	�H;��H;�H;��H;��H;��H;��H;�H;�qH;�SH;,/H;�H;V�G;��G;"G;�XF;�D;J#B;��=;�6;],;�Y;x�	;d�:��:V�@: <9(���lp���ܺ�Z�9)��9�      ��	�p����i���Z���5u9�:k~:T��:�[�:��;��;%;u0;��8;��>;.�B;��D;�XF;iG;��G;��G;��G;/&H;BKH;�iH;"�H;ȗH;u�H;��H;E�H;��H;��H;��H;n�H;��H;�H;��H;�H;��H;m�H;��H;��H;��H;B�H;��H;u�H;ŗH;#�H;�iH;@KH;+&H;��G;��G;��G;kG;�XF;��D;0�B;��>;��8;u0;%;��;��;�[�:P��:k~:�:@6u9�Z���i��h���      �Y�:�o�:�W�:\�:Y&�:���:���:W�	;2Q;�M#;�n-;v�5;�;;�A@;�PC;JGE;vF;"G;��G;
�G;P�G;� H;JEH;�cH;z}H;��H;��H;ޱH;�H;��H;��H;f�H;��H;��H;��H;��H;*�H;��H;��H;��H;��H;g�H;��H;��H;��H;ܱH;�H;��H;z}H;�cH;FEH;� H;N�G;�G;��G;"G;vF;JGE;�PC;�A@;�;;w�5;�n-;�M#;4Q;X�	;���:���:o&�:\�:�W�:~o�:      ���:Q% ;p�;�;*�;Q;Fm;\d';!�.;�=5;�:;��>;B;6BD;��E;{�F;!7G;��G;��G;Q�G;�H;%BH;F`H;�yH;��H;`�H;��H;�H;��H;�H;��H;j�H;��H;|�H;.�H;�H;��H;�H;.�H;|�H;��H;l�H;��H;�H;��H;�H;��H;a�H;��H;�yH;E`H;%BH;�H;S�G;��G;��G;!7G;z�F;��E;6BD;B;��>;�:;�=5;$�.;\d';Fm;Q;-�;�;m�;A% ;      ��";�M#;/%;{�';L�+;c�/;��3;� 8;�;;B?;#�A;ջC;$:E;�@F;*�F;�UG;��G;X�G;��G;� H;$BH;�^H;�wH;X�H;ÝH;�H;̷H;j�H;<�H;d�H;]�H;&�H;��H;�H;��H;��H;��H;��H;��H;�H;��H;&�H;]�H;`�H;8�H;j�H;ɷH;�H;ĝH;V�H;�wH;�^H;"BH;� H;��G;Y�G;��G;�UG;,�F;�@F;$:E;ջC;"�A;B?;�;;� 8;��3;c�/;b�+;{�';-%;�M#;      �46;��6;#l7;Q�8;��:;q�<;V�>;v�@;�tB;��C;�,E;�F;�F;�,G;�xG;X�G;��G;�H;/&H;LEH;F`H;�wH;n�H;r�H;��H;'�H;׿H;��H;�H;9�H;g�H;{�H;��H;��H;��H;��H;��H;��H;��H;��H;��H;{�H;h�H;7�H;�H;��H;ԿH;(�H;��H;p�H;m�H;�wH;B`H;MEH;0&H;�H;��G;W�G;�xG;�,G;�F;�F;�,E;��C;�tB;u�@;V�>;t�<;��:;Q�8;%l7;s�6;      @;gA@;>�@;,RA;�"B;C;_�C;��D;?�E;�@F;��F;�!G;.hG;��G;b�G;�G;�H;0/H;AKH;�cH;�yH;W�H;p�H;�H;C�H;��H;��H;�H;M�H;��H;��H;��H;x�H;��H;�H;��H;��H;��H;�H;��H;u�H;��H;��H;��H;K�H;�H;��H;��H;D�H;��H;p�H;W�H;�yH;�cH;AKH;3/H;�H;�G;b�G;��G;0hG;�!G;��F;�@F;A�E;��D;^�C;C;�"B;.RA;>�@;]A@;      ��D;&�D;�D;�9E;��E;Q�E;rPF;�F;��F;>:G;aoG;ښG;�G;��G;�H;�H;�:H;�SH;�iH;�}H;ÎH;ǝH;��H;L�H;w�H; �H;k�H;��H;��H;j�H;�H;D�H;��H;'�H;��H;\�H;��H;\�H;��H;$�H;��H;F�H;�H;j�H;��H;��H;k�H; �H;w�H;I�H;��H;ɝH;��H;�}H;�iH;�SH;�:H;�H;�H;��G;�G;ۚG;doG;=:G;��F;�F;tPF;Q�E;��E;�9E;�D;&�D;      �F;�F;�F;��F;�F;�!G;�FG;VjG;f�G;+�G;+�G;�G;C�G;�H;�1H;�HH;N^H;�qH;�H;��H;]�H;�H;$�H;��H;�H;L�H;Z�H;��H;��H;��H;��H;��H;+�H;�H;��H;�H;G�H;�H;��H;�H;(�H;��H;��H;��H;��H;��H;[�H;L�H;�H;��H;$�H;�H;Z�H;��H;�H;�qH;M^H;�HH;�1H;�H;D�G;�G;-�G;)�G;g�G;VjG;�FG;�!G;#�F;��F;�F;دF;      �nG;2qG;xG;�G;��G;]�G;|�G;��G;)�G;O�G;�H;}H;�0H;	EH;QXH;OjH;�zH;�H;ȗH;��H;��H;̷H;ֿH;��H;e�H;_�H;}�H;��H;��H;��H;��H;�H;�H;��H;q�H;��H;��H;��H;o�H;��H;�H;�H;��H;��H;��H;��H;{�H;^�H;g�H;��H;ԿH;ͷH;��H;��H;ȗH;�H;�zH;NjH;QXH;	EH;�0H;}H;�H;O�G;,�G;��G;|�G;\�G;��G;�G;	xG;0qG;      �G;�G;��G; �G;�G;7�G;(�G;�H;H;q'H;
8H;�HH;�XH;]hH;>wH;5�H;6�H;�H;r�H;�H;�H;j�H;��H;�H;��H;��H;��H;x�H;��H;��H;��H;�H;��H;��H;�H;?�H;P�H;?�H;�H;��H;��H;�H;��H;�H;��H;x�H;��H;��H;��H;�H;��H;j�H;�H;�H;u�H;�H;5�H;5�H;@wH;[hH;�XH;�HH;
8H;q'H;H;�H;(�G;7�G;)�G;�G;��G;��G;      [H;VH;{H;�H;tH;�%H;�/H;�:H;�FH;�RH;{_H;lH;hxH;o�H;�H;��H;��H;��H;��H;�H;��H;;�H;�H;R�H;��H; �H;��H;��H;^�H;��H;�H;��H;��H;�H;��H;��H;��H;��H;��H;�H;��H;��H;�H;��H;^�H;��H;��H;��H;��H;R�H;�H;;�H;��H;�H;��H;��H;��H;��H;�H;o�H;ixH;lH;y_H;�RH;�FH;�:H;�/H;�%H;zH;�H;zH;MH;      I@H;AH;rCH;9GH;sLH;�RH;6ZH;ubH;]kH;�tH;F~H;�H;a�H;��H;U�H;��H;�H;��H;A�H;��H;�H;a�H;6�H;��H;b�H;��H;��H;�H;��H;�H;��H;��H;7�H;��H;��H;�H;�H;�H;��H;��H;3�H;��H;��H;�H;��H;�H;��H;��H;c�H;��H;4�H;a�H;�H;��H;C�H;��H;�H;��H;U�H;��H;a�H;�H;G~H;�tH;`kH;wbH;6ZH;�RH;oLH;9GH;mCH;AH;      #gH;�gH;piH;VlH;ApH;uH;�zH;��H;ƇH;�H;.�H;��H;��H;��H;C�H;v�H;M�H;��H;��H;��H;��H;]�H;h�H;��H;�H;��H;��H;��H;�H;��H;��H;B�H;��H;��H;�H;I�H;c�H;I�H;�H;��H;��H;C�H;��H;��H;�H;��H;��H;��H;�H;��H;e�H;]�H;��H;��H;��H;��H;K�H;v�H;C�H;��H;��H;��H;/�H;�H;ȇH;��H;�zH;uH;>pH;WlH;piH;�gH;      ��H; �H;]�H;��H;��H;:�H;��H;M�H;b�H;��H;C�H;׭H;B�H;��H;��H;��H;�H;�H;��H;p�H;s�H;*�H;~�H;��H;A�H;��H;�H;�H;��H;��H;?�H;��H;��H;;�H;c�H;��H;�H;��H;c�H;;�H;��H;��H;?�H;��H;��H;�H;�H;��H;D�H;��H;{�H;*�H;p�H;p�H;��H;!�H;�H;��H;��H;��H;B�H;׭H;E�H;��H;c�H;J�H;��H;=�H;��H;��H;_�H;��H;      k�H;њH;ӛH;w�H;��H;~�H;��H;s�H;M�H;c�H;��H;�H;7�H;c�H;X�H;�H;��H;��H;��H;��H;��H;��H;��H;�H;��H;.�H;"�H;��H;��H;>�H;��H;��H;=�H;v�H;��H;��H;��H;��H;��H;v�H;;�H;��H;��H;?�H;��H;��H;�H;-�H;��H;�H;��H;��H;��H;��H;��H;��H;��H;�H;U�H;c�H;6�H;�H;��H;e�H;M�H;q�H;��H;��H;��H;w�H;ӛH;ʚH;      שH;'�H;֪H;%�H;�H;�H;��H;��H;��H;�H;R�H;��H; �H;_�H;��H;��H;_�H;	�H;q�H;��H;��H;�H;��H;��H;�H;�H;��H;��H;�H;��H;��H;;�H;o�H;��H;��H;��H;��H;��H;��H;��H;m�H;=�H;��H;��H;�H;��H;��H;�H;!�H;��H;��H;�H;��H;��H;q�H;�H;]�H;��H;��H;_�H; �H;��H;P�H;�H;��H;��H;��H;�H;ܭH;%�H;تH;�H;      �H;g�H; �H;�H;��H;?�H;e�H;ʽH;Q�H;��H;��H;��H;U�H; �H;��H;R�H;��H;��H;��H;��H;8�H;��H;��H;�H;��H;��H;m�H;�H;��H;��H;�H;f�H;��H;��H;��H;��H;��H;��H;��H;��H;��H;i�H;�H;��H;��H;�H;k�H;��H;��H;	�H;��H;��H;5�H;��H;��H;��H;��H;R�H;��H; �H;U�H;��H;��H;��H;Q�H;ǽH;e�H;C�H;��H;	�H;�H;^�H;      �H;6�H;ӺH;ͻH; �H;��H;l�H;{�H;��H;	�H;}�H;��H;j�H;��H;(�H;a�H;n�H;Q�H;�H;��H;'�H;��H;��H;��H;X�H;�H;��H;?�H;��H;�H;G�H;��H;��H;��H;��H;��H;��H;��H;��H;��H;��H;��H;G�H;�H;��H;?�H;��H;�H;Y�H;��H;��H;��H;%�H;��H;�H;S�H;m�H;a�H;(�H;��H;j�H;��H;{�H;�H;��H;x�H;k�H;��H;�H;ͻH;ֺH;.�H;      ��H;�H;��H;��H;̾H;?�H;�H;�H;:�H;}�H;��H;$�H;v�H;��H;��H;�H;��H;��H;��H;1�H;��H;��H;��H;��H;��H;B�H;��H;V�H;��H;�H;f�H;��H;��H;��H;��H;��H;��H;��H;��H;��H;��H;��H;f�H;�H;��H;V�H;��H;D�H;��H;��H;��H;��H;��H;1�H;��H;��H;��H;�H;��H;��H;v�H;$�H;��H;��H;:�H;�H;�H;C�H;��H;��H;��H;�H;      �H;7�H;ӺH;ͻH;!�H;��H;l�H;{�H;��H;
�H;}�H;��H;j�H;��H;(�H;a�H;n�H;Q�H;�H;��H;(�H;��H;��H;��H;Y�H;�H;��H;?�H;��H;�H;G�H;��H;��H;��H;��H;��H;��H;��H;��H;��H;��H;��H;G�H;�H;��H;?�H;��H;�H;X�H;��H;��H;��H;%�H;��H;�H;S�H;m�H;a�H;(�H;��H;j�H;��H;}�H;
�H;��H;x�H;l�H;��H;�H;ͻH;ҺH;+�H;      �H;g�H;��H;	�H;��H;?�H;e�H;ʽH;Q�H;��H;��H;��H;V�H; �H;��H;R�H;��H;��H;��H;��H;9�H;��H;��H;�H;��H;��H;m�H;�H;��H;��H;�H;f�H;��H;��H;��H;��H;��H;��H;��H;��H;��H;j�H;�H;��H;��H;�H;k�H;��H;��H;�H;��H;��H;5�H;��H;��H;��H;��H;R�H;��H; �H;U�H;��H;��H;��H;Q�H;ǽH;e�H;C�H;��H;	�H; �H;^�H;      ةH;'�H;تH;%�H;�H;�H;��H;��H;��H;�H;R�H;��H; �H;_�H;��H;��H;_�H;�H;q�H;��H;��H;�H;��H;��H;!�H;�H;��H;��H;�H;��H;��H;;�H;o�H;��H;��H;��H;��H;��H;��H;��H;m�H;=�H;��H;��H;�H;��H;��H;�H;�H;��H;��H;�H;��H;��H;q�H;�H;]�H;��H;��H;_�H; �H;��H;R�H;�H;��H;��H;��H;�H;ۭH;%�H;تH;�H;      n�H;њH;ӛH;x�H;��H;~�H;��H;q�H;M�H;c�H;��H;�H;6�H;c�H;U�H;�H;��H;��H;��H;��H;��H;��H;��H;�H;��H;.�H;!�H;��H;��H;>�H;��H;��H;<�H;t�H;��H;��H;��H;��H;��H;t�H;;�H;��H;��H;?�H;��H;��H; �H;-�H;��H;~�H;��H;��H;��H;��H;��H;��H;��H;�H;V�H;c�H;6�H;�H;��H;e�H;M�H;o�H;��H;��H;��H;x�H;қH;̚H;      ��H;�H;_�H;��H;��H;:�H;��H;M�H;b�H;��H;C�H;׭H;B�H;��H;��H;��H;�H;�H;��H;q�H;v�H;*�H;~�H;��H;D�H;��H;�H;�H;��H;��H;?�H;��H;��H;;�H;c�H;��H;�H;��H;c�H;;�H;��H;��H;?�H;��H;��H;�H;�H;��H;A�H;��H;|�H;*�H;q�H;p�H;��H;�H;�H;��H;��H;��H;B�H;׭H;C�H;��H;c�H;J�H;��H;;�H;��H;��H;`�H;��H;      #gH;�gH;piH;WlH;ApH;uH;�zH;��H;ȇH;�H;/�H;��H;��H;��H;C�H;w�H;K�H;��H;��H;��H;��H;]�H;h�H;��H;�H;��H;��H;��H;�H;��H;��H;B�H;��H;��H;�H;I�H;c�H;I�H;�H;��H;��H;C�H;��H;��H;�H;��H;��H;��H;�H;��H;e�H;]�H;��H;��H;��H;��H;K�H;v�H;C�H;��H;��H;��H;,�H;�H;ȇH;��H;�zH;uH;>pH;VlH;piH;�gH;      C@H;AH;qCH;9GH;oLH;�RH;9ZH;xbH;^kH;�tH;F~H;�H;_�H;��H;U�H;��H;�H;��H;B�H;��H;�H;a�H;6�H;��H;c�H;��H;��H;�H;��H;�H;��H;��H;5�H;��H;��H;�H;�H;�H;��H;��H;5�H;��H;��H;�H;��H;�H;��H;��H;b�H;��H;4�H;a�H;�H;��H;A�H;��H;�H;��H;U�H;��H;a�H;�H;F~H;�tH;akH;xbH;9ZH;�RH;nLH;:GH;oCH;AH;      TH;RH;�H;�H;xH;�%H;�/H;�:H;�FH;�RH;{_H;lH;hxH;o�H;�H;��H;��H;��H;��H;�H;��H;;�H;�H;Q�H;��H; �H;��H;��H;^�H;��H;�H;��H;��H;�H;��H;��H;��H;��H;��H;�H;��H;��H;�H;��H;^�H;��H;��H;��H;��H;R�H;�H;;�H;��H;�H;��H;��H;��H;��H;�H;o�H;hxH;lH;{_H;�RH;�FH;�:H;�/H;�%H;vH;�H;�H;TH;      �G;�G;��G;�G;�G;7�G;(�G;�H;H;q'H;8H;�HH;�XH;]hH;@wH;5�H;6�H;�H;u�H;�H;$�H;j�H;��H;�H;��H;��H;��H;x�H;��H;��H;��H;�H;��H;��H;�H;A�H;P�H;?�H;�H;��H;��H;�H;��H;�H;��H;x�H;��H;��H;��H;�H;��H;j�H;�H;�H;r�H;�H;5�H;6�H;>wH;ZhH;�XH;�HH;8H;q'H;H;�H;(�G;4�G;)�G; �G;��G;��G;      �nG;3qG;	xG;݂G;��G;Y�G;{�G;��G;)�G;P�G;�H;}H;�0H;	EH;QXH;OjH;�zH;�H;ȗH;��H;��H;ͷH;ֿH;��H;g�H;_�H;~�H;��H;��H;��H;��H;�H;�H;��H;o�H;��H;��H;��H;q�H;��H;�H;�H;��H;��H;��H;��H;{�H;_�H;e�H;��H;ԿH;̷H;��H;��H;ȗH;�H;�zH;NjH;QXH;	EH;�0H;}H;�H;P�G;)�G;��G;{�G;W�G;��G;݂G;	xG;)qG;      �F;ޯF;�F;��F;�F;�!G;�FG;YjG;e�G;+�G;-�G;�G;D�G;�H;�1H;�HH;N^H;�qH;�H;��H;`�H;�H;$�H;��H;�H;L�H;\�H;��H;��H;��H;��H;��H;*�H;�H;��H;�H;G�H;�H;��H;�H;(�H;��H;��H;��H;��H;��H;Z�H;L�H;�H;��H;$�H;�H;X�H;��H;�H;�qH;M^H;�HH;�1H;�H;C�G;�G;-�G;)�G;f�G;VjG;�FG;�!G;!�F;��F;�F;ԯF;      ��D;&�D;�D;�9E;��E;Q�E;tPF;�F;��F;>:G;foG;ۚG;�G;��G;�H;�H;�:H;�SH;�iH;�}H;ĎH;ɝH;��H;L�H;w�H;�H;l�H;��H;��H;l�H;�H;D�H;��H;$�H;��H;\�H;��H;\�H;��H;&�H;��H;G�H;�H;i�H;��H;��H;k�H; �H;w�H;J�H;��H;ǝH;��H;�}H;�iH;�SH;�:H;�H;�H;��G;�G;ښG;aoG;=:G;��F;�F;rPF;Q�E;��E;�9E;�D;&�D;      �@;dA@;C�@;+RA;�"B;C;\�C;��D;A�E;�@F;��F;�!G;1hG;��G;b�G;�G;�H;0/H;AKH;�cH;�yH;W�H;r�H;�H;D�H;��H;��H;�H;N�H;��H;��H;��H;w�H;��H;�H;��H;��H;��H;�H;��H;w�H;��H;��H;��H;J�H;�H;��H;��H;C�H;��H;o�H;W�H;�yH;�cH;AKH;2/H;�H;�G;b�G;��G;.hG;�!G;��F;�@F;A�E;��D;\�C;!C;�"B;+RA;A�@;[A@;      �46;��6;4l7;Q�8;��:;w�<;Z�>;v�@;�tB;��C;�,E;�F;�F;�,G;�xG;X�G;��G;�H;0&H;LEH;H`H;�wH;n�H;s�H;��H;'�H;׿H;��H;�H;:�H;h�H;{�H;��H;��H;��H;��H;��H;��H;��H;��H;��H;{�H;g�H;6�H;�H;��H;ԿH;(�H;��H;p�H;n�H;�wH;C`H;MEH;/&H;�H;��G;X�G;�xG;�,G;�F;�F;�,E;�C;�tB;u�@;[�>;w�<;��:;P�8;)l7;�6;      ��";�M#;1%;{�';N�+;c�/;��3;� 8;�;;B?;#�A;ջC;$:E;�@F;*�F;�UG;��G;V�G;��G;� H;%BH;�^H;�wH;Z�H;ĝH;�H;̷H;j�H;<�H;d�H;]�H;&�H;��H;�H;��H;��H;��H;��H;��H;�H;��H;&�H;]�H;`�H;8�H;j�H;ɷH;�H;ÝH;V�H;�wH;�^H;$BH;� H;��G;Y�G;��G;�UG;,�F;�@F;$:E;׻C;"�A;B?;�;;� 8;��3;c�/;b�+;{�';.%;�M#;      ���:L% ;t�;�;*�;Q;Jm;_d';!�.;�=5;�:;��>;B;6BD;��E;z�F;#7G;��G;��G;Q�G;�H;%BH;F`H;�yH;��H;a�H;��H;�H;��H;�H;��H;j�H;��H;{�H;.�H;�H;��H;�H;.�H;|�H;��H;m�H;��H;�H;��H;�H;��H;`�H;��H;�yH;E`H;%BH;�H;Q�G;��G;��G;7G;z�F;��E;6BD;B;��>;�:;�=5;"�.;]d';Hm;Q;1�;�;r�;A% ;      �Y�:�o�:�W�:X�:c&�:���:���:Y�	;4Q;�M#;�n-;w�5;�;;�A@;�PC;JGE;vF;"G;��G;
�G;Q�G;� H;JEH;�cH;z}H;��H;��H;ܱH;�H;��H;��H;f�H;��H;��H;��H;��H;*�H;��H;��H;��H;��H;g�H;��H;��H;��H;ޱH;�H;��H;z}H;�cH;GEH;� H;M�G;�G;��G;"G;vF;JGE;�PC;�A@;�;;u�5;�n-;�M#;4Q;X�	;���:���:o&�:X�:�W�:~o�:      ��	�p����i���Z���5u9�:k~:T��:�[�:��;��;%;u0;��8;��>;0�B;��D;�XF;kG;��G;��G;��G;/&H;BKH;�iH;!�H;ȗH;u�H;��H;E�H;��H;��H;��H;m�H;��H;�H;��H;�H;��H;n�H;��H;��H;��H;B�H;��H;u�H;ƗH;#�H;�iH;@KH;+&H;��G;��G;��G;iG;�XF;��D;.�B;��>;��8;u0;%;��;��;�[�:T��:k~:�:@6u9�Z���i��h���      �A?�ܡ9�9)��Z��ܺvp��(��� <9J�@:��:d�:x�	;�Y;Z,;�6;��=;L#B;�D;�XF;"G;��G;V�G;�H;0/H;�SH;�qH;�H;��H;��H;��H;��H;�H;��H;	�H;��H;U�H;��H;U�H;��H;	�H;��H;�H;��H;��H;��H;��H;�H;�qH;�SH;,/H;�H;V�G;��G;"G;�XF;�D;I#B;��=;�6;Z,;�Y;x�	;d�:��:V�@: <9(���lp���ܺ�Z�9)��9�      �EֻN�ѻ��ĻlT���񕻳.o�ȝ.�#ܺP�B� ��8\:�&�:���:^Q;);�=5;;=;L#B;��D;vF;!7G;��G;��G;�H;�:H;O^H;�zH;6�H;��H;�H;G�H;�H;��H;X�H;��H;g�H;��H;g�H;��H;Y�H;��H;�H;G�H;�H;��H;7�H;�zH;Q^H;�:H;�H;��G;��G;!7G;vF;��D;O#B;;=;�=5;);\Q;���:�&�:\:���8L�B�'ܺɝ.��.o���lT����ĻS�ѻ      ZFB�?�>���4�X�$�u��[�����ݎ�YA?�OӺ����P4�9�q�:�X�:w;��';�=5;��=;0�B;PGE;z�F;�UG;X�G;�G;�H;�HH;NjH;5�H;��H;��H;p�H;��H;�H;{�H;I�H;Z�H;�H;Z�H;I�H;}�H;�H;��H;p�H;��H;��H;5�H;MjH; IH;�H;�G;W�G;�UG;z�F;PGE;0�B;��=;�=5;��';u;�X�:�q�:@4�9����TӺYA?��ݎ����[�u��X�$���4�A�>�      my��Dݜ��A���I����s���P��%+������Ļ����2|���o��;u9~X�:",�:t;);�6;��>;�PC;��E;)�F;�xG;e�G;�H;�1H;SXH;=wH;�H;R�H;@�H;��H;U�H;}�H;��H;#�H;��H;#�H;��H;��H;U�H;��H;@�H;P�H;�H;>wH;QXH;�1H;�H;a�G;�xG;)�F;��E;�PC;��>;��6;);u;",�:~X�:�;u9��o�2|�������Ļ����%+���P���s��I���A��Eݜ�      u�����W�Жռ�վ�.Ϥ��I����[�	(��Z����9��{���<9�X�:�X�:_Q;^,;��8;�A@;6BD;�@F;�,G;��G;��G;�H;EH;ZhH;o�H;��H;��H;��H;`�H;[�H;�H;��H;��H;��H;�H;[�H;]�H;��H;��H;��H;o�H;]hH;EH;�H;��G;��G;�,G;�@F;9BD;�A@;��8;`,;\Q;�X�:~X�:�<9�{����9���Z�	(���[��I��-Ϥ� ־�Жռ�W���      6�6�J�3���+�	��d�o�����μ���}���UFB�hs�?T���D��{���;u9�q�:���:�Y;u0;�;;B;":E;�F;4hG;�G;D�G;�0H;�XH;hxH;[�H;��H;>�H;5�H;�H;O�H;g�H;u�H;g�H;P�H;�H;3�H;@�H;��H;[�H;gxH;�XH;�0H;G�G;�G;0hG;�F;":E;B;�;;u0;�Y;���:�q�:�;u9�{���D�?T��hs�UFB�}��������μo���d�	����+�K�3�      r₽�؀���u��Xc���K�|1�������վ��]����P����>T����9���o�H4�9�&�:x�	;~%;y�5;��>;ԻC;�F;�!G;՚G;�G;{H;�HH;lH;هH;��H;έH;�H;��H;��H;��H;�H;��H;��H;��H;�H;ЭH;��H;هH;
lH;�HH;{H;�G;ۚG;�!G;�F;ջC;��>;y�5;~%;z�	;�&�:84�9��o���9�?T�������P��]���վ�����|1���K��Xc���u��؀�      <S���r��v�����ԓ����u���N���(��i�͌˼�A����P�hs��1|�����\:b�:��;�n-;�:;�A;�,E;��F;doG;.�G;�H;8H;}_H;?~H;)�H;<�H;��H;K�H;��H;w�H;��H;w�H;��H;L�H;��H;A�H;)�H;?~H;{_H;8H;�H;.�G;goG;��F;�,E;�A;�:;�n-;��;d�:\:����1|��hs���P��A��Ό˼�i���(���N���u�ԓ�����v���r��      �o��s��置�ս9@��tĥ�{^���Xc�G�3���	�Ό˼�]��UFB��Z򻬜��QӺ ��8��:��;�M#;�=5;>?;��C;�@F;>:G;+�G;Q�G;k'H;�RH;�tH;�H;��H;c�H;�H;��H;
�H;~�H;
�H;��H;�H;b�H;��H;�H;�tH;�RH;k'H;P�G;,�G;A:G;�@F;��C;>?;�=5;�M#;��;��:���8SӺ�����Z�UFB��]��Ό˼��	�G�3��Xc�{^��tĥ�9@����ս���s�      �#�X� �b'������gٽ:S��*l��S�j�G�3��i��վ�}���
(���ĻYA?�H�B�N�@:�[�:6Q;!�.;�;;�tB;A�E;��F;i�G;*�G;H;�FH;VkH;H;^�H;I�H;��H;I�H;��H;2�H;��H;I�H;��H;F�H;_�H;H;VkH;�FH;H;'�G;i�G;��F;>�E;�tB;�;;$�.;5Q;�[�:V�@:T�B�YA?���Ļ
(�}����վ��i�F�3�S�j�+l��:S���gٽ����b'�X� �      �S�*�O��E��5�X� �Z�
���罨9��*l���Xc���(��������[�����ݎ�!ܺP<9V��:[�	;\d';� 8;u�@;��D;�F;YjG;��G;�H;�:H;qbH;�H;E�H;j�H;�H;��H;q�H;�H;r�H;��H;�H;h�H;F�H;�H;qbH;�:H;�H;��G;XjG;�F;��D;u�@;� 8;_d';Y�	;V��:`<9'ܺ�ݎ������[��������(��Xc�*l���9�����Z�
�X� ��5��E�*�O�      �~��*��,�v��9b�}�H�#,�OZ����:S��z^����N������μ�I���%+����̝.����
k~:���:Am;��3;R�>;[�C;tPF;�FG;x�G;#�G;�/H;0ZH;�zH;��H;��H;��H;]�H;a�H;�H;b�H;]�H;��H;��H;��H;�zH;/ZH;�/H;#�G;v�G;�FG;vPF;W�C;R�>;��3;Dm;���:
k~:���Ν.�����%+��I����μ�����N�z^��:S�����OZ�#,�}�H��9b�,�v�*��      ����*����:���M��H�r�*�O�#,�Z�
��gٽsĥ���u�|1�o���.Ϥ���P�[�.o�Zp���:���:
Q;[�/;q�<;!C;O�E;�!G;Y�G;7�G;�%H;�RH;uH;7�H;~�H;�H;@�H;��H;>�H;��H;@�H;�H;|�H;:�H;uH;�RH;�%H;7�G;W�G;�!G;P�E;C;s�<;[�/;Q;���:�:Vp���.o�[򻮎P�.Ϥ�o���|1���u�sĥ��gٽZ�
�#,�*�O�H�r��M���:��*���      :���v��O;������UP��H�r�}�H�X� ���8@��ԓ����K�d� ־���s�t���񕻒ܺ 6u9_&�:.�;J�+;��:;�"B;��E;�F;��G;�G;vH;bLH;4pH;}�H;��H;ܭH;t�H;�H;��H;�H;r�H;ۭH;��H;��H;5pH;`LH;sH;�G;��G;�F;��E;�"B;��:;J�+;1�;_&�:06u9�ܺ��t����s� ־�d���K�ԓ��8@����X� �}�H�H�r�UP������O;���v��      YVھ�*־25ʾu��������M���9b��5�����ս����Xc�	��Жռ�I��X�$�iT���Z�`Z��`�:�;��';X�8;0RA;�9E;��F;��G;!�G;�H;4GH;JlH;��H;q�H;�H;�H;˻H;��H;˻H;�H;�H;p�H;��H;JlH;2GH;�H;!�G;��G;��F;�9E;+RA;\�8;��';�;\�:`Z���Z�jT��W�$��I��Жռ	���Xc������ս���5��9b��M������u���25ʾ�*־      ���쾶�޾25ʾO;���:��+�v��E�b'����u����u���+��W��A����4���Ļ9)��i���W�:h�; %;"l7;5�@;$�D;�F;xG;��G;{H;hCH;ciH;R�H;ɛH;ܪH;��H;˺H;��H;˺H;��H;ܪH;țH;R�H;ciH;eCH;xH;��G;xG;�F;$�D;1�@;%l7; %;j�;�W�:�i��9)���Ļ��4��A���W缇�+���u�u�����b'��E�+�v��:��O;��25ʾ��޾��      Yh���b���쾪*־�v��*���*��*�O�X� �s��r���؀�K�3���Cݜ�?�>�Q�ѻۡ9�P���po�:E% ;�M#;�6;]A@;"�D;կF;/qG;|�G;YH;	AH;�gH;�H;ŚH;�H;Q�H;.�H;�H;.�H;S�H;�H;ĚH;��H;�gH;AH;VH;|�G;.qG;կF;"�D;XA@;��6;�M#;F% ;lo�:P���ڡ9�R�ѻ?�>�Cݜ���J�3��؀��r��s�X� �*�O�*��*����v���*־���b��      ���	^�X_ݾ��ɾl*���{x�)G�R,�����b��c@{���/�����䙼�J;�M�ͻ��4��V�T��:<;��#;V�6;[@;_�D;ޱF;�lG;��G;�H;�:H;�bH;!�H;c�H;j�H;�H;,�H;�H;,�H;�H;j�H;a�H;$�H;�bH;�:H;}H;��G;�lG;ޱF;_�D;[@;Y�6;��#;=;P��:�V���4�O�ͻ�J;��䙼����/�c@{��b�����R,�)G�{x��l*����ɾX_ݾ	^�      	^�6���:پ~�žj�����9t�s�C������誫�\`w�K-����.`����7�6Sɻ�K/�pxƹ���:�/;�f$;�7;�~@;z�D;��F;�nG;'�G;iH;�;H;�cH;��H;��H;��H;H�H;b�H;[�H;b�H;J�H;��H;��H;��H;�cH;�;H;gH;'�G;�nG;��F;z�D;�~@;�7;�f$;�/;���:pxƹ�K/�6Sɻ��7�.`�����K-�\`w�誫������s�C�9t���j���~�ž�:پ7��      X_ݾ�:پ�V;+���Ƥ�Na����g��$:��Z�sݽ�ƣ��l�j.%��߼k���9.�ʴ��NV��0p�?A�:x;b(&;m�7;J�@;/E;1�F;�uG;U�G;�H;>H;�eH;	�H;��H;��H;�H;�H;�H;�H;�H;��H;��H;
�H;�eH;>H;�H;U�G;�uG;1�F;/E;D�@;o�7;`(&;x;9A�:�0p�MV�˴���9.�l���߼j.%��l��ƣ�sݽ�Z��$:���g�Na���Ƥ�+���V;�:پ      ��ɾ~�ž+��sת��#�����T��J+�=��2̽�s���yZ����Rμjy����[Ϩ�J,� 8�6a��:�
;u�(;�N9;�A;�NE;w�F;�G;�G;�H;�AH;lhH;+�H;w�H;�H;�H;޹H;��H;޹H;�H;�H;u�H;+�H;khH;�AH;�H;�G;�G;w�F;�NE;�A;�N9;s�(;�
;]��: 8�6I,�[Ϩ���jy��Rμ����yZ��s���2̽=��J+���T�#����sת�+��~�ž      l*��j����Ƥ���/��B�c��G=����zｔж��ɇ�V�C���("��w;k��&��-��f�˺�Y�9���:9;i,;�	;;QB;��E;G;��G;�G;�H;9GH;�lH;A�H;ӜH;ЫH;x�H;=�H;�H;=�H;w�H;ϫH;ќH;B�H;�lH;6GH;�H;�G;��G;G;��E;QB;�	;;i,;9;���:�Y�9d�˺�-���&�w;k�("����V�C��ɇ��ж��z����G=�B�c��/����Ƥ�j���      ����Na��#���B�c�s�C�}#� ��VvϽ�����l�hg*����
���I���軷\c��쀺u,:@��:�;�_0;��<;�1C;�E;�#G;v�G;C�G;P H;�MH;qqH;�H;��H;�H;j�H;׼H;��H;׼H;k�H;�H;��H;�H;qqH;�MH;L H;C�G;t�G;�#G;�E;�1C;��<;�_0;�;<��:u,:�쀺�\c�����I��
�����hg*��l�����VvϽ ��}#�s�C�B�c�#���Na����      {x�9t���g���T��G=�}#�6�sݽ�b������GG�����Ǽky��N�$�e����$�xuƹz��:$'�:ɡ ;j4;��>;mD;\F;�FG;��G;:�G;A*H;�UH;3wH;;�H;"�H;��H;��H;��H;g�H;��H;��H;��H;"�H;<�H;3wH;�UH;?*H;:�G;��G;�FG;�[F;gD;��>;j4;ɡ ;'�:z��:huƹ�$�e���N�$�ky���Ǽ���GG������b��sݽ6�}#��G=���T���g�9t�      )G�s�C��$:��J+��� ��sݽ`���0I���yZ���"����֫��hT��� �M����˺Pm9lٶ:��; `(;0�8;��@;��D;�F;�hG;��G;�H;q5H;(^H;�}H;(�H;��H;��H;�H;��H;t�H;��H;�H;��H;��H;+�H;�}H;(^H;m5H;�H;��G;�hG;�F;��D;��@;0�8;"`(;��;lٶ:`m9��˺M���� �hT�֫�������"��yZ�0I��`���sݽ �����J+��$:�s�C�      R,����Z�=��z�VvϽ�b��0I��k]a�J-�k� �%"��}�{�H�!�������4�XP(�FoQ:�L�:(�;�/;�'<;�B;"�E;�F;ʇG;��G;mH;}AH;HgH;��H;r�H;�H;ӶH;��H;4�H;��H;4�H;��H;ӶH;�H;t�H;��H;GgH;xAH;jH;��G;ʇG;�F;�E;�B;�'<;�/;&�;�L�:JoQ:XP(���4�����H�!�}�{�%"��k� �J-�j]a�0I���b��VvϽ�z�=��Z���      ������tݽ�2̽�ж����������yZ�K-�ط�3aļ\O���J;����w�|�y�º�O@9킬:\�;�f$;��5;�N?;qD;�LF;3;G;ܤG;(�G;�!H;NH;�pH;ȋH;�H;e�H;+�H;�H;��H;��H;��H;�H;+�H;d�H;�H;ƋH;�pH;NH;�!H;'�G;ޤG;1;G;�LF;pD;�N?;��5;�f$;\�;:�O@9y�ºw�|�����J;�[O��3aļط�J-��yZ����������ж��2̽tݽ���      �b��誫��ƣ��s���ɇ��l�GG���"�k� �2aļe���I��C��ۙ�;��tƹ��k:���:/�;n>.;=
;;��A;BE;��F;HmG;��G;��G;�2H;&[H;�zH;�H;ʥH;ϳH;��H;l�H;:�H;P�H;:�H;l�H;��H;ͳH;ͥH;�H;�zH;"[H;�2H;��G;��G;DmG;��F;BE;��A;;
;;l>.;/�;���:��k:�tƹ:��ۙ��C��I�e��2aļk� ���"�GG��l��ɇ��s���ƣ�誫�      d@{�]`w��l��yZ�V�C�ig*�������&"��[O���I�@|�8Ϩ�fK/�D$T�zQ:���:��;�(&;$6;�%?;��C;�#F;-$G;Z�G;��G;�H;dCH; hH;��H;��H;��H;#�H;.�H;^�H;��H;��H;��H;`�H;+�H;"�H;��H;��H;��H;hH;dCH;�H;��G;U�G;*$G;�#F;��C;�%?;$6;�(&;��;���:zQ:D$T�fK/�8Ϩ�?|��I�[O��&"����鼱��hg*�V�C��yZ��l�]`w�      ��/�K-�j.%����������Ǽ׫��}�{��J;��C�9Ϩ�BO:������[�9���:�;��;a.1;0(<;�5B;OE;F�F;ffG;�G;o�G;/+H;TH;uH;Y�H;��H;[�H;��H;��H;%�H;8�H;]�H;8�H;"�H;��H;��H;\�H;��H;Y�H;uH;TH;,+H;p�G;�G;afG;B�F;OE;�5B;.(<;a.1;��;�;���:�[�9����BO:�9Ϩ��C��J;�|�{�׫���Ǽ��������i.%�K-�      ������߼Rμ("���
��ky��hT�G�!���軼ۙ�dK/������m9B�:���:P�;^�,;�N9;r@;�^D;�LF;�.G;�G;��G;H;�?H;VdH;T�H;��H;F�H;ֶH;��H;�H;�H;��H;��H;��H;�H;�H;��H;ضH;D�H;��H;S�H;VdH;�?H;H;��G;�G;�.G;�LF;�^D;r@;�N9;a�,;P�;���:B�: m9����dK/��ۙ����G�!�hT�ky���
��("��Rμ�߼���      �䙼/`��l��jy��y;k��I�N�$��� �����w�|�<�H$T��[�9B�:���:=�;;�);H7;�>;�tC;F�E; �F;vG;T�G;��G;>,H;�SH;�sH;ÌH;��H;L�H;�H;��H;r�H;��H;/�H;�H;/�H;��H;t�H;��H;�H;J�H;��H;��H;�sH;�SH;?,H;��G;N�G;vG; �F;E�E;�tC;�>;J7;:�);=�;���:B�:�[�9H$T�;�v�|������� �N�$��I�x;k�ky��l��0`��      �J;���7��9.����&����d���M����4�z�º�tƹzQ:���:���:=�;��(;��5;��=;��B;�[E;s�F;UG;�G;��G;�H;�CH;OfH;�H;��H;/�H;ȶH; �H;��H;��H;5�H;v�H;^�H;v�H;5�H;��H;��H;�H;ȶH;.�H;��H;�H;MfH;�CH;�H;��G;ܩG;UG;q�F;�[E;��B;��=;��5;��(;=�;���:���:zQ:�tƹz�º��4�M��d�����軫&����9.���7�      N�ͻ1Sɻ˴��^Ϩ��-���\c��$���˺`P(��O@9��k:���:�;P�;=�);��5;q�=;IQB;�E;#�F;Y8G;v�G;��G;�	H;�5H;�YH;�wH;�H;�H;�H;μH;��H;��H;^�H;��H;��H;`�H;��H;��H;_�H;��H;��H;μH;�H;�H;�H;|wH;�YH;�5H;�	H;}�G;v�G;X8G;$�F;�E;LQB;q�=;��5;=�);P�;�;���:��k:�O@9XP(���˺�$��\c��-��^Ϩ�̴��7Sɻ      ��4��K/�MV�H,�o�˺퀺�uƹ0m9>oQ:킬:���:��;��;[�,;H7;��=;GQB;��D;�cF;T$G;�G;�G;�G;�)H;�NH;nH;�H;�H;d�H;P�H;N�H;�H;��H;�H;�H;��H;P�H;��H;�H;�H;��H;�H;N�H;M�H;a�H; �H;�H;nH;�NH;�)H;�G;�G;��G;U$G;�cF;��D;GQB;��=;H7;^�,;��;��;���:킬:JoQ:m9�uƹ퀺a�˺H,�NV��K/�      xVṐxƹ�/p� 8�6�Y�9u,:���:hٶ:�L�:[�;/�;�(&;a.1;�N9;�>;��B;�E;�cF;G;e�G;��G;�G;� H;(FH;�eH;�H;��H;�H;��H;žH;L�H;�H;��H;��H;*�H;��H;��H;��H;*�H;��H;��H;�H;K�H;þH;�H;�H;�H;�H;�eH;$FH;� H;�G;�G;g�G;G;�cF;�E;��B;�>;�N9;a.1;�(&;/�;[�;�L�:fٶ:���:.u,:�Y�9 6�6�/p��xƹ      T��:��:=A�:_��:���:8��:'�:��;$�;�f$;k>.;$6;,(<;k@;�tC;�[E;�F;P$G;a�G;�G;S�G;�H;@H;�_H;/zH;��H;\�H;��H;q�H;��H;��H;��H;��H;��H;�H;7�H;��H;8�H;�H;��H;��H;��H;��H;��H;k�H;�H;Z�H;��H;0zH;�_H;@H;�H;P�G;�G;a�G;Q$G;�F;�[E;�tC;k@;,(<;$6;l>.;�f$;$�;��;'�:>��:���:_��:9A�:
��:      F;�/;"x;��
;9;�;̡ ; `(;�/;��5;:
;;�%?;�5B;�^D;C�E;r�F;X8G;�G;��G;V�G;	H;�<H;�[H;'vH;ċH;��H;w�H;|�H;��H;��H;��H;��H;H�H;��H;��H;��H;�H;��H;��H;��H;H�H;��H;��H;��H;��H;z�H;v�H;��H;ċH;$vH;�[H;�<H;H;V�G;��G;�G;W8G;r�F;C�E;�^D;�5B;�%?;8
;;��5;�/;`(;Ρ ;�;9;��
;x;�/;      ��#;�f$;s(&;n�(;i,;�_0;x4;9�8;�'<;�N?;��A;��C;OE;�LF; �F;UG;v�G;�G;�G;�H;�<H;�ZH;tH;6�H;ݚH;ɩH;�H;�H;��H;U�H;{�H;n�H;��H;��H;(�H;�H;P�H;�H;(�H;��H;��H;n�H;|�H;Q�H;��H;�H;�H;ʩH;ߚH;2�H;tH;�ZH;�<H;�H;�G;!�G;t�G;UG;!�F;�LF;OE;��C;��A;�N?;�'<;7�8;x4;�_0;i,;n�(;p(&;�f$;      ^�6;�7;o�7;�N9;�	;;��<;��>;��@;�B;pD;BE;�#F;C�F;�.G;vG;ߩG;~�G;�G;� H;@H;�[H;tH;s�H;��H;.�H;h�H;?�H;c�H;8�H;`�H;��H;��H;��H;i�H;v�H;-�H;n�H;-�H;u�H;i�H;~�H;��H;��H;_�H;6�H;b�H;<�H;h�H;.�H;��H;s�H;tH;�[H;@H;� H;�G;~�G;ݩG;vG;�.G;E�F;�#F;BE;pD;�B;��@;��>;��<;�	;;�N9;o�7;�7;      2[@;�~@;T�@;�A;QB;�1C;sD;��D;�E;�LF;��F;-$G;`fG;�G;O�G;��G;�	H;�)H;'FH;�_H;"vH;4�H;��H;��H;x�H;Z�H;h�H; �H;��H;��H;I�H;�H;�H;��H;��H;6�H;�H;6�H;��H;��H;�H;�H;I�H;��H;��H;�H;h�H;Z�H;x�H;��H;��H;5�H;!vH;�_H;'FH;�)H;�	H;��G;Q�G;�G;`fG;-$G;��F;�LF;!�E;��D;qD;�1C;QB;�A;R�@;�~@;      q�D;��D;E;�NE;��E;�E;�[F;�F;�F;0;G;DmG;Z�G;�G;��G;��G;�H;�5H;�NH;�eH;6zH;ƋH;�H;4�H;��H;�H;��H;g�H;��H;5�H;��H;��H;��H;��H;��H;��H;.�H;K�H;,�H;��H;��H;��H;��H;��H;��H;4�H;��H;e�H;��H;�H;}�H;3�H;�H;ƋH;9zH;�eH;�NH;�5H;�H;��G;��G;�G;[�G;DmG;.;G;�F;�F;�[F;�E;��E;�NE;E;��D;      �F;��F;#�F;w�F;G;�#G;�FG;�hG;ɇG;ܤG;��G;��G;l�G;H;;,H;�CH;�YH;nH;�H;��H;��H;ǩH;e�H;X�H;��H;2�H;s�H;��H;Q�H;\�H;��H;B�H;��H;��H;��H;��H;��H;��H;��H;��H;��H;D�H;��H;Z�H;Q�H;��H;u�H;2�H;��H;W�H;d�H;ƩH;��H;��H;�H;nH;�YH;�CH;;,H;H;o�G;��G;��G;ۤG;ʇG;hG;�FG;�#G;G;w�F;!�F;��F;      �lG;�nG;�uG;�G;��G;z�G;��G;��G;��G;%�G;��G;�H;-+H;�?H;�SH;OfH;�wH;�H;��H;_�H;y�H;�H;?�H;l�H;a�H;v�H;��H;�H;�H;h�H;Z�H;��H;��H;��H;;�H;��H;��H;��H;;�H;��H;��H;��H;Z�H;f�H; �H;�H;��H;v�H;c�H;j�H;=�H;�H;w�H;a�H;��H;�H;�wH;OfH;�SH;�?H;-+H;�H;��G;%�G;��G;��G;��G;x�G;�G;�G;�uG;�nG;      ��G;(�G;]�G;�G;�G;C�G;>�G;�H;mH;�!H;�2H;hCH;TH;XdH;�sH;�H;�H;��H;�H;��H;|�H;�H;c�H;�H;��H;��H;�H;��H;M�H;�H;��H;��H;��H;v�H;��H;�H;T�H;�H;��H;x�H;��H;��H;��H;�H;L�H;��H;�H;��H;��H;�H;b�H;�H;y�H;��H;�H;��H;�H;�H;�sH;VdH;TH;hCH;�2H;�!H;oH;�H;>�G;C�G;�G;�G;\�G;3�G;      �H;hH;�H;�H;�H;Q H;F*H;q5H;{AH;NH;%[H;#hH;uH;S�H;��H;��H;�H;a�H;��H;r�H;��H;��H;8�H;��H;/�H;S�H;��H;M�H;�H;��H;��H;��H;q�H;��H;P�H;��H;��H;��H;P�H;��H;o�H;��H;��H;��H;�H;M�H;�H;S�H;1�H;��H;6�H;��H;��H;r�H;��H;c�H;�H;��H;H;S�H;uH;"hH;#[H;NH;~AH;p5H;D*H;Q H;�H;�H;�H;^H;      �:H;�;H;>H;�AH;IGH;�MH;�UH;.^H;PgH; qH;�zH;��H;_�H;��H;��H;1�H;�H;J�H;þH;��H;��H;R�H;_�H;��H;��H;Y�H;f�H;�H;��H;��H;��H;h�H;��H;p�H;��H;��H;��H;��H;��H;p�H;��H;h�H;��H;��H;��H;�H;f�H;Y�H;��H;��H;]�H;R�H;��H;��H;þH;L�H;�H;1�H;��H;��H;_�H;��H;�zH; qH;SgH;0^H;�UH;�MH;EGH;�AH;>H;�;H;      �bH;�cH;�eH;vhH;�lH;sqH;:wH;�}H;��H;̋H;�H;��H;��H;J�H;M�H;϶H;ԼH;M�H;L�H;��H;��H;|�H;��H;M�H;��H;��H;Y�H;��H;��H;��H;}�H;��H;d�H;��H;�H;+�H;M�H;-�H;�H;��H;b�H;��H;|�H;��H;��H;��H;Y�H;��H;��H;M�H;��H;|�H;��H;��H;L�H;M�H;ӼH;ζH;M�H;I�H;��H;��H;�H;͋H;��H;�}H;:wH;tqH;�lH;whH;�eH;�cH;      5�H;��H;�H;1�H;F�H;�H;>�H;1�H;w�H;�H;ХH;��H;^�H;ܶH;
�H;�H;��H;�H;�H;��H;��H;r�H;��H;�H;��H;B�H;��H;��H;��H;j�H;��H;|�H;��H;*�H;P�H;}�H;l�H;{�H;P�H;*�H;��H;|�H;��H;k�H;��H;��H;��H;A�H;��H;�H;��H;r�H;��H;��H;�H;�H;��H;�H;
�H;ܶH;^�H;��H;ХH;�H;w�H;.�H;>�H;�H;E�H;/�H;�H;��H;      h�H;ėH;��H;|�H;ۜH;��H;#�H;��H;	�H;d�H;ϳH;)�H;��H;��H;��H;��H;��H;��H;��H;��H;P�H;��H;��H;�H;��H;��H;��H;��H;v�H;�H;g�H;��H;8�H;Q�H;��H;��H;o�H;��H;��H;Q�H;5�H;��H;g�H;�H;x�H;��H;��H;��H;��H;�H;��H;��H;O�H;��H;��H;��H;��H;��H;��H;��H;��H;'�H;ϳH;e�H;
�H;��H;#�H;��H;ԜH;|�H;��H;��H;      x�H;��H;��H;�H;٫H;�H;ðH;��H;ضH;,�H;��H;1�H;��H;�H;v�H;��H;e�H;�H;��H;��H;��H;��H;j�H;��H;��H;��H;��H;v�H;��H;r�H;��H;*�H;J�H;��H;��H;��H;��H;��H;��H;��H;I�H;+�H;��H;s�H;��H;v�H;��H;��H;��H;��H;j�H;��H;��H;��H;��H;�H;c�H;��H;v�H;�H;��H;1�H;��H;,�H;ضH;��H;ðH;�H;ϫH;�H;��H;��H;      �H;]�H;��H;�H;��H;h�H;��H;�H;žH;��H;r�H;g�H;(�H;�H;��H;=�H;��H;��H;-�H;�H;��H;,�H;v�H;��H;��H;��H;9�H;��H;Q�H;��H;�H;S�H;��H;��H;��H;��H;��H;��H;��H;��H;��H;U�H;�H;��H;S�H;��H;7�H;��H;��H;��H;v�H;,�H;��H;�H;-�H;��H;��H;=�H;��H;�H;(�H;g�H;p�H;��H;žH;�H;��H;m�H;��H;�H;��H;U�H;      '�H;h�H;��H;߹H;L�H;ӼH;ľH;��H;>�H;��H;?�H;��H;=�H;��H;3�H;}�H;��H;��H;��H;B�H;��H;�H;0�H;<�H;'�H;��H;��H;�H;��H;��H;+�H;~�H;��H;��H;��H;��H;��H;��H;��H;��H;��H;��H;+�H;��H;��H;�H;��H;��H;(�H;;�H;0�H;�H;��H;B�H;��H;��H;��H;}�H;2�H;��H;=�H;��H;?�H;��H;>�H;��H;ľH;׼H;@�H;�H;��H;`�H;      �H;b�H;��H;��H;�H;��H;k�H;x�H;��H;��H;U�H;��H;`�H;��H;�H;f�H;e�H;G�H;��H;��H;�H;U�H;n�H;��H;F�H;��H;��H;Z�H;��H;��H;P�H;q�H;m�H;��H;��H;��H;��H;��H;��H;��H;j�H;s�H;P�H;��H;��H;Z�H;��H;��H;F�H;��H;n�H;U�H;�H;��H;��H;I�H;d�H;f�H;�H;��H;`�H;��H;U�H;��H;��H;u�H;k�H;��H;�H;��H; �H;Y�H;      '�H;i�H;��H;�H;L�H;ӼH;ľH;��H;>�H;��H;?�H;��H;=�H;��H;2�H;}�H;��H;��H;��H;B�H;��H;�H;0�H;<�H;(�H;��H;��H;�H;��H;��H;+�H;~�H;��H;��H;��H;��H;��H;��H;��H;��H;��H;��H;+�H;��H;��H;�H;��H;��H;'�H;;�H;0�H;�H;��H;B�H;��H;��H;��H;}�H;2�H;��H;=�H;��H;A�H;��H;@�H;��H;ľH;׼H;@�H;�H;��H;^�H;      �H;]�H;�H;�H;��H;h�H;��H;�H;žH;��H;o�H;g�H;(�H;�H;��H;=�H;��H;��H;-�H;�H;��H;,�H;v�H;��H;��H;��H;9�H;��H;Q�H;��H;�H;S�H;��H;��H;��H;��H;��H;��H;��H;��H;��H;W�H;�H;��H;S�H;��H;7�H;��H;��H;��H;v�H;,�H;��H;�H;-�H;��H;��H;=�H;��H;�H;(�H;g�H;p�H;��H;žH;�H;��H;k�H;��H;�H;��H;U�H;      y�H;��H;��H;�H;٫H;�H;ðH;��H;ضH;,�H;��H;1�H;��H;�H;v�H;��H;e�H;�H;��H;��H;��H;��H;j�H;��H;��H;��H;��H;v�H;��H;r�H;��H;(�H;J�H;��H;��H;��H;��H;��H;��H;��H;I�H;-�H;��H;s�H;��H;v�H;��H;��H;��H;��H;j�H;��H;��H;��H;��H;�H;c�H;��H;v�H;�H;��H;1�H;��H;,�H;ٶH;��H;ðH;�H;ͫH;�H;��H;��H;      k�H;H;��H;~�H;ڜH;��H;#�H;��H;
�H;d�H;ϳH;'�H;��H;��H;��H;��H;��H;��H;��H;��H;Q�H;��H;��H;�H;��H;��H;��H;��H;v�H;�H;g�H;��H;6�H;P�H;��H;��H;o�H;��H;��H;P�H;5�H;��H;g�H;�H;x�H;��H;��H;��H;��H;�H;��H;��H;O�H;��H;��H;��H;��H;��H;��H;��H;��H;)�H;ϳH;e�H;	�H;��H;#�H;��H;ќH;~�H;��H;��H;      5�H;��H;�H;.�H;F�H;�H;A�H;1�H;u�H;�H;ХH;��H;^�H;ܶH;
�H;�H;��H;�H;�H;��H;��H;r�H;��H;�H;��H;B�H;��H;��H;��H;j�H;��H;|�H;��H;*�H;P�H;}�H;l�H;{�H;P�H;*�H;��H;}�H;��H;k�H;��H;��H;��H;A�H;��H;�H;��H;r�H;��H;��H;�H;�H;��H;�H;
�H;ܶH;\�H;��H;ХH;�H;x�H;.�H;A�H;�H;C�H;.�H;�H;��H;      �bH;�cH;�eH;whH;�lH;sqH;:wH;�}H;��H;̋H;�H;��H;��H;J�H;M�H;϶H;ӼH;K�H;L�H;��H;��H;|�H;��H;N�H;��H;��H;Y�H;��H;��H;��H;|�H;��H;d�H;��H;�H;-�H;M�H;+�H;�H;��H;a�H;��H;}�H;��H;��H;��H;Y�H;��H;��H;M�H;��H;|�H;��H;��H;L�H;M�H;ӼH;϶H;M�H;J�H;��H;��H;�H;͋H;��H;�}H;:wH;vqH;�lH;vhH;�eH;�cH;      �:H;�;H;>H;�AH;DGH;�MH;�UH;0^H;RgH;�pH;�zH;��H;_�H;��H;��H;1�H;�H;J�H;þH;��H;��H;R�H;_�H;��H;��H;Z�H;h�H;�H;��H;��H;��H;g�H;��H;o�H;��H;��H;��H;��H;��H;p�H;��H;j�H;��H;��H;��H;�H;e�H;W�H;��H;��H;]�H;R�H;��H;��H;þH;L�H;�H;2�H;��H;��H;_�H;��H;�zH;�pH;SgH;0^H;�UH;�MH;BGH;�AH;>H;�;H;      �H;eH;�H;�H;�H;L H;G*H;s5H;}AH;NH;%[H;#hH;uH;S�H;ÌH;��H;�H;a�H;��H;t�H;��H;��H;8�H;��H;1�H;T�H; �H;M�H;�H;��H;��H;��H;q�H;��H;O�H;��H;��H;��H;P�H;��H;o�H;��H;��H;��H;�H;M�H; �H;Q�H;/�H;��H;6�H;��H;��H;r�H;��H;c�H;�H;��H;��H;S�H;uH;#hH;%[H;NH;~AH;q5H;H*H;P H;�H;�H;�H;eH;      ��G;(�G;]�G;�G;�G;C�G;>�G;�H;mH;�!H;�2H;hCH;TH;XdH;�sH;�H;�H;��H;�H;��H;~�H;�H;c�H;�H;��H;��H;�H;��H;M�H;�H;��H;��H;��H;v�H;��H;�H;T�H;�H;��H;v�H;��H;��H;��H;�H;L�H;��H;�H;��H;��H;�H;b�H;�H;y�H;��H;�H;��H;�H;�H;�sH;VdH;TH;hCH;�2H;�!H;oH;�H;>�G;@�G;�G;�G;]�G;5�G;      �lG;�nG;�uG;�G;��G;v�G;��G;��G;��G;'�G;��G;�H;-+H;�?H;�SH;QfH;�wH;�H;��H;b�H;}�H;�H;?�H;l�H;c�H;w�H;��H;�H; �H;h�H;Z�H;��H;��H;��H;;�H;��H;��H;��H;;�H;��H;��H;��H;Z�H;f�H;��H;�H;��H;v�H;a�H;j�H;=�H;�H;v�H;_�H;��H;�H;wH;OfH;�SH;�?H;-+H;�H;��G;'�G;��G;��G;��G;t�G;��G;�G;�uG;�nG;      ��F;��F;-�F;x�F;G;�#G;�FG;�hG;ȇG;ܤG;��G;��G;o�G;H;;,H;�CH;�YH;nH;�H;��H;��H;ƩH;e�H;X�H;��H;3�H;u�H;��H;S�H;\�H;��H;B�H;��H;��H;��H;��H;��H;��H;��H;��H;��H;D�H;��H;Y�H;P�H;��H;r�H;2�H;��H;X�H;e�H;ǩH;��H;��H;�H;nH;�YH;�CH;;,H;H;l�G;��G;��G;ۤG;ɇG;hG;�FG;�#G;G;x�F;-�F;��F;      q�D;��D;E;�NE;��E;�E;�[F;�F;�F;0;G;FmG;[�G;�G;��G;��G;�H;�5H;�NH;�eH;9zH;ˋH;�H;5�H;��H;�H;��H;g�H;��H;6�H;��H;��H;��H;��H;��H;��H;,�H;K�H;.�H;��H;��H;��H;��H;��H;��H;2�H;��H;d�H;��H;�H;�H;1�H;�H;ƋH;7zH;�eH;�NH;�5H;�H;��G;��G;�G;Z�G;DmG;.;G;�F;�F;�[F;�E;��E;�NE;E;��D;      :[@;�~@;W�@;�A;QB;�1C;pD;��D;!�E;�LF;��F;-$G;afG;�G;Q�G;��G;�	H;�)H;'FH;�_H;%vH;5�H;��H;��H;x�H;Z�H;i�H;�H;��H;��H;I�H;�H;�H;��H;��H;6�H;�H;6�H;��H;��H;�H;�H;I�H;��H;��H; �H;h�H;Z�H;x�H;��H;��H;4�H; vH;�_H;'FH;�)H;�	H;��G;O�G;�G;`fG;-$G;��F;�LF;"�E;��D;pD;�1C;QB;�A;U�@;�~@;      Y�6;�7;�7;�N9;�	;;��<;��>;��@;�B;pD;BE;�#F;C�F;�.G;vG;ߩG;�G;�G;� H;@H;�[H;tH;u�H;��H;.�H;g�H;?�H;b�H;8�H;b�H;��H;��H;��H;i�H;u�H;-�H;n�H;-�H;v�H;i�H;~�H;��H;��H;]�H;5�H;c�H;=�H;h�H;.�H;��H;r�H;tH;�[H;@H;� H;�G;~�G;ߩG;vG;�.G;B�F;�#F;BE;mD;�B;��@;��>;��<;�	;;�N9;t�7;�7;      ��#;�f$;s(&;n�(;i,;�_0;x4;9�8;�'<;�N?;��A;��C;OE;�LF; �F;UG;t�G;�G;�G;�H;�<H;�ZH;tH;6�H;ߚH;ɩH;�H;�H;��H;U�H;|�H;o�H;��H;��H;(�H;�H;P�H;�H;(�H;��H;��H;n�H;{�H;Q�H;��H;�H;�H;ʩH;ݚH;4�H;tH;�ZH;�<H;�H;�G;�G;t�G;UG;!�F;�LF;OE;��C;��A;�N?;�'<;9�8;x4;�_0;i,;n�(;q(&;�f$;      >;�/;&x;��
;9;�;С ;#`(;�/;��5;;
;;�%?;�5B;�^D;C�E;r�F;X8G;�G;��G;U�G;	H;�<H;�[H;(vH;ċH;��H;w�H;z�H;��H;��H;��H;��H;I�H;��H;��H;��H;�H;��H;��H;��H;H�H;��H;��H;��H;��H;|�H;v�H;��H;ċH;$vH;�[H;�<H;H;V�G;��G;�G;W8G;r�F;C�E;�^D;�5B;�%?;:
;;��5;�/;"`(;С ;
�;9;��
;$x;�/;      P��:��:EA�:Y��:���:6��:'�:��;$�;�f$;l>.;$6;,(<;k@;�tC;�[E;�F;P$G;a�G;�G;U�G;�H;@H;�_H;0zH;��H;\�H;�H;q�H;��H;��H;��H;��H;��H;�H;:�H;��H;8�H;�H;��H;��H;��H;��H;��H;k�H;��H;[�H;��H;/zH;�_H;@H;�H;R�G;�G;a�G;Q$G;�F;�[E;�tC;k@;*(<;$6;i>.;�f$;$�;��; '�:<��:���:[��:?A�:��:      xVṐxƹ�/p� 6�6�Y�9u,:���:hٶ:�L�:[�;/�;�(&;a.1;�N9;�>;��B;�E;�cF;G;e�G;��G;�G;� H;(FH;�eH;�H;��H;�H;��H;žH;K�H;�H;��H;��H;(�H;��H;��H;��H;*�H;��H;��H;�H;L�H;þH;�H;�H;�H;�H;�eH;%FH;� H;�G;�G;g�G;G;�cF;�E;��B;�>;�N9;a.1;�(&;/�;[�;�L�:fٶ:���:.u,:�Y�9 8�6�/p��xƹ      ��4��K/�LV�H,�q�˺퀺�uƹ m9>oQ::���:��;��;[�,;H7;��=;GQB;��D;�cF;T$G;�G;�G;�G;�)H;�NH;nH;�H; �H;d�H;O�H;N�H;�H;��H;�H;�H;��H;P�H;��H;�H;�H;��H;�H;N�H;O�H;c�H;�H;�H;nH;�NH;�)H;�G;�G; �G;U$G;�cF;��D;EQB;��=;H7;[�,;��;��;���:킬:JoQ: m9�uƹ퀺d�˺I,�NV��K/�      N�ͻ2Sɻ˴��^Ϩ��-���\c��$���˺`P(��O@9��k:���:�;P�;=�);��5;r�=;HQB;�E;#�F;Y8G;v�G;��G;�	H;�5H;�YH;�wH;�H;�H;�H;μH;��H;��H;_�H;��H;��H;`�H;��H;��H;_�H;��H;��H;μH;�H;�H;�H;}wH;�YH;�5H;�	H;}�G;v�G;X8G;$�F;�E;KQB;q�=;��5;=�);P�;�;���:��k:�O@9XP(���˺�$��\c��-��^Ϩ�̴��8Sɻ      �J;���7��9.����&����d���M����4�y�º�tƹzQ:���:���:=�;��(;��5;��=;��B;�[E;r�F;UG;ݩG;��G;�H;�CH;OfH;�H;��H;.�H;ȶH; �H;��H;��H;5�H;v�H;^�H;v�H;5�H;��H;��H;�H;ȶH;/�H;��H;�H;MfH;�CH;�H;��G;ݩG;UG;r�F;�[E;��B;��=;��5;��(;=�;���:���:zQ:�tƹ|�º��4�M��d�����軫&����9.���7�      �䙼/`��l��jy��x;k��I�O�$��� �����v�|�<�H$T��[�9B�:���:=�;;�);H7;�>;�tC;E�E; �F;vG;R�G;��G;>,H;�SH;�sH;ŌH;��H;J�H;�H;��H;t�H;��H;/�H;�H;/�H;��H;t�H;��H;�H;L�H;��H;��H;�sH;�SH;?,H;��G;O�G;vG; �F;F�E;�tC;�>;J7;:�);=�;���:B�:�[�9L$T�<�x�|������� �N�$��I�x;k�jy��l��0`��      ������߼Rμ("���
��ky��hT�G�!���軼ۙ�fK/������m9B�:���:P�;_�,;�N9;q@;�^D;�LF;�.G;�G;��G;H;�?H;VdH;T�H;��H;D�H;նH;��H;�H;�H;��H;��H;��H;�H;�H;��H;ضH;F�H;��H;S�H;VdH;�?H;H;��G;�G;�.G;�LF;�^D;q@;�N9;a�,;P�;���:B�:�m9����fK/��ۙ����G�!�hT�ky���
��("��Rμ�߼���      ��/�K-�j.%����������Ǽ׫��|�{��J;��C�9Ϩ�BO:������[�9���:�;��;a.1;.(<;�5B;OE;F�F;ffG;�G;n�G;/+H;TH;uH;Y�H;��H;[�H;��H;��H;"�H;8�H;]�H;8�H;$�H;��H;��H;[�H;��H;Y�H;uH;TH;,+H;s�G;�G;`fG;B�F;OE;�5B;.(<;a.1;��;�;���:�[�9����BO:�9Ϩ��C��J;�}�{�׫���Ǽ��������i.%�K-�      d@{�]`w��l��yZ�V�C�hg*�������&"��[O���I�?|�8Ϩ�fK/�D$T�zQ:���:��;�(&;$6;�%?;��C;�#F;-$G;U�G;��G;�H;dCH;hH;��H;��H;��H;%�H;-�H;`�H;��H;��H;��H;^�H;.�H;"�H;��H;��H;��H;hH;dCH;�H;��G;Z�G;($G;�#F;��C;�%?;$6;�(&;��;���:vQ:D$T�fK/�8Ϩ�?|��I�[O��&"����鼱��hg*�V�C��yZ��l�]`w�      �b��誫��ƣ��s���ɇ��l�GG���"�k� �2aļe���I��C��ۙ�:��tƹ��k:���:/�;n>.;:
;;��A;BE;��F;DmG;��G;��G;�2H;%[H;�zH;�H;ʥH;ϳH;��H;l�H;:�H;P�H;:�H;l�H;��H;ͳH;ͥH;�H;�zH;#[H;�2H;��G;��G;HmG;��F;BE;��A;;
;;l>.;/�;���:��k:�tƹ;��ۙ��C��I�e��2aļk� ���"�GG��l��ɇ��s���ƣ�誫�      ������tݽ�2̽�ж����������yZ�K-�ط�3aļ\O���J;����w�|�y�º�O@9킬:\�;�f$;��5;�N?;qD;�LF;1;G;ܤG;(�G;�!H;NH;�pH;ƋH;�H;e�H;+�H;�H;��H;��H;��H;�H;+�H;d�H;�H;ȋH;�pH;NH;�!H;'�G;ޤG;3;G;�LF;pD;�N?;��5;�f$;\�;:�O@9|�ºw�|�����J;�\O��3aļط�K-��yZ����������ж��2̽tݽ���      R,����Z�=��z�VvϽ�b��0I��k]a�J-�k� �%"��}�{�H�!�������4�TP(�FoQ:�L�:(�;�/;�'<;�B;"�E;�F;ʇG;��G;jH;{AH;GgH;��H;r�H;�H;ӶH;��H;4�H;��H;4�H;��H;ӶH;�H;r�H;��H;GgH;zAH;mH;��G;ʇG;�F;�E;�B;�'<;�/;&�;�L�:JoQ:`P(���4�����H�!�}�{�%"��k� �J-�j]a�0I���b��VvϽ�z�=��Z���      )G�s�C��$:��J+��� ��sݽ`���0I���yZ���"����֫��hT��� �M����˺Pm9lٶ:��;`(;0�8;��@;��D;�F;�hG;��G;�H;q5H;(^H;�}H;(�H;��H;��H;�H;��H;t�H;��H;�H;��H;��H;*�H;�}H;(^H;o5H;�H;��G;�hG;�F;��D;��@;0�8;"`(;��;lٶ:`m9��˺M���� �hT�֫�������"��yZ�0I��`���sݽ �����J+��$:�s�C�      {x�9t���g���T��G=�}#�6�sݽ�b������GG�����Ǽky��N�$�e����$�puƹz��:'�:ǡ ;j4;��>;mD;�[F;�FG;��G;:�G;A*H;�UH;3wH;;�H;#�H;��H;��H;��H;g�H;��H;��H;��H;!�H;;�H;3wH;�UH;@*H;:�G;��G;�FG;\F;iD;��>;j4;̡ ;'�:z��:huƹ�$�f���N�$�ky���Ǽ���GG������b��sݽ6�}#��G=���T���g�9t�      ����Na��#���B�c�s�C�}#� ��VvϽ�����l�hg*����
���I���軸\c��쀺u,:<��: �;�_0;��<;�1C;�E;�#G;v�G;C�G;P H;�MH;qqH;�H;��H;�H;k�H;׼H;��H;ڼH;j�H;�H;��H;�H;qqH;�MH;L H;C�G;t�G;�#G;�E;�1C;��<;�_0;�;<��:u,:�쀺�\c�����I��
�����hg*��l�����VvϽ ��}#�s�C�B�c�#���Na����      l*��j����Ƥ���/��B�c��G=����zｔж��ɇ�V�C���("��w;k��&��-��f�˺�Y�9���:9;i,;�	;;QB;��E;G;��G;�G;�H;9GH;�lH;A�H;ӜH;ϫH;x�H;=�H;�H;=�H;w�H;ЫH;ќH;B�H;�lH;6GH;�H;�G;��G;G;��E;QB;�	;;i,;9;���:�Y�9d�˺�-���&�w;k�("����V�C��ɇ��ж��z����G=�B�c��/����Ƥ�j���      ��ɾ~�ž+��sת��#�����T��J+�=��2̽�s���yZ����Rμjy����[Ϩ�I,� 8�6_��:�
;s�(;�N9;�A;�NE;w�F;�G;�G;�H;�AH;khH;+�H;w�H;�H;�H;޹H;��H;޹H;�H;�H;u�H;*�H;lhH;�AH;�H;�G;�G;w�F;�NE;�A;�N9;u�(;�
;_��: 8�6I,�\Ϩ���jy��Rμ����yZ��s���2̽=��J+���T�#����sת�+��~�ž      X_ݾ�:پ�V;+���Ƥ�Na����g��$:��Z�sݽ�ƣ��l�j.%��߼k���9.�ʴ��NV��0p�9A�:x;`(&;k�7;J�@;/E;/�F;�uG;U�G;�H;>H;�eH;
�H;��H;��H;�H;�H;�H;�H;�H;��H;��H;	�H;�eH;>H;�H;U�G;�uG;/�F;/E;F�@;o�7;b(&;x;;A�:�0p�LV�˴���9.�l���߼j.%��l��ƣ�sݽ�Z��$:���g�Na���Ƥ�+���V;�:پ      	^�6���:پ~�žj�����9t�s�C������誫�\`w�K-����.`����7�6Sɻ�K/�pxƹ���:�/;�f$;�7;�~@;z�D;��F;�nG;'�G;iH;�;H;�cH;��H;��H;��H;H�H;b�H;[�H;b�H;J�H;��H;��H;��H;�cH;�;H;gH;'�G;�nG;��F;z�D;�~@;�7;�f$;�/;���:pxƹ�K/�6Sɻ��7�.`�����K-�\`w�誫������s�C�9t���j���~�ž�:پ6��      IF�Zh����XVھ:�������~���S��#��o��<S��r₽6�6�u���my��ZFB��Eֻ�A?���	��Y�:���:{�";�46;j@;��D;کF;�nG; �G;@H;<@H;gH;��H;d�H;ĩH;�H;�H;��H;�H;�H;ĩH;c�H;��H;gH;;@H;=H; �G;�nG;۩F;��D;g@;�46;{�";���:�Y�:��	��A?��EֻZFB�my��u���6�6�r₽<S���o���#��S��~������:��XVھ��Zh��      Zh���b���쾪*־�v��+���*��*�O�X� �s��r���؀�K�3���Cݜ�@�>�R�ѻ�9�`���lo�:A% ;�M#;}�6;[A@;�D;ԯF;,qG;|�G;UH;AH;�gH;�H;ĚH;�H;P�H;,�H;�H;,�H;Q�H;�H;ÚH;�H;�gH;AH;RH;|�G;,qG;ԯF;�D;VA@;��6;�M#;A% ;ho�:h���ޡ9�S�ѻ@�>�Cݜ���K�3��؀��r��s�X� �*�O�*��+����v���*־���b��      ���쾶�޾25ʾO;���:��,�v��E�b'����t����u���+��W��A����4���Ļ9)� j���W�:h�;%;!l7;5�@; �D;�F;xG;��G;xH;hCH;biH;Q�H;ƛH;٪H;��H;ʺH;��H;ʺH;��H;٪H;śH;Q�H;biH;eCH;vH;��G;xG;�F; �D;0�@;#l7;%;g�;�W�: j��9)���Ļ��4��A���W缇�+���u�t�����b'��E�,�v��:��O;��25ʾ��޾��      XVھ�*־25ʾu��������M���9b��5�����ս����Xc�	��Жռ�I��X�$�jT���Z��Z��V�:�;��';X�8;.RA;�9E;��F;݂G;!�G;�H;3GH;IlH;��H;o�H;�H;��H;ɻH;��H;ɻH;��H;�H;m�H;��H;JlH;0GH;�H; �G;݂G;��F;�9E;(RA;[�8;��';�;T�:�Z���Z�kT��X�$��I��Жռ	���Xc������ս���5��9b��M������u���25ʾ�*־      :���v��O;������UP��I�r�~�H�X� ���8@��ԓ����K�d� ־���s�u���񕻗ܺ�5u9[&�:-�;H�+;��:;�"B;��E;�F;�G;�G;qH;bLH;3pH;|�H;��H;ۭH;t�H;�H;��H;�H;q�H;٭H;��H;�H;3pH;`LH;pH;�G;��G;�F;��E;�"B;��:;H�+;.�;Y&�: 6u9�ܺ��u����s� ־�d���K�ԓ��8@����X� �~�H�I�r�UP������O;���v��      ����+����:���M��I�r�*�O�#,�Z�
��gٽtĥ���u�|1�o���.Ϥ���P�[�.o�`p���:���:
Q;Y�/;p�<;C;M�E;�!G;U�G;5�G;�%H;�RH;uH;7�H;|�H;�H;?�H;��H;<�H;��H;?�H;�H;{�H;7�H;uH;�RH;�%H;5�G;S�G;�!G;L�E;C;p�<;X�/;Q;���:�:^p���.o�[򻯎P�.Ϥ�o���{1���u�tĥ��gٽZ�
�#,�*�O�I�r��M���:��+���      �~��*��,�v��9b�~�H�#,�OZ����:S��z^����N������μ�I���%+����ѝ.�8���k~:���:Am;��3;P�>;X�C;uPF;�FG;u�G;!�G;�/H;/ZH;�zH;��H;��H;��H;\�H;a�H;�H;a�H;\�H;��H;��H;��H;�zH;.ZH;�/H;!�G;t�G;�FG;rPF;R�C;O�>;��3;Am;���:k~:(���ҝ.�����%+��I����μ�����N�z^��:S�����OZ�#,�~�H��9b�,�v�*��      �S�*�O��E��5�X� �Z�
���罨9��+l���Xc���(��������[�����ݎ�)ܺ0<9R��:X�	;\d';� 8;r�@;��D;�F;XjG;��G;�H;�:H;nbH;�H;C�H;i�H;�H;��H;p�H;�H;p�H;��H;~�H;f�H;E�H;�H;nbH;�:H;�H;��G;XjG;�F;��D;r�@;� 8;]d';W�	;R��:P<9+ܺ�ݎ������[��������(��Xc�+l���9�����Z�
�X� ��5��E�*�O�      �#�X� �b'������gٽ:S��+l��T�j�G�3��i��վ�}���
(���Ļ\A?�\�B�J�@:�[�:5Q;!�.;�;;�tB;>�E;��F;f�G;'�G;H;�FH;VkH;��H;^�H;F�H;��H;H�H;��H;0�H;��H;H�H;��H;F�H;^�H;��H;SkH;�FH;H;%�G;f�G;��F;;�E;�tB;�;;"�.;4Q;�[�:N�@:X�B�\A?���Ļ
(�}����վ��i�G�3�T�j�+l��:S���gٽ����b'�X� �      �o��s��置�ս9@��tĥ�{^���Xc�G�3���	�Ό˼�]��VFB��Z򻭜��XӺ���8��:��;�M#;�=5;;?;��C;�@F;@:G;)�G;P�G;k'H;�RH;�tH;�H;��H;a�H;�H;��H;	�H;}�H;	�H;��H;�H;_�H;��H;�H;�tH;�RH;k'H;M�G;+�G;<:G;�@F;��C;;?;�=5;�M#;��;��:���8XӺ�����Z�VFB��]��Ό˼��	�G�3��Xc�{^��tĥ�9@����ս���s�      <S���r��t�����ԓ����u���N���(��i�Ό˼�A����P�hs��4|�����\:Z�:��;�n-;	�:;�A;�,E;��F;doG;-�G;�H;8H;|_H;=~H;)�H;>�H;��H;K�H;��H;t�H;��H;t�H;��H;I�H;��H;?�H;(�H;=~H;y_H;8H;�H;.�G;coG;��F;�,E;�A;�:;�n-;��;`�:\:����5|��hs���P��A��Ό˼�i���(���N���u�ԓ�����t���r��      s₽�؀���u��Xc���K�|1�������վ��]����P����@T����9���o�<4�9�&�:t�	;}%;w�5;��>;һC;�F;�!G;ؚG;	�G;yH;�HH;
lH;هH;��H;˭H;�H;��H;��H;��H;�H;��H;��H;��H;�H;έH;��H;ׇH;lH;�HH;xH;�G;՚G;�!G;�F;һC;��>;v�5;}%;w�	;�&�:<4�9��o���9�@T�������P��]���վ�����|1���K��Xc���u��؀�      6�6�K�3���+�	��e�o�����μ���}���VFB�hs�AT��#�D��{���;u9�q�:���:�Y;u0;�;;B;":E;�F;2hG;�G;C�G;�0H;�XH;hxH;[�H;��H;=�H;3�H;�H;N�H;f�H;t�H;f�H;N�H;�H;3�H;>�H;��H;Z�H;exH;�XH;�0H;F�G;�G;.hG;�F;":E;B;�;;u0;�Y;���:�q�:�;u9�{��"�D�@T��hs�VFB�}��������μo���e�	����+�K�3�      u�����W�Жռ ־�.Ϥ��I����[�
(��Z����9��{���<9vX�:�X�:[Q;Z,;��8;�A@;6BD;�@F;�,G;��G;��G;�H;EH;[hH;n�H;��H;��H;��H;]�H;[�H;�H;��H;��H;��H;�H;X�H;]�H;��H;��H;��H;l�H;XhH;	EH;�H;��G;��G;�,G;�@F;6BD;�A@;��8;],;[Q;�X�:zX�:�<9�{����9���Z�	(���[��I��.Ϥ� ־�Жռ�W���      my��Dݜ��A���I����s���P��%+������Ļ����6|���o��;u9tX�:,�:q;�);��6;��>;�PC;��E;'�F;�xG;d�G;�H;�1H;SXH;=wH;�H;R�H;?�H;��H;U�H;}�H;��H;#�H;��H;#�H;��H;~�H;T�H;��H;?�H;O�H;�H;=wH;PXH;�1H;�H;a�G;�xG;'�F;��E;�PC;��>;�6;�);q;,�:tX�:�;u9��o�5|�������Ļ����%+���P���s��I���A��Eݜ�      ZFB�A�>���4�Y�$�v��[�����ݎ�^A?�XӺ����44�9�q�:�X�:s;��';�=5;��=;.�B;QGE;z�F;�UG;Z�G;�G;�H;�HH;NjH;4�H;��H;��H;o�H;��H;�H;|�H;I�H;Z�H;�H;Z�H;I�H;{�H;�H;��H;o�H;��H;��H;4�H;KjH;�HH;�H;�G;V�G;�UG;w�F;NGE;.�B;��=;�=5;��';s;�X�:�q�:<4�9����ZӺ\A?��ݎ����[�v��Y�$���4�B�>�      �EֻM�ѻ��ĻnT���񕻴.o�̝.�+ܺ`�B����8\:�&�:���:ZQ;);�=5;;=;J#B;��D;vF; 7G;��G;��G;�H;�:H;N^H;�zH;6�H;��H;�H;F�H;�H;��H;X�H;��H;e�H;��H;e�H;��H;Y�H;��H;�H;F�H;��H;��H;6�H;�zH;O^H;�:H;�H;��G;��G;7G;vF;��D;M#B;;=;�=5;);ZQ;���:�&�:\:���8X�B�+̝ܺ.��.o���mT����ĻS�ѻ      �A?��9�9)��Z��ܺzp��H��� <9B�@:��:\�:t�	;�Y;W,;��6;��=;I#B;�D;�XF;"G;��G;U�G;�H;//H;�SH;�qH;�H;�H;��H;��H;��H;�H;��H;�H;��H;U�H;��H;T�H;��H;�H;��H;�H;��H;��H;��H;�H;�H;�qH;�SH;,/H;�H;U�G;��G;"G;�XF;�D;H#B;��=;��6;Z,;�Y;t�	;^�:��:N�@:�;9H���tp���ܺ�Z�9)��9�      ��	������i���Z���5u9�:k~:L��:�[�:��;��;~%;u0;��8;��>;.�B;��D;�XF;gG;��G;��G;��G;.&H;BKH;�iH;!�H;ƗH;u�H;��H;E�H;��H;��H;��H;m�H;��H;�H;��H;�H;��H;m�H;��H;��H;��H;B�H;��H;u�H;ėH;"�H;�iH;>KH;+&H;��G;��G;��G;gG;�XF;��D;.�B;��>;��8;u0;~%;��;��;�[�:J��:k~:�:06u9�Z���i��x���      �Y�:�o�:�W�:V�:U&�:���:���:T�	;/Q;�M#;�n-;u�5;�;;�A@;�PC;IGE;
vF; "G;��G;�G;P�G;� H;GEH;�cH;x}H;��H;�H;ޱH;�H;��H;��H;f�H;��H;��H;��H;��H;(�H;��H;��H;��H;��H;i�H;��H;��H;��H;ܱH;�H;��H;x}H;�cH;DEH;� H;M�G;
�G;��G;"G;
vF;JGE;�PC;�A@;�;;u�5;�n-;�M#;1Q;U�	;���:���:m&�:V�:�W�:vo�:      ���:N% ;n�; �;)�;Q;Cm;\d';�.;�=5;�:;��>;B;5BD;��E;w�F;7G;��G;��G;P�G;�H;$BH;F`H;�yH;��H;`�H;��H; �H;��H;�H;��H;l�H;��H;y�H;-�H;�H;��H;�H;-�H;y�H;��H;o�H;��H;
�H;��H;�H;��H;`�H;��H;�yH;C`H;$BH;�H;S�G;��G;��G;7G;w�F;��E;5BD;B;��>;�:;�=5;"�.;[d';Dm;Q;+�;�;l�;>% ;      ��";�M#;.%;z�';J�+;b�/;��3;� 8;�;;>?; �A;ԻC;":E;�@F;'�F;�UG;��G;V�G;��G;� H;"BH;�^H;�wH;X�H;ÝH;�H;̷H;j�H;<�H;c�H;[�H;%�H;��H;�H;��H;��H;��H;��H;��H;�H;��H;%�H;[�H;`�H;8�H;j�H;ɷH;�H;ĝH;T�H;�wH;�^H;!BH;� H;��G;X�G;��G;�UG;)�F;�@F;":E;ԻC;�A;??;�;;� 8;��3;c�/;`�+;z�';+%;�M#;      �46;��6;#l7;N�8;��:;q�<;S�>;s�@;�tB;��C;�,E;�F;�F;�,G;�xG;W�G;��G;�H;,&H;JEH;E`H;�wH;m�H;r�H;��H;'�H;׿H;��H;�H;9�H;g�H;{�H;��H;��H;��H;��H;��H;��H;��H;��H;��H;{�H;g�H;7�H;�H;��H;ԿH;(�H;��H;p�H;k�H;�wH;A`H;LEH;.&H;�H;��G;V�G;�xG;�,G;�F;�F;�,E;��C;�tB;s�@;S�>;s�<;��:;N�8;#l7;v�6;      }@;iA@;>�@;+RA;�"B;C;^�C;��D;>�E;�@F;��F;�!G;.hG;��G;a�G;�G;�H;//H;@KH;�cH;�yH;W�H;p�H;�H;C�H;��H;��H;�H;M�H;��H;��H;��H;x�H;��H;�H;��H;��H;��H;�H;��H;u�H;��H;��H;��H;K�H;�H;��H;��H;D�H;��H;o�H;V�H;�yH;�cH;AKH;2/H;�H;�G;a�G;��G;.hG;�!G;��F;�@F;?�E;��D;\�C;C;�"B;)RA;<�@;]A@;      ��D;%�D;�D;�9E;��E;Q�E;rPF;�F;��F;=:G;coG;ؚG;�G;��G;�H;�H;�:H;�SH;�iH;�}H;��H;ǝH;��H;L�H;w�H; �H;h�H;��H;��H;j�H;�H;D�H;��H;'�H;��H;[�H;��H;\�H;��H;$�H;��H;D�H;�H;i�H;��H;��H;i�H; �H;x�H;I�H;��H;ǝH;��H;�}H;�iH;�SH;�:H;�H;�H;��G;�G;ښG;aoG;<:G;��F;�F;rPF;P�E;��E;�9E;�D;%�D;      �F;�F;�F;��F;�F;�!G;�FG;XjG;c�G;(�G;*�G;�G;A�G;�H;�1H;�HH;M^H;�qH;�H;��H;]�H;�H;$�H;��H;�H;J�H;Z�H;��H;��H;��H;��H;��H;+�H;�H;��H;�H;G�H;�H;��H;�H;*�H;��H;��H;��H;��H;��H;[�H;L�H;�H;��H;$�H;�H;X�H;��H;�H;�qH;M^H;�HH;�1H;�H;A�G;�G;+�G;(�G;e�G;UjG;�FG;�!G;!�F;��F;�F;ٯF;      �nG;0qG;xG;�G;��G;\�G;{�G;��G;&�G;M�G;�H;|H;�0H;	EH;PXH;NjH;�zH;�H;ƗH;��H;��H;̷H;ֿH;��H;d�H;\�H;{�H;��H;��H;��H;��H;�H;�H;��H;o�H;��H;��H;��H;n�H;��H;�H;�H;��H;��H;��H;��H;{�H;\�H;g�H;��H;ԿH;̷H;��H;��H;ƗH;�H;�zH;NjH;QXH;	EH;�0H;|H;�H;M�G;)�G;��G;{�G;W�G;��G;�G;xG;/qG;      �G;�G;��G;�G;�G;5�G;'�G;�H;H;m'H;
8H;�HH;�XH;[hH;=wH;4�H;5�H;�H;r�H;�H;�H;j�H;��H;�H;��H;��H;��H;x�H;��H;��H;��H;��H;��H;��H;�H;>�H;Q�H;>�H;�H;��H;��H;�H;��H;}�H;��H;x�H;��H;��H;��H;�H;��H;i�H;�H;�H;r�H;�H;3�H;4�H;>wH;ZhH;�XH;�HH;
8H;m'H;H;�H;&�G;7�G;*�G;�G;��G;��G;      ZH;UH;zH;�H;qH;�%H;�/H;�:H;�FH;�RH;{_H;lH;gxH;n�H;�H;��H;��H;��H;��H;�H;��H;;�H;�H;R�H;��H;��H;��H;��H;^�H;��H;�H;��H;��H;�H;��H;��H;��H;��H;��H;�H;��H;��H;�H;��H;^�H;��H;��H;��H;��H;R�H;�H;;�H;��H;�H;��H;��H;��H;��H;�H;n�H;hxH;
lH;y_H;�RH;�FH;�:H;�/H;�%H;xH;�H;xH;JH;      I@H;AH;qCH;9GH;rLH;�RH;3ZH;ubH;]kH;�tH;D~H;�H;_�H;��H;S�H;��H;�H;�H;A�H;��H;�H;a�H;6�H;��H;a�H;��H;��H;�H;��H;�H;��H;��H;4�H;��H;��H;�H;�H;�H;��H;��H;3�H;��H;��H;�H;��H;�H;��H;��H;c�H;��H;4�H;a�H;�H;��H;A�H;��H;�H;��H;S�H;��H;_�H;�H;F~H;�tH;`kH;wbH;3ZH;�RH;oLH;7GH;mCH;AH;      "gH;�gH;piH;SlH;?pH;uH;�zH;��H;ŇH;�H;,�H;��H;��H;��H;A�H;v�H;K�H;��H;��H;��H;��H;]�H;j�H;��H;�H;��H;��H;��H;�H;��H;��H;A�H;��H;��H;�H;G�H;c�H;G�H;�H;��H;��H;C�H;��H;��H;�H;��H;��H;��H;�H;��H;e�H;[�H;��H;��H;��H;��H;J�H;u�H;A�H;��H;��H;��H;.�H;�H;ƇH;��H;�zH;	uH;<pH;TlH;piH;�gH;      ��H;�H;_�H;��H;��H;9�H;��H;L�H;a�H;��H;B�H;խH;A�H;��H;��H;��H;�H;�H;��H;p�H;t�H;*�H;~�H;��H;@�H;��H;�H;�H;��H;��H;?�H;��H;��H;9�H;b�H;��H;~�H;��H;b�H;;�H;��H;��H;A�H;��H;��H;�H;�H;��H;C�H;��H;|�H;*�H;s�H;p�H;��H;�H;�H;��H;��H;��H;A�H;ԭH;B�H;��H;b�H;I�H;��H;;�H;��H;��H;_�H;��H;      j�H;ϚH;ЛH;v�H;��H;|�H;��H;q�H;L�H;b�H;��H;�H;6�H;c�H;X�H;�H;��H;��H;��H;��H;��H;��H;��H;~�H;��H;-�H; �H;��H;��H;>�H;��H;��H;=�H;t�H;��H;��H;��H;��H;��H;t�H;;�H;��H;��H;>�H;��H;��H;�H;+�H;��H;�H;��H;��H;��H;��H;��H;��H;��H;�H;U�H;b�H;5�H;�H;��H;c�H;L�H;p�H;��H;�H;��H;v�H;ЛH;ȚH;      ԩH;$�H;֪H;#�H;�H;�H;��H;��H;��H;�H;P�H;��H; �H;_�H;��H;��H;_�H;	�H;q�H;��H;��H;�H;��H;��H;�H;�H;��H;��H;�H;��H;��H;9�H;m�H;��H;��H;��H;��H;��H;��H;��H;m�H;<�H;��H;��H;�H;��H;��H;�H; �H;��H;��H;�H;��H;��H;q�H;�H;]�H;��H;��H;_�H; �H;��H;O�H;�H;��H;��H;��H;�H;ۭH;#�H;تH;�H;      �H;e�H;��H;�H;��H;=�H;c�H;ǽH;O�H;��H;��H;��H;S�H; �H;��H;R�H;��H;��H;��H;��H;8�H;��H;��H;	�H;��H;��H;m�H;�H;��H;��H;�H;f�H;��H;��H;��H;��H;��H;��H;��H;��H;��H;h�H;�H;��H;��H;�H;k�H;��H;��H;	�H;��H;��H;5�H;��H;��H;��H;��H;R�H;��H; �H;S�H;��H;��H;��H;P�H;ĽH;c�H;B�H;��H;�H; �H;]�H;      ��H;5�H;ӺH;̻H;�H;��H;i�H;z�H;��H;�H;}�H;��H;j�H;��H;(�H;a�H;n�H;Q�H;�H;��H;'�H;��H;��H;��H;V�H;�H;��H;?�H;��H;�H;G�H;��H;��H;��H;��H;��H;��H;��H;��H;��H;��H;��H;G�H;�H;��H;?�H;��H;�H;X�H;��H;��H;��H;%�H;��H;�H;S�H;m�H;a�H;(�H;��H;k�H;��H;{�H;�H;��H;x�H;i�H;��H;�H;̻H;ֺH;,�H;      ��H;�H;��H;��H;˾H;<�H;�H;�H;9�H;}�H;��H;$�H;v�H;��H;��H;�H;��H;��H;��H;1�H;��H;��H;��H;��H;��H;B�H;��H;W�H;��H;�H;f�H;��H;��H;��H;��H;��H;��H;��H;��H;��H;��H;��H;f�H;�H;��H;W�H;��H;D�H;��H;��H;��H;��H;��H;1�H;��H;��H;��H;�H;��H;��H;v�H;$�H;��H;��H;:�H;�H;�H;A�H;��H;��H;��H;�H;      ��H;5�H;ӺH;̻H;�H;��H;i�H;z�H;��H;�H;}�H;��H;k�H;��H;(�H;a�H;n�H;Q�H;�H;��H;(�H;��H;��H;��H;X�H;�H;��H;?�H;��H;�H;G�H;��H;��H;��H;��H;��H;��H;��H;��H;��H;��H;��H;G�H;�H;��H;?�H;��H;�H;V�H;��H;��H;��H;%�H;��H;�H;S�H;m�H;a�H;(�H;��H;j�H;��H;}�H;
�H;��H;w�H;i�H;��H;�H;̻H;ҺH;)�H;      �H;e�H;��H;�H;��H;=�H;c�H;ɽH;O�H;��H;��H;��H;S�H; �H;��H;R�H;��H;��H;��H;��H;9�H;��H;��H;�H;��H;��H;m�H;�H;��H;��H;�H;e�H;��H;��H;��H;��H;��H;��H;��H;��H;��H;j�H;�H;��H;��H;�H;k�H;��H;��H;�H;��H;��H;5�H;��H;��H;��H;��H;R�H;��H; �H;S�H;��H;��H;��H;O�H;ĽH;d�H;B�H;��H;�H;��H;]�H;      թH;$�H;֪H;#�H;�H;�H;��H;��H;��H;�H;P�H;��H; �H;_�H;��H;��H;_�H;	�H;q�H;��H;��H;�H;��H;��H; �H;�H;��H;��H;�H;��H;��H;9�H;o�H;��H;��H;��H;��H;��H;��H;��H;l�H;<�H;��H;��H;�H;��H;��H;�H;�H;��H;��H;�H;��H;��H;q�H;�H;]�H;��H;��H;_�H; �H;��H;P�H;�H;��H;��H;��H;�H;٭H;#�H;تH;�H;      m�H;ϚH;қH;w�H;��H;|�H;��H;p�H;L�H;b�H;��H;�H;5�H;c�H;V�H;�H;��H;��H;��H;��H;��H;��H;��H;�H;��H;-�H; �H;��H;��H;<�H;��H;��H;<�H;s�H;��H;��H;��H;��H;��H;s�H;;�H;��H;��H;>�H;��H;��H;�H;+�H;��H;|�H;��H;��H;��H;��H;��H;��H;��H;�H;X�H;b�H;5�H;�H;��H;c�H;L�H;m�H;��H;��H;��H;w�H;ϛH;̚H;      ��H;�H;_�H;��H;��H;9�H;��H;J�H;a�H;��H;B�H;խH;A�H;��H;��H;��H;�H;�H;��H;q�H;w�H;*�H;~�H;��H;C�H;��H;�H;�H;��H;��H;A�H;��H;��H;;�H;b�H;��H;~�H;��H;b�H;9�H;��H;��H;?�H;��H;��H;�H;�H;��H;@�H;��H;|�H;*�H;s�H;p�H;��H;�H;�H;��H;��H;��H;@�H;ԭH;B�H;��H;b�H;H�H;��H;:�H;}�H;��H;`�H;��H;      "gH;�gH;oiH;TlH;?pH;uH;�zH;��H;ŇH;�H;.�H;��H;��H;��H;A�H;v�H;J�H;��H;��H;��H;��H;[�H;j�H;��H;�H;��H;��H;��H;�H;��H;��H;B�H;��H;��H;�H;G�H;c�H;G�H;�H;��H;��H;B�H;��H;��H;�H;��H;��H;��H;�H;��H;g�H;]�H;��H;��H;��H;��H;J�H;v�H;A�H;��H;��H;��H;+�H;�H;ŇH;��H;�zH;	uH;<pH;SlH;piH;�gH;      C@H;AH;oCH;9GH;nLH;�RH;6ZH;wbH;^kH;�tH;D~H;�H;^�H;��H;S�H;��H;�H;�H;A�H;��H;�H;a�H;6�H;��H;c�H;��H;��H;�H;��H;�H;��H;��H;4�H;��H;��H;�H;�H;�H;��H;��H;3�H;��H;��H;�H;��H;�H;��H;��H;a�H;��H;4�H;a�H;�H;��H;A�H;��H;�H;��H;S�H;��H;_�H;�H;D~H;�tH;`kH;wbH;6ZH;�RH;lLH;9GH;oCH;AH;      QH;QH;H;�H;wH;�%H;�/H;�:H;�FH;�RH;{_H;lH;gxH;n�H;�H;��H;��H;��H;��H;�H;��H;;�H;�H;R�H;��H; �H;��H;��H;^�H;��H;�H;��H;��H;�H;~�H;��H;��H;��H;��H;�H;��H;��H;�H;��H;^�H;��H;��H;��H;��H;R�H;�H;;�H;��H;�H;��H;��H;��H;��H;�H;n�H;gxH;lH;|_H;�RH;�FH;�:H;�/H;�%H;sH;�H;}H;OH;      �G;��G;��G;�G;�G;7�G;&�G;�H;H;m'H;8H;�HH;�XH;[hH;>wH;4�H;5�H;�H;r�H;�H;!�H;i�H;��H;�H;��H;��H;��H;x�H;��H;��H;��H;�H;��H;��H;�H;>�H;Q�H;>�H;�H;��H;��H;�H;��H;}�H;��H;x�H;��H;��H;��H;�H;��H;j�H;�H;�H;r�H;�H;3�H;5�H;=wH;XhH;�XH;�HH;8H;m'H;H;�H;'�G;3�G;)�G;�G;��G;��G;      �nG;0qG;xG;܂G;��G;V�G;y�G;��G;&�G;O�G;�H;|H;�0H;	EH;QXH;OjH;�zH;�H;ƗH;��H;��H;̷H;ֿH;��H;g�H;^�H;}�H;��H;��H;��H;��H;�H;�H;��H;n�H;��H;��H;��H;o�H;��H;�H;�H;��H;��H;��H;��H;z�H;\�H;d�H;��H;ԿH;̷H;��H;��H;ƗH;�H;�zH;MjH;PXH;	EH;�0H;|H;�H;M�G;&�G;��G;y�G;W�G;��G;܂G;xG;%qG;      �F;ۯF;�F;��F;�F;�!G;�FG;VjG;c�G;)�G;+�G;	�G;A�G;�H;�1H;�HH;N^H;�qH;�H;��H;^�H;�H;$�H;��H;�H;L�H;[�H;��H;��H;��H;��H;��H;+�H;�H;��H;�H;G�H;�H;��H;�H;(�H;��H;��H;��H;��H;��H;Z�H;J�H;�H;��H;$�H;�H;X�H;��H;�H;�qH;K^H;�HH;�1H;�H;A�G;�G;+�G;(�G;c�G;VjG;�FG;�!G; �F;��F;�F;ԯF;      ��D;%�D;�D;�9E;��E;Q�E;rPF;�F;��F;=:G;coG;ښG;�G;��G;�H;�H;�:H;�SH;�iH;�}H;ÎH;ǝH;��H;L�H;x�H; �H;k�H;��H;��H;j�H;�H;C�H;��H;$�H;��H;\�H;��H;[�H;��H;&�H;��H;G�H;�H;i�H;��H;��H;h�H; �H;w�H;J�H;��H;ǝH;��H;�}H;�iH;�SH;�:H;�H;�H;��G;�G;ؚG;coG;<:G;��F;�F;rPF;Q�E;��E;�9E;�D;&�D;      �@;dA@;A�@;'RA;�"B;C;[�C;��D;?�E;�@F;��F;�!G;0hG;��G;a�G;�G;�H;//H;AKH;�cH;�yH;V�H;p�H;�H;D�H;��H;��H;�H;N�H;��H;��H;��H;w�H;��H;�H;��H;��H;��H;�H;��H;w�H;��H;��H;��H;J�H;�H;��H;��H;C�H;��H;o�H;W�H;�yH;�cH;@KH;0/H;�H;�G;a�G;��G;-hG;�!G;��F;�@F;?�E;��D;[�C;C;�"B;(RA;?�@;[A@;      �46;��6;1l7;N�8;��:;t�<;W�>;s�@;�tB;��C;�,E;�F;�F;�,G;�xG;W�G;��G;�H;.&H;JEH;F`H;�wH;m�H;r�H;��H;'�H;׿H;��H;�H;:�H;g�H;{�H;��H;��H;��H;��H;��H;��H;��H;��H;��H;{�H;g�H;6�H;�H;��H;ԿH;(�H;��H;p�H;k�H;�wH;B`H;LEH;,&H;�H;��G;W�G;�xG;�,G;�F;�F;�,E;�C;�tB;s�@;W�>;v�<;��:;N�8;(l7;}�6;      ��";�M#;/%;z�';J�+;b�/;��3;� 8;�;;??; �A;ԻC;":E;�@F;'�F;�UG;��G;U�G;��G;� H;$BH;�^H;�wH;X�H;ĝH;�H;̷H;j�H;<�H;d�H;[�H;%�H;��H;�H;��H;��H;��H;��H;��H;�H;��H;%�H;[�H;^�H;8�H;j�H;ɷH;�H;ÝH;W�H;�wH;�^H;"BH;� H;��G;X�G;��G;�UG;)�F;�@F;":E;ջC;�A;>?;�;;� 8;��3;b�/;^�+;z�';-%;�M#;      ���:H% ;r�;�;)�;Q;Hm;_d';�.;�=5;�:;��>;B;5BD;��E;w�F;7G;��G;��G;Q�G;�H;$BH;E`H;�yH;��H;`�H;��H;�H;��H;�H;��H;m�H;��H;x�H;-�H;�H;��H;�H;-�H;y�H;��H;m�H;��H;	�H;��H; �H;��H;`�H;��H;�yH;E`H;$BH;�H;Q�G;��G;��G;7G;w�F;��E;5BD;B;��>;�:;�=5;!�.;]d';Gm;Q;.�;�;p�;?% ;      �Y�:�o�:�W�:R�:]&�:���:���:U�	;1Q;�M#;�n-;u�5;�;;�A@;�PC;JGE;
vF; "G;��G;�G;Q�G;� H;GEH;�cH;x}H;��H;�H;ܱH;�H;��H;��H;g�H;��H;��H;��H;��H;(�H;��H;��H;��H;��H;g�H;��H;��H;��H;ޱH;�H;��H;x}H;�cH;DEH;� H;M�G;
�G;��G;"G;
vF;IGE;�PC;�A@;�;;s�5;�n-;�M#;1Q;U�	;���:���:g&�:P�:�W�:vo�:      ��	������i���Z���5u9�:k~:L��:�[�:��;��;~%;u0;��8;��>;.�B;��D;�XF;gG;��G;��G;��G;/&H;BKH;�iH;!�H;ƗH;u�H;��H;E�H;��H;��H;��H;m�H;��H;�H;��H;�H;��H;m�H;��H;��H;��H;B�H;��H;u�H;ėH;"�H;�iH;>KH;)&H;��G;��G;��G;gG;�XF;��D;.�B;��>;��8;u0;~%;��;��;�[�:J��:k~:�: 6u9�Z���i������      �A?��9�9)��Z��ܺ�p��H����;9B�@:��:^�:t�	;�Y;Y,;��6;��=;I#B;��D;�XF;"G;��G;U�G;�H;0/H;�SH;�qH;�H;�H;��H;��H;��H;�H;��H;�H;��H;T�H;��H;U�H;��H;�H;��H;�H;��H;��H;��H;�H;�H;�qH;�SH;*/H;�H;U�G;��G;"G;�XF;�D;H#B;��=;��6;W,;�Y;t�	;\�:��:N�@:�;9H���tp���ܺ�Z�9)��9�      �EֻN�ѻ��ĻnT���񕻶.o�̝.�)ܺ`�B����8\:�&�:���:[Q;);�=5;;=;J#B;��D;vF; 7G;��G;��G;�H;�:H;N^H;�zH;6�H;��H;�H;F�H;�H;��H;Y�H;��H;e�H;��H;e�H;��H;Y�H;��H;�H;F�H; �H;��H;6�H;�zH;O^H;�:H;�H;��G;��G;7G;vF;��D;M#B;;=;�=5;);ZQ;���:�&�:\:���8X�B�-̝ܺ.��.o���nT����ĻS�ѻ      [FB�@�>���4�Y�$�v��[�����ݎ�^A?�XӺ����<4�9�q�:�X�:s;��';�=5;��=;.�B;NGE;x�F;�UG;X�G;�G;�H;�HH;NjH;4�H;��H;��H;o�H;��H;�H;{�H;I�H;Z�H;�H;Z�H;I�H;|�H;�H;��H;o�H;��H;��H;4�H;KjH;�HH;�H;�G;V�G;�UG;x�F;NGE;.�B;��=;�=5;��';s;�X�:�q�:44�9����ZӺ\A?��ݎ����[�v��Y�$���4�C�>�      my��Dݜ��A���I����s���P��%+������Ļ����6|���o��;u9tX�:,�:q;�);��6;��>;�PC;��E;'�F;�xG;d�G;�H;�1H;QXH;=wH;�H;R�H;?�H;��H;V�H;~�H;��H;#�H;��H;#�H;��H;~�H;U�H;��H;?�H;O�H;�H;=wH;QXH;�1H;�H;a�G;�xG;'�F;��E;�PC;��>;�6;�);q;,�:tX�:�;u9��o�6|�������Ļ����%+���P���s��I���A��Eݜ�      u�����W�Жռ ־�.Ϥ��I����[�
(��Z����9��{���<9zX�:�X�:\Q;\,;��8;�A@;5BD;�@F;�,G;��G;��G;�H;EH;XhH;n�H;��H;��H;��H;_�H;Z�H;�H;��H;��H;��H;�H;Z�H;\�H;��H;��H;��H;n�H;[hH;	EH;�H;��G;��G;�,G;�@F;6BD;�A@;��8;],;ZQ;�X�:xX�:�<9�{����9���Z�
(���[��I��.Ϥ� ־�Жռ�W���      6�6�K�3���+�	��e�o�����μ���}���VFB�hs�@T��"�D��{���;u9�q�:���:�Y;u0;�;;B;":E;�F;2hG;�G;C�G;�0H;�XH;gxH;Z�H;��H;=�H;3�H;�H;N�H;f�H;t�H;g�H;N�H;�H;2�H;=�H;��H;[�H;gxH;�XH;�0H;G�G;�G;-hG;�F;":E;B;�;;u0;�Y;���:�q�:�;u9�{��#�D�AT��hs�VFB�}��������μo���e�	����+�K�3�      s₽�؀���u��Xc���K�|1�������վ��]����P����@T����9���o�<4�9�&�:v�	;}%;v�5;��>;һC;�F;�!G;՚G;	�G;yH;�HH;lH;ׇH;��H;˭H;�H;��H;��H;��H;�H;��H;��H;��H;�H;έH;��H;هH;lH;�HH;xH;�G;ؚG;�!G;�F;һC;��>;v�5;}%;w�	;�&�:,4�9��o���9�@T�������P��]���վ�����|1���K��Xc���u��؀�      <S���r��t�����ԓ����u���N���(��i�Ό˼�A����P�hs��4|�����\:^�:��;�n-;�:;�A;�,E;��F;coG;-�G;�H;8H;|_H;=~H;(�H;<�H;��H;I�H;��H;t�H;��H;t�H;��H;K�H;��H;?�H;)�H;=~H;y_H;8H;�H;.�G;doG;��F;�,E;�A;�:;�n-;��;`�:�\:����5|��hs���P��A��Ό˼�i���(���N���u�ԓ�����t���r��      �o��s��置�ս9@��tĥ�{^���Xc�G�3���	�Ό˼�]��VFB��Z򻬜��XӺ���8��:��;�M#;�=5;;?;��C;�@F;<:G;)�G;O�G;k'H;�RH;�tH;�H;��H;b�H;�H;��H;�H;}�H;	�H;��H;�H;a�H;��H;�H;�tH;�RH;k'H;M�G;+�G;@:G;�@F;��C;;?;�=5;�M#;��;��:���8ZӺ�����Z�VFB��]��Ό˼��	�G�3��Xc�{^��tĥ�9@����ս���s�      �#�X� �b'������gٽ:S��+l��T�j�G�3��i��վ�}���
(���Ļ]A?�T�B�J�@:�[�:5Q;�.;�;;�tB;>�E;��F;f�G;'�G;H;�FH;UkH;��H;\�H;G�H;��H;H�H;��H;0�H;��H;H�H;��H;D�H;^�H;��H;UkH;�FH;H;%�G;f�G;��F;;�E;�tB;�;;"�.;4Q;�[�:N�@:`�B�\A?���Ļ
(�}����վ��i�G�3�T�j�+l��:S���gٽ����b'�X� �      �S�*�O��E��5�X� �Z�
���罨9��*l���Xc���(��������[�����ݎ�(ܺ0<9R��:X�	;[d';� 8;r�@;��D;�F;XjG;��G;�H;�:H;nbH;�H;C�H;i�H;�H;��H;p�H;�H;q�H;��H;��H;h�H;E�H;�H;nbH;�:H;�H;��G;VjG;�F;��D;r�@;� 8;]d';W�	;R��:@<9-ܺ�ݎ������[��������(��Xc�*l���9�����Z�
�X� ��5��E�*�O�      �~��*��,�v��9b�~�H�#,�OZ����:S��z^����N������μ�I���%+����Н.�0���k~:���:?m;��3;O�>;X�C;rPF;�FG;u�G;!�G;�/H;/ZH;�zH;��H;��H;��H;\�H;a�H;�H;a�H;\�H;��H;��H;��H;�zH;.ZH;�/H;!�G;t�G;�FG;uPF;T�C;O�>;��3;Cm;���:k~:(���ҝ.�����%+��I����μ�����N�z^��:S�����OZ�#,�~�H��9b�,�v�*��      ����+����:���M��H�r�*�O�#,�Z�
��gٽtĥ���u�|1�o���.Ϥ���P�[�.o�`p���:���:Q;X�/;o�<;C;L�E;�!G;U�G;5�G;�%H;�RH;uH;6�H;|�H;�H;?�H;��H;<�H;��H;?�H;�H;{�H;9�H;uH;�RH;�%H;5�G;S�G;�!G;M�E;C;p�<;Y�/;Q;���:�:^p���.o�[򻯎P�.Ϥ�o���|1���u�tĥ��gٽZ�
�#,�*�O�I�r��M���:��+���      :���v��O;������UP��I�r�~�H�X� ���8@��ԓ����K�d� ־���s�u���񕻗ܺ 6u9Y&�:+�;H�+;��:;�"B;��E;�F;�G;�G;sH;bLH;3pH;|�H;��H;٭H;r�H;�H;��H;�H;q�H;ۭH;��H;�H;3pH;`LH;pH;�G;��G;�F;��E;�"B;��:;H�+;.�;Y&�:�5u9�ܺ��u����s� ־�d���K�ԓ��8@����X� �~�H�I�r�UP������O;���v��      XVھ�*־25ʾu��������M���9b��5�����ս����Xc�	��Жռ�I��X�$�jT���Z��Z��V�:�;��';X�8;.RA;�9E;��F;݂G; �G;�H;4GH;JlH;��H;o�H;�H;��H;ɻH;��H;ɻH;��H;�H;m�H;��H;IlH;2GH;�H;!�G;݂G;��F;�9E;)RA;[�8;��';�;T�:�Z���Z�lT��X�$��I��Жռ	���Xc������ս���5��9b��M������u���25ʾ�*־      ���쾶�޾25ʾO;���:��,�v��E�b'����t����u���+��W��A����4���Ļ9)� j���W�:f�;%;!l7;5�@; �D;�F;xG;��G;xH;hCH;biH;Q�H;țH;٪H;��H;ʺH;��H;ʺH;��H;٪H;śH;Q�H;biH;eCH;vH;��G;xG;�F; �D;0�@;#l7;%;h�;�W�: j��9)���Ļ��4��A���W缇�+���u�t�����b'��E�,�v��:��O;��25ʾ��޾��      Zh���b���쾪*־�v��+���*��*�O�X� �s��r���؀�K�3���Cݜ�@�>�R�ѻ�9�h���jo�:A% ;�M#;}�6;[A@;�D;ԯF;,qG;|�G;UH;AH;�gH;�H;ĚH;�H;P�H;,�H;�H;,�H;Q�H;�H;ÚH;�H;�gH;AH;RH;|�G;+qG;ԯF;�D;XA@;��6;�M#;A% ;ho�:h���ޡ9�R�ѻ@�>�Dݜ���K�3��؀��r��s�X� �*�O�*��+����v���*־���b��      3�$��� ����%��D��*�þ�*��6Dx���=�����Pν	���''K��c�"��s�V����E^�`�S� x[:���:&e;g�4;R`?;�mD;��F;avG;J�G;�H;�OH;�sH;�H;��H;��H;,�H;��H;[�H;��H;+�H;��H;��H;��H;�sH;�OH;�H;J�G;`vG;��F;�mD;O`?;j�4;&e;���:x[:`�S�E^����t�V�#���c�''K�	����Pν�����=�6Dx��*��*�þD��%������� �      �� ����T��P��2��
����0��8�s�ڀ:�i9� �ʽ4Z���G��8�.���5S�����/X�@�D�Cd:�B�: ;/�4;ֈ?;D;Z�F;$yG;��G;� H;SPH;OtH;H�H;�H;�H;i�H;��H;l�H;��H;j�H;�H;��H;I�H;OtH;PPH;� H;��G;$yG;\�F;D;ш?;4�4; ;�B�:Cd:@�D��/X���껱5S�.���8��G�4Z�� �ʽi9�ڀ:�8�s��0��
���2��P��T�����      ���T��;�
������Yؾ"���॒���f���0�\[�R8��Ґ����>�����NȤ��6H�`�ܻrF������}: ��:z";i�5;�?;��D;�F; �G;��G;x#H;�RH;�uH;��H;��H;��H;�H;&�H;��H;&�H;�H;��H;��H;��H;�uH;�RH;u#H;��G; �G;�F;��D;�?;l�5;z"; ��:��}:���rF�a�ܻ�6H�NȤ�������>�Ґ��R8��\[���0���f�॒�"����Yؾ����:�
�T��      %��P������AI�*�þ�R��=���xS��Q"��s������}��0��켋�����6�E�ƻ3}*�����'�:�x;o%;m7;�@;��D;�F;��G;��G;:(H;VH;�xH;��H;{�H;ٲH;�H;��H;��H;��H;�H;ٲH;z�H;��H;�xH;VH;7(H;��G;��G;�F;��D;�@;m7;o%;�x;%�:����2}*�F�ƻ��6��������0���}�����s��Q"�xS�=����R��*�þAIᾦ���P��      C��2�很Yؾ*�þĪ�~쏾�k�ڀ:���~�ؽ�����c�`y���Ҽ ���E� �f�%�� 2(7��:��
;�(;�_9;ɘA;�\E;��F;ڝG;��G;�.H;�ZH;#|H;*�H;�H;��H;I�H;�H;��H;�H;G�H;��H;|�H;-�H;#|H;�ZH;�.H;��G;۝G;��F;�\E;ĘA;�_9;�(;��
;��: 2(7$��g�E� � �����Ҽ`y��c�����~�ؽ��ڀ:��k�~쏾Ī�*�þ�Yؾ2��      *�þ
���"����R��~쏾9�s��H�����������ѐ����D��c�����B�f�U,�����P����9��:�;?j-;��;;��B;�E;�G;��G;��G;�6H;�`H;��H;��H;	�H;��H;ݾH;��H;�H;��H;ݾH;��H;�H;��H;��H;�`H;�6H;��G;��G;�G;�E;��B;��;;?j-;�;��:��9�P�����U,�A�f������c���D�ѐ�������������H�8�s�~쏾�R��"���
���      �*���0��॒�=����k��H��#%�\[��Pν
t��e�f�6/%���伈���x�=��?ػ�FL���D���R:H�:E�;S2;��=;ךC;�0F;�GG;��G;YH;@H;�gH;��H;i�H;�H;θH;��H;(�H;��H;(�H;��H;͸H;�H;k�H;��H;�gH;@H;VH;��G;�GG;�0F;ӚC;��=;R2;F�;@�:��R:x�D��FL��?ػx�=��������6/%�e�f�
t���Pν\[��#%��H��k�=���॒��0��      6Dx�8�s���f�xS�ڀ:����\[��7ս�榽��}���;��8�X�����r����9G������ˬ�R��:5�;�}$;�6;5�?;�D;��F;�pG;��G;H;`JH;moH;v�H;��H;4�H;r�H;��H;��H;a�H;��H;��H;r�H;3�H;��H;v�H;moH;_JH;H;��G;�pG;��F;�D;5�?;�6;�}$;4�;T��:@ˬ����9G�������r�X����8���;���}��榽�7ս\[����ڀ:�xS���f�8�s�      ��=�ڀ:���0��Q"��������Pν�榽B�� �G�4����Ҽ ��LE:�>�ܻ�D^������i:v��:�;Q|,;ԡ:;��A;diE;��F;X�G;��G;�(H;qUH;�wH;��H;a�H;ɳH;.�H;�H;��H;M�H;��H;�H;.�H;ɳH;b�H;��H;�wH;oUH;�(H;��G;Z�G;��F;aiE;��A;ԡ:;S|,;�;x��:�i:�����D^�=�ܻKE:� ����Ҽ4�� �G�B���榽�Pν�������Q"���0�ڀ:�      ���j9�][��s��ؽ���t����}� �G������3c��Z�V�G,��*����������:N��:| ;��3;�0>;��C;F;9G;k�G;�H;&8H;�`H;7�H;'�H;5�H;�H;$�H;��H;�H;M�H;�H;��H;$�H;}�H;6�H;'�H;7�H;�`H;%8H;�H;m�G;9G;F;��C;�0>;��3;{ ;N��:��:�������*��G,�Z�V�3c������� �G���}�t������ؽ�s�][�j9�      �Pν �ʽR8���������ѐ��e�f���;�5�����FȤ�8�f�+��Mߵ�No5���D���-:q��:�>;�+;�_9;�A;��D;K�F;�vG;�G;OH;�GH;�lH;�H;ΞH;0�H;c�H;0�H;��H;=�H;`�H;<�H;��H;0�H;a�H;3�H;ΞH;�H;�lH;�GH;LH;�G;�vG;G�F;��D;�A;�_9;�+;�>;u��:��-:��D�No5�Lߵ�+��7�f�FȤ����5����;�e�f�ѐ���������R8�� �ʽ      	���4Z��Ґ����}��c���D�6/%��8���Ҽ2c��7�f�����ƻx/X�@���(��9:�:T�;�";��3;`>;mYC;��E;G;$�G;��G;�,H;;WH;LxH;��H;l�H;#�H;I�H;(�H;l�H;{�H;k�H;{�H;n�H;&�H;I�H;&�H;l�H;��H;JxH;;WH;�,H;��G;!�G;G;��E;mYC;`>;��3;�";W�;6�:(��9@���x/X��ƻ���7�f�2c����Ҽ�8�6/%���D��c���}�Ґ��4Z��      ('K��G���>��0�ay��c����X��� ��Z�V�+���ƻ�od�n�º �(7�4�:���:��;Q.;�:;8zA;Z�D;��F;~nG;t�G;*H;�@H;\fH;��H;d�H;�H;�H;#�H;'�H;��H;��H;t�H;��H;��H;'�H;!�H;�H;�H;d�H;��H;\fH;�@H;*H;p�G;znG;��F;Z�D;8zA;�:;Q.;¡;���:�4�: �(7n�º�od��ƻ*��Z�V� ��X�����优c�ay��0���>��G�      �c��8���������Ҽ����������r�KE:�F,�Lߵ�v/X�l�º Ŭ���}:5�:;c�);Jm7;@�?;��C;5F;�)G;B�G;��G;=*H;�SH;�tH;��H;��H;,�H;�H;��H;�H;J�H;��H;��H;��H;J�H;�H;��H;�H;,�H;��H;��H;�tH;�SH;@*H;�G;A�G;�)G;5F;��C;?�?;Jm7;f�);
;5�:��}:�Ĭ�l�ºv/X�Lߵ�F,�KE:���r�����������Ҽ�켼����8�      "��.��NȤ��������B�f�y�=����?�ܻ�*��Po5�D��� �(7��}:�n�:E�;�>&;��4;�=;��B;�E;C�F;ȁG;&�G;hH;�AH;�eH;w�H;�H;��H;�H;��H;[�H;��H;��H;��H;��H;��H;��H;��H;Y�H;��H;�H;��H;�H;w�H;�eH;�AH;gH;$�G;ÁG;C�F;�E;��B;�=;��4;�>&;E�;�n�:��}: �(7D���Po5��*��>�ܻ���y�=�B�f��������NȤ�.��      s�V��5S��6H���6�F� �V,��?ػ;G���D^������D� ��9�4�:/�:G�;%;��3;;�<;~B;�E;/�F;�XG;8�G;} H;�0H;�WH;�vH;*�H;��H;��H;ͽH;�H;��H;��H;��H;��H;u�H;��H;��H;��H;��H;�H;ͽH;��H;��H;*�H;�vH;�WH;�0H;y H;5�G;�XG;,�F;�E;~B;=�<;��3;%;G�;3�:�4�: ��9��D�����D^�;G���?ػU,�F� ���6��6H��5S�      ��ﻬ��b�ܻH�ƻh󩻶��{FL�������������-:8�:���:
;�>&;��3;x9<;6�A;�D;xZF;Q5G;/�G;�G;�!H;kJH;kkH;ޅH;��H;��H;׸H;%�H;��H;��H;�H;��H;��H;.�H;��H;��H;�H;��H;��H;%�H;ָH;��H;��H;مH;mkH;kJH;�!H;�G;/�G;P5G;xZF;�D;9�A;z9<;��3;�>&;
;���:8�:��-:����������{FL����g�H�ƻb�ܻ���      E^� 0X�rF�2}*�*���P����D��ˬ��i:��:s��:Q�;��;`�);��4;8�<;5�A;I�D;�9F;G;��G;y�G;uH;S?H;�aH;M}H;��H;��H;ԳH;�H;��H;��H;��H;V�H;��H;]�H;��H;]�H;��H;V�H;��H;��H;��H;�H;ҳH;��H;��H;P}H;�aH;O?H;rH;y�G;��G;G;�9F;K�D;3�A;8�<;��4;c�);��;S�;s��:��:�i: ̬���D��P��$��2}*�rF�0X�      T�S�P�D�d������ .(7��9ƍR:N��:t��:J��:�>;�";Q.;Im7;�=;|B;�D;�9F;NG;Q�G;��G;�H;�6H;�YH;vH;Z�H;*�H;:�H;=�H;��H;]�H;��H;T�H;q�H;��H;��H;/�H;��H;��H;q�H;R�H;��H;^�H;��H;:�H;9�H;'�H;\�H;vH;�YH;�6H;�H;��G;R�G;NG;�9F;�D;|B;�=;Im7;Q.;�";�>;J��:z��:L��:ʍR:(�9 4(7����d��L�D�      $x[:DCd:��}:%�:��:��:>�:0�;�;| ;�+;��3;��:;8�?;��B;�E;rZF;�G;M�G;��G;wH;�1H;TH;�pH;�H;��H;"�H;��H;��H;��H;:�H;�H;��H;\�H;1�H;O�H;��H;Q�H;1�H;\�H;��H;�H;:�H;��H;��H;��H;�H;��H;�H;�pH;TH;�1H;tH;��G;M�G; G;rZF;�E;��B;8�?;��:;��3;�+;{ ;�;1�;>�:��:��:'�:��}:$Cd:       ��:�B�:��:x;��
;�;G�;�}$;P|,;��3;�_9;^>;6zA;��C;�E;,�F;N5G;��G;��G;xH;�/H;+QH;=mH;��H;ٗH;ϧH;��H;7�H;��H;R�H;��H;��H;��H;�H;��H;��H;��H;�H;��H;�H;��H;��H;��H;O�H;��H;7�H;��H;ϧH;ٗH;��H;<mH;+QH;�/H;zH;��G;��G;M5G;,�F;�E;��C;6zA;\>;�_9;��3;S|,;�}$;I�;�;��
;�x;��:�B�:      .e;7 ;�";h%;
�(;Gj-;]2;�6;֡:;�0>;�A;nYC;Z�D;4F;E�F;�XG;-�G;y�G;�H;�1H;+QH;lH;��H;��H;s�H;j�H;�H;��H;��H;J�H;��H;�H;��H;��H;��H;��H;��H;��H;��H;��H;��H;�H;��H;F�H;��H;��H;�H;k�H;t�H;��H;��H;lH;*QH;�1H;�H;{�G;,�G;�XG;F�F;4F;Z�D;nYC;�A;�0>;ء:;�6;\2;Jj-;�(;i%;�";2 ;      m�4;6�4;l�5;m7;�_9;��;;��=;8�?;��A;��C;��D;��E;��F;�)G;ƁG;5�G;�G;sH;�6H;TH;<mH;��H;�H;F�H;��H;��H;b�H;n�H;�H;��H;S�H;'�H;p�H;��H;��H;��H;��H;��H;��H;��H;m�H;&�H;S�H;��H;�H;o�H;a�H;��H;��H;C�H;�H;��H;8mH;TH;�6H;uH;�G;4�G;ƁG;�)G;��F;��E;��D;��C;��A;5�?;��=;��;;�_9;m7;m�5;(�4;      f`?;�?;�?;�@;˘A;��B;ޚC;�D;diE;F;I�F;G;znG;C�G;$�G;y H;�!H;R?H;�YH;�pH;��H;��H;E�H;��H;ʺH;g�H;��H;C�H;��H;��H;��H;��H;��H;�H;��H;q�H;��H;p�H;��H;	�H;��H;��H;��H;��H;��H;C�H;��H;e�H;̺H;~�H;C�H;��H;��H;�pH;�YH;S?H;�!H;y H;%�G;C�G;znG;G;I�F;F;eiE;�D;ۚC;��B;ҘA;�@;�?;؈?;      �mD;	D;v�D;�D;�\E;�E;�0F;��F;��F;9G;�vG;$�G;t�G;��G;jH;�0H;qJH;�aH;!vH;�H;ۗH;w�H;��H;ҺH;)�H;�H;��H;O�H;#�H;4�H;��H;y�H;��H;�H;��H;!�H;d�H;�H;��H;�H;��H;|�H;��H;3�H;"�H;O�H;��H;�H;*�H;ѺH;��H;w�H;ڗH; �H;!vH;�aH;nJH;�0H;jH;��G;r�G;%�G;�vG;9G;��F;��F;�0F;�E;�\E;�D;u�D;	D;      ��F;j�F;ܮF;�F;��F;�G;�GG;�pG;W�G;j�G;�G;��G;(H;=*H;�AH;�WH;jkH;L}H;W�H;��H;̧H;g�H;��H;e�H;��H;r�H;��H;��H;��H;N�H;L�H;��H;��H;��H;r�H;��H;�H;��H;t�H;��H;��H;��H;L�H;N�H;��H;��H;��H;t�H;�H;d�H;��H;g�H;ȧH;��H;W�H;M}H;hkH;�WH;�AH;=*H;'H;��G;�G;i�G;X�G;�pG;�GG;�G;��F;�F;ٮF;`�F;      uvG;(yG;#�G;��G;�G;��G;�G;��G;��G;�H;OH;�,H;�@H;�SH;�eH;�vH;ޅH;��H;)�H;%�H;��H;�H;b�H;��H;��H;��H;��H;��H;�H;�H;��H;��H;��H;�H;�H;`�H;`�H;^�H;�H;}�H;��H;��H;��H;�H;�H;��H;��H;��H;��H;��H;a�H;�H;��H;%�H;)�H;��H;܅H;�vH;�eH;�SH;�@H;�,H;OH;�H;��G;��G;�G;��G;�G;��G;!�G;(yG;      ?�G;��G;��G;��G;��G;��G;]H;%H;�(H;*8H;�GH;@WH;]fH;�tH;x�H;*�H;��H;��H;7�H;��H;7�H;��H;q�H;F�H;I�H;��H;��H;��H;��H;��H;��H;��H;��H;�H;��H;��H;��H;��H;��H;�H;��H;��H;��H;��H;��H;��H;��H;��H;L�H;H�H;o�H;��H;4�H;��H;7�H;��H;�H;*�H;x�H;�tH;\fH;AWH;�GH;)8H;�(H;%H;]H;��G;��G;��G;��G;��G;      �H;� H;y#H;>(H;�.H;�6H;"@H;dJH;qUH;�`H;�lH;PxH;��H;��H;�H;��H;��H;гH;=�H;��H;��H;��H;�H;��H;�H;��H;�H;��H;p�H;��H;��H;��H;*�H;��H;��H;�H;-�H;�H;��H;��H;'�H;��H;��H;��H;o�H;��H;�H;��H; �H;��H;�H;��H;��H;��H;=�H;ӳH;��H;��H;�H;��H;��H;MxH;�lH;�`H;sUH;bJH;"@H;�6H;�.H;>(H;x#H;� H;      �OH;ZPH;�RH;VH;�ZH;�`H;�gH;toH;�wH;?�H;��H;͑H;j�H;��H;��H;��H;ظH;�H;��H;��H;T�H;H�H;��H;��H;,�H;L�H;�H;��H;��H;��H;��H;&�H;��H;�H;8�H;\�H;q�H;\�H;8�H;�H;��H;)�H;��H;��H;��H;��H;�H;J�H;-�H;��H;��H;H�H;R�H;��H;��H;�H;׸H;��H;��H;��H;j�H;ˑH;��H;?�H;�wH;uoH;�gH;�`H;�ZH;VH;�RH;WPH;      �sH;atH;�uH;�xH;1|H;��H;ƅH;��H;��H;,�H;ҞH;v�H;�H;2�H;�H;ԽH;*�H;��H;^�H;A�H;��H;��H;T�H;��H;��H;N�H;��H;��H;��H;��H;�H;��H;�H;N�H;��H;��H;��H;��H;��H;P�H;�H;��H;�H;��H;��H;��H;��H;L�H;��H;��H;Q�H;��H;��H;A�H;^�H;��H;)�H;ҽH;�H;0�H;�H;t�H;ӞH;.�H;��H;��H;ƅH;��H;-|H;�xH;�uH;atH;      �H;W�H;��H;��H;1�H;��H;n�H;��H;f�H;7�H;7�H;-�H;�H;�H;��H;�H;�H;��H;��H;�H;��H;"�H;)�H;��H;v�H;��H;��H;��H;��H;*�H;��H;�H;J�H;��H;��H;��H;��H;��H;��H;��H;I�H;�H;��H;,�H;��H;��H;��H;��H;y�H;��H;)�H;"�H;��H;�H;��H;��H;�H;�H;��H;�H;�H;*�H;6�H;7�H;h�H;��H;n�H;��H;/�H;��H;��H;S�H;      ��H;�H;�H;��H;��H;	�H;�H;<�H;ϳH;��H;d�H;P�H;%�H;��H;\�H;��H;��H;��H;X�H;��H;��H;��H;p�H;��H;��H;��H;��H;��H;0�H;��H;�H;N�H;��H;��H;��H;��H;�H;��H;��H;��H;��H;P�H;�H;��H;1�H;��H;��H;��H;��H;��H;p�H;��H;��H;��H;X�H;��H;��H;��H;\�H;��H;#�H;O�H;e�H;��H;ϳH;;�H;�H;�H;�H;��H;�H;�H;      ɰH;�H;��H;�H;��H;��H;ѸH;|�H;2�H;&�H;4�H;,�H;(�H;�H;��H;��H;�H;V�H;v�H;e�H;'�H;��H;��H;�H;�H;��H;|�H;�H;��H;�H;L�H;��H;��H;��H;��H;�H;	�H;�H;��H;��H;��H;��H;L�H;�H;��H;�H;|�H;��H;�H;�H;��H;��H;&�H;d�H;v�H;W�H;�H;��H;��H;�H;(�H;,�H;3�H;&�H;2�H;{�H;ѸH;��H;��H;�H;��H;�H;      )�H;�H;�H;��H;a�H;ھH;��H;��H;�H;��H;��H;w�H;��H;Q�H;��H;��H;��H;��H;��H;;�H;��H;��H;��H;��H;��H;q�H;�H;��H;��H;<�H;��H;��H;��H;��H;�H;�H;�H;�H;�H;��H;��H;��H;��H;=�H;��H;��H;�H;q�H;��H;��H;��H;��H;��H;9�H;��H;��H;��H;��H;��H;P�H;��H;w�H;��H;��H;�H;��H;��H;߾H;W�H;�H;�H;w�H;      ��H;��H;.�H;��H;(�H;��H;/�H;�H;��H;�H;D�H;��H;��H;��H;��H;��H;��H;Y�H;��H;[�H;��H;��H;��H;w�H;�H;��H;^�H;��H;�H;_�H;��H;��H;��H;�H;�H;/�H;%�H;/�H;�H;�H;��H;��H;��H;_�H;�H;��H;]�H;��H;�H;u�H;��H;��H;��H;[�H;��H;Z�H;��H;��H;��H;��H;��H;��H;C�H;�H;��H;��H;/�H;��H;�H;��H;0�H;��H;      \�H;s�H;��H;��H;��H;�H;��H;g�H;T�H;M�H;g�H;s�H;x�H;��H;��H;}�H;5�H;��H;1�H;��H;��H;��H;��H;��H;`�H;
�H;^�H;��H;/�H;x�H;��H;��H;�H;�H;�H;(�H;2�H;(�H;�H;�H;�H;��H;��H;z�H;2�H;��H;]�H;�H;`�H;��H;��H;��H;��H;��H;1�H;��H;3�H;}�H;��H;��H;x�H;s�H;g�H;P�H;U�H;d�H;��H;�H;��H;��H;��H;i�H;      ��H;��H;.�H;��H;(�H;��H;/�H;�H;��H;�H;D�H;��H;��H;��H;��H;��H;��H;Y�H;��H;[�H;��H;��H;��H;w�H;�H;��H;^�H;��H;�H;_�H;��H;��H;��H;�H;�H;/�H;%�H;/�H;�H;�H;��H;��H;��H;_�H;�H;��H;]�H;��H;�H;u�H;��H;��H;��H;[�H;��H;Z�H;��H;��H;��H;��H;��H;��H;D�H;�H;��H;��H;/�H;��H;�H;��H;-�H;��H;      (�H;�H;
�H;��H;a�H;ھH;��H;��H;�H;��H;��H;w�H;��H;Q�H;��H;��H;��H;��H;��H;;�H;��H;��H;��H;�H;��H;q�H;�H;��H;��H;<�H;��H;��H;��H;��H;�H;�H;�H;�H;�H;��H;��H;��H;��H;=�H;��H;��H;�H;q�H;��H;��H;��H;��H;��H;9�H;��H;��H;��H;��H;��H;Q�H;��H;w�H;��H;��H;�H;��H;��H;߾H;W�H;��H;�H;u�H;      ʰH;�H;��H;�H;��H;��H;ѸH;{�H;0�H;&�H;4�H;,�H;(�H;�H;��H;��H;�H;V�H;v�H;e�H;*�H;��H;��H;�H;�H;��H;|�H;�H;��H;�H;L�H;��H;��H;��H;��H;�H;	�H;�H;��H;��H;��H;��H;L�H;�H;��H;�H;|�H;��H;�H;�H;��H;��H;&�H;d�H;v�H;W�H;�H;��H;��H;�H;(�H;,�H;4�H;&�H;2�H;y�H;ѸH;��H;��H;�H;��H;�H;      ��H;�H;�H;��H;��H;�H;�H;;�H;ϳH;��H;e�H;O�H;#�H;��H;\�H;��H;��H;��H;X�H;��H;��H;��H;q�H;��H;��H;��H;��H;��H;0�H;��H;�H;N�H;��H;��H;��H;��H;�H;��H;��H;��H;��H;Q�H;�H;��H;1�H;��H;��H;��H;��H;��H;n�H;��H;��H;��H;X�H;��H;��H;��H;]�H;��H;#�H;P�H;d�H;��H;ͳH;:�H;�H;�H;}�H;��H; �H;
�H;      	�H;W�H;��H;��H;1�H;��H;p�H;��H;f�H;7�H;6�H;,�H;�H;�H;��H;�H;�H;��H;��H;�H;��H;"�H;*�H;��H;y�H;��H;��H;��H;��H;*�H;��H;�H;J�H;��H;��H;��H;��H;��H;��H;��H;G�H;�H;��H;,�H;��H;��H;��H;��H;v�H;��H;'�H;"�H;��H;�H;��H;��H;�H;�H;��H;�H;�H;,�H;7�H;7�H;h�H;��H;p�H;��H;.�H;��H;��H;R�H;      �sH;atH;�uH;�xH;0|H;��H;ƅH;��H;��H;-�H;ҞH;t�H;�H;3�H;�H;ԽH;)�H;��H;^�H;A�H;��H;��H;T�H;��H;��H;N�H;��H;��H;��H;��H;�H;��H;�H;P�H;��H;��H;��H;��H;��H;N�H;�H;��H;�H;��H;��H;��H;��H;L�H;��H;��H;Q�H;��H;��H;A�H;^�H;��H;)�H;ԽH;�H;2�H;�H;v�H;ўH;-�H;��H;��H;ƅH;��H;-|H;�xH;�uH;atH;      �OH;ZPH;�RH;VH;�ZH;�`H;�gH;uoH;�wH;?�H;��H;͑H;j�H;��H;��H;��H;ظH;�H;��H;��H;V�H;H�H;��H;��H;/�H;L�H;�H;��H;��H;��H;��H;'�H;��H;�H;8�H;\�H;q�H;\�H;8�H;�H;��H;'�H;��H;��H;��H;��H;�H;J�H;,�H;��H;��H;H�H;R�H;��H;��H;�H;׸H;��H;��H;��H;j�H;͑H;��H;>�H;�wH;uoH;�gH;�`H;�ZH;VH;�RH;XPH;      �H;� H;#H;<(H;�.H;�6H;%@H;fJH;qUH;�`H;�lH;PxH;��H;��H;�H;��H;��H;гH;=�H;��H;��H;��H;�H;��H; �H;��H;�H;��H;p�H;��H;��H;��H;*�H;��H;��H;�H;-�H;�H;��H;��H;)�H;��H;��H;��H;p�H;��H;�H;��H;�H;��H;�H;��H;��H;��H;=�H;ҳH;��H;��H;�H;��H;��H;PxH;�lH;�`H;sUH;dJH;%@H;�6H;�.H;8(H;|#H;� H;      ?�G;��G;��G;��G;��G;��G;]H;(H;�(H;)8H;�GH;AWH;\fH;�tH;x�H;*�H;��H;��H;7�H;��H;:�H;��H;q�H;H�H;L�H;��H;��H;��H;��H;��H;��H;��H;��H;�H;��H;��H;��H;��H;��H;�H;��H;��H;��H;��H;��H;��H;��H;��H;I�H;F�H;o�H;��H;6�H;��H;7�H;��H;�H;,�H;x�H;�tH;]fH;@WH;�GH;*8H;�(H;%H;]H;��G;��G;��G;��G;��G;      ovG;(yG; �G;��G;ݝG;��G; �G;��G;��G;�H;OH;�,H;�@H;�SH;�eH;�vH;ޅH;��H;)�H;&�H;��H;�H;b�H;��H;��H; �H;��H;��H;�H;�H;��H;��H;��H;}�H;�H;^�H;`�H;^�H;�H;}�H;��H;��H;��H;�H;�H;��H;��H;��H;��H;��H;a�H;�H;��H;#�H;)�H;��H;܅H;�vH;�eH;�SH;�@H;�,H;PH;�H;��G;��G; �G;��G;��G;��G; �G;yG;      ��F;b�F;�F;�F;��F;�G;�GG;�pG;W�G;j�G;�G;��G;'H;=*H;�AH;�WH;jkH;L}H;W�H;��H;ͧH;g�H;��H;e�H;�H;t�H;��H;��H;��H;P�H;L�H;��H;��H;��H;q�H;��H;�H;��H;t�H;��H;��H;��H;L�H;M�H;��H;��H;��H;r�H;��H;d�H;��H;g�H;ȧH;��H;W�H;M}H;hkH;�WH;�AH;=*H;(H;��G;�G;i�G;W�G;�pG;�GG;�G;��F;�F;�F;Z�F;      �mD;	D;v�D;�D;�\E;�E;�0F;��F;��F;9G;�vG;%�G;r�G;��G;jH;�0H;pJH;�aH;!vH; �H;ݗH;w�H;��H;ӺH;*�H;�H;��H;O�H;#�H;4�H;��H;{�H;��H;�H;��H;�H;d�H;�H;��H;�H;��H;|�H;��H;3�H; �H;O�H;��H;�H;)�H;ѺH;��H;w�H;ۗH; �H;!vH;�aH;nJH;�0H;jH;��G;t�G;$�G;�vG;9G;��F;��F;�0F;�E;�\E;�D;u�D;	D;      k`?;�?;�?;�@;ĘA;��B;ښC;�D;eiE;F;K�F;G;{nG;C�G;%�G;y H;�!H;P?H;�YH;�pH;��H;��H;E�H;��H;̺H;g�H;��H;C�H;��H;��H;��H;��H;��H;�H;��H;q�H;��H;q�H;��H;�H;��H;��H;��H;��H;��H;C�H;�H;g�H;ʺH;��H;C�H;��H;��H;�pH;�YH;S?H;�!H;y H;%�G;C�G;znG;G;H�F;F;eiE;�D;ښC;��B;ԘA;�@;�?;ֈ?;      j�4;@�4;z�5;m7;�_9;��;;��=;7�?;��A;��C;��D;��E;��F;�)G;ƁG;5�G;�G;rH;�6H;TH;?mH;��H;�H;F�H;��H;��H;d�H;o�H;�H;��H;S�H;'�H;p�H;��H;��H;��H;��H;��H;��H;��H;n�H;'�H;S�H;��H;�H;n�H;`�H;��H;��H;C�H;�H;��H;9mH;TH;�6H;uH;�G;5�G;ǁG;�)G;��F;��E;��D;��C;��A;7�?;��=;��;;�_9;m7;p�5;0�4;      .e;7 ;�";i%;�(;Hj-;\2;�6;֡:;�0>;�A;nYC;Z�D;4F;E�F;�XG;,�G;y�G;�H;�1H;-QH;lH;��H;��H;t�H;j�H;�H;��H;��H;J�H;��H;�H;��H;��H;��H;��H;��H;��H;��H;��H;��H;�H;��H;F�H;��H;��H;�H;k�H;s�H;��H;��H;lH;*QH;�1H;�H;{�G;,�G;�XG;F�F;4F;Z�D;oYC;�A;�0>;١:;�6;]2;Gj-;�(;h%;�";2 ;      ���:�B�:��:�x;��
;�;L�;�}$;P|,;��3;�_9;\>;6zA;��C;�E;,�F;N5G;��G;��G;xH;�/H;+QH;=mH;��H;ٗH;ϧH;��H;7�H;��H;R�H;��H;��H;��H;�H;��H;�H;��H;��H;��H;�H;��H;��H;��H;O�H;��H;7�H;��H;ϧH;ٗH;��H;<mH;+QH;�/H;zH;��G;��G;M5G;,�F;�E;��C;6zA;\>;�_9;��3;S|,;�}$;L�;�;��
;�x;��:�B�:       x[:HCd:��}:#�:��:��:@�:1�;�;| ;�+;��3;��:;8�?;��B;�E;rZF;�G;M�G;��G;zH;�1H;TH;�pH;�H;��H;"�H;��H;��H;��H;:�H;�H;��H;\�H;1�H;Q�H;��H;Q�H;1�H;\�H;��H;�H;:�H;��H;��H;��H;�H;��H;�H;�pH;TH;�1H;vH;��G;M�G; G;rZF;�E;��B;8�?;��:;��3;�+;{ ;�;2�;@�:��:��:!�:��}: Cd:      T�S�P�D�d������ -(7��9ʍR:N��:v��:J��:�>;�";Q.;Im7;�=;|B;�D;�9F;NG;Q�G;��G;�H;�6H;�YH;vH;[�H;*�H;9�H;=�H;��H;^�H;��H;U�H;q�H;��H;��H;/�H;��H;��H;q�H;R�H;��H;]�H;��H;:�H;:�H;'�H;\�H;vH;�YH;�6H;�H;��G;R�G;NG;�9F;�D;|B;�=;Im7;Q.;�";�>;J��:z��:L��:ƍR: �9 3(7����d��P�D�      E^�0X�rF�3}*�,���P����D� ̬��i:��:s��:Q�;��;b�);��4;8�<;5�A;I�D;�9F;G;��G;y�G;uH;S?H;�aH;N}H;��H;��H;ԳH;�H;��H;��H;��H;V�H;��H;]�H;��H;]�H;��H;V�H;��H;��H;��H;�H;ҳH;��H;��H;P}H;�aH;O?H;rH;y�G;��G;G;�9F;I�D;3�A;8�<;��4;`�);��;Q�;s��:��:�i:`̬���D��P��&��3}*�rF�0X�      ��ﻭ��b�ܻH�ƻh󩻷��|FL�������������-::�:���:
;�>&;��3;z9<;6�A;�D;wZF;Q5G;/�G;�G;�!H;kJH;kkH;ޅH;��H;��H;׸H;%�H;��H;��H;�H;��H;��H;.�H;��H;��H;�H;��H;��H;%�H;ָH;��H;��H;مH;mkH;kJH;�!H;�G;/�G;P5G;xZF;�D;9�A;x9<;��3;�>&;
;���:8�:��-:����������|FL����g�H�ƻb�ܻ���      t�V��5S��6H���6�F� �V,��?ػ;G���D^������D� ��9�4�:/�:G�;%;��3;;�<;~B;�E;/�F;�XG;7�G;} H;�0H;�WH;�vH;*�H;��H;��H;ͽH; �H;��H;��H;��H;��H;u�H;��H;��H;��H;��H;�H;ͽH;��H;��H;*�H;�vH;�WH;�0H;y H;5�G;�XG;.�F;�E;~B;=�<;��3;%;H�;/�:�4�: ��9��D�����D^�<G���?ػU,�F� ���6��6H��5S�      "��.��NȤ��������B�f�y�=����?�ܻ�*��Po5�D��� �(7��}:�n�:E�;�>&;��4;�=;��B;�E;C�F;ǁG;(�G;gH;�AH;�eH;w�H;�H;��H;�H;��H;\�H;��H;��H;��H;��H;��H;��H;��H;[�H;��H;�H;��H;�H;w�H;�eH;�AH;hH;$�G;��G;C�F;�E;��B;�=;��4;�>&;E�;�n�:��}: �(7D���Po5��*��?�ܻ���y�=�A�f��������NȤ�.��      �c��8���������Ҽ����������r�KE:�F,�Lߵ�v/X�l�º Ŭ���}:5�:;e�);Jm7;>�?;��C;5F;�)G;C�G;�G;=*H;�SH;�tH;��H;��H;,�H;�H;��H;�H;J�H;��H;��H;��H;J�H;�H;��H;�H;,�H;��H;��H;�tH;�SH;@*H;��G;A�G;�)G;5F;��C;?�?;Jm7;f�);
;3�:��}: Ŭ�l�ºv/X�Lߵ�F,�KE:���r�����������Ҽ�켼����8�      ('K��G���>��0�ay��c����X��� ��Z�V�*���ƻ�od�n�º �(7�4�:���:��;Q.;�:;6zA;Z�D;��F;~nG;p�G;(H;�@H;\fH;��H;d�H;�H;�H;!�H;'�H;��H;��H;t�H;��H;��H;'�H;"�H;�H;�H;d�H;��H;\fH;�@H;+H;t�G;znG;��F;Z�D;8zA;�:;Q.;��;���:�4�: �(7p�º�od��ƻ+��Z�V� ��Y�����众c�ay��0���>��G�      	���4Z��Ґ����}��c���D�6/%��8���Ҽ2c��7�f�����ƻx/X�@���(��9:�:U�;�";��3;^>;mYC;��E;G;!�G;��G;�,H;;WH;LxH;��H;l�H;#�H;K�H;(�H;n�H;|�H;k�H;|�H;l�H;(�H;H�H;%�H;l�H;��H;JxH;;WH;�,H;��G;$�G;G;��E;mYC;b>;��3;�";U�;6�: ��9@���x/X��ƻ���7�f�2c����Ҽ�8�6/%���D��c���}�Ґ��4Z��      �Pν �ʽR8���������ѐ��e�f���;�5�����FȤ�7�f�*��Mߵ�No5���D���-:s��:�>;�+;�_9;�A;��D;K�F;�vG;�G;OH;�GH;�lH;�H;ΞH;0�H;d�H;0�H;��H;<�H;`�H;=�H;��H;0�H;a�H;2�H;ΞH;�H;�lH;�GH;LH;�G;�vG;G�F;��D;�A;�_9;�+;�>;u��:��-:��D�No5�Mߵ�+��8�f�FȤ����5����;�e�f�ѐ���������R8�� �ʽ      ���j9�][��s��ؽ���t����}� �G������3c��Z�V�G,��*����������:N��:| ;��3;�0>;��C;F;9G;k�G;�H;%8H;�`H;7�H;'�H;5�H;��H;$�H;��H;�H;M�H;�H;��H;$�H;}�H;5�H;'�H;7�H;�`H;&8H;�H;m�G;9G;F;��C;�0>;��3;{ ;N��:��:�������*��G,�Z�V�3c������� �G���}�t������ؽ�s�][�j9�      ��=�ڀ:���0��Q"��������Pν�榽B�� �G�4����Ҽ ��KE:�=�ܻ�D^������i:x��:�;P|,;ԡ:;��A;diE;��F;X�G;��G;�(H;qUH;�wH;��H;a�H;̳H;.�H;�H;��H;M�H;��H;�H;.�H;ȳH;a�H;��H;�wH;oUH;�(H;��G;Z�G;��F;aiE;��A;ԡ:;S|,;�;v��:�i:�����D^�>�ܻLE:� ����Ҽ5����G�B���榽�Pν�������Q"���0�ڀ:�      6Dx�8�s���f�xS�ڀ:����\[��7ս�榽��}���;��8�X�����r����9G������ˬ�T��:5�;�}$;�6;5�?;�D;��F;�pG;��G;H;bJH;moH;v�H;��H;4�H;t�H;��H;��H;a�H;��H;��H;t�H;3�H;��H;v�H;moH;_JH;H;��G;�pG;��F;�D;5�?;�6;�}$;4�;R��:@ˬ����9G�������r�X����8���;���}��榽�7ս\[����ڀ:�xS���f�8�s�      �*���0��॒�=����k��H��#%�\[��Pν
t��e�f�6/%���伈���x�=��?ػ�FL�|�D���R:D�:C�;R2;��=;ךC;�0F;�GG;��G;VH;@H;�gH;��H;i�H;�H;θH;��H;(�H;��H;(�H;��H;θH;�H;i�H;��H;�gH;@H;YH;��G;�GG;�0F;ԚC;��=;S2;F�;B�:��R:|�D��FL��?ػx�=��������6/%�e�f�
t���Pν\[��#%��H��k�=���॒��0��      *�þ
���"����R��~쏾8�s��H�����������ѐ����D��c�����A�f�U,�����P����9��:�;?j-;��;;��B;�E;�G;��G;��G;�6H;�`H;��H;��H;�H;��H;ݾH;��H;�H;��H;ݾH;��H;�H;��H;��H;�`H;�6H;��G;��G;�G;�E;��B;��;;?j-;�;��:��9�P�����U,�A�f������c���D�ѐ�������������H�8�s�~쏾�R��"���
���      C��2�很Yؾ*�þĪ�~쏾�k�ڀ:���~�ؽ�����c�`y���Ҽ ���E� �f�%�� 1(7��:��
;�(;�_9;ʘA;�\E;��F;ڝG;��G;�.H;�ZH;#|H;*�H;�H;��H;I�H;�H;��H;�H;G�H;��H;|�H;-�H;#|H;�ZH;�.H;��G;۝G;��F;�\E;ƘA;�_9;�(;��
;��: 2(7$��g�E� � �����Ҽ`y��c�����~�ؽ��ڀ:��k�~쏾Ī�*�þ�Yؾ2��      %��P������AI�*�þ�R��=���xS��Q"��s������}��0��켋�����6�E�ƻ2}*�����'�:�x;o%;m7;�@;��D;�F;��G;��G;:(H;VH;�xH;��H;{�H;ٲH;�H;��H;��H;��H;�H;ٲH;z�H;��H;�xH;VH;7(H;��G;��G;�F;��D;�@;m7;o%;�x;%�:����2}*�F�ƻ��6��������0���}�����s��Q"�xS�=����R��*�þAIᾦ���P��      ���T��:�
������Yؾ"���॒���f���0�\[�R8��Ґ����>�����NȤ��6H�`�ܻrF������}:���:z";i�5;�?;��D;�F; �G;��G;x#H;�RH;�uH;��H;��H;��H;�H;&�H;��H;&�H;�H;��H;��H;��H;�uH;�RH;u#H;��G; �G;�F;��D;�?;l�5;z"; ��:��}:���rF�a�ܻ�6H�NȤ�������>�Ґ��R8��\[���0���f�॒�"����Yؾ����:�
�T��      �� ����T��P��2��
����0��8�s�ڀ:�i9� �ʽ4Z���G��8�.���5S�����/X�@�D�Cd:�B�: ;/�4;׈?;D;Z�F;$yG;��G;� H;SPH;OtH;H�H;�H;�H;i�H;��H;l�H;��H;j�H;�H;��H;I�H;OtH;PPH;� H;��G;#yG;\�F;D;ӈ?;4�4; ;�B�:Cd:@�D��/X���껱5S�.���8��G�4Z�� �ʽi9�ڀ:�8�s��0��
���2��P��T�����      HEb�c]��N���7����u� ���˾��,�j��!,�t���O��Hm�.��;,˼��x�Z���1����:�:�;T�1;C,>;��C;�wF;�G;� H;?H;�hH;b�H;��H;M�H;.�H;��H;<�H;��H;<�H;��H;.�H;L�H;��H;b�H;�hH;?H;� H;�G;�wF;��C;@,>;W�1;�;�:��:��1��Z��ªx�;,˼.��Hm�O��t����!,�,�j�����˾u� ������7��N�c]�      c]�g�W��TI�v3� E�������Ǿx����f�;)�(��u;���Fi��k���Ǽ�[t�L�	�(Ȅ� X��|�:��:��;kJ2;`Z>;W	D;�F;Q�G;(H;�?H;�iH;��H;�H;��H;J�H;��H;h�H;��H;h�H;��H;J�H;��H;�H;��H;�iH;�?H;(H;Q�G;�F;W	D;\Z>;qJ2;��;��:t�: X��'Ȅ�L�	��[t���Ǽ�k��Fi�u;��(��;)��f�x�����Ǿ���� E�v3��TI�g�W�      �N��TI���;�1�'�l��쾂���{󐾷Z��K ��s�C����&^���"����g����̨u�� ��~3<:-��:;xg3;�>;�BD;ĖF;��G;�H;YBH;�kH;f�H;�H;;�H;�H;~�H;��H;V�H;��H;}�H;�H;9�H;�H;f�H;�kH;VBH;�H;��G;ƖF;�BD;��>;{g3;;-��:v3<:� ��ʨu������g��"����&^�C����s潧K ��Z�{󐾂�����l�1�'���;��TI�      ��7�v3�1�'����u� ��{Ծ!���J���|�F�����ӽ���b�L�Lv��뮼ST����PV�X�=�*i:���:�z ;�$5;��?;�D;޺F;�G;�H;�FH;�nH;��H;��H;~�H;�H;F�H;e�H;�H;e�H;F�H;�H;|�H;��H;��H;�nH;�FH;�H;�G;޺F;�D;��?;�$5;�z ;���:*i:X�=��PV���ST��뮼Lv�b�L�����ӽ���|�F�J���!����{Ծu� ����1�'�v3�      ��� E�l�u� �Y�ݾm���X͓��f��>/�����'���섽R�6��t�w��_�:�!Tʻr.��ڷ��t�:�;��$;�Y7;h�@;	
E;-�F;G�G;�H;JLH;�rH;H;ؤH;1�H;/�H;@�H;X�H;��H;X�H;?�H;/�H;.�H;ڤH;��H;�rH;ILH;�H;I�G;,�F;
E;d�@;�Y7;��$;�;�t�:�ڷ�q.�"Tʻ_�:�w���t�R�6��섽�'������>/��f�X͓�m���Y�ݾu� �l� E�      u� ��������{Ծm���x���^�x��SC��^��޽B���|�e�*��F�Ѽ'G������R�����@�8��:�Y;c�);�9;�A;΄E;�G;-�G;v!H;OSH;�wH;��H;��H;N�H;��H;��H;��H;��H;��H;��H;��H;N�H;��H;��H;�wH;KSH;u!H;+�G;�G;˄E;�A;�9;c�);�Y;��:@�8����R�����'G��F�Ѽ*��|�e�B����޽�^��SC�^�x�x���m����{Ծ�쾣���      ��˾��Ǿ����!���X͓�^�x���J��K �r��� ������?����뮼-�[����3|�~W����:��:�';�/;xg<;�C;}F;�NG;��G;<-H;|[H;�}H;ӗH;ӪH;ɸH;��H;�H;��H;�H;��H;�H;��H;ɸH;ժH;ӗH;�}H;x[H;<-H;��G;�NG;yF;�C;vg<;�/;�';��:��:xW��3|����-�[��뮼���?���� ��r����K ���J�^�x�X͓�!���������Ǿ      ��x���{�J����f��SC��K �rn���Ž����Z��k�"}ռ.X��by-�)���].� ���P�:�+�:��;14;I�>;D;�wF;C�G;��G;�9H;gdH;��H;��H;m�H;{�H;��H;��H;`�H;}�H;`�H;��H;��H;y�H;p�H;��H;~�H;bdH;�9H;��G;C�G;�wF;	D;I�>;14;��;�+�:�P�:���_.�)���by-�.X��"}ռ�k��Z�����Žrn���K ��SC��f�J���{�x���      ,�j��f��Z�|�F��>/��^�r����ŽI ���Fi��Q+�~t�qT��q�W�����1��Ⱥ�X�9�P�:�Y;��(;�8;A;�E;�F;y�G;�H;�FH;�mH;��H;ΡH;K�H;z�H;��H;��H;�H;�H;�H;��H;��H;z�H;M�H;ΡH;��H;�mH;�FH;�H;{�G;�F;�E;A;�8;��(;�Y;�P�:�X�9Ⱥ�1�����q�W�qT��~t�Q+��Fi�I ���Žr����^��>/�|�F��Z��f�      �!,�;)��K ��������޽ ������Fi��0����鷼��x�����.��F�(����X+i:���:Q�;��0;`�<;�C;��E;=G;�G;%H;sTH;�wH;��H;%�H;Y�H;��H;L�H;��H;��H;��H;��H;��H;L�H;��H;[�H;%�H;��H;�wH;sTH;%H;�G;=G;��E;�C;`�<;��0;P�;���:\+i:���E�(��.�������x�鷼����0��Fi���� ���޽�������K �;)�      t���(��s��ӽ�'��B�������Z��Q+�����"��G��»0���׻b�W���Y�9 ��:>`;�*';�Y7; $@;;�D;�F;'�G;��G;H8H;bH;�H;f�H;��H;�H;��H;��H;��H;\�H;H�H;\�H;��H;��H;��H;��H;��H;d�H;�H;bH;G8H;��G;"�G;�F;8�D; $@;�Y7;�*';>`;��:�Y�9W��b���׻��0�G���"������Q+��Z����B����'���ӽ�s�(��      P��u;��C�������섽|�e��?��k�t�鷼G���e7�����Ǆ�T0���t�Vu�:1,�:�;�1;h�<;w�B;9�E;G;�G;pH;�JH;moH;�H;��H;"�H;��H;��H;+�H;��H;�H;��H;�H;��H;,�H;��H;��H;"�H;��H;�H;moH;�JH;rH;�G;G;6�E;w�B;h�<;�1;�;3,�:Ru�:��t�T0��Ǆ���껅e7�G��鷼t��k��?�|�e��섽���C���u;��      Hm��Fi��&^�b�L�R�6�*����#}ռqT����x���0�������
���׷�Ho`:��:0�;>�*;N�8;%�@;K�D;z�F;~G;��G;�1H;�[H;~|H;ΕH;�H;��H;��H;��H;��H;��H;��H;��H;��H;��H;��H;��H;��H;��H;�H;˕H;~|H;�[H;�1H;��G;~G;v�F;K�D;#�@;N�8;>�*;4�;��:Po`:�׷�����������0���x�qT��#}ռ��*��S�6�b�L��&^��Fi�      .���k��Lv��t�F�Ѽ�뮼.X��p�W������׻�Ǆ�
�����^5<:���:�Y;�t%;%5;�Z>;aC;��E;G*G;v�G;'H;HH;}lH;�H;�H;үH;߼H;��H;��H;�H;��H;}�H;=�H;}�H;��H;�H;��H;��H;߼H;ЯH;�H;�H;|lH;HH;&H;t�G;C*G;��E;aC;�Z>;%5;�t%;�Y;���:b5<:���
���Ǆ���׻���p�W�/X���뮼F�Ѽ�t�Lv���k�      ;,˼��Ǽ�"���뮼w��'G��.�[�cy-�����.��ĕb�Z0�ط�V5<:M�:�\;��!;�J2;�g<;d0B;?CE;=�F;a�G;�G;�4H;�\H;|H;��H;��H;i�H;��H;O�H;��H;^�H;`�H;�H;��H;�H;a�H;a�H;��H;Q�H;��H;f�H;��H;��H;|H;�\H;�4H;�G;\�G;=�F;=CE;f0B;�g<;�J2;��!;�\;M�:V5<:ط�Z0�b��.�����cy-�.�[�'G��w���뮼�"����Ǽ      ªx��[t���g�ST�`�:�������+����1��F�(�W��@�t�Do`:���: ];!{ ;��0;r;;=A;,�D;�wF;�cG;g�G;�!H;�MH;�oH;��H;��H;ӯH;��H;u�H;��H;h�H;}�H;�H;��H;3�H;��H;�H;}�H;g�H;��H;u�H;��H;ϯH;��H;��H;�oH;�MH;�!H;d�G;�cG;�wF;*�D;=A;s;;��0;!{ ; ];���:Do`:@�t�W��H�(��1��+���������`�:�ST���g��[t�      Z��J�	������#Tʻ�R��3|�_.�Ⱥ����Y�9Ru�:��:�Y;��!;��0;��:;ĵ@;CD;�2F;�8G;��G;�H;{@H;8dH;րH;��H;W�H;Y�H;]�H;��H;��H;��H;}�H;��H;�H;��H;�H;��H;~�H;��H; �H;��H;[�H;V�H;W�H;��H;׀H;7dH;w@H;�H;��G;�8G;�2F;CD;Ƶ@;��:;��0;��!;�Y;��:Ru�:�Y�9���Ⱥ_.�3|��R��"Tʻ�����M�	�      �1��*Ȅ�̨u��PV�x.�����W����X�9T+i: ��:+,�:0�;�t%;�J2;o;;ĵ@;D;F;:G;��G;�H;�5H;�ZH;FxH;P�H;:�H;'�H;$�H;k�H;~�H;*�H;?�H;9�H;M�H;g�H;��H;g�H;M�H;9�H;>�H;,�H;~�H;j�H;!�H;(�H;9�H;S�H;FxH;�ZH;�5H;�H;��G;<G;F;�D;µ@;m;;�J2;�t%;0�;-,�: ��:P+i:�X�9(��W�����r.��PV�̨u�.Ȅ�      ꥥ�X��� ��T�=��ڷ���8��:�P�:�P�:���:>`;�;<�*;%5;�g<;=A;CD;F;�G;��G;y�G;�-H;*SH;jqH;��H;НH;��H;%�H;J�H;�H;�H;��H;d�H;��H;��H;��H;��H;��H;��H;��H;c�H;��H;�H; �H;H�H;%�H;��H;ҝH;��H;fqH;)SH;�-H;v�G;��G;�G; F;CD;=A;�g<;%5;<�*;�;>`;���:�P�:�P�:��:`�8�ڷ�X�=�� ��X��      �:��:z3<: *i:�t�:��:��:�+�:�Y;Q�;�*';�1;J�8;�Z>;a0B;%�D;�2F;6G;��G;.�G;�)H;�NH;�lH;^�H;x�H;��H;��H;@�H;��H;�H;I�H;9�H;C�H;j�H;��H;��H;��H;��H;��H;j�H;A�H;;�H;I�H;�H;��H;?�H;��H;��H;z�H;Z�H;�lH;�NH;�)H;.�G;��G;7G;�2F;%�D;a0B;�Z>;L�8;�1;�*';N�;�Y;�+�:��:��:�t�:*i:z3<:��:      ��:2��:5��:z��:�;�Y;�';��;��(;��0;�Y7;d�<;!�@;aC;=CE;�wF;�8G;��G;v�G;�)H;�LH;jH;G�H;m�H;��H;�H;̾H;u�H;6�H;��H;&�H;e�H;��H;��H;��H;��H;��H;��H;��H;��H;��H;g�H;&�H;��H;3�H;t�H;̾H;�H;��H;j�H;F�H;jH;�LH;�)H;w�G;��G;�8G;�wF;=CE;aC;!�@;d�<;�Y7;��0;��(;��;�';�Y;�;~��:5��:��:      �;��;$;�z ;��$;l�);�/;84;"�8;a�<;$$@;v�B;K�D;��E;>�F;�cG;��G;�H;�-H;�NH;jH;Z�H;ƔH;¤H;�H;ѼH;��H;��H;\�H;�H;��H;B�H;Z�H;��H;��H;{�H;��H;{�H;��H;��H;Y�H;B�H;��H;��H;X�H;��H;��H;ԼH;�H;��H;ŔH;Z�H;jH;�NH;�-H;�H;��G;�cG;@�F;��E;K�D;v�B;"$@;a�<;"�8;84;�/;o�);��$;�z ;#;��;      X�1;oJ2;yg3;�$5;�Y7;�9;zg<;K�>;A;�C;;�D;<�E;x�F;F*G;^�G;d�G;�H;�5H;)SH;�lH;F�H;ƔH;<�H;�H;��H;}�H;t�H;F�H;�H;��H;��H;��H;��H;��H;��H;;�H;��H;;�H;��H;��H;��H;��H;��H;��H;�H;G�H;r�H;~�H;��H;�H;<�H;ǔH;C�H;�lH;)SH;�5H;�H;c�G;^�G;F*G;x�F;:�E;;�D;�C;A;I�>;zg<;�9;�Y7;�$5;{g3;dJ2;      V,>;qZ>;�>;��?;j�@;�A;�C;D;�E;��E;�F;G;~G;v�G;�G;�!H;w@H;�ZH;fqH;[�H;i�H;��H;�H;0�H;��H;��H;]�H;(�H;�H;�H;|�H;J�H;��H;��H;v�H;��H;�H;��H;v�H;��H;��H;L�H;{�H;�H;�H;(�H;]�H;��H;��H;-�H;�H;��H;g�H;\�H;hqH;�ZH;u@H;�!H;�G;v�G;�}G;G;	�F;��E;�E;D;�C;�A;r�@;��?;�>;cZ>;      ��C;`	D;vBD;�D;	
E;τE;zF;�wF;�F;=G;$�G;�G;��G;*H;�4H;�MH;;dH;FxH;��H;�H;��H;�H;��H;��H;]�H;�H;��H;��H;��H;��H;��H;��H;��H;n�H;�H;r�H;y�H;p�H;�H;m�H;��H;��H;��H;��H;��H;��H;��H;�H;_�H;��H;��H;�H;��H;��H;��H;JxH;:dH;�MH;�4H;(H;��G;�G;$�G;=G;�F;�wF;zF;τE;
E;�D;uBD;^	D;      �wF;�F;��F;ݺF;,�F;�G;�NG;B�G;x�G;
�G;��G;rH;�1H;HH;�\H;�oH;ԀH;M�H;˝H;��H;޳H;мH;z�H;��H;�H;��H;O�H;L�H;��H;��H;G�H;��H;d�H;'�H;��H;��H;��H;��H;��H;'�H;a�H;��H;G�H;��H;��H;K�H;P�H;��H;�H;��H;|�H;ѼH;۳H;��H;͝H;P�H;ӀH;�oH;�\H;HH;�1H;rH;��G;�G;y�G;@�G;�NG;�G;3�F;ݺF;��F;�F;      �G;U�G;��G;�G;N�G;2�G;��G;��G;�H;%H;H8H;�JH;�[H;}lH;|H;��H;��H;7�H;��H;��H;ξH;��H;r�H;a�H;��H;S�H;3�H;��H;{�H;'�H;g�H;@�H;�H;��H;�H;6�H;D�H;6�H;��H;��H;�H;A�H;g�H;&�H;y�H;��H;3�H;Q�H;��H;a�H;r�H;��H;̾H;��H;��H;9�H;��H;��H;|H;}lH;�[H;�JH;I8H;%H;�H;��G;��G;/�G;T�G;
�G;��G;T�G;      � H;-H;�H;�H;�H;w!H;A-H;�9H;�FH;wTH;bH;roH;�|H;�H;��H;��H;U�H;$�H;"�H;C�H;t�H;��H;G�H;+�H;��H;L�H;��H;��H;�H;6�H;7�H;
�H;��H;�H;J�H;��H;��H;��H;J�H;�H;��H;
�H;9�H;5�H;	�H;��H;��H;L�H;��H;-�H;G�H;��H;r�H;C�H;$�H;$�H;T�H;��H;��H;�H;~|H;roH;bH;wTH;GH;�9H;A-H;w!H;�H;�H;�H;9H;      ?H;�?H;ZBH;�FH;LLH;OSH;�[H;idH;�mH;�wH;�H;�H;ЕH;�H;��H;ԯH;Z�H;!�H;I�H;��H;7�H;Y�H;�H;�H;��H;��H;v�H;�H;U�H;#�H;��H;��H;�H;i�H;��H;��H;��H;��H;��H;i�H;�H;��H;��H;%�H;U�H;�H;y�H;��H;��H;�H;�H;[�H;6�H;��H;J�H;"�H;Y�H;ԯH;��H;�H;ЕH;�H;�H;�wH;�mH;idH;�[H;NSH;SLH;�FH;ZBH;�?H;      iH;�iH;�kH;�nH;�rH; xH;�}H;��H;��H; �H;p�H;ˡH;�H;گH;j�H;��H;`�H;e�H;��H; �H;��H;��H;��H;�H;��H;��H;$�H;7�H;%�H;��H;��H;�H;U�H;��H;��H;��H;��H;��H;��H;��H;S�H;�H;��H; �H;#�H;6�H;#�H;��H;��H;�H;��H;��H;��H;�H;��H;g�H;]�H;��H;j�H;ׯH;�H;ɡH;p�H;��H;��H;��H;�}H; xH;�rH;�nH;�kH;�iH;      h�H;�H;u�H;��H;ЏH;��H;ۗH;ŜH;աH;)�H;��H;.�H;��H;�H;��H;|�H;��H;|�H;�H;P�H;*�H;��H;��H;�H;��H;I�H;d�H;:�H;��H;��H;�H;c�H;��H;��H;�H;�H;�H;�H;�H;��H;��H;e�H;�H;��H;��H;:�H;f�H;G�H;��H;�H;��H;��H;)�H;P�H;�H;|�H;��H;{�H;��H;�H;��H;,�H;��H;,�H;աH;ŜH;ۗH;��H;̏H;��H;r�H;�H;      ��H;�H;��H;��H;�H;��H;تH;x�H;Q�H;\�H;��H;��H;��H;��H;U�H;��H;�H;*�H;��H;B�H;m�H;D�H;��H;P�H;��H;��H;@�H;�H;��H;�H;b�H;��H;��H;�H;�H;9�H;U�H;9�H;�H;�H;��H;��H;b�H;�H;��H;�H;@�H;��H;��H;P�H;��H;D�H;m�H;B�H;��H;-�H;�H;��H;U�H;��H;��H;��H;��H;]�H;T�H;u�H;٪H;��H;ߤH;��H;��H;��H;      Q�H;��H;D�H;��H;;�H;N�H;̸H;��H;�H;��H;��H;��H;��H;��H;��H;n�H;��H;;�H;f�H;I�H;��H;\�H;��H;��H;��H;e�H;�H;��H;	�H;[�H;��H;��H;�H;.�H;R�H;G�H;:�H;G�H;Q�H;.�H;�H;��H;��H;\�H;�H;��H;�H;d�H;��H;��H;��H;\�H;��H;J�H;f�H;<�H;��H;n�H;��H;��H;��H;��H;��H;��H;��H;��H;̸H;R�H;4�H;��H;D�H;��H;      ;�H;W�H;�H;��H;7�H;��H;��H;��H;��H;N�H;��H;2�H;��H;�H;c�H;��H;��H;9�H;��H;r�H;��H;��H;��H;��H;h�H;&�H;��H;�H;h�H;��H;��H;�H;'�H;:�H;f�H;q�H;R�H;q�H;f�H;<�H;%�H;�H;��H;��H;j�H;�H;��H;&�H;j�H;��H;��H;��H;��H;r�H;��H;:�H;��H;��H;c�H;�H;��H;2�H;��H;N�H;��H;��H;��H;��H;-�H;��H;�H;P�H;      ��H;�H;��H;N�H;[�H;��H;�H;��H;��H;��H;��H;��H;��H;��H;e�H;�H;��H;J�H;��H;��H;��H;��H;��H;|�H;�H;��H;��H;J�H;��H;��H;�H;�H;Q�H;i�H;K�H;i�H;��H;i�H;K�H;i�H;N�H;�H;�H;��H;��H;J�H;��H;��H;�H;{�H;��H;��H;��H;��H;��H;L�H;��H;�H;e�H;��H;��H;��H;��H;��H;��H;��H;�H;��H;Q�H;M�H;��H;�H;      8�H;r�H;��H;j�H;j�H;��H;��H;k�H;�H;��H;d�H;&�H;��H;��H; �H;��H;�H;d�H;��H;��H;��H;~�H;=�H;��H;l�H;��H;5�H;��H;��H;��H;�H;=�H;G�H;w�H;i�H;_�H;p�H;_�H;i�H;t�H;D�H;@�H;�H;��H;��H;��H;5�H;��H;n�H;��H;=�H;~�H;��H;��H;��H;f�H;�H;��H; �H;��H;��H;&�H;c�H;��H;�H;i�H;��H;��H;_�H;j�H;��H;i�H;      ��H;��H;g�H;�H;��H;��H;�H;��H;	�H;��H;O�H;��H;��H;F�H;��H;<�H;��H;��H;��H;��H;��H;��H;��H;�H;s�H;��H;B�H;��H;��H;�H;�H;\�H;:�H;V�H;��H;q�H;]�H;q�H;��H;V�H;7�H;]�H;�H;�H;��H;��H;B�H;��H;s�H;
�H;��H;��H;��H;��H;��H;��H;��H;<�H;��H;F�H;��H;��H;O�H;��H;	�H;��H;�H;��H;��H;�H;g�H;��H;      8�H;r�H;��H;j�H;j�H;��H;��H;k�H;�H;��H;d�H;&�H;��H;��H;!�H;��H;�H;d�H;��H;��H;��H;~�H;=�H;��H;n�H;��H;5�H;��H;��H;��H;�H;=�H;G�H;w�H;i�H;_�H;p�H;_�H;i�H;t�H;D�H;@�H;�H;��H;��H;��H;5�H;��H;l�H;��H;=�H;~�H;��H;��H;��H;f�H;�H;��H; �H;��H;��H;&�H;d�H;��H;�H;i�H;��H;��H;_�H;j�H;��H;h�H;      ��H;�H;��H;N�H;[�H;��H;�H;��H;��H;��H;��H;��H;��H;��H;e�H;�H;��H;J�H;��H;��H;��H;��H;��H;|�H;�H;��H;��H;J�H;��H;��H;�H;�H;Q�H;i�H;K�H;i�H;��H;i�H;K�H;i�H;N�H;�H;�H;��H;��H;J�H;��H;��H;�H;y�H;��H;��H;��H;��H;��H;L�H;��H;�H;e�H;��H;��H;��H;��H;��H;��H;��H;�H;��H;Q�H;N�H;��H;�H;      <�H;W�H;�H;��H;7�H;��H;��H;��H;��H;N�H;��H;2�H;��H;�H;c�H;��H;��H;9�H;��H;r�H;��H;��H;��H;��H;j�H;'�H;��H;�H;h�H;��H;��H;�H;'�H;<�H;f�H;r�H;R�H;q�H;f�H;:�H;%�H;�H;��H;��H;j�H;�H;��H;'�H;h�H;��H;��H;��H;��H;r�H;��H;:�H;��H;��H;c�H;�H;��H;2�H;��H;N�H;��H;��H;��H;��H;-�H;��H;�H;P�H;      T�H;��H;F�H;��H;8�H;O�H;̸H;��H;��H;��H;��H;��H;��H;��H;��H;n�H;��H;:�H;f�H;I�H;��H;\�H;��H;��H;��H;e�H;�H;��H;	�H;[�H;��H;��H;�H;,�H;Q�H;G�H;:�H;G�H;R�H;,�H;�H;��H;��H;\�H;�H;��H;�H;d�H;��H;��H;��H;\�H;��H;J�H;f�H;;�H;��H;n�H;��H;��H;��H;��H;��H;��H;�H;��H;ʸH;R�H;1�H;��H;D�H;��H;      ��H;�H;��H;��H;ߤH;��H;ڪH;w�H;Q�H;]�H;��H;��H;��H;��H;U�H;��H;�H;*�H;��H;C�H;q�H;D�H;��H;P�H;��H;��H;@�H;�H;��H;�H;b�H;��H;��H;�H;�H;9�H;U�H;9�H;�H;�H;��H;��H;b�H;�H;��H;�H;@�H;��H;��H;P�H;��H;D�H;k�H;B�H;��H;,�H;�H;��H;U�H;��H;��H;��H;��H;]�H;R�H;u�H;ڪH;��H;ݤH;��H;��H;��H;      h�H;�H;r�H;��H;ϏH;��H;ۗH;ŜH;աH;*�H;��H;,�H;��H;�H;��H;|�H;��H;{�H;�H;Q�H;-�H;��H;��H;��H;��H;I�H;f�H;:�H;��H;��H;�H;c�H;��H;��H;�H;�H;�H;�H;�H;��H;��H;e�H;�H;��H;��H;:�H;f�H;G�H;��H;�H;��H;��H;'�H;P�H;�H;|�H;��H;|�H;��H;�H;��H;.�H;��H;*�H;աH;ŜH;ۗH;��H;͏H;��H;u�H;�H;      iH;�iH;�kH;�nH;�rH;�wH;�}H;��H;��H;��H;n�H;ɡH;�H;گH;j�H;��H;_�H;e�H;��H;"�H;��H;��H;��H;�H;��H;��H;$�H;6�H;%�H;�H;��H;�H;T�H;��H;��H;��H;��H;��H;��H;��H;T�H;�H;��H;��H;%�H;7�H;#�H;��H;��H;�H;��H;��H;��H;�H;��H;g�H;_�H;��H;j�H;ٯH;�H;ʡH;p�H;��H;��H;��H;�}H;�wH;�rH;�nH;�kH;�iH;      ?H;�?H;`BH;�FH;PLH;KSH;�[H;ldH;�mH;�wH;�H;�H;ЕH;�H;��H;ԯH;Z�H;!�H;J�H;��H;<�H;[�H;�H;�H;��H;��H;v�H;�H;U�H;&�H;��H;��H;�H;i�H;��H;��H;��H;��H;��H;i�H;�H;��H;��H;"�H;U�H;�H;y�H;��H;��H;	�H;�H;Y�H;5�H;��H;I�H;"�H;Y�H;֯H;��H;�H;ЕH;�H;�H;�wH;�mH;kdH;�[H;NSH;MLH;�FH;]BH;�?H;      � H;-H;�H;�H;�H;w!H;A-H;�9H; GH;wTH;bH;roH;~|H;�H;��H;��H;U�H;"�H;$�H;D�H;x�H;��H;I�H;-�H;��H;L�H;��H;��H;�H;7�H;9�H;
�H;��H;�H;I�H;��H;��H;��H;J�H;�H;��H;�H;7�H;3�H;	�H;��H;��H;L�H;��H;+�H;F�H;��H;q�H;B�H;"�H;$�H;T�H;��H;��H;�H;�|H;roH;bH;wTH;GH;�9H;A-H;u!H;�H;�H;�H;8H;      �G;T�G;��G;�G;J�G;.�G;��G;��G;�H;%H;I8H;�JH;�[H;}lH;|H;��H;��H;7�H;��H;��H;ҾH;��H;t�H;b�H;��H;T�H;4�H;��H;{�H;'�H;g�H;A�H;�H;��H;��H;6�H;D�H;5�H;�H;��H;�H;A�H;g�H;&�H;y�H;��H;3�H;Q�H;��H;`�H;q�H;��H;˾H;��H;��H;9�H;��H;��H;|H;}lH;�[H;�JH;I8H;%H;�H;��G;��G;-�G;M�G;�G;��G;I�G;      �wF;�F;F;ݺF;-�F;�G;�NG;B�G;v�G;
�G;��G;pH;�1H;HH;�\H;�oH;րH;O�H;͝H;��H;�H;ѼH;z�H;��H;�H;��H;P�H;K�H;��H;��H;G�H;��H;c�H;'�H;��H;��H;��H;��H;��H;'�H;a�H;��H;G�H;��H;��H;L�H;O�H;��H;�H;��H;z�H;мH;۳H;��H;˝H;O�H;рH;�oH;�\H;HH;�1H;rH;��G;�G;x�G;?�G;�NG;�G;2�F;�F;ÖF;�F;      ��C;`	D;uBD;�D;
E;τE;zF;�wF;�F;=G;%�G;�G;��G;(H;�4H;�MH;;dH;HxH;��H;��H;��H;�H;��H;��H;_�H;�H;��H;��H;��H;��H;��H;��H;��H;m�H;�H;p�H;y�H;r�H;�H;m�H;��H;��H;��H;��H;��H;��H;��H;�H;]�H;��H;��H;�H;��H;�H;��H;IxH;8dH;�MH;�4H;(H;��G;�G;$�G;=G;�F;�wF;zF;τE;
E;�D;uBD;`	D;      \,>;mZ>;�>;��?;d�@;�A;�C;D;�E;��E;�F;G;~G;v�G;�G;�!H;w@H;�ZH;hqH;\�H;k�H;��H;�H;2�H;��H;��H;^�H;(�H;�H;�H;{�H;J�H;��H;��H;t�H;��H;�H;��H;x�H;��H;��H;L�H;|�H;�H;�H;(�H;]�H;��H;��H;/�H;�H;��H;f�H;[�H;fqH;�ZH;u@H;�!H;�G;v�G;�}G;G;�F;��E;�E;D;�C;�A;t�@;��?;�>;_Z>;      U�1;|J2;�g3;�$5;�Y7;�9;~g<;I�>;A;�C;9�D;:�E;w�F;F*G;^�G;d�G;�H;�5H;)SH;�lH;H�H;ǔH;>�H;�H;��H;~�H;u�H;G�H;�H;��H;��H;��H;��H;��H;��H;;�H;��H;;�H;��H;��H;��H;��H;��H;��H;�H;F�H;q�H;}�H;��H;�H;;�H;ƔH;A�H;�lH;)SH;�5H;�H;d�G;`�G;F*G;w�F;<�E;;�D;�C;A;I�>;�g<;�9;�Y7;�$5;}g3;jJ2;      �;��;$;�z ;��$;m�);�/;84;"�8;a�<;#$@;v�B;K�D;��E;>�F;�cG;��G;�H;�-H;�NH;jH;Z�H;ǔH;äH;�H;ӼH;��H;��H;\�H; �H;��H;B�H;Z�H;��H;��H;{�H;��H;{�H;��H;��H;Y�H;B�H;��H;��H;X�H;��H;��H;ӼH;�H;��H;ÔH;Z�H;jH;�NH;�-H;�H;��G;�cG;@�F;��E;K�D;w�B;"$@;a�<;"�8;64;�/;l�);��$;�z ;$;��;      ��:(��:;��:~��:�;�Y;�';��;��(;��0;�Y7;d�<;"�@;aC;=CE;�wF;�8G;��G;w�G;�)H;�LH;jH;G�H;n�H;��H;�H;ξH;t�H;6�H;��H;&�H;e�H;��H;��H;��H;��H;��H;��H;��H;��H;��H;g�H;&�H;��H;3�H;u�H;˾H;�H;��H;i�H;F�H;jH;�LH;�)H;v�G;��G;�8G;�wF;=CE;aC;!�@;d�<;�Y7;��0;��(;��;�';�Y;�;~��:;��:��:      ��:��:�3<:�)i:�t�:��:��:�+�:�Y;P�;�*';�1;J�8;�Z>;a0B;%�D;�2F;6G;��G;.�G;�)H;�NH;�lH;^�H;z�H;��H;��H;?�H;��H;�H;I�H;9�H;C�H;j�H;��H;��H;��H;��H;��H;j�H;B�H;;�H;I�H;�H;��H;@�H;��H;��H;x�H;Z�H;�lH;�NH;�)H;.�G;��G;7G;�2F;%�D;a0B;�Z>;J�8;�1;�*';P�;�Y;�+�:��:��:�t�:�)i:�3<:��:      ꥥ�X��� ��X�=��ڷ���8��:�P�:�P�:���:>`;�;<�*;%5;�g<;=A;CD;F;�G;��G;y�G;�-H;,SH;jqH;��H;ѝH;��H;%�H;J�H;�H;�H;��H;d�H;��H;��H;��H;��H;��H;��H;��H;c�H;��H;�H; �H;H�H;%�H;��H;ѝH;��H;fqH;(SH;�-H;v�G;��G;�G; F;CD;=A;�g<;%5;<�*;�;>`;���:�P�:�P�:��:@�8�ڷ�T�=�� ��X��      �1��*Ȅ�˨u��PV�z.�����W��(��X�9P+i: ��:-,�:0�;�t%;�J2;m;;ĵ@;D;F;:G;��G;�H;�5H;�ZH;FxH;P�H;;�H;(�H;$�H;k�H;~�H;*�H;?�H;9�H;M�H;g�H;��H;g�H;M�H;9�H;>�H;,�H;~�H;j�H;!�H;'�H;7�H;S�H;FxH;�ZH;�5H;�H;��G;<G;F;�D;µ@;o;;�J2;�t%;0�;+,�: ��:X+i:�X�98��W�����s.��PV�˨u�.Ȅ�      Z��J�	������$Tʻ�R��3|�_.�Ⱥ����Y�9Ru�:��:�Y;��!;��0; �:;ĵ@;CD;�2F;�8G;��G;�H;{@H;7dH;րH;��H;W�H;Y�H;]�H;��H; �H;��H;~�H;��H;�H;��H;�H;��H;~�H;��H; �H;��H;[�H;V�H;W�H;��H;׀H;8dH;x@H;�H;��G;�8G;�2F;CD;Ƶ@;��:;��0;��!;�Y;��:Ru�:�Y�9���Ⱥ`.�3|��R��#Tʻ�����M�	�      ªx��[t���g�ST�`�:�������+����1��G�(�W��@�t�Do`:���: ];!{ ;��0;r;;=A;*�D;�wF;�cG;f�G;�!H;�MH;�oH;��H;��H;ԯH;��H;u�H;��H;h�H;}�H;�H;��H;3�H;��H;�H;}�H;g�H;��H;u�H;��H;ϯH;��H;��H;�oH;�MH;�!H;d�G;�cG;�wF;*�D;=A;s;;��0;!{ ; ];���:Do`:@�t�W��G�(��1��,���������`�:�ST���g��[t�      ;,˼��Ǽ�"���뮼w��'G��.�[�cy-�����.��ĕb�X0�ط�V5<:M�:�\;��!;�J2;�g<;d0B;?CE;=�F;a�G;�G;�4H;�\H;|H;��H;��H;i�H;��H;O�H;��H;a�H;a�H;�H;��H;�H;`�H;_�H;��H;R�H;��H;g�H;��H;��H;|H;�\H;�4H;�G;\�G;=�F;?CE;f0B;�g<;�J2;��!;�\;M�:V5<:ط�Z0�ĕb��.�����dy-�.�[�'G��w���뮼�"����Ǽ      .���k��Lv��t�F�Ѽ�뮼.X��p�W������׻�Ǆ�
�����b5<:���:�Y;�t%;%5;�Z>;aC;��E;G*G;v�G;&H;HH;~lH;�H;�H;үH;߼H;��H;��H;�H;��H;}�H;=�H;}�H;��H;�H;��H;��H;߼H;үH;�H;�H;|lH;HH;'H;t�G;C*G;��E;aC;�Z>;%5;�t%;�Y;���:^5<:���	���Ǆ���׻���p�W�/X���뮼F�Ѽ�t�Lv���k�      Hm��Fi��&^�b�L�S�6�*����#}ռqT����x���0����������׷�Ho`:��:2�;>�*;L�8;"�@;K�D;z�F;~G;��G;�1H;�[H;~|H;͕H;�H;��H;��H;��H;��H;��H;��H;��H;��H;��H;��H;��H;��H;��H;�H;˕H;~|H;�[H;�1H;��G;�}G;v�F;K�D;%�@;N�8;>�*;4�;��:Ho`:�׷�
����������0���x�qT��#}ռ��*��S�6�b�L��&^��Fi�      P��u;��C�������섽|�e��?��k�t�鷼G���e7�����Ǆ�T0���t�Tu�:1,�:�;�1;f�<;w�B;9�E;G;�G;pH;�JH;moH;�H;��H;"�H;��H;��H;.�H;��H;�H;��H;�H;��H;+�H;��H;��H;"�H;��H;�H;moH;�JH;rH;�G;G;6�E;w�B;h�<;�1;�;7,�:Ru�:@�t�T0��Ǆ���껅e7�G��鷼t��k��?�|�e��섽���C���u;��      t���(��s��ӽ�'��B�������Z��Q+�����"��G����0���׻b�W���Y�9��:>`;�*';�Y7; $@;;�D;�F;"�G;��G;H8H;bH;�H;f�H;��H;�H;��H;��H;��H;\�H;H�H;\�H;��H;��H;��H;��H;��H;f�H;	�H;bH;G8H;��G;'�G;�F;8�D; $@;�Y7;�*';>`;��:�Y�9W��b���׻»0�G���"������Q+��Z����B����'���ӽ�s�(��      �!,�;)��K ��������޽ ������Fi��0����鷼��x�����.��E�(����X+i:���:Q�;��0;`�<;�C;��E;=G;�G;%H;sTH;�wH;��H;%�H;Y�H;��H;L�H;��H;��H;��H;��H;��H;L�H;��H;Y�H;%�H;��H;�wH;sTH;%H;�G;=G;��E;�C;`�<;��0;P�;���:\+i:���F�(��.�������x�鷼����0��Fi���� ���޽�������K �;)�      ,�j��f��Z�|�F��>/��^�r����ŽI ���Fi��Q+�~t�qT��q�W�����1�� Ⱥ�X�9�P�:�Y;��(;�8;A;�E;�F;y�G;�H;�FH;�mH;��H;ΡH;K�H;{�H;��H;��H;�H;�H;�H;��H;��H;x�H;K�H;ΡH;��H;�mH;�FH;�H;{�G;�F;�E;A;�8;��(;�Y;�P�:�X�9Ⱥ�1�����p�W�qT��~t�Q+��Fi�I ���Žr����^��>/�|�F��Z��f�      ��x���{�J����f��SC��K �rn���Ž����Z��k�"}ռ.X��by-�)���].� ���P�:�+�:��;14;I�>;D;�wF;C�G;��G;�9H;edH;��H;��H;n�H;|�H;��H;��H;`�H;}�H;b�H;��H;��H;y�H;n�H;��H;��H;ddH;�9H;��G;B�G;�wF;	D;I�>;14;��;�+�:�P�:���_.�*���by-�.X��"}ռ�k��Z�����Žrn���K ��SC��f�J���{�x���      ��˾��Ǿ����!���X͓�^�x���J��K �r��� ������?����뮼-�[����3|�|W����:��:�';�/;xg<;�C;yF;�NG;��G;<-H;{[H;�}H;ӗH;ӪH;ʸH;��H;�H;��H;�H;��H;�H;��H;ǸH;ӪH;ӗH;�}H;{[H;<-H;��G;�NG;}F;�C;vg<;�/;�';��:��:xW��3|����-�[��뮼���?���� ��r����K ���J�^�x�X͓�!���������Ǿ      u� ��������{Ծm���x���^�x��SC��^��޽B���|�e�*��F�Ѽ'G������R�����@�8��:�Y;c�); �9;�A;˄E;�G;-�G;u!H;OSH;�wH;��H;��H;O�H;��H;��H;��H;��H;��H;��H;��H;M�H;��H;��H;�wH;KSH;v!H;+�G;�G;΄E;
�A;�9;c�);�Y;��:@�8����R�����'G��F�Ѽ*��|�e�B����޽�^��SC�^�x�x���m����{Ծ�쾣���      ��� E�l�u� �Y�ݾm���X͓��f��>/�����'���섽R�6��t�w��_�:�!Tʻr.��ڷ��t�:�;��$;�Y7;h�@;
E;-�F;G�G;�H;LLH;�rH;��H;ؤH;1�H;/�H;@�H;X�H;��H;X�H;?�H;/�H;.�H;ڤH;H;�rH;ILH;�H;I�G;,�F;	
E;f�@;�Y7;��$;�;�t�:�ڷ�q.�"Tʻ_�:�w���t�R�6��섽�'������>/��f�X͓�m���Y�ݾu� �l� E�      ��7�v3�1�'����u� ��{Ծ!���J���|�F�����ӽ���b�L�Lv��뮼ST����PV�X�=�*i:���:�z ;�$5;��?;�D;޺F;�G;�H;�FH;�nH;��H;��H;~�H;�H;F�H;e�H;�H;e�H;F�H;�H;|�H;��H;��H;�nH;�FH;�H;�G;޺F;�D;��?;�$5;�z ;���:*i:X�=��PV���ST��뮼Lv�b�L�����ӽ���|�F�J���!����{Ծu� ����1�'�v3�      �N��TI���;�1�'�l��쾂���{󐾷Z��K ��s�C����&^���"����g����̨u�� ��v3<:)��:;xg3;�>;�BD;ĖF;��G;�H;YBH;�kH;f�H;�H;;�H;�H;~�H;��H;V�H;��H;~�H;�H;9�H;�H;f�H;�kH;VBH;�H;��G;ƖF;�BD;��>;{g3;;-��:z3<:� ��˨u������g��"����&^�C����s潧K ��Z�{󐾂�����l�1�'���;��TI�      c]�g�W��TI�v3� E�������Ǿx����f�;)�(��u;���Fi��k���Ǽ�[t�L�	�(Ȅ� X��|�:��:��;kJ2;`Z>;W	D;�F;Q�G;(H;�?H;�iH;��H;�H;��H;J�H;��H;h�H;��H;h�H;��H;J�H;��H;�H;��H;�iH;�?H;(H;P�G;�F;W	D;]Z>;qJ2;��;��:t�: X��'Ȅ�L�	��[t���Ǽ�k��Fi�u;��(��;)��f�x�����Ǿ���� E�v3��TI�g�W�      �?��~h��?v��� ��9�X��O/�2y�C�;Ⱆ��+X����ѽ����bn;�^�������B(�՚��0��p�e9.�:;�Y.;`�<;�WC;0[F;�G;50H;|jH;^�H;}�H;��H;Y�H;��H;��H;��H;��H;��H;��H;��H;X�H;õH;}�H;]�H;yjH;50H;�G;2[F;�WC;^�<;�Y.;;0�:`�e90��Ԛ���B(�����^��bn;������ѽ���+X�Ⱆ�C�;2y��O/�9�X�� ��?v��~h��      ~h��1���c�����y�YvS�rM+��v�9ɾ�����T�"]�\ν����{\8�����x��%�H���N����9�-�:��;��.;)�<;oC;�dF;��G;�1H;)kH;ьH;ۤH;�H;��H;�H;��H;�H;��H;�H;��H;�H;��H;�H;ۤH;ΌH;%kH;�1H;��G;�dF;oC;%�<;��.;��;�-�:��9N��H���%��x�����{\8�����\ν"]��T�����9ɾ�v�rM+�YvS���y�c���1���      ?v��c���X ��c�h�9E�Z��m���~㼾~���nH�Ո�|�ý�Ȅ��s/��o��#�����J�� к�
�9ng�:m;d0;/]=;�C;*�F;��G;R6H;emH;Q�H;٥H;��H;0�H;x�H;�H;:�H;�H;:�H;�H;x�H;-�H;��H;٥H;M�H;bmH;R6H;��G;+�F;�C;,]=;f0;m;jg�:�
�9 кJ������#���o��s/��Ȅ�|�ýՈ��nH�~��~㼾m���Z��9E�c�h�X ��c���      � ����y�c�h��N��O/����E�߾B���*|��6�r}�䳽mSt�?�!�rrμAF{��_��X������ :G��:[;�2;�O>;�D;w�F;��G;M=H;�pH;��H;�H;�H;�H;�H;��H;��H;��H;��H;��H;�H;�H;�H;�H;��H;�pH;M=H;��G;v�F;�D;�O>;�2;[;G��: :�����X���_�AF{�rrμ?�!�mSt�䳽r}��6��*|�B��E�߾����O/��N�c�h���y�      9�X�YvS�9E��O/��S�KW����������OS\��� ���<����Y�|��҃����]�}����b�@�Y��Y:��:�`;r�4;�?;n�D;�F;*�G;7FH;�uH;�H;ĩH;��H;G�H;��H;X�H;M�H;.�H;M�H;V�H; �H;F�H;��H;ĩH;�H;�uH;7FH;,�G;�F;m�D;��?;v�4;�`;��:��Y:D�Y��b�~�����]�҃��|���Y�<����当� �OS\���������KW���S��O/�9E�YvS�      �O/�rM+�Y�����KW��9ɾB���Mw�� :�k��z�ý�L��_n;�a���uv���E<��˻��-�`���y�:�^;�%;��7;��@;I5E;�"G;)�G;mPH;={H;�H;��H;��H;��H;,�H;E�H;�H;��H;�H;E�H;,�H;��H;��H;��H;�H;9{H;lPH;'�G;�"G;H5E;��@;��7;�%;�^;�y�:`����-��˻�E<�uv��a���_n;��L��z�ýk��� :��Mw�B��9ɾKW�����Y��rM+�      2y��v�m���E�߾����B��@����nH���FὟu����d�1O�lrμJ"������������s89�;�:u�;�+;�|:;�7B;�E;?bG;�H;![H;��H;T�H;ЯH;,�H;z�H;{�H;>�H;�H;��H;�H;>�H;|�H;y�H;.�H;ЯH;S�H;��H;![H;�H;@bG;�E;�7B;�|:;�+;w�;�;�:�s89|��������J"��lrμ1O���d��u��F����nH�@���B������E�߾m����v�      C�;9ɾ~㼾B�������Mw��nH�����Z�䳽̕��t\8�r#������^N�H���b��Hx��5:@��:H�;�0;T]=;b�C;�[F;�G;	*H;fH;��H;N�H;t�H;��H;N�H;�H;c�H;�H;��H;�H;c�H;�H;M�H;��H;u�H;N�H;��H;fH;*H;�G;�[F;_�C;T]=;�0;H�;>��:�5:�Hx��b�H��^N�����r#��t\8�̕��䳽�Z񽲯��nH��Mw�����B��~㼾9ɾ      Ⱆ�����~���*|�OS\�� :����Z�n$�������K�w���Oļ����������(&�p���/�:�^;��#;�G6;o�?;�D;~�F;��G;+@H;�pH;�H;��H;G�H;��H;`�H;��H;��H;	�H;��H;	�H;��H;��H;`�H;��H;G�H;��H;�H;�pH;)@H;��G;{�F;�D;n�?;�G6;��#;�^;�/�:p��(&������������Oļw���K�����n$���Z���� :�OS\��*|�~������      �+X��T��nH��6��� �k��F�䳽�����mR����ټ�����E<��?ݻ%d\�����T!:�d�:��;H�,;��:;�7B;��E;�LG;lH;�SH;�{H;��H;�H;H�H;r�H;��H;B�H;��H;%�H;��H;'�H;��H;C�H;��H;u�H;I�H;�H;��H;�{H;�SH;lH;�LG;��E;�7B;��:;H�,;��;�d�:T!:����%d\��?ݻ�E<�����ټ����mR�����䳽F�k���� ��6��nH��T�      ��"]�Ո�r}���z�ý�u��̕���K�����o�kv���&R���N^��R�� >�0��:�B;k";��4;��>;vD;��F;*�G;*H;�dH;��H;G�H;��H;`�H;b�H;��H;��H;U�H;A�H;�H;A�H;U�H;��H;��H;e�H;`�H;��H;D�H;��H;�dH;*H;'�G;��F;sD;��>;��4;i";�B;6��: $>�R��N^�����&R�kv���o�����K�̕���u��z�ý��r}�Ո�"]�      �ѽ\ν|�ý䳽=����L����d�t\8�w��ټkv����Y��_�����*��P[��Y:���:om;�r-;0�:;��A;doE;�"G;��G;�GH;�sH;�H;��H;�H;^�H;L�H;��H;��H;��H;[�H;�H;[�H;��H;��H;��H;O�H;^�H;�H;��H;�H;�sH;�GH;��G;�"G;boE;��A;0�:;�r-;qm;���:�Y:T[�+�������_���Y�kv��ټw��t\8���d��L��=���䳽|�ý\ν      ���������Ȅ�mSt��Y�_n;�2O�r#���Oļ�����&R��_������N3�|�Y�T4:J�:�;	@&;H6;�X?;�D;_xF;�G;f!H;�^H;��H;"�H;�H;s�H;9�H;/�H;�H;C�H;�H;��H;A�H;��H;�H;C�H;�H;0�H;9�H;s�H;�H;"�H;��H;�^H;d!H;�G;[xF;�D;�X?;H6;	@&;�;F�:\4:|�Y��N3������_��&R������Oļs#��2O�_n;��Y�mSt��Ȅ�����      bn;�z\8��s/�?�!�|��a���lrμ��������E<��������N3��Gx���9*�:_;r ;R2;��<;�B;ٲE;d5G;5�G;dFH;�qH;ӎH;|�H;�H;~�H;��H;��H;0�H;��H;L�H;��H;;�H;��H;L�H;��H;/�H;��H;��H;~�H;�H;|�H;ҎH;�qH;cFH;2�G;^5G;ٲE;�B;��<;R2;t ;_;.�:��9�Gx��N3��������E<��������lrμ`���|��?�!��s/�{\8�      ^������o�srμӃ��vv��K"��^N�����?ݻO^��/����Y�x�9$�:��:�;p�.;�|:;?A;��D;Y�F;�G;*H;MaH;G�H;��H;�H;k�H;N�H;k�H;��H;+�H;J�H;��H;��H;�H;��H;��H;L�H;*�H;��H;k�H;M�H;h�H;�H;��H;J�H;LaH;*H;޶G;X�F;��D;?A;�|:;s�.;�;��:$�:p�9��Y�/��O^���?ݻ���^N�K"��uv��Ӄ��srμ�o����      �����x���#��AF{���]��E<����J�뻢���&d\�V��X[�P4:(�:��:�[;��,;
�8;E!@; 1D;�[F;O{G;$H;tPH;HvH;�H;q�H;.�H;_�H;��H;��H;
�H;�H;��H;��H;��H;��H;��H;��H;��H;
�H;�H;��H;��H;[�H;.�H;o�H;�H;GvH;pPH; H;M{G;�[F; 1D;D!@;�8;��,;�[;��:*�:P4:X[�V��(d\�����J�뻢���E<���]�AF{��#���x��      �B(� %�����_�����˻�����b�*&�����  >��Y:D�:_;�;��,;4`8;��?;�C;�F;GG;x�G;"@H;YkH;1�H;6�H;#�H;��H;��H;��H;��H;L�H;��H;�H;��H;��H;��H;��H;��H;�H;��H;M�H;��H;��H;��H;��H;!�H;9�H;1�H;TkH;@H;x�G;GG;�F;�C;��?;3`8;��,;�;_;D�:�Y: $>�����(&���b�����˻~����_����%�      ٚ��L���J���X���b���-�����Hx����T!:0��:���:�;p ;q�.;�8;��?; �C;��E;f#G;�G;2H;bH;y�H;��H;��H;ݷH;�H;��H;J�H;h�H;j�H;�H;H�H;��H;j�H;��H;j�H;��H;H�H;�H;k�H;h�H;H�H;��H;�H;ڷH;��H;��H;v�H;bH;2H;�G;g#G;��E;"�C;��?;�8;p�.;p ;�;���:0��:L!:p���Hx������-��b��X��J��P���      ,��T���к����X�Y�P�� t89�5:~/�:�d�:�B;om;@&;R2;�|:;C!@;�C;��E;�G;	�G;�(H;+[H;�zH;n�H;�H;ҳH;��H;��H;��H;��H;��H;-�H;�H;_�H;~�H;-�H;��H;/�H;~�H;_�H;}�H;.�H;��H;��H;��H;��H;��H;ԳH;�H;k�H;�zH;+[H;�(H;
�G;�G;��E;�C;C!@;�|:;R2;@&;qm;�B;�d�:�/�:�5: t89 ��D�Y������кT��      `�e9@�9�
�9�:��Y:�y�:�;�:2��:�^;��;h";�r-;�G6;��<;?A;�0D;�F;b#G;�G;%H;�WH;�vH;��H;s�H;y�H;��H;A�H;��H;��H;l�H;�H;��H;��H;\�H;@�H;��H;,�H;��H;@�H;\�H;��H;��H;�H;i�H;��H;��H;@�H;��H;y�H;o�H;��H;�vH;�WH;%H;�G;c#G;�F;�0D;?A;��<;�G6;�r-;h";��;�^;8��:�;�:�y�:(�Y:  :�
�9�9      <�:�-�:pg�:3��:��:�^;x�;D�;��#;H�,;��4;,�:;�X?;�B;��D;�[F;GG;�G;�(H;�WH;�uH;��H;G�H;.�H;V�H;-�H;��H;!�H;�H;��H;��H;�H;��H;"�H; �H;��H;��H;��H; �H;"�H;��H;�H;��H;��H;�H;!�H;��H;-�H;U�H;)�H;G�H;��H;�uH;�WH;�(H;�G;GG;�[F;��D;�B;�X?;,�:;��4;H�,;��#;D�;x�;�^;��:9��:rg�:�-�:      ;��;m;[;�`;�%;�+;�0;�G6;��:;��>;��A;�D;زE;Y�F;L{G;x�G;2H;*[H;�vH;��H;�H;��H;�H;��H;��H;��H;��H;��H;�H;r�H;l�H;��H;��H;��H;��H;�H;��H;��H;��H;��H;l�H;r�H;�H;��H;��H;��H;��H;��H;��H;��H;�H;��H;�vH;*[H;2H;v�G;L{G;[�F;زE;�D;��A;��>;��:;�G6;�0;�+;�%;�`;[;m;��;      �Y.;��.;e0;�2;n�4;��7;�|:;U]=;q�?;�7B;tD;foE;\xF;a5G;߶G; H; @H;bH;�zH;��H;G�H;��H;~�H;�H;��H;��H;��H;-�H;T�H;��H;��H;��H;��H;z�H;!�H;T�H;~�H;T�H;!�H;|�H;��H;��H;��H;��H;Q�H;-�H;��H;��H;��H;��H;~�H;��H;B�H;��H;�zH;bH;@H;H;߶G;a5G;\xF;foE;vD;�7B;r�?;U]=;�|:;��7;v�4;�2;e0;��.;      r�<;9�<;7]=;�O>;�?;��@;�7B;`�C;�D;��E;��F;�"G;�G;6�G;*H;qPH;VkH;z�H;k�H;q�H;)�H;��H;�H;m�H;j�H;n�H;��H;��H;X�H;p�H;0�H;D�H;A�H;�H;w�H;��H;��H;��H;x�H;�H;>�H;E�H;2�H;o�H;U�H;��H;~�H;n�H;k�H;j�H;�H; �H;'�H;q�H;k�H;|�H;TkH;qPH;*H;5�G;�G;�"G;��F;��E;�D;b�C;�7B;��@;�?;�O>;7]=;)�<;      �WC;oC;��C;�D;o�D;L5E;�E;�[F;~�F;�LG;*�G;��G;f!H;iFH;OaH;JvH;8�H;��H;�H;��H;Y�H;��H;��H;q�H;-�H;?�H;x�H;��H; �H;��H;�H;��H;��H;l�H;��H;�H;�H;�H;��H;j�H;��H;��H;�H;��H;�H;��H;x�H;?�H;0�H;o�H;��H;��H;X�H;��H;�H;��H;4�H;HvH;OaH;fFH;f!H;��G;*�G;�LG;��F;�[F;�E;L5E;r�D;�D;��C;oC;      <[F;�dF; �F;t�F;�F;�"G;@bG;�G;��G;lH;*H;�GH;�^H;�qH;F�H;�H;6�H;��H;ϳH;��H;*�H;��H;��H;n�H;8�H;c�H;��H;��H;��H;��H;��H;��H;[�H;��H;	�H;J�H;J�H;J�H;�H;��H;X�H;��H;��H;��H;��H;��H;��H;d�H;<�H;n�H;��H;��H;&�H;��H;ϳH;��H;5�H;�H;F�H;�qH;�^H;�GH;*H;lH;��G;�G;@bG;�"G;�F;t�F;�F;�dF;      �G;�G;��G;��G;0�G;0�G;�H;*H;.@H;�SH;�dH;�sH;��H;ՎH;��H;q�H;%�H;ڷH;��H;D�H;��H;��H;��H;��H;r�H;��H;��H;z�H;��H;��H;��H;/�H;��H;�H;<�H;m�H;��H;m�H;:�H;�H;��H;.�H;��H;��H;��H;x�H;��H;��H;v�H;��H;��H;��H;��H;C�H;��H;۷H;#�H;p�H;��H;ӎH;��H;�sH;�dH;�SH;0@H;*H;�H;+�G;6�G;��G;��G;�G;      ,0H;�1H;Z6H;F=H;=FH;oPH;&[H;fH;�pH;�{H;��H;#�H;%�H;~�H;�H;.�H;��H;�H;��H;��H;!�H;��H;-�H;��H;��H;��H;w�H;��H;��H;��H;6�H;��H;��H;F�H;z�H;��H;~�H;��H;z�H;F�H;��H;��H;8�H;��H;��H;��H;w�H;��H;��H;��H;-�H;��H;�H;��H;��H;�H;��H;.�H;�H;}�H;"�H;!�H;��H;�{H;�pH; fH;&[H;pPH;HFH;G=H;Y6H;�1H;      �jH;,kH;emH;�pH;�uH;<{H;��H;��H;�H;��H;H�H;ŦH;�H;�H;k�H;_�H;��H;��H;��H;��H;�H;��H;Q�H;[�H;�H;��H;��H;��H;��H;$�H;��H;��H;,�H;i�H;��H;��H;��H;��H;��H;i�H;)�H;��H;��H;$�H;��H;��H;��H;��H;�H;[�H;P�H;��H;�H;��H;��H;��H;��H;_�H;k�H;�H;�H;ĦH;G�H;��H;�H;��H;��H;<{H;�uH;�pH;emH; kH;      l�H;،H;[�H;��H;��H;�H;[�H;U�H;��H;�H;��H;(�H;z�H;��H;Q�H;��H;��H;F�H;��H;o�H;��H;�H;��H;s�H;��H;��H;��H;��H;#�H;�H;��H;2�H;i�H;��H;��H;��H;��H;��H;��H;��H;f�H;3�H;��H;�H;#�H;��H;��H;��H;��H;r�H;��H;�H;��H;o�H;��H;G�H;��H;��H;Q�H;��H;z�H;&�H;��H;�H;��H;W�H;[�H;�H;��H;��H;V�H;ԌH;      ��H;�H;�H;��H;ԩH;��H;گH;��H;O�H;N�H;g�H;j�H;>�H;��H;n�H;��H;��H;h�H;��H;�H;��H;r�H;��H;5�H;�H;��H;��H;9�H;��H;��H;.�H;_�H;��H;��H;��H;��H;��H;��H;��H;��H;��H;`�H;.�H;��H;��H;;�H;��H;��H;�H;5�H;��H;r�H;��H;�H;��H;h�H;��H;��H;n�H;��H;=�H;g�H;g�H;P�H;P�H;��H;گH;��H;ѩH;��H;�H;�H;      ԵH; �H;˶H;�H;ǹH;��H;0�H;��H;��H;w�H;j�H;W�H;4�H;��H;��H;�H;T�H;k�H;1�H;��H;�H;q�H;��H;I�H;��H;��H;.�H;��H;��H;3�H;]�H;x�H;��H;��H;��H;��H;��H;��H;��H;��H;��H;z�H;]�H;6�H;��H;��H;/�H;��H;��H;I�H;��H;q�H;�H;��H;1�H;m�H;S�H;�H;��H;��H;3�H;T�H;i�H;u�H;��H;��H;2�H;��H;ƹH;�H;ʶH;�H;      _�H;��H;:�H;�H;S�H;��H;}�H;V�H;e�H;��H;��H;��H;�H;6�H;/�H;�H;��H;�H;��H;��H;��H;��H;��H;H�H;��H;[�H;��H;��H;/�H;m�H;��H;��H;��H;��H;��H;��H;��H;��H;��H;��H;��H;��H;��H;p�H;0�H;��H;��H;[�H;��H;H�H;��H;��H;��H;��H;��H;�H;��H;�H;-�H;6�H;�H;��H;��H;��H;g�H;U�H;|�H;��H;L�H;�H;9�H;��H;      ��H;�H;t�H;�H;�H;(�H;��H;�H;��H;E�H;�H;��H;F�H;��H;P�H;��H;�H;I�H;c�H;d�H;)�H;��H;z�H;�H;e�H;��H;�H;F�H;i�H;��H;��H;��H;��H;��H;��H;��H;��H;��H;��H;��H;��H;��H;��H;��H;k�H;F�H;�H;��H;f�H;�H;z�H;��H;(�H;d�H;c�H;J�H;�H;��H;O�H;��H;F�H;��H;�H;E�H;��H;�H;��H;.�H;��H;�H;t�H;�H;      ��H;��H;�H;��H;q�H;@�H;F�H;p�H;��H; �H;\�H;��H;�H;T�H;��H;��H;��H;��H;��H;H�H;�H;��H; �H;}�H;��H;�H;6�H;z�H;��H;��H;��H;��H;��H;��H;��H;��H;��H;��H;��H;��H;��H;��H;��H;��H;��H;z�H;6�H;�H;��H;{�H;!�H;��H;�H;H�H;��H;��H;��H;��H;��H;T�H;�H;��H;[�H;�H;��H;m�H;E�H;D�H;g�H;��H;�H;��H;      ��H;�H;C�H;��H;\�H;�H;�H;�H;�H;%�H;I�H;e�H;��H;��H;��H;��H;��H;g�H;3�H;��H;��H;��H;T�H;��H;�H;G�H;j�H;��H;��H;��H;��H;��H;��H;��H;��H;��H;��H;��H;��H;��H;��H;��H;��H;��H;��H;��H;j�H;F�H;�H;��H;T�H;��H;��H;��H;3�H;i�H;��H;��H;��H;��H;��H;e�H;H�H;)�H;�H;
�H;�H;�H;Q�H;��H;C�H;�H;      ��H;��H;&�H;��H;?�H;��H;��H;��H;��H;��H;
�H;*�H;G�H;D�H;�H;��H;��H;��H;��H;3�H;��H;�H;}�H;��H;�H;F�H;��H;��H;��H;��H;��H;��H;��H;��H;��H;��H;��H;��H;��H;��H;��H;��H;��H;��H;��H;��H;��H;G�H;�H;��H;}�H;�H;��H;3�H;��H;��H;��H;��H;�H;D�H;G�H;*�H;
�H;��H;��H;��H;��H;��H;2�H;��H;&�H;��H;      ��H;�H;C�H;��H;\�H;�H;�H;�H;�H;%�H;I�H;e�H;��H;��H;��H;��H;��H;g�H;3�H;��H;��H;��H;T�H;��H;�H;G�H;k�H;��H;��H;��H;��H;��H;��H;��H;��H;��H;��H;��H;��H;��H;��H;��H;��H;��H;��H;��H;j�H;F�H;�H;��H;T�H;��H;��H;��H;3�H;i�H;��H;��H;��H;��H;��H;e�H;I�H;'�H;�H;
�H;�H;�H;Q�H;��H;?�H;�H;      ��H;��H;�H;��H;r�H;@�H;F�H;p�H;��H; �H;[�H;��H;�H;T�H;��H;��H;��H;��H;��H;H�H;�H;��H; �H;}�H;��H;�H;6�H;z�H;��H;��H;��H;��H;��H;��H;��H;��H;��H;��H;��H;��H;��H;��H;��H;��H;��H;z�H;6�H;�H;��H;z�H;!�H;��H;�H;H�H;��H;��H;��H;��H;��H;T�H;�H;��H;[�H;�H;��H;m�H;F�H;D�H;g�H;��H;�H;��H;      ��H;�H;t�H;�H;�H;(�H;��H;�H;��H;E�H;�H;��H;F�H;��H;O�H;��H;�H;I�H;c�H;d�H;-�H;��H;z�H;�H;f�H;��H;�H;F�H;i�H;��H;��H;��H;��H;��H;��H;��H;��H;��H;��H;��H;��H;��H;��H;��H;k�H;F�H;�H;��H;e�H;�H;z�H;��H;)�H;d�H;c�H;J�H;�H;��H;Q�H;��H;F�H;��H;�H;E�H;��H;�H;��H;,�H;��H;�H;t�H;�H;      b�H;��H;;�H;�H;P�H;��H;|�H;U�H;e�H;��H;��H;��H;�H;6�H;-�H;�H;��H;�H;��H;��H;��H;��H;��H;H�H;��H;\�H;��H;��H;/�H;n�H;��H;��H;��H;��H;��H;��H;��H;��H;��H;��H;��H;��H;��H;n�H;0�H;��H;��H;[�H;��H;F�H;��H;��H;��H;��H;��H;�H;��H;�H;/�H;6�H;�H;��H;��H;��H;e�H;T�H;}�H;��H;J�H;�H;9�H;��H;      յH; �H;̶H;�H;ƹH;��H;3�H;��H;��H;w�H;i�H;V�H;3�H;��H;��H;�H;U�H;k�H;1�H;��H;�H;q�H;��H;K�H;��H;��H;.�H;��H;��H;5�H;]�H;x�H;��H;��H;��H;��H;��H;��H;��H;��H;��H;z�H;]�H;5�H;��H;��H;/�H;��H;��H;I�H;��H;q�H;�H;��H;1�H;m�H;S�H;�H;��H;��H;4�H;V�H;j�H;x�H;��H;��H;3�H;��H;ùH;�H;̶H;�H;      ��H;�H;�H;��H;ԩH;��H;گH;��H;O�H;O�H;g�H;g�H;=�H;��H;p�H;��H;��H;g�H;��H;�H;��H;r�H;��H;6�H;�H;��H;��H;;�H;��H;��H;.�H;_�H;��H;��H;��H;��H;��H;��H;��H;��H;��H;`�H;.�H;��H;��H;9�H;��H;��H;�H;5�H;��H;r�H;��H;�H;��H;h�H;��H;��H;n�H;��H;>�H;j�H;e�H;O�H;O�H;��H;گH;��H;ЩH;��H;�H;�H;      e�H;،H;Y�H;��H;��H;�H;]�H;W�H;��H;�H;��H;(�H;y�H;��H;Q�H;��H;��H;F�H;��H;p�H;��H;�H;��H;s�H;��H;��H;��H;��H;$�H;��H;��H;2�H;g�H;��H;��H;��H;��H;��H;��H;��H;g�H;3�H;��H;~�H;#�H;��H;��H;��H;��H;r�H;��H;�H;��H;o�H;��H;G�H;��H;��H;Q�H;��H;y�H;(�H;��H;�H;��H;W�H;]�H;�H;��H;��H;[�H;׌H;      �jH;(kH;kmH;�pH;�uH;8{H;��H;��H;�H;��H;H�H;ŦH;�H;�H;k�H;_�H;��H;��H;��H;��H;�H;��H;Q�H;[�H;�H;��H;��H;��H;��H;&�H;��H;��H;+�H;i�H;��H;��H;��H;��H;��H;i�H;+�H;��H;��H;#�H;��H;��H;��H;��H;�H;[�H;P�H;��H;�H;��H;��H;��H;��H;a�H;k�H;�H;�H;ŦH;H�H;��H;�H;��H;��H;9{H;�uH;�pH;imH;(kH;      ,0H;�1H;Y6H;G=H;<FH;pPH;&[H;"fH;�pH;�{H;��H;!�H;"�H;~�H;�H;.�H;��H;�H;��H;��H;$�H;��H;.�H;��H;��H;��H;w�H;��H;��H;��H;8�H;��H;��H;D�H;x�H;��H;~�H;��H;z�H;F�H;��H;��H;6�H;��H;��H;��H;w�H;��H;��H;��H;+�H;��H;�H;��H;��H;�H;��H;/�H;�H;}�H;%�H;#�H;��H;�{H;�pH;fH;&[H;lPH;EFH;F=H;Y6H;�1H;      �G;�G;��G;��G;,�G;*�G;�H;*H;.@H;�SH;�dH;�sH;��H;ӎH;��H;q�H;%�H;ڷH;��H;F�H;��H;��H;��H;��H;v�H;��H;��H;x�H;��H;��H;��H;/�H;��H;�H;:�H;m�H;��H;k�H;<�H;�H;��H;1�H;��H;��H;��H;z�H;��H;��H;r�H;��H;��H;��H;��H;C�H;��H;۷H;#�H;p�H;��H;ՎH;��H;�sH;�dH;�SH;.@H;
*H;�H;*�G;0�G;��G;��G;��G;      C[F;�dF;'�F;t�F;�F;�"G;BbG;�G;��G;nH;*H;�GH;�^H;�qH;D�H;�H;6�H;��H;ϳH;��H;,�H;��H;��H;o�H;<�H;d�H;��H;��H;��H;��H;��H;��H;Z�H;��H;�H;J�H;J�H;J�H;�H;��H;X�H;��H;��H;��H;��H;��H;��H;c�H;8�H;l�H;��H;��H;&�H;��H;ϳH;��H;5�H;�H;F�H;�qH;�^H;�GH;*H;lH;��G;�G;CbG;�"G;�F;w�F;*�F;�dF;      �WC;oC;��C;�D;o�D;L5E;�E;�[F;��F;�LG;,�G;��G;f!H;fFH;OaH;JvH;7�H;��H;�H;��H;[�H;��H;��H;r�H;0�H;?�H;x�H;��H; �H;��H;�H;��H;��H;j�H;��H;�H;�H;�H;��H;j�H;��H;��H;�H;��H;�H;��H;x�H;?�H;-�H;o�H;��H;��H;X�H;��H;�H;��H;4�H;JvH;OaH;gFH;f!H;��G;*�G;�LG;~�F;�[F;�E;L5E;n�D;�D;��C;oC;      v�<;6�<;=]=;�O>;��?;��@;�7B;`�C;�D;²E;��F;�"G;�G;5�G;*H;qPH;VkH;y�H;k�H;q�H;+�H; �H;�H;o�H;k�H;n�H;��H;��H;X�H;r�H;2�H;D�H;?�H;�H;v�H;��H;��H;��H;x�H;�H;?�H;E�H;0�H;n�H;U�H;��H;~�H;n�H;j�H;j�H;�H;��H;'�H;q�H;k�H;|�H;TkH;qPH;*H;6�G;�G;�"G;��F;��E;�D;`�C;�7B;��@;�?;�O>;@]=;(�<;      �Y.;��.;r0;�2;j�4;��7;�|:;U]=;q�?;�7B;vD;foE;[xF;a5G;߶G; H; @H;bH;�zH;��H;H�H;��H;~�H;�H;��H;��H;��H;-�H;T�H;��H;��H;��H;��H;|�H;!�H;T�H;~�H;T�H;!�H;z�H;��H;��H;��H;��H;Q�H;-�H;��H;��H;��H;��H;~�H;��H;B�H;��H;�zH;bH; @H; H;�G;a5G;[xF;doE;tD;�7B;r�?;T]=;�|:;��7;p�4;�2;i0;��.;      ;��;m;[;�`;�%;�+;�0;�G6;��:;��>;��A;�D;زE;Y�F;M{G;v�G;2H;*[H;�vH;��H;�H;��H;�H;��H;��H;��H;��H;��H;�H;r�H;l�H;��H;��H;��H;��H;�H;��H;��H;��H;��H;l�H;r�H;�H;��H;��H;��H;��H;��H;��H;��H;�H;��H;�vH;*[H;2H;v�G;L{G;[�F;زE;�D;��A;��>;��:;�G6;
�0;�+;�%;�`;[;m;��;      0�:�-�:vg�:9��:��:�^;{�;H�;��#;H�,;��4;,�:;�X?;�B;��D;�[F;GG;�G;�(H;�WH;�uH;��H;G�H;/�H;U�H;-�H;��H;!�H;�H;��H;��H;�H;��H;!�H;��H;��H;��H;��H; �H;"�H;��H;�H;��H;��H;�H;!�H;��H;-�H;V�H;)�H;G�H;��H;�uH;�WH;�(H;�G;GG;�[F;��D;�B;�X?;,�:;��4;D�,;��#;H�;{�;�^;��:9��:xg�:�-�:      @�e9P�9�9�:�Y:�y�:�;�:4��:�^;��;h";�r-;�G6;��<;?A;�0D;�F;b#G;�G;%H;�WH;�vH;��H;t�H;y�H;��H;C�H;��H;��H;l�H;�H;��H;��H;\�H;@�H;��H;,�H;��H;@�H;\�H;��H;��H;�H;i�H;��H;��H;@�H;��H;y�H;o�H;��H;�vH;�WH;%H;�G;c#G;�F;�0D;?A;��<;�G6;�r-;f";��;�^;8��:�;�:�y�:�Y:�:�
�9��9      ,��T���к����`�Y�P�� t89�5:~/�:�d�:�B;qm;@&;R2;�|:;C!@;�C;��E;�G;	�G;�(H;+[H;�zH;p�H;�H;ӳH;��H;��H;��H;��H;��H;-�H;��H;_�H;~�H;-�H;��H;-�H;~�H;_�H;}�H;.�H;��H;��H;��H;��H;��H;ԳH;�H;j�H;�zH;+[H;�(H;
�G;�G;��E;�C;C!@;�|:;R2;@&;om;�B;�d�:�/�:�5: t89 ��H�Y������кT��      ؚ��L���J���X���b���-�����Hx����L!:0��:���:�;n ;p�.;�8;��?; �C;��E;f#G;�G;2H;bH;y�H;��H;��H;ݷH;�H;��H;J�H;h�H;j�H;�H;H�H;��H;j�H;��H;j�H;��H;H�H;�H;k�H;h�H;H�H;��H;�H;ڷH;��H;��H;v�H;bH;2H;�G;f#G;��E;!�C;��?;�8;q�.;p ;�;���:2��:T!:p���Hx������-��b��X��J��P���      �B(� %�����_������˻����b�)&����� >��Y:D�:_;�;��,;4`8;��?;�C;�F;GG;x�G;"@H;YkH;1�H;7�H;#�H;��H;��H;��H;��H;M�H;��H;�H;��H;��H;��H;��H;��H;�H;��H;M�H;��H;��H;��H;��H;�H;9�H;1�H;TkH;@H;x�G;GG;�F;�C;��?;4`8;��,;�;_;D�:�Y:  >�����(&���b�����˻����_����%�      �����x���#��AF{���]��E<����J�뻢���(d\�V��X[�P4:(�:��:�[;��,;
�8;D!@; 1D;�[F;M{G;#H;tPH;GvH;�H;q�H;.�H;_�H;��H;��H;
�H;�H;��H;��H;��H;��H;��H;��H;��H;�H;�H;��H;��H;[�H;.�H;o�H;�H;HvH;qPH; H;O{G;�[F; 1D;E!@;�8;��,;�[;��:(�:P4:X[�V��&d\�����J�뻢���E<���]�AF{��#���x��      ^������o�srμӃ��vv��K"��^N�����?ݻP^��.����Y�x�9$�:��:�;p�.;�|:;?A;��D;X�F;�G;*H;LaH;H�H;��H;�H;n�H;N�H;k�H;��H;+�H;L�H;��H;��H;�H;��H;��H;L�H;+�H;��H;k�H;M�H;h�H;�H;��H;J�H;MaH;*H;ݶG;Y�F;��D;?A;�|:;s�.;�;��:$�:x�9��Y�/��O^���?ݻ���^N�K"��uv��Ӄ��srμ�o����      bn;�z\8��s/�?�!�|��a���lrμ��������E<��������N3��Gx���9.�:_;r ;R2;��<;�B;ٲE;b5G;5�G;cFH;�qH;ӎH;|�H;�H;~�H;��H;��H;0�H;��H;L�H;��H;;�H;��H;L�H;��H;/�H;��H;��H;~�H;�H;|�H;ҎH;�qH;dFH;3�G;`5G;ٲE;�B;��<;R2;t ;_;*�:��9�Gx��N3��������E<��������lrμ`���|��?�!��s/�{\8�      ���������Ȅ�mSt��Y�_n;�2O�r#���Oļ�����&R��_������N3�|�Y�T4:J�:�;	@&;H6;�X?;�D;_xF;�G;d!H;�^H;��H;"�H;�H;s�H;9�H;0�H;�H;C�H;
�H;��H;A�H;��H;�H;C�H;�H;0�H;9�H;s�H;��H;"�H;��H;�^H;f!H;�G;[xF;�D;�X?;H6;	@&;�;F�:T4:|�Y��N3������_��&R������Oļs#��2O�_n;��Y�mSt��Ȅ�����      �ѽ\ν|�ý䳽=����L����d�t\8�w��ټkv����Y��_�����+��T[��Y:���:qm;�r-;.�:;��A;doE;�"G;��G;�GH;�sH;�H;��H;�H;^�H;L�H;��H;��H;��H;]�H;�H;]�H;��H;��H;��H;M�H;^�H;�H;��H;�H;�sH;�GH;��G;�"G;boE;��A;0�:;�r-;om;���:�Y:X[�*�������_���Y�kv��ټw��t\8���d��L��=���䳽|�ý\ν      ��"]�Ո�r}���z�ý�u��̕���K�����o�kv���&R���N^��R�� >�2��:�B;k";��4;��>;vD;��F;'�G;*H;�dH;��H;G�H;��H;`�H;b�H;��H;��H;U�H;A�H;�H;A�H;U�H;��H;��H;c�H;`�H;��H;D�H;��H;�dH;*H;*�G;��F;sD;��>;��4;i";�B;2��: $>�V��N^�����&R�kv���o�����K�̕���u��z�ý��r}�Ո�"]�      �+X��T��nH��6��� �k��F�䳽�����mR����ټ�����E<��?ݻ%d\�����L!:�d�:��;F�,;��:;�7B;��E;�LG;lH;�SH;�{H;��H;�H;I�H;t�H;��H;C�H;��H;%�H;��H;'�H;��H;B�H;��H;r�H;H�H;�H;��H;�{H;�SH;lH;�LG;��E;�7B;��:;H�,;��;�d�:X!:����&d\��?ݻ�E<�����ټ����mR�����䳽F�k���� ��6��nH��T�      Ⱆ�����~���*|�OS\�� :����Z�n$�������K�w���Oļ����������'&�����/�:�^;��#;�G6;o�?;�D;{�F;��G;+@H;�pH;�H;��H;G�H;��H;a�H;��H;��H;	�H;��H;	�H;��H;��H;^�H;��H;G�H;��H;�H;�pH;)@H;��G;~�F;�D;n�?;�G6;��#;�^;�/�:`��*&������������Oļw���K�����n$���Z���� :�OS\��*|�~������      C�;9ɾ~㼾B�������Mw��nH�����Z�䳽̕��t\8�r#������^N�H���b��Hx��5:>��:F�;�0;T]=;`�C;�[F;�G;	*H;fH;��H;N�H;u�H;��H;N�H;�H;e�H;�H;��H;�H;c�H;�H;M�H;��H;t�H;N�H;��H;fH;*H;�G;�[F;_�C;T]=;�0;H�;>��:�5:�Hx���b�H��^N�����r#��t\8�̕��䳽�Z񽲯��nH��Mw�����B��~㼾9ɾ      2y��v�m���E�߾����B��@����nH���FὟu����d�1O�lrμJ"������������s89�;�:u�;�+;�|:;�7B;�E;@bG;�H;![H;��H;T�H;ЯH;,�H;z�H;}�H;>�H;�H;��H;�H;>�H;{�H;y�H;,�H;ЯH;S�H;��H;![H;�H;@bG;�E;�7B;�|:;�+;w�;�;�:�s89~��������J"��lrμ1O���d��u��F����nH�@���B������E�߾m����v�      �O/�rM+�Y�����KW��9ɾB���Mw�� :�k��z�ý�L��_n;�a���uv���E<��˻��-�`���y�:�^;�%;��7;��@;H5E;�"G;*�G;lPH;={H;�H;��H;��H;��H;,�H;E�H;�H;��H;�H;E�H;,�H;��H;��H;��H;�H;9{H;mPH;'�G;�"G;I5E;��@;��7;�%;�^;�y�:`����-��˻�E<�uv��a���_n;��L��z�ýk��� :��Mw�B��9ɾKW�����Y��rM+�      9�X�YvS�9E��O/��S�KW����������OS\��� ���<����Y�|��҃����]�}����b�D�Y���Y:��:�`;r�4;�?;m�D;�F;*�G;7FH;�uH;�H;ĩH;��H;G�H; �H;X�H;M�H;.�H;M�H;U�H;��H;F�H;��H;ĩH;�H;�uH;7FH;,�G;�F;n�D;��?;v�4;�`;��:��Y:@�Y��b�~�����]�҃��|���Y�<����当� �OS\���������KW���S��O/�9E�YvS�      � ����y�c�h��N��O/����E�߾B���*|��6�r}�䳽mSt�?�!�rrμAF{��_��X������ :C��:[;�2;�O>;�D;v�F;��G;M=H;�pH;��H;�H;�H;�H;�H;��H;��H;��H;��H;��H;�H;�H;�H;�H;��H;�pH;M=H;��G;w�F;�D;�O>;�2;[;G��: :�����X���_�AF{�rrμ?�!�mSt�䳽r}��6��*|�B��E�߾����O/��N�c�h���y�      ?v��c���X ��c�h�9E�Y��m���~㼾~���nH�Ո�|�ý�Ȅ��s/��o��#�����J�� к�
�9jg�:m;d0;/]=;�C;*�F;��G;R6H;emH;O�H;٥H;��H;0�H;x�H;�H;:�H;�H;:�H;�H;x�H;-�H;��H;٥H;N�H;bmH;R6H;��G;+�F;�C;+]=;f0;m;jg�:�
�9 кJ������#���o��s/��Ȅ�|�ýՈ��nH�~��~㼾m���Y��9E�c�h�X ��c���      ~h��1���c�����y�YvS�rM+��v�9ɾ�����T�"]�\ν����{\8�����x��%�H���N����9�-�:��;��.;)�<;oC;�dF;��G;�1H;)kH;ьH;ۤH;�H;��H;�H;��H;�H;��H;�H;��H;�H;��H;�H;ۤH;ΌH;%kH;�1H;��G;�dF;oC;&�<;��.;��;�-�:��9N��H���%��x�����{\8�����\ν"]��T�����9ɾ�v�rM+�YvS���y�c���1���      gܿ5�ֿ�aǿ?^��1���[o���7����iþ�(���-=��` �A���_�2]�/p���I�K�ѻl�)�0�R���:L�
;�*;,�:;�B;NIF;:�G;�lH;>�H;��H;u�H;��H;��H;��H;��H;=�H;��H;=�H;��H;��H;��H;��H;u�H;��H;;�H;�lH;:�G;OIF;�B;)�:;�*;L�
;��:@�R�l�)�J�ѻ��I�/p��2]��_�A���` ��-=��(���iþ����7�[o�1���?^���aǿ5�ֿ      5�ֿFpѿ�¿������bXi�ѕ3��
�XD��Gl��D�9��.���R��#\� �ex��.�E��ͻ�$�����:Z�;��*;C�:;!�B;,UF;��G;^nH;ءH;�H;��H;��H;��H;��H;��H;Q�H;��H;Q�H;��H;��H;��H;��H;��H;�H;աH;^nH;��G;-UF;!�B;A�:;��*;Z�;�: ���$��ͻ.�E�ex�� �#\��R���.��D�9�Gl��XD���
�ѕ3�bXi��������¿Fpѿ      �aǿ�¿����������"Y��f'�����9o���.}��k/����'ڟ�%<Q�/#�ע��(;�&��� �� 07��:�;�,;��;;�C;LwF;-�G;�rH;e�H;ʸH;I�H;.�H;*�H;��H;��H;~�H;�H;~�H;��H;��H;)�H;/�H;I�H;ǸH;b�H;�rH;-�G;LwF;�C;��;;�,;�;�: 17� ��%����(;�ע�/#�%<Q�'ڟ�����k/��.}�9o�������f'��"Y�����������¿      ?^������m���[o���@�*�&�޾����<ce�2����ڽ����g@������R���O*�@G������F^9L��:$;�d.;�<;̐C;@�F;��G;�yH;ϥH;A�H;W�H;��H;��H;�H;%�H;��H;K�H;��H;%�H;	�H;��H;��H;V�H;@�H;̥H;�yH;��G;@�F;ʐC;�<;�d.;$;N��:�F^9���@G���O*��R������g@�������ڽ2��<ce�����&�޾*���@�[o�m�������      1����������[o��!J�M�#��\��XD������|PH�����b��!C��� +���ټ)����俐�欷�<�:K��:h�;�Y1;>;�0D;��F;H;y�H;�H;5�H;��H;��H;<�H;��H;��H;��H;��H;��H;��H;��H;;�H;��H;��H;1�H;�H;y�H;�H;��F;�0D;>;�Y1;h�;M��:8�:䬷�⿐���(����ټ� +�!C���b�����|PH�����XD���\��M�#��!J�[o��������      [o�bXi��"Y���@�M�#��
��о�A���i���(����xr���_��5��ɺ�o�`��<��R�d� �\��X:�P�:a;�4;ԧ?;��D;�8G;�0H;͋H;��H;��H;:�H;��H;��H;.�H;��H;A�H;��H;A�H;��H;.�H;��H;��H;:�H;��H;��H;͋H;�0H;�8G;��D;ҧ?;�4;a;�P�:�X:��\�Q�d��<��o�`��ɺ��5��_�xr�������(��i��A���о�
�M�#���@��"Y�bXi�      ��7�ѕ3��f'�*��\���о�����.}��-=�}
���Ľ]��-:�����������7�GĻ��$�8N��%��:�{;�D&;+,8;4JA;,�E;��G;�LH;�H;��H;\�H;�H;;�H;��H;��H;S�H;��H;K�H;��H;S�H;��H;��H;<�H;�H;[�H;��H;�H;�LH;��G;)�E;1JA;*,8;�D&;�{;��:8N����$�GĻ��7���������-:�]����Ľ}
��-=��.}������о�\��*��f'�ѕ3�      ���
�����&�޾XD���A���.}�+�D�jt���ڽ�!��\����]�ļ�
v�:�������Iɺ�S�9#��:8(;�-;��;;��B;�IF;��G;DfH;ϝH;$�H;W�H;��H;��H;��H;��H;��H;#�H;��H;%�H;��H;��H;��H;��H;��H;W�H;!�H;ϝH;CfH;��G;�IF;��B;��;;�-;8(;!��:�S�9�Iɺ����:���
v�]�ļ���\��!����ڽjt�+�D��.}��A��XD��&�޾�����
�      �iþXD��9o�����������i��-=�jt����R��kys�| +����y񗼒(;�#�ѻ�s@�t�!��4j:Q�:
�;�D3;k�>;;FD;��F;�	H;e|H;ťH;��H;a�H;'�H;)�H;��H;P�H;f�H;��H;�H;��H;g�H;P�H;��H;*�H;(�H;`�H;��H;ťH;b|H;�	H;��F;8FD;j�>;�D3;�;Q�:�4j:h�!��s@�"�ѻ�(;�y����| +�kys��R����jt��-=��i���������9o��XD��      �(��Gl���.}�<ce�}PH���(�}
���ڽ�R���{�E�6�� �-p��]�`�ʨ��,��IҺN^9ׇ�:�;�~(;[�8;JA;,|E;FjG;�=H;q�H;�H;X�H;��H;\�H;��H;��H;�H;��H;&�H;��H;&�H;��H;�H;��H;��H;]�H;��H;U�H;�H;q�H;�=H;DjG;+|E;JA;Y�8;�~(;�;ׇ�:0N^9
IҺ�,��ʨ�]�`�-p��� �E�6��{��R����ڽ}
���(�}PH�<ce��.}�Hl��      �-=�D�9��k/�2��������Ľ�!��kys�E�6�'#��ɺ��vz����7^��R�$��}�r:J��:�;�Y1;*I=;_xC;SwF;V�G;8fH;v�H;��H;��H;��H;��H;�H;�H;��H;��H;��H;��H;��H;��H;��H;�H;�H;��H;��H;��H;��H;t�H;9fH;S�G;OwF;\xC;)I=;�Y1;�;J��:��r:�}�Q�$�8^������vz��ɺ�&#�E�6�kys��!����Ľ����2���k/�D�9�      �` ��.�������ڽ�b��xr��]��\�| +�� ��ɺ�@��O*�<ͻ�5R��ƅ�X�:i��:��;�); u8;��@;�*E;�8G;x$H;|�H;r�H;)�H;]�H;��H;��H;��H;4�H;��H;&�H;�H;W�H;�H;'�H;��H;4�H;��H;��H;��H;\�H;)�H;p�H;|�H;w$H;�8G;�*E;��@; u8;�);��;o��:P�:�ƅ��5R�<ͻ�O*�@��ɺ�� �| +�\�]��xr���b����ڽ��.��      A���R��'ڟ�����"C���_�-:�������-p���vz��O*��4ֻ�k����� �09��:(1;{� ;�D3;q�=;ؐC;lF;��G;�\H;ЗH;��H;7�H;v�H;��H;��H;�H;1�H;A�H;��H;��H;��H;��H;��H;A�H;1�H;�H;��H;��H;u�H;7�H;}�H;ӗH;�\H;��G;lF;ؐC;q�=;�D3;{� ;,1;~�:0�09�����k��4ֻ�O*��vz�-p����輦��-:��_�"C������'ڟ��R��      �_�"\�$<Q�g@�� +��5�����]�ļy�]�`����<ͻ�k��Hɺ j6��:$Q�:L�;e.;}�:;M�A;\|E;�NG;x'H;8�H;�H;��H;��H;c�H;��H;��H;j�H;/�H;��H;F�H;��H;6�H;��H;F�H;��H;/�H;m�H;��H;��H;a�H;��H;��H;�H;7�H;w'H;�NG;\|E;M�A;}�:;e.;N�; Q�:�: g6��Hɺ�k�<ͻ���]�`�y�]�ļ�����5�� +�g@�$<Q�#\�      2]� �/#�������ټ�ɺ������
v��(;�ʨ�8^���5R����� k6���:)��: �;J�*;,8;�!@;��D;��F;.�G;fH;��H;ǰH;ٿH;��H;�H;��H;Z�H;��H;�H;��H;��H;`�H;��H;`�H;��H;��H;�H;��H;[�H;��H;�H;��H;ٿH;ɰH;��H;	fH;*�G;��F;��D;�!@;,8;L�*; �;%��:��: m6������5R�8^��ʨ��(;��
v������ɺ���ټ����/#� �      /p��dx��ע��R��)��q�`���7�:��"�ѻ�,��R�$��ƅ� �09y�:/��:�;�~(;�Z6;��>;��C;%IF;�G;"EH;��H;�H;�H;J�H;d�H;N�H;2�H;�H;��H;��H;I�H;$�H;��H;��H;��H;$�H;I�H;��H;��H;�H;2�H;J�H;d�H;H�H;�H;�H;~�H;EH;�G;"IF;��C;��>;�Z6;�~(;�;+��:}�:��09�ƅ�S�$��,��"�ѻ:����7�o�`�)���R��ע�ex��      ��I�,�E��(;��O*����<��GĻ�����s@�
IҺ�}�L�:z�:Q�:"�;�~(;8�5;�>;gC;k�E;�cG;s$H;2|H;s�H;X�H;��H;��H;v�H;�H;Z�H;��H;��H;��H;��H;{�H;�H;,�H;�H;{�H;��H;��H;��H;��H;X�H;�H;v�H;��H;��H;X�H;n�H;,|H;s$H;�cG;m�E;gC;�>;6�5;�~(; �;Q�:x�:L�:�}�
IҺ�s@�����GĻ�<�����O*��(;�/�E�      N�ѻ�ͻ$���@G��濐�`�d���$��Iɺl�!�N^9��r:g��:(1;I�;K�*;�Z6;�>;d�B;��E;9G;�	H;8nH;R�H;��H;�H;��H;��H;�H;��H;:�H;��H;��H;9�H;5�H;��H;>�H;`�H;>�H;��H;6�H;8�H;��H;��H;:�H;��H;�H;��H;��H;�H;~�H;O�H;9nH;�	H;9G;��E;f�B;�>;�Z6;J�*;I�;(1;e��:��r:�M^9h�!��Iɺ��$�\�d�⿐�@G��$����ͻ      h�)�
�$�������𬷺��\�N���S�9�4j:Ӈ�:F��:��;z� ;e.;	,8;��>;gC;��E;�)G;��G;JdH;��H;ҫH;��H;��H;r�H;�H;�H;��H;��H;��H;��H;��H;��H;:�H;n�H;��H;n�H;:�H;��H;��H;��H;��H;��H;��H;�H;�H;u�H;��H;��H;ΫH;��H;HdH;��G;�)G;��E;dC;��>;	,8;e.;x� ;��;J��:͇�:�4j:�S�9N����\�䬷������
�$�      0�R�0�� ,7��F^90�:��X:��:��:
Q�:�;�;�);�D3;v�:;�!@;��C;g�E;9G;��G;�`H;��H;Q�H;X�H;��H;|�H;q�H;��H;��H;��H;�H;��H;F�H;%�H;��H;j�H;��H;��H;��H;j�H;��H;$�H;G�H;��H;�H;��H;��H;��H;r�H;|�H;��H;V�H;R�H;��H;�`H;��G;9G;g�E;��C;�!@;v�:;�D3;�);�;
�;
Q�:��:��:�X:\�:�F^9 -7����      ��:��:�:8��:9��:�P�:�{;5(;�;�~(;�Y1;u8;p�=;K�A;��D;IF;�cG;�	H;HdH;��H;��H;�H;n�H;2�H;	�H;|�H;��H;��H;c�H;!�H;��H;��H;��H;#�H;��H;��H;��H;��H;��H;#�H;��H;��H;��H;�H;a�H;��H;��H;|�H;	�H;-�H;m�H;�H;��H;��H;HdH;�	H;�cG;IF;��D;L�A;p�=;u8;�Y1;�~(;
�;7(;�{;�P�:=��:>��:�:퍨:      S�
;v�;�;;h�;a;�D&;�-;�D3;\�8;-I=;��@;ؐC;\|E;��F;�G;q$H;6nH;��H;R�H;�H;��H;w�H;\�H;��H;��H;!�H;��H;��H;E�H;^�H;2�H;��H;\�H;��H;��H;��H;��H;��H;\�H;��H;2�H;^�H;B�H;��H;��H; �H;��H;��H;X�H;t�H;��H;�H;U�H;��H;8nH;p$H;�G;��F;[|E;ؐC;��@;+I=;[�8;�D3;�-;�D&;a;~�;; �;r�;      �*;��*;�,;�d.;�Y1;�4;,,8;��;;m�>;JA;]xC;�*E;lF;�NG;-�G;EH;/|H;P�H;ϫH;W�H;m�H;x�H;��H;7�H;6�H;��H;J�H;(�H;��H;�H;��H;��H;"�H;v�H;��H;��H;��H;��H;��H;v�H;�H;��H;��H;�H;��H;(�H;H�H;��H;7�H;5�H;��H;x�H;j�H;Z�H;ϫH;R�H;,|H;EH;-�G;�NG;lF;�*E;_xC;JA;m�>;��;;,,8;�4;�Y1;�d.;�,;��*;      >�:;Q�:;��;;�<;">;ӧ?;=JA;��B;<FD;.|E;SwF;�8G;��G;x'H;fH;~�H;q�H;��H;��H;��H;-�H;Z�H;6�H;!�H;W�H;��H;��H;r�H;��H;��H;U�H;��H;Y�H;��H;��H;��H;��H;��H;��H;��H;V�H;��H;U�H;��H;��H;r�H;��H;��H;X�H;�H;5�H;Z�H;*�H;��H;��H;��H;p�H;}�H;	fH;x'H;��G;�8G;RwF;,|E;<FD;��B;;JA;ԧ?;*>;�<;��;;B�:;      �B;*�B;�C;АC;�0D;��D;,�E;�IF;��F;DjG;V�G;{$H;�\H;;�H;��H;�H;^�H;�H;��H;��H;�H;��H;<�H;^�H;��H;��H;9�H;��H;h�H;5�H;��H;�H;m�H;��H;��H;��H;��H;��H;��H;��H;j�H;�H;��H;3�H;e�H;��H;7�H;��H;��H;[�H;:�H;��H;�H;��H;��H;�H;Z�H;�H;��H;9�H;�\H;{$H;V�G;DjG;��F;�IF;,�E;��D;�0D;АC;�C;*�B;      WIF;:UF;AwF;>�F;��F;�8G;��G;��G;�	H;�=H;8fH;~�H;ЗH;�H;İH;�H;��H;��H;p�H;q�H;y�H;��H;��H;��H;��H;6�H;e�H;I�H;��H;��H;�H;]�H;r�H;��H;��H;��H;��H;��H;��H;��H;o�H;^�H;�H;��H;��H;I�H;d�H;7�H;��H;��H;��H;��H;u�H;o�H;p�H;��H;��H;�H;İH;�H;ЗH;~�H;9fH;�=H;�	H;��G;��G;�8G;��F;@�F;AwF;/UF;      G�G;��G;.�G;��G;�H;�0H;�LH;GfH;i|H;r�H;z�H;w�H;��H;��H;ٿH;J�H;��H;��H;�H;��H;��H;!�H;I�H;��H;3�H;h�H;;�H;��H;��H;��H;�H;k�H;��H;��H;��H;��H;��H;��H;��H;��H;��H;k�H;�H;��H;��H;��H;9�H;g�H;9�H;��H;H�H;!�H;��H;��H;�H;��H;��H;J�H;ٿH;��H;��H;w�H;z�H;r�H;j|H;GfH;�LH;�0H;�H;��G;-�G;��G;      �lH;bnH;�rH;�yH;}�H;ҋH;�H;ٝH;˥H;�H;��H;0�H;;�H;��H;��H;e�H;u�H;�H;�H;��H;��H;��H;(�H;u�H;z�H;J�H;��H;r�H;��H;(�H;G�H;u�H;��H;��H;��H;��H;��H;��H;��H;��H;��H;t�H;E�H;%�H;��H;r�H;��H;J�H;|�H;t�H;(�H;��H;��H;��H;�H;�H;t�H;d�H;��H;��H;8�H;2�H;��H;�H;̥H;۝H;�H;ҋH;��H;�yH;�rH;onH;      Q�H;ܡH;c�H;ӥH;�H;��H;��H;(�H;��H;[�H;��H;d�H;y�H;d�H;�H;O�H;�H;��H;��H;��H;b�H;��H;��H;��H;a�H;��H;��H;��H;	�H;L�H;j�H;��H;��H;��H;��H;��H;��H;��H;��H;��H;��H;��H;h�H;L�H;	�H;��H;��H;��H;c�H;��H;��H;��H;_�H;��H;��H;��H;�H;N�H;�H;c�H;y�H;c�H;��H;[�H;��H;*�H;��H;��H;�H;ԥH;c�H;ѡH;      ��H;�H;ԸH;C�H;C�H;��H;c�H;^�H;k�H;��H;��H;��H;��H;��H; �H;6�H;\�H;9�H;��H;�H;"�H;B�H;�H;��H;,�H;��H;��H;(�H;K�H;`�H;�H;}�H;��H;��H;��H;��H;��H;��H;��H;��H;��H;�H;�H;^�H;I�H;(�H;��H;��H;.�H;��H;�H;B�H;"�H;�H;��H;:�H;[�H;4�H;��H;��H;��H;��H;��H;��H;m�H;`�H;b�H;��H;C�H;D�H;иH;�H;      z�H;��H;V�H;b�H;��H;:�H;�H;�H;1�H;c�H;��H;��H;��H;��H;_�H;�H;��H;��H;��H;��H;��H;^�H;��H;Y�H;��H;�H;�H;H�H;g�H;��H;��H;��H;{�H;}�H;��H;��H;k�H;��H;��H;}�H;x�H;��H;��H;��H;h�H;H�H;�H;�H;��H;Y�H;��H;^�H;��H;��H;��H;��H;��H;�H;^�H;��H;��H;��H;��H;e�H;1�H;
�H;�H;:�H;��H;b�H;U�H;��H;      ��H;��H;6�H;��H;��H;��H;?�H;��H;.�H;��H;�H;��H;�H;r�H;��H;��H;��H;��H;��H;P�H;��H;7�H;��H;��H;�H;^�H;h�H;v�H;��H;�H;��H;��H;{�H;u�H;��H;m�H;c�H;k�H;��H;u�H;v�H;��H;��H;��H;��H;v�H;j�H;]�H;�H;��H;��H;7�H;��H;P�H;��H;��H;��H;��H;��H;r�H;�H;��H;�H;��H;1�H;��H;@�H;��H;��H;��H;6�H;��H;      ��H;��H;4�H;��H;I�H;��H;��H;��H;��H;��H;�H;A�H;6�H;6�H;	�H;��H;��H;8�H;��H;,�H;��H;��H;!�H;^�H;g�H;r�H;��H;��H;��H;��H;|�H;|�H;�H;}�H;\�H;Z�H;��H;Z�H;\�H;}�H;{�H;}�H;|�H;��H;��H;��H;��H;q�H;h�H;^�H;�H;��H;��H;.�H;��H;9�H;��H;��H;�H;6�H;5�H;?�H;�H;��H;��H;��H;��H;��H;B�H;��H;4�H;��H;      ��H;��H;��H;�H;��H;)�H;��H;��H;V�H;�H;��H;��H;E�H;�H;��H;S�H;��H;7�H;��H;��H;*�H;]�H;v�H;��H;��H;��H;��H;��H;��H;��H;{�H;u�H;x�H;g�H;V�H;]�H;a�H;]�H;V�H;g�H;v�H;x�H;{�H;��H;��H;��H;��H;��H;��H;��H;x�H;]�H;)�H;��H;��H;9�H;��H;S�H;��H;�H;E�H;��H;��H;�H;W�H;��H;��H;.�H;��H;�H;��H;��H;      ��H;��H;��H;0�H;��H;��H;\�H;��H;p�H;��H;��H;5�H;��H;N�H;��H;.�H;��H;��H;=�H;o�H;��H;��H;��H;��H;��H;��H;��H;��H;��H;��H;��H;��H;Z�H;W�H;a�H;W�H;:�H;W�H;a�H;W�H;W�H;��H;��H;��H;��H;��H;��H;��H;��H;��H;��H;��H;��H;o�H;=�H;��H;��H;.�H;��H;M�H;��H;5�H;��H;��H;q�H;��H;\�H;��H;��H;.�H;��H;��H;      6�H;\�H;��H;��H;��H;=�H;��H;0�H;��H;'�H;��H;&�H;��H;��H;f�H;��H;�H;;�H;t�H;��H;��H;��H;��H;��H;��H;��H;��H;��H;��H;��H;��H;o�H;Z�H;a�H;W�H;S�H;D�H;S�H;W�H;^�H;Y�H;r�H;��H;��H;��H;��H;��H;��H;��H;��H;��H;��H;��H;��H;t�H;=�H;�H;��H;f�H;��H;��H;&�H;��H;*�H;��H;/�H;��H;A�H;��H;��H;��H;U�H;      ��H;�H;�H;N�H;��H;��H;P�H;��H;"�H;��H;��H;b�H;��H;@�H;��H;��H;3�H;]�H;��H;��H;��H;��H;��H;�H;��H;��H;��H;��H;��H;��H;n�H;h�H;��H;d�H;:�H;D�H;>�H;D�H;:�H;d�H;��H;j�H;n�H;��H;��H;��H;��H;��H;��H;�H;��H;��H;��H;��H;��H;^�H;2�H;��H;��H;@�H;��H;b�H;��H;��H;#�H;��H;P�H;��H;��H;N�H;�H;��H;      6�H;\�H;��H;��H;��H;=�H;��H;0�H;��H;'�H;��H;&�H;��H;��H;f�H;��H;�H;;�H;t�H;��H;��H;��H;��H;��H;��H;��H;��H;��H;��H;��H;��H;o�H;Z�H;a�H;W�H;S�H;D�H;S�H;W�H;^�H;Y�H;r�H;��H;��H;��H;��H;��H;��H;��H;��H;��H;��H;��H;��H;t�H;=�H;�H;��H;f�H;��H;��H;&�H;��H;)�H;��H;/�H;��H;A�H;��H;��H;��H;T�H;      ��H;��H;��H;0�H;��H;��H;\�H;��H;p�H;��H;��H;5�H;��H;N�H;��H;.�H;��H;��H;=�H;q�H;��H;��H;��H;��H;��H;��H;��H;��H;��H;��H;��H;��H;Z�H;W�H;a�H;W�H;:�H;W�H;a�H;W�H;W�H;��H;��H;��H;��H;��H;��H;��H;��H;��H;��H;��H;��H;o�H;=�H;��H;��H;.�H;��H;N�H;��H;5�H;��H;��H;p�H;��H;\�H;��H;��H;.�H;��H;��H;      ��H;��H;��H;�H;��H;)�H;��H;��H;V�H;�H;��H;��H;E�H;�H;��H;S�H;��H;7�H;��H;��H;-�H;]�H;v�H;��H;��H;��H;��H;��H;��H;��H;{�H;u�H;x�H;g�H;V�H;]�H;a�H;]�H;V�H;g�H;v�H;x�H;{�H;��H;��H;��H;��H;��H;��H;��H;x�H;]�H;)�H;��H;��H;9�H;��H;S�H;��H;�H;E�H;��H;��H;�H;W�H;��H;��H;.�H;��H;�H;��H;��H;      ��H;��H;5�H;��H;G�H;��H;��H;��H;��H;��H;�H;?�H;5�H;6�H;�H;��H;��H;8�H;��H;,�H;��H;��H;!�H;^�H;h�H;r�H;��H;��H;��H;��H;|�H;|�H;}�H;|�H;\�H;Z�H;��H;Z�H;\�H;|�H;{�H;�H;|�H;��H;��H;��H;��H;q�H;g�H;]�H;�H;��H;��H;,�H;��H;8�H;��H;��H;	�H;6�H;5�H;?�H;�H;��H;��H;��H;��H;��H;@�H;��H;3�H;��H;      ��H;��H;9�H;��H;��H;��H;B�H;��H;.�H;��H;�H;��H;�H;r�H;��H;��H;��H;��H;��H;Q�H;��H;7�H;��H;��H;�H;^�H;j�H;v�H;��H;�H;��H;��H;y�H;u�H;��H;k�H;c�H;k�H;��H;u�H;v�H;��H;��H;��H;��H;v�H;j�H;]�H;�H;��H;��H;7�H;��H;P�H;��H;��H;��H;��H;��H;r�H;�H;��H;�H;��H;0�H;��H;@�H;��H;��H;��H;8�H;��H;      z�H;��H;V�H;b�H;��H;9�H;�H;
�H;1�H;d�H;��H;��H;��H;��H;^�H;�H;��H;��H;��H;��H;��H;^�H;��H;[�H;��H;�H;�H;H�H;h�H;��H;��H;��H;y�H;}�H;��H;��H;k�H;��H;��H;}�H;x�H;��H;��H;��H;h�H;H�H;�H;�H;��H;X�H;��H;^�H;��H;��H;��H;��H;��H;�H;_�H;��H;��H;��H;��H;d�H;1�H;
�H;�H;;�H;��H;b�H;V�H;��H;      ��H;�H;ѸH;D�H;A�H;��H;c�H;^�H;m�H;��H;��H;��H;��H;��H;��H;4�H;\�H;7�H;��H;�H;&�H;B�H;�H;��H;.�H;��H;��H;(�H;K�H;`�H;�H;}�H;��H;��H;��H;��H;��H;��H;��H;��H;��H;�H;�H;^�H;K�H;(�H;��H;��H;,�H;��H;�H;B�H;!�H;�H;��H;9�H;[�H;7�H; �H;��H;��H;��H;��H;��H;n�H;`�H;e�H;��H;A�H;C�H;ԸH;�H;      I�H;ءH;i�H;ҥH;�H;��H;��H;+�H;��H;[�H;��H;d�H;y�H;c�H;�H;N�H;�H;��H;��H;��H;e�H;��H;��H;��H;c�H;��H;��H;��H;	�H;N�H;h�H;��H;��H;��H;��H;��H;��H;��H;��H;��H;��H;��H;j�H;I�H;	�H;��H;��H;��H;a�H;��H;��H;��H;_�H;��H;��H;��H;�H;Q�H;�H;d�H;y�H;d�H;��H;Y�H;��H;*�H;��H;��H;	�H;ϥH;g�H;١H;      �lH;bnH;�rH;�yH;{�H;ҋH;�H;ܝH;˥H;�H;��H;2�H;8�H;��H;��H;d�H;u�H;�H;�H;��H;��H;��H;(�H;u�H;|�H;J�H;��H;r�H;��H;(�H;E�H;t�H;��H;��H;��H;��H;��H;��H;��H;��H;��H;v�H;G�H;%�H;��H;r�H;��H;J�H;z�H;t�H;(�H;��H;��H;��H;�H;�H;t�H;g�H;��H;��H;;�H;2�H;��H;�H;̥H;ٝH;�H;ϋH;��H;�yH;�rH;mnH;      A�G;��G;-�G;��G;�H;�0H;�LH;GfH;i|H;t�H;z�H;w�H;��H;��H;ٿH;K�H;��H;��H;�H;��H;��H;!�H;I�H;��H;9�H;h�H;;�H;��H;��H;��H;�H;k�H;��H;��H;��H;��H;��H;��H;��H;��H;��H;m�H;�H;��H;��H;��H;9�H;h�H;3�H;��H;H�H;!�H;��H;��H;�H;��H;��H;H�H;ٿH;��H;��H;w�H;{�H;t�H;i|H;FfH;�LH;�0H;�H;��G;+�G;��G;      ^IF;3UF;JwF;A�F;��F;�8G;��G;��G;�	H;�=H;8fH;|�H;ЗH;�H;ðH;�H;��H;��H;p�H;o�H;{�H;��H;��H;��H;��H;7�H;e�H;I�H;��H;��H;�H;]�H;q�H;��H;��H;��H;��H;��H;��H;��H;o�H;^�H;�H;��H;��H;I�H;d�H;7�H;��H;��H;��H;��H;u�H;o�H;p�H;��H;��H;�H;İH;�H;ЗH;~�H;8fH;�=H;�	H;��G;��G;�8G;��F;A�F;KwF;*UF;      �B;*�B;�C;АC;�0D;��D;,�E;�IF;��F;EjG;X�G;{$H;�\H;9�H;��H;�H;[�H;�H;��H;��H;�H;��H;:�H;^�H;��H;��H;9�H;��H;i�H;5�H;��H;�H;k�H;��H;��H;��H;��H;��H;��H;��H;k�H;�H;��H;3�H;e�H;��H;7�H;��H;��H;\�H;:�H;��H;�H;��H;��H;�H;Z�H;�H;��H;9�H;�\H;{$H;V�G;BjG;��F;�IF;,�E;��D;�0D;АC;�C;*�B;      A�:;O�:;��;;�<;>;٧?;8JA;��B;>FD;/|E;UwF;�8G;��G;y'H;	fH;}�H;q�H;��H;��H;��H;/�H;Z�H;6�H;!�H;X�H;��H;��H;r�H;��H;��H;U�H;��H;W�H;��H;��H;��H;��H;��H;��H;��H;W�H;��H;U�H;��H;��H;r�H;��H;��H;W�H; �H;5�H;Z�H;*�H;��H;��H;��H;p�H;~�H;fH;y'H;��G;�8G;RwF;.|E;>FD;��B;8JA;٧?;*>;�<;��;;A�:;      �*;��*;�,;�d.;�Y1;	�4;1,8;��;;m�>;JA;_xC;�*E;lF;�NG;-�G;EH;/|H;O�H;ϫH;X�H;p�H;x�H;��H;7�H;7�H;��H;J�H;(�H;��H;�H;��H;��H;"�H;v�H;��H;��H;��H;��H;��H;v�H;�H;��H;��H;�H;��H;(�H;H�H;��H;6�H;5�H;��H;x�H;i�H;X�H;ϫH;P�H;.|H;EH;.�G;�NG;lF;�*E;]xC;JA;m�>;��;;1,8;	�4;�Y1;�d.;�,;��*;      S�
;x�;�;;f�;a;�D&;�-;�D3;[�8;-I=;��@;ؐC;[|E;��F;�G;p$H;6nH;��H;T�H;�H;��H;w�H;\�H;��H;��H;"�H;��H;��H;F�H;^�H;2�H;��H;\�H;��H;��H;��H;��H;��H;\�H;��H;2�H;^�H;A�H;��H;��H; �H;��H;��H;X�H;t�H;��H;�H;T�H;��H;8nH;p$H;�G;��F;\|E;ؐC;��@;+I=;\�8;�D3;�-;�D&;a;z�;; �;p�;      ��:��:�:<��:9��:�P�:�{;9(;	�;�~(;�Y1;u8;p�=;L�A;��D;IF;�cG;�	H;HdH;��H;��H;�H;n�H;2�H;	�H;|�H;��H;��H;c�H;"�H;��H;��H;��H;"�H;��H;��H;��H;��H;��H;#�H;��H;��H;��H;�H;_�H;��H;��H;|�H;	�H;-�H;m�H;�H;~�H;��H;HdH;�	H;�cG;IF;��D;L�A;p�=;u8;�Y1;�~(;
�;8(;�{;�P�:A��:<��:�:퍨:      @�R��� )7��F^9<�:�X:��:��:
Q�:�;�;�);�D3;v�:;�!@;��C;g�E;9G;��G;�`H;��H;R�H;X�H;��H;|�H;r�H;��H;��H;��H;�H;��H;F�H;%�H;��H;j�H;��H;��H;��H;j�H;��H;$�H;G�H;��H;	�H;��H;��H;��H;q�H;|�H;��H;V�H;Q�H;��H;�`H;��G;9G;g�E;��C;�!@;v�:;�D3;�);�;
�;Q�:��:��:�X:L�:�F^9 -7����      h�)�
�$������򬷺��\�N���S�9�4j:͇�:J��:��;x� ;e.;,8;��>;fC;��E;�)G;��G;KdH;��H;ҫH;��H;��H;t�H;�H;�H;��H;��H;��H;��H;��H;��H;:�H;m�H;��H;n�H;:�H;��H;��H;��H;��H;��H;��H;�H;�H;t�H;��H;��H;ΫH;��H;GdH;��G;�)G;��E;fC;��>;,8;e.;z� ;��;F��:Ӈ�:�4j:�S�9N����\�欷�������
�$�      M�ѻ�ͻ$���@G��濐�a�d���$��Iɺl�!��M^9��r:e��:(1;I�;J�*;�Z6;�>;d�B;��E;9G;�	H;9nH;R�H;��H;�H;��H;��H;�H;��H;;�H;��H;��H;9�H;6�H;��H;>�H;`�H;>�H;��H;5�H;8�H;��H;��H;9�H;��H;�H;��H;��H;�H;}�H;O�H;8nH;�	H;9G;��E;d�B;�>;�Z6;K�*;I�;(1;g��:��r:N^9l�!��Iɺ��$�[�d�俐�@G��$����ͻ      ��I�,�E��(;��O*����<��GĻ�����s@�
IҺ�}�L�:x�:Q�: �;�~(;9�5;�>;gC;k�E;�cG;s$H;2|H;s�H;X�H;��H;��H;v�H;�H;Z�H;��H;��H;��H;��H;{�H;�H;,�H;�H;{�H;��H;��H;��H;��H;W�H;�H;v�H;��H;��H;X�H;n�H;,|H;s$H;�cG;m�E;gC;�>;8�5;�~(;"�;Q�:z�:P�:�}�
IҺ�s@�����GĻ�<�����O*��(;�.�E�      /p��dx��ע��R��)��p�`���7�:��"�ѻ�,��S�$��ƅ���09y�:+��:�;�~(;�Z6;��>;��C;%IF;�G;!EH;��H;�H;�H;K�H;d�H;N�H;2�H;�H;��H;��H;I�H;$�H;��H;��H;��H;$�H;I�H;��H;��H;�H;2�H;J�H;d�H;H�H;�H;�H;~�H;EH;�G;"IF;��C;��>;�Z6;�~(;�;/��:}�: �09�ƅ�R�$��,��"�ѻ;����7�p�`�)���R��ע�ex��      2]� �/#�������ټ�ɺ������
v��(;�ʨ�8^���5R����� m6���:%��: �;J�*;,8;�!@;��D;��F;/�G;fH;��H;ǰH;ٿH;��H;�H;��H;[�H;��H;�H;��H;��H;`�H;��H;`�H;��H;��H;�H;��H;Z�H;��H;�H;��H;׿H;ɰH;��H;	fH;(�G;��F;��D;�!@;,8;L�*; �;)��:��: k6������5R�8^��ʨ��(;��
v������ɺ���ټ����/#� �      �_�"\�$<Q�g@�� +��5�����]�ļy�]�`����<ͻ�k��Hɺ h6��:$Q�:M�;e.;z�:;M�A;\|E;�NG;x'H;7�H;�H;��H;��H;c�H;��H;��H;j�H;0�H;��H;F�H;��H;6�H;��H;F�H;��H;.�H;k�H;��H;��H;`�H;��H;��H;�H;8�H;w'H;�NG;\|E;M�A;{�:;e.;N�; Q�:�: j6��Hɺ�k�<ͻ���]�`�x�]�ļ�����5�� +�g@�$<Q�#\�      A���R��'ڟ�����"C���_�-:�������-p���vz��O*��4ֻ�k������09��:*1;{� ;�D3;q�=;ؐC;lF;��G;�\H;їH;��H;7�H;v�H;��H;��H;�H;1�H;A�H;��H;��H;��H;��H;��H;A�H;/�H;�H;��H;��H;t�H;7�H;}�H;ԗH;�\H;��G;lF;ؐC;q�=;�D3;{� ;,1;~�: �09�����k��4ֻ�O*��vz�-p����輦��-:��_�"C������'ڟ��R��      �` ��.�������ڽ�b��xr��]��\�| +�� ��ɺ�@��O*�<ͻ�5R��ƅ�X�:m��:��;�);u8;��@;�*E;�8G;w$H;|�H;r�H;)�H;]�H;��H;��H;��H;5�H;��H;'�H;�H;W�H;�H;&�H;��H;3�H;��H;��H;��H;\�H;)�H;p�H;|�H;x$H;�8G;�*E;��@; u8;�);��;o��:P�:�ƅ��5R�<ͻ�O*�@��ɺ�� �| +�\�]��xr���b��¯ڽ��.��      �-=�D�9��k/�2��������Ľ�!��kys�E�6�&#��ɺ��vz����8^��Q�$��}�r:J��:�;�Y1;)I=;_xC;SwF;S�G;8fH;v�H;��H;��H;��H;��H;�H;�H;��H;��H;��H;��H;��H;��H;��H;�H;�H;��H;��H;��H;��H;t�H;8fH;V�G;QwF;\xC;*I=;�Y1;�;J��:��r:�}�S�$�7^������vz��ɺ�'#�E�6�kys��!����Ľ����2���k/�D�9�      �(��Gl���.}�<ce�}PH���(�}
���ڽ�R���{�E�6�� �-p��]�`�ʨ��,��IҺN^9ׇ�:�;�~(;Y�8;JA;.|E;DjG;�=H;q�H;�H;X�H;��H;]�H;��H;��H;�H;��H;&�H;��H;&�H;��H;�H;��H;��H;\�H;��H;U�H;�H;p�H;�=H;FjG;+|E;JA;[�8;�~(;�;ׇ�:0N^9
IҺ�,��ʨ�]�`�-p��� �E�6��{��R����ڽ}
���(�}PH�<ce��.}�Hl��      �iþXD��9o�����������i��-=�jt����R��kys�| +����y񗼒(;�#�ѻ�s@�l�!��4j:Q�:	�;�D3;k�>;;FD;��F;�	H;e|H;ťH;��H;`�H;(�H;)�H;��H;P�H;g�H;��H;�H;��H;f�H;P�H;��H;)�H;'�H;`�H;��H;ťH;b|H;�	H;��F;9FD;j�>;�D3;�;Q�:�4j:l�!��s@�#�ѻ�(;�y����| +�kys��R����jt��-=��i���������9o��XD��      ���
�����&�޾XD���A���.}�+�D�jt���ڽ�!��\����]�ļ�
v�:�������Iɺ�S�9!��:7(;�-;��;;��B;�IF;��G;DfH;ϝH;$�H;W�H;��H;��H;��H;��H;��H;#�H;��H;%�H;��H;��H;��H;��H;��H;W�H;!�H;ϝH;CfH;��G;�IF;��B;��;;�-;9(;��:�S�9�Iɺ����:���
v�]�ļ���\��!����ڽjt�+�D��.}��A��XD��&�޾�����
�      ��7�ѕ3��f'�*��\���о�����.}��-=�}
���Ľ]��-:�����������7�GĻ��$�8N����:�{;�D&;+,8;6JA;)�E;��G;�LH;�H;��H;\�H;�H;;�H;��H;��H;S�H;��H;K�H;��H;S�H;��H;��H;;�H;�H;[�H;��H;�H;�LH;��G;,�E;3JA;*,8;�D&;�{;��:8N����$�GĻ��7���������-:�]����Ľ}
��-=��.}������о�\��*��f'�ѕ3�      [o�bXi��"Y���@�M�#��
��о�A���i���(����xr���_��5��ɺ�o�`��<��R�d���\��X:�P�:a;�4;ԧ?;��D;�8G;�0H;͋H;��H;��H;:�H;��H;��H;.�H;��H;A�H;��H;C�H;��H;.�H;��H;��H;:�H;��H;��H;͋H;�0H;�8G;��D;ҧ?;�4;a;�P�:�X: �\�Q�d��<��o�`��ɺ��5��_�xr�������(��i��A���о�
�M�#���@��"Y�bXi�      1����������[o��!J�M�#��\��XD������|PH�����b��!C��� +���ټ)����㿐�欷�8�:K��:h�;�Y1;>;�0D;��F;H;y�H;	�H;4�H;��H;��H;<�H;��H;��H;��H;��H;��H;��H;��H;;�H;��H;��H;3�H;�H;y�H;�H;��F;�0D;>;�Y1;h�;M��:8�:欷�㿐���)����ټ� +�!C���b�����|PH�����XD���\��M�#��!J�[o��������      ?^������m���[o���@�*�&�޾����<ce�2����ڽ����g@������R���O*�@G������F^9J��:$;�d.;�<;ʐC;@�F;��G;�yH;ϥH;C�H;V�H;��H;��H;	�H;%�H;��H;K�H;��H;%�H;�H;��H;��H;W�H;@�H;̥H;�yH;��G;@�F;̐C;�<;�d.;$;N��:�F^9���@G���O*��R������g@�������ڽ2��<ce�����&�޾*���@�[o�m�������      �aǿ�¿����������"Y��f'�����9o���.}��k/����'ڟ�%<Q�/#�ע��(;�&��� �� 17��:�;�,;��;;�C;LwF;-�G;�rH;e�H;ʸH;I�H;/�H;*�H;��H;��H;~�H;�H;~�H;��H;��H;)�H;.�H;I�H;ǸH;b�H;�rH;-�G;LwF;�C;��;;�,;�;�: 17� ��%����(;�ע�/#�%<Q�'ڟ�����k/��.}�9o�������f'��"Y�����������¿      5�ֿFpѿ�¿������bXi�ѕ3��
�XD��Gl��D�9��.���R��#\� �dx��.�E��ͻ�$�����:Z�;��*;C�:;!�B;,UF;��G;^nH;ءH;�H;��H;��H;��H;��H;��H;Q�H;��H;Q�H;��H;��H;��H;��H;��H;�H;աH;^nH;��G;-UF;!�B;A�:;��*;Z�;�: ���$��ͻ.�E�ex�� �#\��R���.��D�9�Gl��XD���
�ѕ3�bXi��������¿Fpѿ      ��"$������꿱�ſ�ޞ�(3s��2�A����� j���|HͽǸ����'�C<ͼn�n�\���+Q^�-.����:�W;�S%;qo8;��A;lDF;�H;��H;��H;�H;[�H;O�H;Z�H;��H;�H;��H;?�H;��H;�H;��H;Y�H;Q�H;[�H;�H;��H;��H;�H;lDF;��A;oo8;�S%;�W;���:-.�+Q^�\���n�n�C<ͼ��'�Ǹ��|Hͽ�� j���A����2�(3s��ޞ���ſ������"$�      "$�������忊�����!cm�W�-�����Rh��Yde�#-�ڪɽ�v��)�$���ɼumj�0����X�<��
Ɔ:�x;P�%;?�8;{B;{RF;H;<�H;b�H;�H;~�H;T�H;K�H;��H;��H;��H;:�H;��H;��H;��H;I�H;T�H;~�H;�H;_�H;<�H;H;zRF;{B;<�8;V�%;�x;
Ɔ:D���X�/���vmj���ɼ)�$��v��ڪɽ#-�Yde�Rh������W�-�!cm��������忞����      ��������� �ԿNw�����<�\�"����m��\0X�����;����w����������]��黲F�(��ʒ:
�;I�';̏9;/pB;�zF;�!H;��H;E�H;-�H;��H;Y�H;O�H;��H;��H;��H;&�H;��H;��H;��H;N�H;Y�H;��H;*�H;B�H;��H;�!H;�zF;/pB;ɏ9;K�';
�;ʒ:0�깲F��黩�]����������w��;�����\0X�m�����"�<�\����Nw�� �Կ��𿞏�      ����� �Կp���ޞ�bF�j�C�.E�%�;�I���D��� "��i�c�}��֯���J��ѻ��)��|K�B��:)�
;�M*;��:;�C;�F;�8H;c�H;��H;��H;��H;R�H;O�H;��H;��H;��H;�H;��H;��H;��H;N�H;R�H;��H;��H;��H;d�H;�8H;�F;�C;~�:; N*;+�
;F��:�|K���)��ѻ��J��֯�}�i�c� "�����D��I��%�;.E�j�C�bF��ޞ�p�� �Կ��      ��ſ���Nw���ޞ�����A�W�7�%�����jɰ��|x�h{+�Ա����J��  �Ͷ��V�1� ���+��#
9�:��;�-;��<;��C;�G;�TH;Y�H;
�H;��H;��H;i�H;G�H;��H;��H;��H;�H;��H;��H;��H;E�H;j�H;��H;��H;	�H;Y�H;�TH;�G;��C;��<;"�-;��; �:�#
9 +����V�1�Ͷ���  ��J���Ա�h{+��|x�jɰ�����7�%�A�W������ޞ�Nw�����      �ޞ�������bF�A�W�Y�-����BKɾ�G����O����ƽɸ��Є-���ۼㄼ/4�ǐ��ζ��]:%��:�;��1;d>;{�D;�\G;QsH;��H;x�H;q�H;4�H;��H;=�H;�H;��H;��H;��H;��H;��H;��H;=�H;��H;4�H;n�H;t�H;��H;OsH;�\G;z�D;�c>;��1;�;'��:�]:�ζ�ǐ�04�ㄼ��ۼЄ-�ɸ��ƽ�����O��G��BKɾ���Y�-�A�W�bF�������      (3s�!cm�<�\�j�C�7�%�����TҾl�� j��C(����`P����[�}������Y�.��MX���<���k:m��:� ;�5;SR@;quE;�G;?�H;T�H;��H;�H;W�H;�H;9�H;x�H;��H;k�H;��H;k�H;��H;x�H;9�H;��H;W�H;�H;��H;U�H;>�H;�G;nuE;OR@;�5;� ;o��:��k:��<�JX�.����Y����}���[�`P����콭C(� j�l���TҾ���7�%�j�C�<�\�!cm�      �2�W�-�"�.E�����BKɾl����s�;�5���x㻽�v��
z0��;��+���*����6��9S��M�:m�	;��(;)�9;�/B;�DF;_H;ޫH;��H;��H;��H;��H;��H;#�H;G�H;U�H;P�H;o�H;P�H;U�H;G�H;#�H;��H;��H;��H;��H;��H;ܫH;_H;�DF;�/B;)�9;��(;n�	;�M�:�9S�6�����*��+���;�
z0��v��x㻽��;�5���s�l��BKɾ����.E�"�W�-�      A����������%�;jɰ��G�� j�;�5��	�Ҫɽ[����J�t���沼��]�����	x�	���n:��:�v;��/;�-=;��C;R�F;*IH;��H;1�H;��H;0�H;��H;��H;��H;�H;"�H;)�H;:�H;)�H;"�H;�H;��H;��H;��H;.�H;��H;1�H;��H;,IH;O�F;��C;�-=;��/;�v;��:�n:	���	x������]��沼t���J�[���Ҫɽ�	�;�5� j��G��jɰ�%�;��徹���      ��Rh��m���I���|x���O��C(���Ҫɽ����TDX�I��'<ͼㄼ�X!��s���W��sK�d��:�y;"�#;I6;CR@;�PE;��G;��H;��H;>�H;��H;��H;��H;��H;��H;��H;��H;��H;��H;��H;��H;��H;��H;��H;��H;��H;��H;>�H;��H;��H;��G;�PE;AR@;I6;"�#;�y;d��:�sK��W��s���X!�ㄼ'<ͼI��TDX�����Ҫɽ���C(���O��|x��I��m��Sh��       j�Yde�\0X��D�h{+�������x㻽[���TDX������ۼ˾����;�<>ۻX���y�d?":���:��;�-;��;;�B;�zF;�H;��H;��H;2�H;��H;�H;��H;��H;��H;��H;��H;��H;��H;��H;��H;��H;��H;��H;��H;�H;��H;2�H;��H;��H;�H;�zF;�B;��;;�-;��;���:t?":��y�X�<>ۻ��;�˾����ۼ���TDX�[���x㻽��콄��h{+��D�\0X�Yde�      ��#-������Ա�ƽ`P���v���J�I����ۼ��`�J�����z+��PrѺ�*
9N�: �;� $;�5;�?;��D;o\G;fH; �H;��H;��H;��H;/�H;�H;i�H;��H;r�H;j�H;x�H;Q�H;z�H;m�H;t�H;��H;k�H;�H;/�H;��H;��H;��H;�H;fH;n\G;��D;�?;�5;� $; �;N�:p*
9NrѺz+������`�J�����ۼI���J��v��`P��ƽԱ轅����$-�      }Hͽڪɽ�;�� "����ɸ����[�z0�t��'<ͼʾ��`�J�����j��]*���:��:wb�:d�;��/;�L<;C;<mF;��G;�H;�H; �H;!�H;W�H;h�H;�H;=�H;H�H;5�H;/�H;�H;�H;�H;.�H;5�H;H�H;=�H;�H;h�H;V�H;!�H;�H;�H;�H;��G;8mF;C;�L<;��/;d�;}b�:8��:��_*��j�����`�J�ʾ��(<ͼt��z0���[�ɸ���� "���;��ڪɽ      Ǹ���v����w�i�c��J�Є-�}��;缆沼ㄼ��;������j���5�p�김?Q:���:ti;�M*;��8;��@;�PE;�uG;OiH;��H;��H;&�H;7�H;��H;��H;��H;�H;��H;��H;��H;��H;��H;��H;��H;��H;��H;�H;��H;��H;��H;7�H;%�H;��H;��H;LiH;�uG;�PE;��@;��8;�M*;wi;���:x?Q:p�깋5��j��������;�ㄼ�沼�;�}�τ-��J�i�c���w��v��      ��'�)�$����}��  ���ۼ����+����]��X!�=>ۻ|+��b*����L�>:��:%�;E�%;��5;��>;�(D;"�F;�!H;G�H;g�H;�H;��H;��H;�H;��H;��H;��H;��H;��H;��H;h�H;��H;i�H;��H;��H;��H;��H;��H;��H; �H;��H;��H;�H;g�H;C�H;�!H;"�F;�(D;��>;��5;I�%;#�;��:L�>:���b*�|+��<>ۻ�X!���]��+�������ۼ�  �}����)�$�      B<ͼ��ɼ�����֯�Ͷ��ㄼ��Y��*�����s��X�TrѺ��t?Q:��:��
;a�#;u�3;�c=;$C;8DF;�G;'�H;��H;'�H;O�H;�H;p�H;=�H;�H;��H;}�H;S�H;l�H;&�H;�H;#�H;�H;&�H;j�H;P�H;~�H;��H;�H;9�H;p�H;�H;Q�H;%�H;��H;#�H;�G;6DF;$C;�c=;w�3;`�#;��
;��:x?Q:��TrѺX��s������*���Y�ㄼͶ���֯�������ɼ      n�n�smj���]���J�V�1�/4�*������	x��W���y�p*
92��:���:%�;]�#;j�2;�<;pB;=�E;ōG;�eH;�H;K�H;��H;�H;��H;��H;W�H;e�H;T�H;+�H;�H;��H;��H;��H;��H;��H;��H;��H;�H;+�H;T�H;c�H;T�H;��H;��H;�H;��H;I�H;�H;�eH;čG;>�E;�pB;�<;h�2;[�#;$�;���:0��:P*
9��y��W��	x����+��.4�V�1���J���]�vmj�      `���0������ѻ!���ǐ�NX�6�	���sK�p?":N�:sb�:qi;H�%;q�3;�<;W0B;��E;�\G;�HH;]�H;��H;v�H;�H;P�H;X�H;��H;4�H;6�H;�H;��H;��H;|�H;o�H;n�H;L�H;n�H;o�H;}�H;��H;��H;�H;5�H;1�H;��H;W�H;S�H;�H;s�H;��H;]�H;�HH;�\G;��E;Z0B;�<;q�3;F�%;ri;ub�:N�:l?": tK�	��6�NX�ǐ�����ѻ��4���      &Q^��X��F���)�+��ζ���<� ;S��n:^��:���: �;b�;�M*;��5;�c=;pB;��E;�JG;k8H;��H;��H;,�H;F�H;��H;��H;��H;�H;�H;��H;��H;��H;u�H; �H;�H;�H;��H;�H;�H; �H;r�H;��H;��H;��H;�H;�H;��H;��H;��H;B�H;'�H;��H;��H;l8H;�JG;��E;|pB;�c=;��5;�M*;`�;��;���:\��:�n:�:S���<��ζ�+���)��F��X�      -.����깐|K��#
9�]:��k:�M�:��:�y;��;� $;��/;��8;��>;$C;;�E;�\G;h8H;ݥH; �H;;�H;��H;R�H;��H;p�H;��H;��H;��H;��H;[�H;1�H;�H;��H;��H;��H;��H;��H;��H;��H; �H;3�H;[�H;��H;��H;��H;��H;r�H;��H;N�H;��H;;�H;�H;ޥH;h8H;�\G;9�E;$C;��>;��8;��/;� $;��;�y;��:�M�:��k:�]: $
9�|K��� ��      ���:(Ɔ:ʒ:2��:
�:/��:m��:i�	;�v;#�#;�-;�5;�L<;��@;�(D;6DF;ōG;�HH;��H;�H;��H;h�H;��H;|�H;?�H;��H;��H;��H;��H;B�H;&�H;��H;��H;��H;R�H;B�H;D�H;D�H;R�H;��H;��H;��H;&�H;?�H;}�H;��H;��H;��H;A�H;y�H;��H;h�H;��H; �H;��H;�HH;čG;4DF;�(D;��@;�L<;�5;�-;"�#;�v;i�	;m��:5��:�::��:ʒ:Ɔ:      �W;�x;�;�
;��;�;� ;��(;��/;I6;��;;�?;C;�PE;#�F;�G;�eH;\�H;��H;=�H;g�H;��H;O�H;�H;��H;��H;��H;��H;�H;��H;��H;h�H;@�H;-�H;��H;��H;��H;��H;��H;-�H;;�H;h�H;��H;��H;�H;��H;��H;��H;��H;�H;N�H;��H;e�H;>�H;��H;]�H;�eH;�G;$�F;�PE;C;�?;��;;I6;��/;��(;� ;�;ԅ;!�
;�;�x;      �S%;R�%;G�';�M*;�-;��1;�5;)�9;�-=;CR@;�B;��D;<mF;�uG;�!H;#�H;�H;��H;*�H;��H;��H;P�H;%�H;��H;��H;��H;]�H;�H;��H;��H;I�H;�H;��H;��H;��H;��H;x�H;��H;��H;��H;��H;�H;H�H;��H;��H;�H;Z�H;��H;��H;��H;%�H;R�H;��H;��H;*�H;��H;
�H;#�H;�!H;�uG;;mF;��D;�B;AR@;�-=;)�9;�5;��1;"�-;�M*;G�';E�%;      �o8;K�8;ӏ9;~�:;��<; d>;[R@;�/B;��C;�PE;�zF;s\G;��G;OiH;F�H;��H;M�H;w�H;E�H;O�H;x�H;�H;��H;��H;��H;o�H;�H;��H;��H;9�H;��H;��H;��H;T�H;N�H;C�H;�H;C�H;Q�H;T�H;��H;��H;��H;6�H;��H;��H;�H;p�H;��H;��H;��H;�H;v�H;O�H;C�H;x�H;J�H;��H;F�H;OiH;��G;p\G;�zF;�PE;��C;�/B;YR@;d>;��<;��:;ԏ9;=�8;      ��A;�B;pB;�C;��C;~�D;quE;�DF;Q�F;��G;�H;fH;�H;��H;j�H;(�H;��H;�H;��H;��H;B�H;��H;��H;��H;P�H;��H;��H;��H;0�H;��H;��H;k�H;:�H;�H;��H;��H;��H;��H;��H;�H;7�H;m�H;��H;��H;-�H;��H;��H;��H;Q�H;��H;��H;��H;A�H;��H;��H;�H;��H;'�H;j�H;��H;�H;fH;�H;��G;R�F;�DF;quE;~�D;��C;�C;pB;�B;      vDF;�RF;�zF;�F;�G;�\G;�G;]H;,IH;��H;��H;�H;�H;��H;�H;M�H;�H;P�H;��H;o�H;��H;��H;��H;o�H;��H;��H;��H;)�H;��H;��H;H�H;�H;��H;��H;��H;��H;��H;��H;��H;��H;��H;	�H;G�H;��H;��H;)�H;��H;��H;��H;l�H;��H;��H;��H;p�H;��H;R�H;�H;M�H;�H;��H;�H;�H;��H;��H;*IH;]H;�G;�\G;�G;�F;�zF;|RF;      �H;H;�!H;�8H;�TH;TsH;G�H;ޫH;��H;��H;��H;��H; �H;&�H;��H;�H;��H;V�H;��H;��H;��H;��H;[�H;�H;��H;��H;�H;��H;x�H;G�H;��H;��H;��H;w�H;Z�H;6�H;J�H;6�H;X�H;v�H;��H;��H;��H;F�H;w�H;��H;�H;��H;��H;�H;[�H;��H;��H;��H;��H;W�H;��H;�H;��H;&�H;�H;��H;��H;��H;��H;߫H;F�H;QsH;�TH;�8H;�!H;H;      ��H;A�H;��H;_�H;^�H;��H;Y�H;��H;6�H;D�H;:�H;��H;%�H;=�H;��H;p�H;��H;��H;�H;��H;��H;��H;�H;��H;��H;)�H;��H;��H;7�H;��H;��H;x�H;S�H; �H;�H;�H;�H;�H;�H; �H;P�H;x�H;��H;��H;6�H;��H;��H;)�H;��H;��H;�H;��H;��H;��H;�H;��H;��H;p�H;��H;:�H;!�H;��H;7�H;C�H;7�H;��H;Y�H;��H;i�H;_�H;��H;L�H;      �H;d�H;B�H;��H;
�H;x�H;��H;��H;��H;��H;��H;��H;Z�H;��H;�H;=�H;[�H;2�H;	�H;��H;��H;�H;��H;��H;)�H;��H;u�H;9�H;��H;��H;l�H;4�H;��H;��H;��H;��H;��H;��H;��H;��H;��H;5�H;j�H;��H;��H;9�H;u�H;��H;,�H;��H;��H;�H;��H;��H;	�H;2�H;X�H;=�H;�H;��H;X�H;��H;��H;��H;��H;��H;��H;w�H;�H;��H;B�H;[�H;      �H;�H;5�H;��H;�H;u�H;�H;��H;:�H;��H;�H;=�H;m�H;��H;��H;��H;h�H;4�H;��H;��H;B�H;��H;��H;;�H;��H;��H;C�H;��H;��H;b�H;2�H;��H;��H;��H;��H;��H;v�H;��H;��H;��H;��H;��H;2�H;a�H;��H;��H;C�H;��H;��H;9�H;��H;��H;A�H;��H;��H;4�H;f�H;��H;��H;��H;o�H;=�H;�H;��H;;�H;��H;�H;w�H;	�H;��H;1�H;�H;      ^�H;��H;��H;��H;�H;2�H;a�H;��H;��H;��H;�H;�H;�H;�H;��H;��H;\�H;�H;��H;a�H;,�H;��H;I�H;��H;��H;J�H;��H;��H;i�H;4�H;��H;��H;��H;v�H;T�H;^�H;]�H;^�H;T�H;v�H;��H;��H;��H;2�H;j�H;��H;��H;J�H;��H;��H;G�H;��H;)�H;a�H;��H;�H;Z�H;��H;��H;�H;�H;�H;�H;��H;��H;��H;a�H;4�H;�H;��H;��H;��H;      \�H;d�H;`�H;\�H;p�H;��H;��H;��H;��H;��H;��H;u�H;A�H;�H;��H;��H;5�H;��H;��H;;�H;��H;n�H;�H;��H;j�H;�H;��H;z�H;2�H;��H;��H;��H;w�H;E�H;0�H;-�H;1�H;-�H;0�H;E�H;s�H;��H;��H;��H;4�H;z�H;��H;�H;m�H;��H;�H;n�H;��H;;�H;��H;��H;4�H;��H;��H;�H;@�H;r�H;��H;��H;��H;��H;��H;��H;n�H;[�H;`�H;`�H;      ]�H;\�H;Y�H;\�H;U�H;=�H;;�H;/�H;�H;��H;��H;��H;N�H;��H;��H;X�H;�H;��H;z�H;�H;��H;A�H;��H;��H;3�H;��H;��H;U�H; �H;��H;��H;y�H;3�H;'�H;'�H;�H;��H;�H;'�H;'�H;0�H;z�H;��H;��H;�H;U�H;��H;��H;5�H;��H;��H;A�H;��H;
�H;z�H;��H;�H;Z�H;��H;��H;M�H;��H;��H;��H;�H;/�H;=�H;@�H;N�H;\�H;Y�H;V�H;      ��H;��H;��H;��H;��H;|�H;|�H;R�H;�H; �H;��H;{�H;7�H;��H;��H;t�H;��H;~�H;&�H;��H;��H;0�H;��H;Y�H;	�H;��H;q�H;�H;��H;��H;v�H;E�H;#�H;�H;�H;��H;��H;��H;�H;�H;"�H;I�H;v�H;��H;��H;�H;q�H;��H;�H;X�H;��H;0�H;��H;��H;%�H;��H;��H;v�H;��H;��H;7�H;{�H;��H;�H;!�H;S�H;|�H;��H;��H;��H;��H;��H;      �H;�H;��H;��H;��H;��H;��H;c�H;*�H;��H;��H;{�H;7�H;��H;��H;1�H;��H;o�H;�H;��H;\�H;��H;��H;T�H;��H;��H;X�H;�H;��H;��H;T�H;3�H;&�H;�H;��H;��H;��H;��H;��H;�H;#�H;5�H;T�H;��H;��H;�H;W�H;��H;��H;R�H;��H;��H;V�H;��H;�H;p�H;��H;1�H;��H;��H;7�H;{�H;��H;��H;*�H;a�H;��H;��H;��H;��H;��H;�H;      ��H;��H;��H;��H;��H;��H;u�H;\�H;4�H;��H;��H;��H;$�H;��H;o�H;�H;��H;l�H;�H;��H;L�H;��H;��H;H�H;��H;��H;5�H;�H;��H;��H;`�H;1�H;�H;��H;��H;��H;��H;��H;��H;��H; �H;4�H;`�H;��H;��H;�H;5�H;��H;��H;G�H;��H;��H;K�H;��H;�H;n�H;��H;�H;m�H;��H;$�H;��H;��H;��H;6�H;Z�H;u�H;��H;��H;��H;��H;��H;      ?�H;C�H;8�H;�H;�H;��H;��H;x�H;A�H;��H;��H;\�H;�H;��H;��H;-�H;��H;F�H;��H;��H;G�H;��H;w�H;"�H;��H;��H;G�H;�H;��H;y�H;`�H;7�H;��H;��H;��H;��H;��H;��H;��H;��H;��H;8�H;`�H;z�H;��H;�H;G�H;��H;��H; �H;w�H;��H;E�H;��H;��H;H�H;��H;-�H;��H;��H;�H;\�H;��H;��H;B�H;v�H;��H;��H;�H;�H;7�H;<�H;      ��H;��H;��H;��H;��H;��H;u�H;\�H;4�H;��H;��H;��H;$�H;��H;o�H;�H;��H;l�H;�H;��H;N�H;��H;��H;H�H;��H;��H;6�H;�H;��H;��H;`�H;1�H;�H;��H;��H;��H;��H;��H;��H;��H; �H;4�H;`�H;��H;��H;�H;5�H;��H;��H;F�H;��H;��H;K�H;��H;�H;n�H;��H;�H;o�H;��H;$�H;��H;��H;��H;4�H;Z�H;u�H;��H;��H;��H;��H;��H;      �H;�H;��H;��H;��H;��H;��H;c�H;*�H;��H;��H;{�H;7�H;��H;��H;1�H;��H;o�H;�H;��H;\�H;��H;��H;T�H;��H;��H;X�H;�H;��H;��H;T�H;3�H;&�H;�H;��H;��H;��H;��H;��H;�H;#�H;7�H;T�H;��H;��H;�H;W�H;��H;��H;Q�H;��H;��H;W�H;��H;�H;p�H;��H;1�H;��H;��H;7�H;{�H;��H;��H;*�H;a�H;��H;��H;��H;��H;��H;�H;      ��H;��H;��H;��H;��H;|�H;|�H;R�H;�H;�H;��H;{�H;7�H;��H;��H;v�H;��H;~�H;%�H;��H;��H;0�H;��H;Y�H;�H;��H;q�H;�H;��H;��H;v�H;F�H;#�H;�H;�H;��H;��H;��H;�H;�H;"�H;I�H;v�H;��H;��H;�H;q�H;��H;	�H;X�H;��H;0�H;��H;��H;&�H;��H;��H;t�H;��H;��H;7�H;{�H;��H; �H;!�H;R�H;|�H;��H;��H;��H;��H;��H;      a�H;]�H;Z�H;]�H;R�H;;�H;;�H;-�H;�H;��H;��H;��H;M�H;��H;��H;Z�H;�H;��H;z�H;�H;��H;A�H;��H;��H;5�H;��H;��H;U�H; �H;��H;��H;y�H;1�H;&�H;'�H;�H;��H;�H;'�H;&�H;0�H;|�H;��H;��H;�H;U�H;��H;��H;3�H;��H;��H;A�H;��H;
�H;z�H;��H;�H;X�H;��H;��H;M�H;��H;��H;��H;�H;,�H;:�H;>�H;K�H;\�H;W�H;\�H;      \�H;d�H;c�H;[�H;n�H;��H;��H;��H;��H;��H;��H;t�H;@�H;�H;��H;��H;5�H;��H;��H;<�H;��H;n�H;�H;��H;m�H;	�H;��H;z�H;2�H;��H;��H;��H;v�H;E�H;0�H;-�H;1�H;-�H;0�H;E�H;s�H;��H;��H;��H;4�H;z�H;��H;�H;j�H;��H;�H;n�H;��H;;�H;��H;��H;4�H;��H;��H;�H;A�H;t�H;��H;��H;��H;��H;��H;��H;k�H;Y�H;c�H;b�H;      ^�H;��H;��H;��H;�H;4�H;a�H;��H;��H;��H;�H;�H;�H;�H;��H;��H;Z�H;�H;��H;a�H;-�H;��H;I�H;��H;��H;K�H;��H;��H;i�H;4�H;��H;��H;��H;v�H;T�H;^�H;]�H;^�H;T�H;v�H;��H;��H;��H;2�H;j�H;��H;��H;H�H;��H;��H;G�H;��H;)�H;a�H;��H;�H;[�H;��H;��H;�H;�H;�H;�H;��H;��H;��H;a�H;4�H;�H;��H;��H;��H;      �H;�H;2�H;��H;�H;t�H;�H;��H;;�H;��H;�H;=�H;o�H;��H;��H;��H;h�H;2�H;��H;��H;F�H;��H;��H;;�H;��H;��H;C�H;��H;��H;b�H;2�H;��H;��H;��H;��H;��H;v�H;��H;��H;��H;��H;��H;2�H;a�H;��H;��H;A�H;��H;��H;:�H;��H;��H;A�H;��H;��H;5�H;f�H;��H;��H;��H;m�H;=�H;�H;��H;;�H;��H;�H;u�H;�H;��H;4�H;�H;      
�H;`�H;F�H;��H;�H;t�H;��H;��H;��H;��H;��H;��H;X�H;��H;�H;=�H;Z�H;1�H;	�H;��H;��H;�H;��H;��H;,�H;��H;t�H;9�H;��H;��H;j�H;2�H;��H;��H;��H;��H;��H;��H;��H;��H;��H;5�H;l�H;��H;��H;9�H;w�H;��H;)�H;��H;��H;�H;��H;��H;	�H;4�H;Z�H;?�H;�H;��H;Z�H;��H;��H;��H;��H;��H;��H;u�H;�H;��H;F�H;`�H;      ��H;?�H;��H;_�H;\�H;��H;Y�H;��H;6�H;C�H;9�H;��H;!�H;;�H;��H;p�H;��H;��H;�H;��H;��H;��H;�H;��H;��H;)�H;��H;��H;9�H;��H;��H;x�H;Q�H;�H;�H;�H;�H;�H;�H; �H;Q�H;z�H;��H;��H;6�H;��H;��H;)�H;��H;��H;�H;��H;��H;��H;�H;��H;��H;r�H;��H;;�H;%�H;��H;9�H;D�H;7�H;��H;Y�H;��H;f�H;_�H;��H;L�H;      �H;H;�!H;�8H;�TH;QsH;E�H;ޫH;��H;��H;��H;��H; �H;&�H;��H;�H;��H;V�H;��H;��H;��H;��H;[�H;�H;��H;��H;�H;��H;x�H;G�H;��H;��H;��H;v�H;X�H;6�H;J�H;5�H;Z�H;v�H;��H;��H;��H;F�H;w�H;��H;�H;��H;��H;�H;[�H;��H;��H;��H;��H;W�H;��H;�H;��H;&�H; �H;��H;��H;��H;��H;ޫH;E�H;NsH;�TH;�8H;�!H;	H;      }DF;�RF;�zF;�F;�G;�\G;�G;]H;)IH;��H;��H;�H;�H;��H;�H;O�H;�H;P�H;��H;p�H;��H;��H;��H;o�H;��H;��H;��H;)�H;��H;��H;G�H;�H;��H;��H;��H;��H;��H;��H;��H;��H;��H;	�H;H�H;��H;��H;)�H;��H;��H;��H;l�H;��H;��H;��H;o�H;��H;R�H;�H;M�H;�H;��H;�H;�H;��H;��H;*IH;[H;�G;�\G;�G;�F;�zF;xRF;      ��A;�B;pB;�C;��C;~�D;quE;�DF;R�F;��G;�H;fH;�H;��H;j�H;(�H;��H;�H;��H;��H;E�H;��H;��H;��H;Q�H;��H;��H;��H;0�H;��H;��H;k�H;9�H;�H;��H;��H;��H;��H;��H;�H;9�H;n�H;��H;��H;-�H;��H;��H;��H;P�H;��H;��H;��H;?�H;��H;��H;�H;��H;(�H;j�H;��H;�H;fH;�H;��G;Q�F;�DF;quE;~�D;��C;�C;pB;�B;      �o8;K�8;ۏ9;}�:;��<;d>;VR@;�/B;��C;�PE;�zF;r\G;��G;OiH;F�H;��H;M�H;v�H;C�H;O�H;{�H;�H;��H;��H;��H;o�H;�H;��H;��H;:�H;��H;��H;��H;R�H;M�H;C�H;�H;C�H;O�H;T�H;��H;��H;��H;6�H;��H;��H;�H;p�H;��H;��H;��H;�H;u�H;O�H;E�H;x�H;J�H;��H;F�H;OiH;��G;s\G;�zF;�PE;��C;�/B;VR@;d>;��<;z�:;ݏ9;<�8;      �S%;`�%;U�';�M*;�-;��1;�5;)�9;�-=;CR@;�B;��D;9mF;�uG;�!H;$�H;�H;��H;*�H;��H;��H;R�H;&�H;��H;��H;��H;]�H;�H;��H;��H;H�H;�H;��H;��H;��H;��H;x�H;��H;��H;��H;��H;�H;I�H;��H;��H;�H;[�H;��H;��H;��H;#�H;P�H;��H;��H;*�H;��H;�H;#�H;�!H;�uG;;mF;��D;�B;@R@;�-=;'�9;�5;��1;�-;�M*;M�';O�%;      �W;�x;�;!�
;��;�;� ;��(;��/;I6;��;;�?;C;�PE;#�F;�G;�eH;\�H;��H;=�H;h�H;��H;P�H;�H;��H;��H;��H;��H;�H;��H;��H;h�H;=�H;-�H;��H;��H;��H;��H;��H;-�H;>�H;h�H;��H;��H;�H;��H;��H;��H;��H;�H;L�H;��H;e�H;>�H;��H;]�H;�eH;�G;$�F;�PE;C;�?;��;;I6;��/;��(;� ;�;Ѕ;�
;�;�x;      ���:$Ɔ:ʒ:8��:�:��:s��:l�	;�v; �#;�-;�5;�L<;��@;�(D;4DF;ōG;�HH;��H;�H;��H;h�H;��H;}�H;A�H;��H;��H;��H;��H;B�H;&�H;��H;��H;��H;R�H;B�H;D�H;B�H;R�H;��H;��H;��H;&�H;?�H;}�H;��H;��H;��H;?�H;x�H;��H;h�H;��H; �H;��H;�HH;čG;6DF;�(D;��@;�L<;�5;�-;�#;�v;l�	;s��:3��:�:4��:ʒ:Ɔ:      -.������깐|K��#
9�]:��k:�M�:��:�y;��;� $;��/;��8;��>;$C;:�E;�\G;h8H;ݥH;!�H;;�H;��H;R�H;��H;r�H;��H;��H;��H;��H;[�H;3�H;�H;��H;��H;��H;��H;��H;��H;��H;�H;3�H;[�H;��H;��H;��H;��H;r�H;��H;M�H;��H;;�H;�H;ޥH;h8H;�\G;:�E;$C;��>;��8;��/;� $;��;�y;��:�M�:��k:�]:�#
9�|K���,��      &Q^��X��F���)�	+��ζ���<� ;S��n:\��:���:��;`�;�M*;��5;�c=;~pB;��E;�JG;k8H;��H;��H;,�H;F�H;��H;��H;��H;�H;	�H;��H;��H;��H;u�H; �H;�H;�H;��H;�H;�H; �H;s�H;��H;��H;��H;�H;�H;��H;��H;��H;B�H;'�H;��H;��H;l8H;�JG;��E;~pB;�c=; �5;�M*;b�; �;���:^��:�n: ;S���<��ζ�+���)��F��X�      ^���0������ѻ"���ǐ�NX� 6�	�� tK�l?":N�:sb�:qi;F�%;q�3;�<;W0B;��E;�\G;�HH;]�H;��H;w�H;�H;R�H;X�H;��H;5�H;6�H;�H;��H;��H;}�H;o�H;n�H;L�H;n�H;o�H;|�H;��H;��H;�H;5�H;1�H;��H;V�H;S�H;�H;q�H;��H;]�H;�HH;�\G;��E;X0B;�<;q�3;H�%;ri;ub�:N�:p?":�sK�	��#6�PX�ǐ�����ѻ��4���      n�n�smj���]���J�W�1�04�+������	x��W���y�P*
90��:���:$�;[�#;j�2;�<;�pB;=�E;ōG;�eH;�H;M�H;��H;�H;��H;��H;W�H;f�H;T�H;+�H;�H;��H;��H;��H;��H;��H;��H;��H;�H;-�H;T�H;c�H;S�H;��H;��H;�H;��H;G�H;�H;�eH;čG;>�E;pB;�<;j�2;]�#;%�;���:2��:p*
9��y��W��	x����+��/4�V�1���J���]�vmj�      B<ͼ��ɼ�����֯�Ͷ��ㄼ��Y��*�����s��X�TrѺ��t?Q:��:��
;a�#;u�3;�c=;$C;8DF;�G;&�H;��H;%�H;P�H;�H;p�H;?�H;�H;��H;~�H;Q�H;j�H;&�H;�H;#�H;�H;&�H;l�H;Q�H;~�H;��H;�H;9�H;p�H;�H;Q�H;'�H;��H;#�H;�G;6DF;$C;�c=;w�3;`�#;��
;��:t?Q:��TrѺX��s������*���Y�ㄼͶ���֯�������ɼ      ��'�)�$����}��  ���ۼ����+����]��X!�=>ۻ|+��b*����L�>:��:%�;F�%;��5;��>;�(D;"�F;�!H;G�H;g�H;�H;��H;��H;�H;��H;��H;��H;��H;��H;��H;h�H;��H;h�H;��H;��H;��H;��H;��H;��H;��H;��H;��H;�H;g�H;C�H;�!H;"�F;�(D;��>;��5;H�%;$�;��:L�>:���b*�|+��=>ۻ�X!���]��+�������ۼ�  �}����)�$�      Ǹ���v����w�i�c��J�Є-�}��;缆沼ㄼ��;������j���5�p��x?Q:���:ui;�M*;��8;��@;�PE;�uG;OiH;��H;��H;&�H;7�H;��H;��H;��H;�H;��H;��H;��H;��H;��H;��H;��H;��H;��H;�H;��H;��H;��H;7�H;%�H;��H;��H;LiH;�uG;�PE;��@;��8;�M*;wi;���:�?Q:p�깋5��j��������;�ㄼ�沼�;�}�τ-��J�i�c���w��v��      }Hͽڪɽ�;�� "����ɸ����[�z0�t��(<ͼʾ��`�J�����j��_*���:��:{b�:d�;��/;�L<;C;<mF;��G;�H;�H; �H;!�H;X�H;h�H;�H;<�H;H�H;5�H;.�H;�H;�H;�H;/�H;5�H;G�H;=�H;�H;h�H;T�H;!�H;�H;�H;�H;��G;8mF;C;�L<;��/;d�;}b�:8��:��]*��j�����`�J�ʾ��'<ͼt��z0���[�ɸ���� "���;��ڪɽ      ��#-������Ա�ƽ`P���v���J�I����ۼ��`�J�����z+��NrѺ�*
9N�: �;� $;�5;�?;��D;o\G;fH;�H;��H;��H;��H;/�H;�H;i�H;��H;u�H;m�H;z�H;Q�H;z�H;j�H;r�H;��H;j�H;�H;/�H;��H;��H;��H;�H;fH;n\G;��D;�?;�5;� $; �;N�:p*
9TrѺz+������`�J�����ۼI���J��v��`P��ƽԱ轅����$-�       j�Yde�\0X��D�h{+�������x㻽[���TDX������ۼ˾����;�<>ۻX���y�p?":���:��;�-;��;;�B;�zF;�H;��H;��H;2�H;��H;�H;��H;��H;��H;��H;��H;��H;��H;��H;��H;��H;��H;��H;��H;�H;��H;2�H;��H;��H;�H;�zF;�B;��;;�-;��;���:p?":��y�X�<>ۻ��;�˾����ۼ���TDX�[���x㻽��콄��h{+��D�\0X�Yde�      ��Rh��m���I���|x���O��C(���Ҫɽ����TDX�I��'<ͼㄼ�X!��s���W��sK�d��:�y; �#;I6;CR@;�PE;��G;��H;��H;>�H;��H;��H;��H;��H;��H;��H;��H;��H;��H;��H;��H;��H;��H;��H;��H;��H;��H;>�H;��H;��H;��G;�PE;AR@;I6;"�#;�y;d��:�sK��W��s���X!�ㄼ'<ͼI��TDX�����Ҫɽ���C(���O��|x��I��m��Sh��      A����������%�;jɰ��G�� j�;�5��	�Ҫɽ[����J�t���沼��]�����	x�	���n:��:�v;��/;�-=;��C;O�F;,IH;��H;1�H;��H;.�H;��H;��H;��H;�H;"�H;)�H;:�H;)�H;"�H;�H;��H;��H;��H;.�H;��H;1�H;��H;*IH;R�F;��C;�-=;��/;�v;��:�n:	���	x������]��沼t���J�[���Ҫɽ�	�;�5� j��G��jɰ�%�;��徹���      �2�W�-�"�.E�����BKɾl����s�;�5���x㻽�v��
z0��;��+���*����6��9S��M�:l�	;��(;)�9;�/B;�DF;_H;ޫH;��H;��H;��H;��H;��H;%�H;H�H;V�H;P�H;o�H;R�H;U�H;H�H;"�H;��H;��H;��H;��H;��H;ܫH;^H;�DF;�/B;)�9;��(;n�	;�M�:�9S�6�����*��+���;�z0��v��x㻽��;�5���s�l��BKɾ����.E�"�W�-�      (3s�!cm�<�\�j�C�7�%�����TҾl�� j��C(����`P����[�}������Y�-��LX���<���k:i��:� ;�5;SR@;nuE;�G;?�H;U�H;��H;�H;W�H;��H;:�H;y�H;��H;k�H;��H;k�H;��H;x�H;7�H;�H;W�H;�H;��H;T�H;>�H;�G;quE;QR@;�5;� ;m��:��k:��<�JX�.����Y����}���[�`P����콭C(� j�l���TҾ���7�%�j�C�<�\�!cm�      �ޞ�������bF�A�W�Y�-����BKɾ�G����O����ƽɸ��Є-���ۼㄼ/4�ǐ��ζ��]:��:�;��1;d>;z�D;�\G;QsH;��H;x�H;q�H;4�H;��H;>�H;��H;��H;��H;��H;��H;��H;�H;;�H;��H;4�H;n�H;t�H;��H;OsH;�\G;{�D;�c>;��1;�;'��:�]:�ζ�ǐ�04�ㄼ��ۼЄ-�ɸ��ƽ�����O��G��BKɾ���Y�-�A�W�bF�������      ��ſ���Nw���ޞ�����A�W�7�%�����jɰ��|x�h{+�Ա����J��  �Ͷ��V�1� ��� +��#
9�:��;�-;��<;��C;�G;�TH;Y�H;�H;��H;��H;i�H;G�H;��H;��H;��H;�H;��H;��H;��H;E�H;i�H;��H;��H;	�H;Y�H;�TH;�G;��C;��<;"�-;��; �:`#
9+� ���V�1�Ͷ���  ��J���Ա�h{+��|x�jɰ�����7�%�A�W������ޞ�Nw�����      ����� �Կp���ޞ�bF�j�C�.E�%�;�I���D��� "��i�c�}��֯���J��ѻ��)��|K�@��:+�
;�M*;��:;�C;�F;�8H;d�H;��H;��H;��H;R�H;O�H;��H;��H;��H;�H;��H;��H;��H;N�H;Q�H;��H;��H;��H;c�H;�8H;�F;�C;}�:;�M*;)�
;F��:�|K���)��ѻ��J��֯�}�i�c� "�����D��I��%�;.E�j�C�bF��ޞ�p�� �Կ��      ��������� �ԿNw�����<�\�"����m��\0X�����;����w����������]��黲F�0��ʒ:
�;I�';̏9;/pB;�zF;�!H;��H;E�H;-�H;��H;Y�H;P�H;��H;��H;��H;&�H;��H;��H;��H;N�H;X�H;��H;(�H;B�H;��H;�!H;�zF;/pB;ɏ9;K�';
�;ʒ:@�깲F��黩�]����������w��;�����\0X�m�����"�<�\����Nw�� �Կ��𿞏�      "$�������忊�����!cm�W�-�����Rh��Yde�#-�ڪɽ�v��)�$���ɼumj�0����X�<��
Ɔ:�x;P�%;?�8;{B;{RF;H;<�H;b�H;�H;~�H;T�H;K�H;��H;��H;��H;:�H;��H;��H;��H;I�H;T�H;~�H;�H;_�H;<�H;H;zRF;{B;=�8;V�%;�x;
Ɔ:D���X�/���vmj���ɼ)�$��v��ڪɽ#-�Yde�Rh������W�-�!cm��������忞����      �>���8���*�O������˿p��G�b�E\�6m־^��S�:��J�*��G�B�=��������#/��ܯ��$�>:�t�:]p ;�J6;EA;�IF;�NH;�H;"I;�I;'I;�I;�I;I;� I;��H;@�H;��H;� I;I;�I;�I;'I;�I;"I;�H;�NH;�IF;EA;�J6;`p ;�t�:(�>:௕�#/���������=��G�B�*���J�S�:�^��6m־E\�G�b�p���˿����O���*���8�      ��8��4��g&�7��>����<ƿ򲗿�>]�î�Q�Ѿ�p���*7����&W��MR?� }�o8�������b�����G:� �:�!;"�6;-lA;�YF;�TH;�H;/"I;�I;I;�I;]I;I;y I;��H;)�H;��H;z I;I;\I;�I;I;�I;,"I;�H;�TH;�YF;-lA;�6;�!;� �:��G:d��������o8�� }�MR?�'W�����*7��p��Q�Ѿî��>]�򲗿�<ƿ>���7���g&��4�      ��*��g&��#�v�V[�sL�������M�s5��>ľ����,��D�뒐��5�2�ݼ���q
���x�@tk��b:ml�:#;ڗ7;��A;��F;�dH;�I;l"I;I;}I;VI;	I;�I;7 I;��H;��H;��H;5 I;�I;I;TI;}I;I;k"I;�I;�dH;��F;��A;֗7;#;ml�:�b:Htk���x��q
���2�ݼ�5�뒐��DὭ�,����>ľs5���M����sL��V[�v��#��g&�      O�7��v����˿B1��:�y�Ŏ6��z �����5�l�+��ͽ$�����&���˼<�k������X�$� ����:[�;!&;�9;��B;!�F;�}H;�	I;x"I;BI;�I;�I;�I;]I;��H;9�H;��H;9�H;��H;]I;�I;�I;�I;AI;u"I;�	I;�}H;!�F;��B;�9;%&;[�;���:(� ���X����<�k���˼��&�$����ͽ+�5�l������z �Ŏ6�:�y�B1���˿���v�7��      ����>���V[忸˿�T���}�R�®��E۾ԗ����M���	������j��3�d����O�0�׻��/����r��:� 
;*;m;;kC;�'G;��H;I;"I;I;�I;�
I;�I;�I;\�H;��H;�H;��H;Z�H;�I;�I;�
I;�I;I;"I;I;��H;�'G;kC;i;;"*;� 
;t��:�����/�.�׻��O�d���3���j������	���M�ԗ���E۾®�}�R���T���˿V[�>���      �˿�<ƿsL��B1����>]���)�%��ֳ���{���,�t��)��S`I��J���,���3/��+���� �`069�4�:��;p.;2.=;vaD;��G;{�H;�I;R!I;nI;bI;�	I;�I; I;��H;'�H;w�H;'�H;��H; I;�I;�	I;bI;kI;O!I;�I;z�H;��G;vaD;/.=;p.;��;�4�:@069�� ��+���3/��,���J��S`I�)��t�齧�,���{�ֳ�%����)��>]��B1��sL���<ƿ      p��򲗿���:�y�}�R���)�ov��>ľ^���I�Zl����������&�ԮҼ�}�+B���������P�!:%+�:Jz;�3;lj?;�\E;��G;��H;�I;�I;�I;�I;�I;�I;. I;��H;w�H;��H;w�H;��H;0 I;�I;�I;�I;�I;�I;�I;��H;��G;�\E;ij?;�3;Jz;'+�:H�!:��������+B��}�ԮҼ��&��������Zl��I�^���>ľov���)�}�R�:�y����򲗿      G�b��>]���M�Ŏ6�®�%���>ľ%q��|�Z�+�T9ݽ"W����L����!F�� �G���׻�;�n��Ȋ:�i;,P$;�7;{�A;#JF;DCH;��H;� I;}I;�I;-I;@I;�I;*�H;��H;��H;%�H;��H;��H;,�H;�I;BI;-I;�I;zI;� I;��H;DCH; JF;w�A;�7;,P$;�i;�Ȋ:n��;���׻ �G�!F�������L�"W��T9ݽ+�|�Z�%q���>ľ%��®�Ŏ6���M��>]�      E\�î�s5��z ��E۾ֳ�^��|�Z�N?#����A����j�&��Dϼ ����������lۺ�:�9�4�:g�;r�,;��;;H�C;�G;]�H;�I;�!I;�I;TI;;I;�I;SI;0�H;�H;��H;7�H;��H;�H;2�H;TI;�I;;I;RI;�I;�!I;�I;`�H;�G;F�C;��;;r�,;i�;�4�:�:�9�lۺ������� ��Eϼ&����j��A�����M?#�|�Z�^��ֳ��E۾�z �s5�î�      6m־Q�Ѿ�>ľ����ԗ����{��I�+�����V���{�?�/�&���,��:=�7�һH�@��� �<�k:)�:b;��3;Cj?;|2E;��G;|�H;FI;� I;�I;�I;4	I;I;��H;�H;��H;��H;m�H;��H;��H;�H;��H;I;5	I;�I;�I;� I;FI;�H;��G;{2E;Bj?;��3;b;)�:<�k:�� �J�@�7�һ:=��,��&��?�/��{��V�����+��I���{�ԗ�������>ľQ�Ѿ      ^���p����5�l���M���,�Zl�T9ݽ�A���{���5��J��;���T[�?�����P�� Q�9��:��;8*;3�9;pkB;�F;�NH;��H;/ I;�I;�I;/I;"I;UI;u�H;��H;��H;��H;��H;��H;��H;��H;t�H;XI;"I;/I;�I;�I;0 I;��H;�NH;�F;nkB;3�9;6*;��;��:8Q�9P������?��T[�;���J����5��{��A��T9ݽZl���,���M�5�l����p��      S�:��*7���,�+���	�t�齄���"W����j�?�/��J���I���k�f� .��F������Ɋ:o�:&;or3;2�>;?�D;~�G;`�H;I;A!I;�I;�I;�
I;I;u I;��H;��H;��H;��H;x�H;��H;��H;��H;��H;w I;I;�
I;�I;�I;A!I;I;^�H;{�G;<�D;2�>;or3;&;o�:Ɋ: ��F�� .��f��k��I���J��?�/���j�"W������t�齄�	�+���,��*7�      �J�����D��ͽ���(�������L�&��&��;���k����^I����/�/�К>:d��:�B;w�,;��:;B�B;�xF;�<H;�H;I;�I;�I;XI;�I;�I;��H;��H;M�H;��H;��H;��H;��H;��H;N�H;��H;��H;�I;�I;XI;�I;�I;I;�H;�<H;�xF;B�B;��:;v�,;�B;l��:Ț>:/���/�^I������k�;��&��&����L����(������ͽ�D����      *��&W��꒐�$�����j�R`I���&����Dϼ�,���T[�f�^I��E;�,nk�:H5�:�;&;�6;�!@;L2E;�G;��H;I;!I;fI;%I;I;NI;� I;��H;�H;��H;z�H;��H;_�H;��H;z�H;��H;�H;��H;� I;PI;I;'I;fI;!I;I;��H;�G;L2E;�!@;�6;&;�;B5�::,nk�E;�^I��f��T[��,��Dϼ�����&�R`I���j�$���꒐�&W��      F�B�MR?��5���&��3��J��ԮҼ!F�� ��;=�?�.����/�8nk���9j׳:��;D!;l3;�=;��C;5�F;*dH;�H;�I;&I;�I;:I;�I;�I;\�H;�H;��H;��H;[�H;��H;Q�H;��H;\�H;��H;��H;�H;\�H;�I;�I;<I;�I;)I;�I;�H;%dH;5�F;��C;�=;l3;I!;��;j׳:��98nk���/�.��?�<=� ��!F��ԮҼ�J���3���&��5�NR?�      <�� }�0�ݼ��˼d���,���}� �G����7�һ����G��/��:r׳:�;�b;ģ0;�<;��B;�IF;�H;=�H;�I;� I;1I;PI;r
I;�I;: I;H�H;l�H;%�H;?�H;;�H;��H;U�H;��H;;�H;@�H;%�H;o�H;H�H;: I;�I;t
I;NI;4I;� I;�I;9�H;�H;�IF;��B;�<;ţ0;�b;�;p׳:�:/�G������8�һ��� �G��}��,��d����˼0�ݼ }�      ����m8����;�k���O��3/�)B���׻����H�@�P�� ��Ě>:B5�:��;}b;��/;?;;R�A;��E;ؿG;�H;�
I;� I;I;I;�I;�I;�I;��H;V�H;��H;��H;�H;/�H;��H;M�H;��H;/�H;�H;��H;��H;V�H;��H;�I;�I;�I;I;I;| I;�
I;�H;ؿG;��E;R�A;B;;��/;|b;��;>5�:��>: ��P��J�@�������׻)B��3/���O�;�k���o8��      ������q
����0�׻�+�������;��lۺĖ �8Q�9Ɋ:d��:�;G!;��0;@;;ғA;�pE;��G;�H;��H;�I;OI;qI;=I;�I;�I;�H;]�H;��H;�H;;�H;�H;�H;}�H;W�H;}�H;�H;�H;:�H;!�H;��H;\�H;�H;�I;�I;>I;qI;NI;�I;��H;��H;��G;�pE;ՓA;?;;��0;F!;�;`��:Ɋ: Q�9Ȗ ��lۺ�;������+��-�׻����q
���       /�������x���X���/��� �����8n칠:�94�k:��:o�:�B;&;l3;�<;R�A;�pE;vtG;}H;A�H;BI;�I;^I;I;�
I;I;n I;k�H;@�H;��H;��H;��H;��H;�H;��H;��H;��H;�H;��H;��H;��H;��H;=�H;i�H;o I;I;�
I;I;ZI;�I;BI;@�H;}H;wtG;�pE;O�A;�<;l3;&;�B;}o�:��:0�k:�:�98n������ ���/���X���x����      ֯��B���8tk�(� ���� 069H�!:�Ȋ:�4�:)�:��;";r�,;�6;�=;��B;��E;��G;}H;��H;�I;. I;�I;uI;�I;FI;�I;e�H;�H;Z�H;�H;/�H;��H;��H;�H;��H;��H;��H;�H;��H;��H;0�H;�H;W�H;�H;e�H;�I;FI;�I;qI;�I;. I;�I;��H;}H;��G;��E;��B;�=;�6;r�,;";��;!�:�4�:�Ȋ:H�!:@069H��(� �8tk�T���      <�>:�G: �b:���:`��:�4�:%+�:�i;f�;b;5*;kr3;��:;�!@;��C;�IF;ؿG;�H;A�H;�I;5 I;^I;VI;�I;0I;{I;=�H;��H;��H;��H;j�H;��H;��H;��H;2�H;��H;��H;��H;2�H;��H;��H;��H;j�H;��H;��H;��H;<�H;|I;0I;�I;VI;^I;4 I;�I;A�H;�H;׿G;�IF;��C;�!@;��:;kr3;3*;b;g�;�i;'+�:�4�:d��:���:,�b:��G:      �t�:� �:�l�:R�;� 
;�;Sz;0P$;v�,;��3;7�9;5�>;B�B;L2E;5�F;�H;�H;��H;AI;. I;]I;�I;UI;�I;I;��H;A�H;l�H;��H;��H;�H;��H;��H;��H;T�H;�H;��H;�H;T�H;��H;��H;��H;��H;��H;��H;l�H;@�H;��H;I;�I;SI;�I;[I;1 I;AI;��H;
�H;�H;6�F;K2E;A�B;4�>;6�9;��3;u�,;3P$;Sz;�;� 
;R�;�l�:� �:      `p ;�!;#;&;*;p.;�3;�7;��;;Dj?;pkB;A�D;�xF;�G;)dH;9�H;�
I;�I;�I;�I;VI;WI;�I;uI;R�H;��H;��H;G�H;�H;5�H;��H;��H;��H;	�H;s�H;9�H;&�H;9�H;s�H;	�H;��H;��H;��H;2�H;�H;G�H;��H;��H;U�H;tI;�I;WI;RI;�I;�I;�I;�
I;8�H;'dH;�G;�xF;A�D;qkB;Bj?;��;;�7;�3;p.;*;&;#;�!;      �J6;-�6;��7;�9;m;;/.=;sj?;w�A;K�C;}2E;�F;��G;�<H;��H;�H;�I;} I;PI;]I;tI;�I;�I;uI;j�H;��H;��H;��H;O�H;\�H;��H;��H;��H;��H;G�H;��H;��H;i�H;��H;��H;I�H;��H;��H;��H;��H;Y�H;O�H;��H;��H;��H;h�H;uI;�I;�I;tI;]I;RI;| I;�I;�H;��H;�<H;�G;�F;|2E;K�C;z�A;qj?;1.=;t;;�9;�7;�6;      !EA;7lA;w�A;��B;	kC;xaD;�\E;!JF;�G;��G;�NH;b�H;�H;I;�I;� I;I;rI;I;�I;3I;I;W�H;��H;�H;��H;X�H;m�H;��H;��H;��H;��H;��H;~�H;�H;��H;��H;��H;�H;}�H;��H;��H;��H;��H;��H;m�H;V�H;��H;�H;��H;W�H;I;2I;�I;I;uI;I;� I;�I;I;�H;b�H;�NH;��G;�G; JF;�\E;yaD;	kC;��B;x�A;7lA;      �IF;�YF;�F;�F;�'G;��G;��G;ACH;`�H;~�H;��H; I;I;!I;&I;/I;I;;I;�
I;CI;zI;��H;��H;��H;��H;��H;��H;��H;��H;��H;��H;��H;W�H;��H;q�H;S�H;B�H;S�H;r�H;��H;S�H;��H;��H;��H;��H;��H;��H;��H;��H;��H;��H;��H;tI;CI;�
I;;I;I;/I;&I;!I;I; I;��H;|�H;`�H;ACH;��G;��G;�'G;�F;�F;�YF;      �NH;�TH;�dH;�}H;��H;|�H;��H;��H;�I;FI;2 I;E!I;�I;gI;�I;QI;�I;�I;I;�I;?�H;B�H;��H;��H;S�H;��H;��H;��H;��H;��H;��H;�H;��H;,�H;��H;��H;��H;��H;��H;*�H;��H;�H;��H;��H;��H;��H;��H;��H;T�H;��H;��H;D�H;:�H;�I;I;�I;�I;PI;�I;gI;�I;E!I;2 I;FI;�I;��H;��H;z�H;�H;�}H;�dH;�TH;      �H;��H;�I;�	I;I;�I;�I;� I;�!I;� I;�I;�I;�I;)I;=I;t
I;�I;�I;l I;h�H;��H;l�H;J�H;Q�H;i�H;��H;��H;��H;��H;��H;�H;n�H;	�H;��H;n�H;?�H;6�H;?�H;n�H;��H;�H;n�H;�H;��H;�H;��H;��H;��H;j�H;Q�H;H�H;n�H;��H;h�H;l I;�I;�I;r
I;:I;'I;�I;�I;�I;� I;�!I;� I;�I;�I;I;�	I;�I;��H;      %"I;/"I;h"I;|"I;"I;O!I;�I;�I;�I;�I;�I;�I;YI;I;�I;�I;�I;�H;l�H;�H;��H;��H;�H;`�H;��H;��H;��H;��H;��H;
�H;c�H;��H;�H;0�H;��H;��H;��H;��H;��H;0�H;|�H;��H;c�H;�H;��H;��H;��H;��H;��H;`�H;�H;��H;��H;�H;k�H;�H;�I;�I;�I;I;XI;�I;�I;�I;�I;�I;�I;N!I;"I;|"I;i"I;'"I;      �I;�I;I;AI;I;rI;�I;�I;\I;�I;9I;�
I;�I;ZI;�I;> I;��H;Z�H;=�H;\�H;��H;��H;0�H;��H;��H;��H;��H;��H;�H;S�H;��H;z�H;�H;��H;��H;��H;o�H;��H;��H;��H;��H;{�H;��H;R�H;�H;��H;��H;��H;��H;��H;/�H;��H;��H;\�H;=�H;\�H;��H;< I;�I;WI;�I;�
I;9I;�I;]I;�I;�I;rI;I;BI;I;�I;      *I;I;�I;�I;�I;`I;�I;6I;EI;;	I;-I;I;�I;� I;b�H;P�H;`�H;��H;��H;�H;o�H;�H;��H;��H;��H;��H;��H;�H;a�H;��H;]�H;��H;��H;s�H;@�H;#�H;�H;#�H;@�H;s�H;��H;��H;\�H;��H;c�H;�H;��H;��H;��H;��H;��H;�H;m�H;	�H;��H;��H;]�H;O�H;`�H;� I;�I;I;,I;=	I;EI;8I;�I;aI;�I;�I;�I;I;      �I;�I;ZI;�I;�
I;�	I;�I;KI;�I;I;\I;� I;��H;��H;�H;w�H;��H;"�H;��H;:�H;��H;��H;��H;��H;��H;��H;�H;o�H;��H;z�H;��H;��H;X�H;1�H;��H;��H;��H;��H;��H;1�H;U�H;��H;��H;{�H;��H;o�H;�H;��H;��H;��H;��H;��H;��H;9�H;��H;$�H;��H;v�H;�H;��H;��H;� I;\I;I;�I;II;�I;�	I;�
I;�I;ZI;�I;      �I;oI;I;�I;�I;�I;�I;�I;\I;��H;|�H;��H;��H;"�H;��H;,�H;��H;:�H;��H;��H;��H;��H;��H;��H;��H;V�H;��H;
�H;��H;�H;��H;Z�H;�H;��H;��H;��H;��H;��H;��H;��H;�H;[�H;��H;�H;��H;
�H;��H;T�H;��H;��H;��H;��H;��H;��H;��H;;�H;��H;,�H;��H;"�H;��H;��H;|�H;��H;\I;�I;�I;�I;�I;�I;I;hI;      #I;I;�I;dI;�I;� I;3 I;7�H;7�H;�H;��H;��H;S�H;��H;��H;J�H;#�H;	�H;��H;��H;��H;��H;�H;L�H;y�H;��H;&�H;��H;.�H;��H;q�H;1�H;��H;��H;��H;��H;p�H;��H;��H;��H;��H;4�H;q�H;��H;0�H;��H;&�H;��H;z�H;J�H;�H;��H;��H;��H;��H;
�H;"�H;I�H;��H;��H;S�H;��H;��H;�H;9�H;9�H;3 I;� I;�I;dI;�I;I;      � I;� I;C I;��H;v�H;��H;��H;�H;#�H;��H;��H;��H;��H;��H;a�H;F�H;:�H;�H;�H;�H;:�H;V�H;q�H;��H;�H;o�H;��H;n�H;��H;��H;@�H;��H;��H;��H;k�H;`�H;a�H;`�H;k�H;��H;��H; �H;@�H;��H;��H;n�H;��H;q�H;�H;��H;s�H;V�H;7�H;�H;	�H;�H;9�H;E�H;b�H;��H;��H;��H;��H;�H;%�H;�H;��H;��H;m�H;��H;B I;� I;      ��H;��H;��H;?�H;��H;#�H;��H;��H;��H;��H;��H;��H;��H;��H;��H;��H;��H;{�H;��H;��H;��H;�H;;�H;��H;��H;P�H;��H;?�H;��H;�H;$�H;��H;��H;��H;`�H;E�H;E�H;E�H;`�H;��H;��H;��H;$�H;��H;��H;?�H;��H;O�H;��H;��H;;�H;�H;��H;��H;��H;}�H;��H;��H;��H;��H;��H;��H;��H;��H;��H;��H;��H;'�H;��H;<�H;��H;��H;      =�H;3�H;�H;��H;'�H;u�H;��H;/�H;?�H;m�H;��H;��H;��H;i�H;W�H;^�H;U�H;S�H;��H;��H;��H;��H;$�H;l�H;��H;@�H;��H;:�H;��H;q�H;�H;��H;��H;s�H;a�H;F�H;B�H;F�H;a�H;s�H;��H;��H;�H;s�H;��H;:�H;��H;A�H;��H;i�H;$�H;��H;��H;��H;��H;T�H;T�H;^�H;W�H;i�H;��H;��H;��H;p�H;@�H;-�H;��H;y�H;�H;��H;�H;+�H;      ��H;��H;��H;<�H;��H;#�H;��H;��H;��H;��H;��H;��H;��H;��H;��H;��H;��H;{�H;��H;��H;��H;�H;;�H;��H;��H;P�H;��H;?�H;��H;�H;$�H;��H;��H;��H;`�H;E�H;E�H;E�H;`�H;��H;��H;��H;$�H;��H;��H;?�H;��H;O�H;��H;��H;;�H;�H;��H;��H;��H;}�H;��H;��H;��H;��H;��H;��H;��H;��H;��H;��H;��H;'�H;��H;?�H;��H;��H;      � I;� I;B I;��H;v�H;��H;��H;�H;%�H; �H;��H;��H;��H;��H;b�H;E�H;:�H;�H;	�H;�H;;�H;V�H;s�H;��H;�H;o�H;��H;n�H;��H;��H;@�H;��H;��H;��H;k�H;`�H;a�H;`�H;k�H;��H;��H;�H;@�H;��H;��H;n�H;��H;o�H;�H;��H;q�H;V�H;7�H;�H;�H;�H;9�H;F�H;b�H;��H;��H;��H;��H; �H;#�H;�H;��H;��H;m�H;��H;A I;� I;      %I;I;�I;dI;�I;� I;3 I;7�H;7�H;�H;��H;��H;S�H;��H;��H;I�H;#�H;	�H;��H;��H;��H;��H;�H;L�H;z�H;��H;&�H;��H;/�H;��H;q�H;1�H;��H;��H;��H;��H;p�H;��H;��H;��H;��H;4�H;q�H;��H;0�H;��H;&�H;��H;y�H;J�H;�H;��H;��H;��H;��H;
�H; �H;J�H;��H;��H;S�H;��H;��H;�H;9�H;7�H;3 I;� I;�I;dI;�I;I;      �I;oI;I;�I;�I;�I;�I;�I;\I;��H;|�H;��H;��H;"�H;��H;,�H;��H;:�H;��H;��H;��H;��H;��H;��H;��H;V�H;��H;
�H;��H;�H;��H;Z�H;�H;��H;��H;��H;��H;��H;��H;��H;�H;\�H;��H;�H;��H;
�H;��H;T�H;��H;��H;��H;��H;��H;��H;��H;:�H;��H;,�H;��H;"�H;��H;��H;|�H;��H;\I;�I;�I;�I;�I;�I;I;nI;      �I;�I;]I;�I;�
I;�	I;�I;II;�I;I;\I;� I;��H;��H;�H;v�H;��H;"�H;��H;:�H;��H;��H;��H;��H;��H;��H;�H;o�H;��H;z�H;��H;��H;W�H;1�H;��H;��H;��H;��H;��H;1�H;U�H;��H;��H;{�H;��H;o�H;�H;��H;��H;��H;��H;��H;��H;:�H;��H;$�H;��H;w�H;�H;��H;��H;� I;\I;I;�I;HI;�I;�	I;�
I;�I;]I;�I;      *I;I;�I;�I;�I;`I;�I;6I;EI;<	I;,I;I;�I;� I;`�H;P�H;_�H;��H;��H;	�H;q�H;�H;��H;��H;��H;��H;��H;�H;a�H;��H;\�H;��H;��H;s�H;@�H;#�H;�H;#�H;@�H;s�H;��H;��H;]�H;��H;c�H;�H;��H;��H;��H;��H;��H;�H;m�H;�H;��H;��H;]�H;P�H;b�H;� I;�I;I;*I;<	I;EI;6I;�I;aI;�I;�I;�I;I;      �I;�I;I;BI;I;oI;�I;�I;_I;�I;9I;�
I;�I;XI;�I;< I;��H;Z�H;=�H;^�H;��H;��H;0�H;��H;��H;��H;��H;��H;�H;S�H;��H;z�H;��H;��H;��H;��H;o�H;��H;��H;��H;��H;{�H;��H;R�H;�H;��H;��H;��H;��H;��H;/�H;��H;��H;\�H;=�H;\�H;��H;? I;�I;XI;�I;�
I;9I;�I;_I;�I;�I;pI;I;AI;I;�I;      "I;+"I;m"I;y"I;"I;K!I;�I;�I;�I;�I;�I;�I;XI;I;�I;�I;�I;�H;k�H;�H;��H;��H;�H;`�H;��H;��H;��H;��H;��H;�H;c�H;��H;~�H;0�H;��H;��H;��H;��H;��H;0�H;~�H;��H;c�H;�H;��H;��H;��H;��H;��H;`�H;�H;��H;��H;�H;l�H;�H;�I;�I;�I;I;YI;�I;�I;�I;�I;�I;�I;M!I;"I;x"I;o"I;,"I;      �H;�H;�I;�	I;I;�I;�I;� I;�!I;� I;�I;�I;�I;(I;<I;r
I;�I;�I;l I;h�H;��H;n�H;J�H;Q�H;j�H;��H;��H;��H;��H;��H;�H;n�H;�H;��H;m�H;?�H;6�H;?�H;n�H;��H;�H;o�H;�H;��H;�H;��H;��H;��H;i�H;Q�H;H�H;l�H;��H;h�H;l I;�I;�I;u
I;=I;(I;�I;�I;�I;� I;�!I;� I;�I;�I;I;�	I;�I;��H;      �NH;�TH;�dH;�}H;��H;x�H;��H;��H;�I;GI;2 I;E!I;�I;fI;�I;QI;�I;�I;I;�I;A�H;D�H;��H;��H;T�H;��H;��H;��H;��H;��H;��H;�H;��H;*�H;��H;��H;��H;��H;��H;*�H;��H;�H;��H;��H;��H;��H;��H;��H;S�H;��H;��H;B�H;:�H;�I;I;�I;�I;PI;�I;gI;�I;E!I;2 I;GI;�I;��H;��H;w�H;��H;�}H;�dH;�TH;      �IF;�YF;�F; �F;�'G;��G;��G;ACH;_�H;~�H;��H;I;I;!I;%I;/I;I;:I;�
I;CI;{I;��H;��H;��H;��H;��H;��H;��H;��H;��H;��H;��H;V�H;��H;o�H;S�H;B�H;S�H;r�H;��H;S�H;��H;��H;��H;��H;��H;��H;��H;��H;��H;��H;��H;tI;CI;�
I;=I;I;/I;&I;!I;I; I;��H;{�H;_�H;@CH;��G;��G;�'G;�F;��F;�YF;      !EA;7lA;w�A;��B;kC;xaD;�\E;JF;�G;��G;�NH;b�H;�H;I;�I;� I;I;rI;I;�I;4I;I;Y�H;��H;�H;��H;W�H;m�H;��H;��H;��H;��H;��H;}�H;�H;��H;��H;��H;�H;}�H;��H;��H;��H;��H;��H;m�H;W�H;��H;�H;��H;V�H;I;2I;�I;I;uI;I;� I;�I;I;�H;b�H;�NH;��G;�G; JF;�\E;xaD;kC;��B;x�A;8lA;      �J6;,�6;�7;�9;f;;5.=;pj?;x�A;M�C;2E;�F;�G;�<H;��H;�H;�I;} I;PI;]I;tI;�I;�I;vI;m�H;��H;��H;��H;O�H;]�H;��H;��H;��H;��H;G�H;��H;��H;i�H;��H;��H;G�H;��H;��H;��H;��H;Y�H;O�H;�H;��H;��H;j�H;tI;�I;�I;tI;]I;RI;| I;�I;�H;��H;�<H;��G;�F;|2E;M�C;x�A;pj?;5.=;t;;�9;�7;�6;      [p ;!;&#;&;*;p.;�3;�7;��;;Cj?;qkB;A�D;�xF;�G;'dH;9�H;�
I;�I;�I;�I;YI;WI;�I;vI;U�H;��H;��H;G�H;�H;5�H;��H;��H;��H;	�H;s�H;9�H;&�H;9�H;s�H;	�H;��H;��H;��H;2�H;�H;G�H;��H;��H;R�H;rI;�I;WI;RI;�I;�I;�I;�
I;9�H;*dH;�G;�xF;A�D;qkB;Bj?;��;;�7;�3;p.;*;&;#;�!;      �t�:� �:�l�:R�;� 
;�;Sz;1P$;u�,;��3;7�9;4�>;A�B;K2E;5�F;�H;
�H;��H;AI;0 I;_I;�I;UI;�I;I;��H;A�H;l�H;��H;��H;��H;��H;��H;��H;T�H;�H;��H;�H;T�H;��H;��H;��H;�H;��H;��H;l�H;>�H;��H;I;�I;SI;�I;[I;0 I;AI;��H;
�H;�H;6�F;L2E;B�B;7�>;6�9;��3;v�,;0P$;Sz;�;� 
;R�;�l�:� �:      $�>:��G:4�b:���:`��:�4�:-+�:�i;f�;b;5*;kr3;��:;�!@;��C;�IF;ؿG;�H;A�H;�I;6 I;^I;VI;�I;0I;|I;=�H;��H;��H;��H;j�H;��H;��H;��H;2�H;��H;��H;��H;2�H;��H;��H;��H;j�H;��H;��H;��H;<�H;{I;0I;�I;UI;^I;2 I;�I;A�H;�H;׿G;�IF;��C;�!@;��:;kr3;6*;b;i�;�i;++�:�4�:h��:���:8�b:��G:      ޯ��@���,tk�,� ����0069H�!:�Ȋ:�4�:#�:��;";p�,;�6;�=;��B;��E;��G;}H;��H;�I;. I;�I;wI;�I;FI;�I;e�H;�H;Z�H;�H;/�H;��H;��H;�H;��H;��H;��H;�H;��H;��H;0�H;�H;W�H;�H;e�H;�I;FI;�I;qI;�I;. I;�I;��H;}H;��G;��E;��B;�=;�6;r�,; ;��;'�:�4�:�Ȋ:H�!:0069p��,� �8tk�T���       /�������x���X���/��� �����8n치:�90�k:��:}o�:�B;&;l3;�<;R�A;�pE;wtG;}H;D�H;BI;�I;^I;I;�
I;I;o I;l�H;@�H;��H;��H;��H;��H;�H;��H;��H;��H;�H;��H;��H;��H;��H;=�H;g�H;n I;I;�
I;I;ZI;�I;BI;>�H;}H;vtG;�pE;O�A;�<;n3;&;�B;o�:��:4�k:�:�9@n������ ���/���X���x����      ������q
����1�׻�+�������;��lۺȖ �0Q�9Ɋ:`��:�;F!;��0;@;;ԓA;�pE;��G;�H;��H;�I;RI;qI;>I;�I;�I;�H;]�H;��H; �H;;�H;�H;�H;}�H;W�H;}�H;�H;�H;:�H;!�H;��H;\�H;�H;�I;�I;>I;qI;KI;�I;��H;ߎH;��G;�pE;ԓA;?;;��0;G!;�;d��:Ɋ:8Q�9Ė ��lۺ�;������+��.�׻����q
���      ����m8����<�k���O��3/�*B���׻����J�@�P�� ����>:>5�:��;|b;��/;?;;R�A;��E;ٿG;�H;�
I;� I;I;I;�I;�I;�I;��H;V�H;��H;��H;�H;/�H;��H;M�H;��H;/�H;�H;��H;��H;V�H;��H;�I;�I;�I;I;I;| I;�
I;�H;տG;��E;R�A;B;;��/;}b;��;B5�:Ě>: ��P��J�@�������׻*B��3/���O�<�k���n8��      =�� }�0�ݼ��˼d���,���}� �G����8�һ����G��/��:l׳:�;�b;ģ0;�<;��B;�IF;�H;<�H;�I;� I;2I;QI;t
I;�I;: I;H�H;m�H;&�H;@�H;;�H;��H;U�H;��H;;�H;?�H;#�H;o�H;H�H;: I;�I;r
I;MI;2I;� I;�I;9�H;�H;�IF;��B;�<;ţ0;b;�;p׳:�:/�G������7�һ����G��}��,��d����˼0�ݼ }�      F�B�MR?��5���&��3��J��ԮҼ!F�� ��<=�?�.����/�8nk���9j׳:��;F!;l3;�=;��C;5�F;*dH;�H;�I;)I;�I;<I;�I;�I;\�H;�H;��H;��H;\�H;��H;Q�H;��H;[�H;��H;��H;�H;\�H;�I;�I;:I;�I;(I;�I;�H;#dH;5�F;��C;�=;l3;G!;��;j׳:��98nk���/�.��?�;=� ��"F��ԮҼ�J���3���&��5�NR?�      *��&W��꒐�$�����j�R`I���&����Dϼ�,���T[�f�^I��E;�,nk�:H5�:�;&;�6;�!@;L2E;�G;��H;I;!I;gI;'I;I;PI;� I;��H;�H;��H;z�H;��H;_�H;��H;z�H;��H;�H;��H;� I;NI;I;%I;fI;!I;I;��H;�G;L2E;�!@;�6;&;�;D5�::,nk�E;�^I��f��T[��,��Dϼ�����&�R`I���j�$���꒐�&W��      �J�����D��ͽ���(�������L�&��&��;���k����^I����/�/�К>:h��:�B;v�,;��:;B�B;�xF;�<H;�H;I;�I;�I;YI;�I;�I;��H;��H;N�H;��H;��H;��H;��H;��H;M�H;��H;��H;�I;�I;UI;�I;�I;I;�H;�<H;�xF;B�B;��:;v�,;�B;l��:Ț>:/���/�^I������k�;��&��&����L����(������ͽ�D����      S�:��*7���,�+���	�t�齄���"W����j�?�/��J���I���k�f� .��F��  ��Ɋ:o�:%;lr3;2�>;?�D;~�G;^�H; I;C!I;�I;�I;�
I;I;u I;��H;��H;��H;��H;x�H;��H;��H;��H;��H;v I;I;�
I;�I;�I;@!I;I;`�H;{�G;<�D;2�>;or3;%;o�:Ɋ:  ��G�� .��f��k��I���J��?�/���j�"W������t�齄�	�+���,��*7�      ^���p����5�l���M���,�Zl�T9ݽ�A���{���5��J��;���T[�?�����P��0Q�9��:��;5*;3�9;pkB;�F;�NH;��H;0 I;�I;�I;/I;"I;TI;u�H;��H;��H;��H;��H;��H;��H;��H;t�H;VI;"I;/I;�I;�I;/ I;��H;�NH;�F;mkB;3�9;5*;��;��:8Q�9P������?��T[�;���J����5��{��A��T9ݽZl���,���M�5�l����p��      6m־Q�Ѿ�>ľ����ԗ����{��I�+�����V���{�?�/�&���,��;=�7�һH�@��� �<�k:)�:b;��3;Cj?;}2E;��G;�H;GI;� I;�I;�I;5	I;I;��H;�H;��H;��H;m�H;��H;��H;�H;��H;I;4	I;�I;�I;� I;DI;|�H;��G;y2E;Bj?;��3;b;'�:<�k:�� �J�@�8�һ;=��,��&��?�/��{��V�����+��I���{�ԗ�������>ľQ�Ѿ      E\�î�s5��z ��E۾ֳ�^��|�Z�M?#����A����j�&��Dϼ ����������lۺ�:�9�4�:f�;r�,;��;;H�C;�G;`�H;�I;�!I;�I;RI;;I;�I;UI;2�H;�H;��H;7�H;��H;�H;0�H;QI;�I;;I;RI;�I;�!I;�I;]�H;�G;F�C;��;;r�,;i�;�4�:�:�9�lۺ������� ��Dϼ&����j��A�����N?#�|�Z�^��ֳ��E۾�z �s5�î�      G�b��>]���M�Ŏ6�®�%���>ľ%q��|�Z�+�T9ݽ"W����L����!F�� �G���׻�;�n��Ȋ:�i;,P$;�7;z�A; JF;DCH;��H;� I;}I;�I;-I;AI;�I;-�H;��H;��H;%�H;��H;��H;,�H;�I;@I;-I;�I;zI;� I;��H;BCH;#JF;w�A;�7;,P$;�i;�Ȋ:n��;� �׻ �G�!F�������L�"W��T9ݽ+�|�Z�%q���>ľ%��®�Ŏ6���M��>]�      p��򲗿���:�y�}�R���)�ov��>ľ^���I�Zl����������&�ԮҼ�}�*B���������L�!:!+�:Jz;�3;mj?;�\E;��G;��H;�I;�I;�I;�I;�I;�I;1 I;��H;w�H;��H;w�H;��H;. I;�I;�I;�I;�I;�I;�I;��H;��G;�\E;jj?;�3;Jz;'+�:H�!:��������+B��}�ԮҼ��&��������Zl��I�^���>ľov���)�}�R�:�y����򲗿      �˿�<ƿsL��B1����>]���)�%��ֳ���{���,�t��)��S`I��J���,���3/��+���� �0069�4�:��;p.;3.=;vaD;��G;{�H;�I;T!I;oI;bI;�	I;�I; I;��H;'�H;w�H;(�H;��H; I;�I;�	I;bI;kI;N!I;�I;z�H;��G;vaD;..=;p.;��;�4�:0069�� ��+���3/��,���J��S`I�)��t�齧�,���{�ֳ�%����)��>]��B1��sL���<ƿ      ����>���V[忸˿�T���}�R�®��E۾ԗ����M���	������j��3�d����O�/�׻��/����n��:� 
;*;m;;kC;�'G;��H;I;"I;I;�I;�
I;�I;�I;\�H;��H;�H;��H;Z�H;�I;�I;�
I;�I;I;"I;I;��H;�'G;kC;j;;*;� 
;t��:�����/�/�׻��O�d���3���j������	���M�ԗ���E۾®�}�R���T���˿V[�>���      O�7��v����˿B1��:�y�Ŏ6��z �����5�l�+��ͽ$�����&���˼<�k������X�$� ����:[�;#&;�9;��B;!�F;�}H;�	I;x"I;DI;�I;�I;�I;]I;��H;9�H;��H;9�H;��H;]I;�I;�I;�I;AI;u"I;�	I;�}H;!�F;��B;�9;$&;[�;���:(� ���X����<�k���˼��&�$����ͽ+�5�l������z �Ŏ6�:�y�B1���˿���v�7��      ��*��g&��#�v�V[�sL�������M�s5��>ľ����,��D�뒐��5�2�ݼ���q
���x�Htk��b:ml�:#;ڗ7;��A;��F;�dH;�I;m"I;I;}I;VI;	I;�I;7 I;��H;��H;��H;7 I;�I;I;TI;}I;I;i"I;�I;�dH;��F;��A;֗7;#;ml�:�b:Htk���x��q
���2�ݼ�5�뒐��DὭ�,����>ľs5���M����sL��V[�v��#��g&�      ��8��4��g&�7��>����<ƿ򲗿�>]�î�Q�Ѿ�p���*7����'W��MR?� }�o8�������b�����G:� �:�!;$�6;-lA;�YF;�TH;�H;/"I;�I;I;�I;]I;I;y I;��H;)�H;��H;z I;I;\I;�I;I;�I;,"I;�H;�TH;�YF;-lA;!�6;�!;� �:��G:d��������o8�� }�MR?�'W�����*7��p��Q�Ѿî��>]�򲗿�<ƿ>���7���g&��4�      �Aq���i���U�H:�@�����>���w���}A�e5�� ���^Z�����A���]�����d��E",��5��B�Ѻ���9��:i�;lY4;}�@;�VF;��H;�GI;�bI;AOI;R:I;*I;TI;�I; I;�I;�I;�I; I;�I;RI;*I;R:I;@OI;�bI;�GI;��H;�VF;}�@;jY4;l�;��:���9F�Ѻ�5��E",��d������]��A������^Z�� ��e5�}A�w���>�������@�H:���U���i�      ��i���b�\�O�.5�2i�������������q<���� f��c
V�HE	�!���IY�j9�B�����(��R����Ⱥ��:���:*�;S�4;w�@;vhF;͗H;CII;�bI;�NI;�9I;�)I;I;�I;�I;�I;�I;�I;�I;�I;I;�)I;�9I;�NI;�bI;CII;͗H;vhF;w�@;O�4;0�;���:��:��Ⱥ�R����(�B���j9��IY�!��HE	�c
V� f������q<������������2i�.5�\�O���b�      ��U�\�O�J-?�/�'���O�ῶ欿d�{�ga/���뾟���I����e���ZN�]5������6H�T ������ܫ":��:��;��5;�`A;�F;h�H;IMI;+bI;�MI;�8I;)I;wI;I;uI;;I;=I;;I;tI;I;vI;)I;�8I;�MI;(bI;KMI;i�H;�F;�`A;��5;��;��:ܫ": ���T ��6H�����]5���ZN�e������I�������ga/�d�{��欿O����/�'�J-?�\�O�      H:�.5�/�'��������lȿ���n$_���Y�Ҿݕ���6�����*���`=�<�漬)��BG�6��H����Q:�:0";#�7;�&B;�F;��H;SI;�`I;�KI;U7I;�'I;pI;OI;�I;�I;�
I;�I;�I;PI;pI;�'I;U7I;�KI;�`I;SI;��H;�F;�&B;�7;!0";�:��Q:J��6��BG��)��<���`=��*������6�ݕ��Y�Ҿ��n$_����lȿ�������/�'�.5�      @�2i�������K�ѿl������q<��:��a����q����Wн轅���'�Tb̼�zl��.��-�X�|��"�:��;�&;�9;\C;�MG;�H;kYI;�^I;�HI;5I;&I;I;>I;�I;�
I;�	I;�
I;�I;>I;I;&I;5I;�HI;�^I;kYI;�H;�MG;ZC;�9;�&;��;(�:���-�X��.���zl�Tb̼��'�轅��Wн����q��a���:��q<���l���K�ѿ������2i�      �������O��lȿl���������O���~]׾|����I�����A��@�d�n�|֮�RH��jλ/�$�@%����:nN;ц+;<;14D;�G;�I;�^I;�[I;EI;X2I;�#I;vI;�I;�I;�	I;�I;�	I;�I;�I;vI;�#I;X2I;EI;�[I;�^I;�I;�G;04D;<;҆+;nN;���:`%�-�$��jλRH�|֮�n�@�d��A������I�|���~]׾����O�����l���lȿO�Ῥ��      >��������欿�������O��x����� ���l���"��ܽ���`=����t���k"�R���ۺh��9�?�:�L;��0;؟>;�ME;�#H;&I;bI;:WI;�@I;)/I;v!I;qI;8I;DI;�I;�I;�I;DI;:I;qI;w!I;)/I;�@I;7WI;bI;�%I;�#H;�ME;ԟ>;��0;�L;�?�:P��9�ۺR���k"�t������`=����ܽ��"��l�� ����뾂x���O�������欿����      w�������c�{�n$_��q<������~��	w���6�����!���h����᷾�~ d�o.��w^e�`H[���Z:���:�, ;��5;�A;WF;ڄH;AI;�bI;�QI; <I;u+I;�I;BI;nI;�	I;I;dI;I;�	I;nI;@I;�I;u+I; <I;�QI;�bI;AI;ڄH;WF;�A;��5;�, ;���:��Z:\H[�v^e�p.��~ d�᷾�����h�!�������6�	w��~��������q<�n$_�c�{�����      }A��q<�ga/����:�~]׾� ��	w��>�EE	�����۽����3�`�꼘���",��W��=���Q�఩:�M
;�f);�:;S@C;*@G;��H;wTI;�_I;_KI;7I;�'I;�I;�I;rI;I;�I;�I;�I;I;sI;�I;�I;�'I;7I;\KI;�_I;vTI;��H;'@G;P@C;�:;�f);�M
;ް�:@Q�:���W��",�����`�꼙�3�۽������EE	�>�	w��� ��~]׾�:���ga/��q<�      e5�������Y�Ҿ�a��|����l��6�EE	���Ƚk���aG����c֮��W����I�k����Xd,:���:&�;Ǔ1;y�>;lE;]�G;SI;Z_I;yZI;oDI;�1I;g#I;yI;.I;9
I;AI;I;UI;I;CI;:
I;-I;yI;e#I;�1I;lDI;yZI;X_I;UI;[�G;iE;w�>;Ǔ1;&�;���:Xd,:���J�k�����W�c֮�����aG�k����ȽEE	��6��l�|����a��Y�Ҿ������      � �� f�����ݕ����q��I���"���������k���ZN�[� ¼L�y��$��Q��c� � �W��:P0;V�&;x8;� B;��F;�H;�@I;*bI;�RI;Q=I;H,I;I;I;�I;I;oI;QI;�I;QI;oI;I;�I;I;I;H,I;N=I;�RI;)bI;�@I;�H;��F;� B;x8;U�&;N0;�: �W�f� ��Q���$�L�y� ¼[��ZN�k������������"��I���q�ݕ����� f��      �^Z�b
V��I��6�������ܽ!��۽���aG�[�	�ȼ�)��w�(�X��+G5���4�Z:r�:DS;<'1;�=;ݠD;a�G;%�H;�XI;N^I;�II;.6I;�&I;�I;�I;�
I;�I;�I;� I;��H;� I;�I;�I;�
I;�I;�I;�&I;,6I;�II;N^I;�XI;$�H;^�G;ڠD;�=;<'1;BS;r�:@�Z:��+G5�X��w�(��)��	�ȼ[��aG�۽��!���ܽ������6��I�c
V�      ���HE	��������Wн�A�����h���3���� ¼�)��,x/��һP�X�*#���9���:�>;if);�`9;�&B;�F;�}H;7I;�aI;�UI;�@I;/I;2!I;I;]I;I;�I;� I;��H;3�H;��H;� I;�I;I;_I;�I;4!I;/I;�@I;�UI;�aI;7I;�}H;�F;�&B;�`9;hf);�>;���:�9(#��P�X��һ,x/��)�� ¼�����3��h��󑽣A���Wн��콻��HE	�      �A��!��e���*��轅�?�d��`=����_��c֮�K�y�w�(��һ|]e�����жf9 ��:^�;v1";R�4;�m?;E;��G;��H;�WI;�^I;AKI;�7I;,(I;�I;_I;�
I;ZI;TI;��H;�H;u�H;�H;��H;TI;ZI;�
I;_I;�I;*(I;�7I;AKI;�^I;�WI;��H;��G;E;�m?;R�4;v1";a�;���:жf9����z]e��һw�(�K�y�c֮�_�꼘���`=�?�d�轅��*��e��!��      �]��IY��ZN��`=���'�n����᷾������W��$�Y��R�X������9���:���:��;ָ0;�<;��C;XG;3�H;�?I;caI;	UI;u@I;I/I;�!I;�I;HI;�I;�I;�H;��H;D�H;��H;D�H;��H;�H;�I;�I;HI;�I;�!I;I/I;u@I;UI;baI;�?I;-�H;XG;��C;�<;ո0;��;���:���:�9����R�X�Z���$��W�����᷾����n���'��`=��ZN��IY�      ���i9�[5��;��Tb̼|֮�s�� d�",�����Q��+G5�.#��жf9���:��:=�;��-;��:;LB;pVF;LKH;I;]I;Z\I;�HI;?6I;W'I;SI;�I;R
I;yI;4 I;��H;��H;��H;$�H;��H;��H;��H;3 I;zI;R
I;�I;PI;Y'I;=6I;�HI;Z\I;]I;I;NKH;mVF;LB;��:;��-;;�;��:���:��f9.#��+G5��Q�����",�~ d�s��|֮�Tb̼;��[5��j9�      �d��@��������)���zl�RH��k"�n.���W��H�k�c� ����9���:���:9�;�-;��9;xaA;�E;]�G;��H;:SI;N`I;!PI;�<I;�,I;�I;lI;II;�I;�I;��H;��H;�H;��H;��H;��H;�H;��H;��H;�I;�I;GI;iI;�I;�,I;�<I;"PI;I`I;6SI;��H;[�G;�E;waA;��9;�-;9�;���:���: �9��d� �I�k��W��n.���k"�RH��zl��)������B���      F",���(�5H�AG��.���jλR��x^e�:����� �W�4�Z:���:\�;��;��-;��9;�A;dE;Y�G;��H;�GI;-aI;�UI;zBI;�1I;%$I;I;&I;�I;-I;��H;��H;�H;D�H;N�H; �H;O�H;D�H;�H;��H;��H;-I;�I;#I;I;#$I;�1I;{BI;�UI;+aI;�GI;��H;Z�G;dE;�A;��9;��-;��;^�;���:,�Z: �W����;��z^e�R���jλ�.��AG�5H���(�      �5���R��P ��6��1�X�)�$��ۺpH[�@Q�Xd,:�:t�:�>;v1";ָ0;��:;waA;dE;,�G;��H;�=I;f`I;�YI;)GI;6I;�'I;'I;�I;4I;�I; I;>�H;Z�H;0�H;��H;��H;y�H;��H;��H;0�H;X�H;?�H; I;�I;3I;�I;%I;�'I;6I;%GI;�YI;f`I;�=I;��H;,�G;dE;taA;��:;ظ0;v1";�>;p�:�:Xd,: Q�lH[��ۺ%�$�,�X�6��P ���R��      @�Ѻx�Ⱥ����J������%�H��9��Z:ܰ�:���:N0;@S;df);K�4;�<;LB;�E;V�G;��H;�:I;�_I;�[I;ZJI;=9I;�*I;�I;/I;;I;�I;JI;$�H;��H;K�H;h�H;3�H;m�H;"�H;n�H;4�H;i�H;K�H;��H;$�H;GI;�I;;I;.I;�I;�*I;<9I;WJI;�[I;�_I;�:I;��H;W�G;�E;LB;�<;K�4;df);@S;N0;���:ذ�:��Z:P��9@%�\��L��������Ⱥ      ��9�:�":p�Q:�:���:�?�:���:�M
;&�;U�&;9'1;�`9;�m?;��C;lVF;^�G;��H;�=I;�_I;J\I;�KI;O;I;	-I;!I;,I;�I;"I;�I;�H;q�H;��H;s�H;��H;��H;�H;��H;�H;��H;��H;q�H;��H;q�H;�H;�I;#I;�I;-I;!I;-I;O;I;�KI;H\I;�_I;�=I;��H;Z�G;lVF;��C;�m?;�`9;7'1;R�&;&�;�M
;���:�?�:���:�:p�Q:�":��:      $��:���:��:��:��;vN;�L;�, ;�f);Ǔ1;x8;�=;�&B;E;XG;KKH;��H;�GI;f`I;�[I;�KI;�;I;'.I;k"I;rI;PI;W	I;�I;��H;(�H;�H;��H;��H;X�H;{�H;��H;��H;��H;{�H;X�H;��H;��H;�H;#�H;��H;�I;T	I;SI;sI;g"I;%.I;�;I;�KI;�[I;f`I;�GI;��H;HKH;XG;E;�&B;�=;x8;Ɠ1;�f);�, ;�L;vN;��;��:��:���:      o�;,�;��;0";
�&;҆+;��0;��5;�:;y�>;� B;�D;�F;��G;1�H;I;8SI;/aI;�YI;\JI;O;I;).I;�"I;;I;�I;9
I;iI;��H;��H;��H;��H;��H;6�H;�H;-�H;��H;��H;��H;.�H;�H;5�H;��H;��H;��H;��H;��H;gI;<
I;�I;8I;�"I;+.I;K;I;]JI;�YI;0aI;7SI;I;1�H;��G;�F;ߠD;� B;w�>;�:;��5;��0;ӆ+;�&;0";��; �;      �Y4;^�4;��5;�7;�9;<;ܟ>;�A;S@C;lE;��F;c�G;�}H;��H;�?I;]I;N`I;�UI;'GI;;9I;-I;j"I;;I;^I;�
I;�I;) I;%�H;��H;%�H;��H;2�H;��H;��H; �H;��H;��H;��H;�H;��H;��H;2�H;��H;"�H;��H;%�H;' I;�I;�
I;[I;9I;k"I;-I;;9I;'GI;�UI;K`I;]I;�?I;��H;�}H;a�G;��F;iE;S@C;�A;ܟ>;<;�9;"�7;��5;P�4;      ��@;~�@;�`A;�&B;\C;14D;�ME;WF;)@G;X�G;�H;(�H;7I;�WI;eaI;\\I;(PI;{BI;!6I;�*I;!I;vI;I;�
I;*I;Z I;o�H;!�H;_�H;�H;?�H;��H;��H;��H;�H;��H;��H;��H;�H;��H;��H;��H;?�H;�H;\�H;!�H;l�H;Z I;+I;�
I;�I;vI;!I;�*I;!6I;~BI;%PI;Z\I;eaI;�WI;7I;'�H;�H;X�G;)@G;WF;�ME;34D;\C;�&B;�`A;~�@;      �VF;�hF;֛F;�F;�MG;�G;�#H;քH;��H;SI;�@I;�XI;�aI;�^I;	UI;�HI;�<I;�1I;�'I;�I;*I;PI;6
I;�I;S I;��H;T�H;��H;*�H;7�H;��H;��H;|�H;��H;@�H;��H;��H;��H;B�H;��H;z�H;��H;��H;6�H;)�H;��H;Q�H;��H;T I;�I;6
I;PI;&I;�I;�'I;�1I;�<I;�HI;	UI;�^I;�aI;�XI;�@I;RI;��H;ׄH;�#H;�G;�MG;�F;כF;xhF;      ��H;̗H;b�H;��H;�H;�I;&I;AI;zTI;Z_I;*bI;S^I;�UI;AKI;v@I;?6I;�,I;#$I;)I;2I;�I;W	I;hI;* I;h�H;U�H;��H;O�H;g�H;��H;h�H;K�H;x�H;��H;u�H;�H;�H;�H;s�H;��H;s�H;K�H;h�H;��H;f�H;O�H;��H;U�H;k�H;) I;gI;W	I;�I;2I;)I;#$I;�,I;=6I;v@I;AKI;�UI;Q^I;*bI;X_I;{TI;AI;&I;�I;�H;��H;b�H;͗H;      �GI;DII;LMI;SI;lYI;�^I;
bI;�bI;`I;|ZI;�RI;�II;�@I;�7I;K/I;W'I;�I;I;�I;=I;#I;�I;��H;&�H;�H;��H;M�H;D�H;��H;h�H;A�H;G�H;��H;�H;��H;|�H;t�H;|�H;��H;�H;��H;G�H;@�H;e�H;��H;D�H;L�H;��H;�H;&�H;��H;�I; I;=I;�I; I;�I;W'I;K/I;�7I;�@I;�II;�RI;}ZI;`I;�bI;
bI;�^I;yYI;SI;OMI;OII;      cI;�bI;&bI;�`I;�^I;�[I;=WI;�QI;`KI;oDI;Q=I;36I;/I;,(I;�!I;SI;pI;%I;7I;�I;�I;��H;��H;��H;X�H;,�H;d�H;��H;\�H;=�H;5�H;w�H;��H;g�H;
�H;��H;��H;��H;
�H;g�H;��H;y�H;5�H;<�H;Z�H;��H;f�H;,�H;[�H;��H;��H;��H;�I;�I;7I;&I;lI;SI;�!I;,(I;/I;26I;P=I;oDI;`KI;�QI;=WI;�[I;�^I;�`I;&bI;�bI;      KOI;�NI;�MI;�KI;�HI;EI;�@I;%<I;7I;�1I;P,I;�&I;9!I;�I;�I;�I;NI;�I;�I;MI;�H;&�H;��H;$�H;�H;5�H;��H;e�H;<�H;=�H;g�H;��H;3�H;��H;�H;]�H;Y�H;_�H;�H;��H;0�H;��H;g�H;<�H;:�H;g�H;��H;5�H;�H;$�H;��H;&�H;�H;MI;�I;�I;JI;�I;�I;�I;9!I;�&I;P,I;�1I;7I;)<I;�@I;EI;�HI;�KI;�MI;�NI;      V:I;�9I;�8I;a7I;(5I;V2I;2/I;}+I;�'I;m#I;I;�I;�I;fI;MI;[
I;�I;0I; I;*�H;x�H;�H;��H;��H;9�H;��H;e�H;A�H;2�H;h�H;��H;,�H;��H;N�H;�H;��H;��H;��H;�H;N�H;��H;-�H;��H;g�H;4�H;A�H;d�H;��H;:�H;��H;��H;�H;u�H;+�H; I;0I;�I;Y
I;NI;dI;�I;�I;I;o#I;�'I;+I;2/I;X2I;&5I;a7I;�8I;�9I;      *I;�)I;)I;�'I;&I;�#I;x!I;�I;�I;|I;#I;�I;bI;�
I;�I;�I;�I;��H;E�H;��H;��H;��H;��H;6�H;��H;��H;J�H;G�H;u�H;��H;*�H;��H;,�H;��H;��H;��H;v�H;��H;��H;��H;)�H;��H;,�H;��H;v�H;G�H;J�H;��H;��H;6�H;��H;��H;��H;��H;E�H;��H;�I;�I;�I;�
I;`I;�I;!I;zI;�I;�I;x!I;�#I;&I;�'I;)I;�)I;      VI;,I;I;}I;#I;vI;rI;GI;�I;0I;�I;�
I;I;_I;�I;: I;��H;��H;_�H;P�H;z�H;��H;6�H;��H;��H;|�H;w�H;��H;��H;6�H;��H;/�H;��H;��H;J�H;@�H;M�H;@�H;J�H;��H;��H;0�H;��H;7�H;��H;��H;t�H;{�H;��H;��H;5�H;��H;x�H;R�H;_�H;��H;��H;: I;�I;_I;I;�
I;�I;0I;�I;II;rI;wI;I;}I;~I;%I;      �I;�I;I;XI;HI;�I;<I;xI;yI;<
I;I;�I;�I;[I;!�H;�H;��H;�H;6�H;p�H;��H;[�H;�H;��H;��H;��H;��H;�H;e�H;��H;K�H;��H;��H;Z�H; �H;�H;��H;�H; �H;Z�H;��H;��H;K�H;��H;h�H;�H;��H;��H;��H;��H;�H;[�H;��H;p�H;6�H;�H;��H;�H;!�H;[I;�I;�I;I;<
I;yI;zI;<I;�I;=I;XI;I;�I;      �I;�I;I;�I;�I;�I;II;�	I;I;FI;wI;�I;� I;��H;��H;��H;�H;D�H;��H;;�H;��H;�H;.�H;�H;�H;@�H;p�H;��H;
�H;�H;�H;��H;J�H;!�H;�H;��H;��H;��H;�H; �H;G�H;��H;�H;��H;�H;��H;o�H;@�H;�H;�H;-�H;�H;��H;;�H;��H;D�H;�H;��H;��H;��H;� I;�I;vI;GI;I;�	I;II;�I;�I;�I;I;�I;      �I;�I;EI;�I;�
I;�	I;�I;*I;�I;
I;[I;� I;��H;�H;I�H;��H;��H;M�H;��H;u�H;�H;��H;��H;��H;��H;��H;�H;|�H;��H;\�H;��H;��H;?�H;	�H;��H;��H;��H;��H;��H;�H;=�H;��H;��H;]�H;��H;|�H;�H;��H;��H;��H;��H;��H;�H;u�H;��H;N�H;��H;��H;I�H;�H;��H;� I;XI;I;�I;*I;�I;�	I;�
I;�I;CI;�I;      �I;�I;KI;�
I;�	I;�I;�I;kI;�I;UI;�I;��H;9�H;}�H;��H;-�H;��H;�H;}�H;)�H;��H;��H;��H;��H;��H;��H;�H;v�H;��H;\�H;��H;z�H;M�H;��H;��H;��H;��H;��H;��H;��H;J�H;{�H;��H;_�H;��H;v�H;�H;��H;��H;��H;��H;��H;��H;)�H;}�H;�H;��H;-�H;��H;}�H;9�H;��H;�I;WI;�I;jI;�I;�I;�	I;�
I;KI;�I;      �I;�I;EI;�I;�
I;�	I;�I;*I;�I;
I;[I;� I;��H;�H;I�H;��H;��H;M�H;��H;u�H;�H;��H;��H;��H;��H;��H;�H;|�H;��H;\�H;��H;��H;?�H;	�H;��H;��H;��H;��H;��H;�H;=�H;��H;��H;_�H;��H;|�H;�H;��H;��H;��H;��H;��H;�H;u�H;��H;N�H;��H;��H;I�H;�H;��H;� I;YI;I;�I;*I;�I;�	I;�
I;�I;AI;�I;      �I;�I;I;�I;�I;�I;II;�	I;I;GI;vI;�I;� I;��H;��H;��H;�H;D�H;��H;;�H;��H;�H;.�H;�H;�H;@�H;r�H;��H;�H;�H;�H;��H;J�H; �H;�H;��H;��H;��H;�H;!�H;G�H;��H;�H;��H;�H;��H;o�H;@�H;�H;�H;-�H;�H;��H;;�H;��H;D�H;�H;��H;��H;��H;� I;�I;vI;GI;I;�	I;II;�I;�I;�I;}I;�I;      �I;�I;I;XI;HI;�I;<I;xI;wI;<
I;I;�I;�I;[I;!�H;�H;��H;�H;6�H;p�H;��H;[�H;�H;��H;��H;��H;��H;�H;e�H;��H;K�H;��H;��H;Z�H; �H;�H;��H;�H; �H;Z�H;��H;��H;K�H;��H;h�H;�H;��H;��H;��H;��H;�H;[�H;��H;p�H;6�H;�H;��H;�H;!�H;[I;�I;�I;I;<
I;zI;xI;<I;�I;=I;XI;I;�I;      YI;.I;�I;~I;"I;tI;qI;FI;�I;.I;�I;�
I;I;_I;�I;: I;��H;��H;_�H;P�H;{�H;��H;7�H;��H;��H;|�H;w�H;��H;��H;6�H;��H;/�H;��H;��H;J�H;@�H;M�H;@�H;J�H;��H;��H;2�H;��H;7�H;��H;��H;s�H;{�H;��H;��H;5�H;��H;w�H;R�H;_�H;��H;��H;: I;�I;_I;I;�
I;�I;1I;�I;FI;rI;wI;I;~I;~I;+I;      *I;�)I;!)I;�'I;&I;�#I;z!I;�I;�I;zI;!I;�I;`I;�
I;�I;�I;�I;��H;E�H;��H;��H;��H;��H;6�H;��H;��H;J�H;G�H;v�H;��H;,�H;��H;,�H;��H;��H;��H;v�H;��H;��H;��H;)�H;��H;*�H;��H;v�H;G�H;H�H;��H;��H;6�H;��H;��H;��H;��H;E�H;��H;�I;�I;�I;�
I;bI;�I;#I;}I;�I;�I;{!I;�#I;&I;�'I; )I;�)I;      V:I;�9I;�8I;a7I;'5I;V2I;2/I;}+I;�'I;n#I;I;�I;�I;fI;NI;[
I;�I;/I; I;*�H;z�H;�H;��H;��H;:�H;��H;d�H;A�H;2�H;h�H;��H;-�H;��H;N�H;�H;��H;��H;��H;�H;N�H;��H;-�H;��H;g�H;4�H;A�H;d�H;��H;9�H;��H;��H;�H;t�H;+�H; I;0I;�I;[
I;NI;fI;�I;�I;I;n#I;�'I;}+I;2/I;X2I;&5I;a7I;�8I;�9I;      AOI;�NI;�MI;�KI;�HI;EI;�@I;&<I;!7I;�1I;P,I;�&I;9!I;�I;�I;�I;LI;�I;�I;NI;�H;&�H;��H;$�H;�H;6�H;��H;g�H;=�H;=�H;g�H;��H;2�H;��H;�H;]�H;Y�H;_�H;�H;��H;2�H;��H;g�H;<�H;<�H;e�H;��H;5�H;�H;$�H;��H;&�H;�H;MI;�I;�I;LI;�I;�I;�I;8!I;�&I;P,I;�1I;!7I;'<I;�@I;EI;�HI;�KI;�MI;�NI;       cI;�bI;,bI;�`I;�^I;�[I;>WI;�QI;`KI;oDI;S=I;36I;/I;,(I;�!I;SI;oI;%I;7I;�I;�I;��H;��H;��H;[�H;,�H;c�H;��H;\�H;=�H;5�H;v�H;��H;g�H;	�H;��H;��H;��H;
�H;g�H;��H;y�H;5�H;<�H;Z�H;��H;d�H;,�H;X�H;��H;��H;��H;�I;�I;7I;&I;mI;UI;�!I;-(I;/I;36I;Q=I;nDI;`KI;�QI;>WI;�[I;�^I;�`I;,bI;�bI;      �GI;CII;OMI;SI;lYI;�^I;
bI;�bI;`I;}ZI;�RI;�II;�@I;�7I;K/I;W'I;�I;�I;�I;=I;&I;�I;��H;&�H;�H;��H;L�H;D�H;��H;g�H;@�H;G�H;��H;�H;��H;|�H;t�H;|�H;��H;�H;��H;I�H;A�H;e�H;��H;D�H;L�H;��H;�H;'�H;��H;�I;I;=I;�I;I;�I;Y'I;K/I;�7I;�@I;�II;�RI;|ZI;`I;�bI;
bI;�^I;vYI;SI;MMI;RII;      ��H;ʗH;g�H;��H;�H;�I;&I;AI;zTI;Z_I;*bI;Q^I;�UI;AKI;v@I;?6I;�,I;#$I;)I;4I;�I;W	I;hI;* I;k�H;U�H;��H;O�H;g�H;��H;h�H;K�H;v�H;��H;s�H;�H;�H;�H;u�H;��H;w�H;M�H;h�H;��H;f�H;O�H;��H;W�H;h�H;* I;gI;W	I;�I;2I;)I;%$I;�,I;=6I;v@I;BKI;�UI;S^I;+bI;Z_I;yTI;AI;&I;�I;�H;��H;d�H;×H;      �VF;hF;��F;�F;�MG;�G;�#H;ׄH;��H;SI;�@I;�XI;�aI;�^I;UI;�HI;�<I;�1I;�'I;�I;,I;PI;6
I;�I;T I;��H;S�H;��H;,�H;7�H;��H;��H;{�H;��H;@�H;��H;��H;��H;B�H;��H;z�H;��H;��H;5�H;)�H;��H;Q�H;��H;S I;�I;7
I;PI;&I;�I;�'I;�1I;�<I;�HI;	UI;�^I;�aI;�XI;�@I;QI;��H;քH;�#H;�G;�MG;�F;�F;uhF;      ��@;�@;�`A;�&B;\C;14D;�ME;WF;*@G;Z�G;�H;'�H;7I;�WI;eaI;\\I;'PI;{BI;!6I;�*I;!I;vI; I;�
I;+I;Z I;n�H;!�H;_�H;�H;?�H;��H;��H;��H;�H;��H;��H;��H;�H;��H;��H;��H;?�H;�H;\�H;!�H;l�H;Z I;*I;�
I; I;vI;!I;�*I;!6I;~BI;%PI;\\I;eaI;�WI;7I;(�H;�H;W�G;)@G;WF;�ME;14D;ZC;�&B;�`A;�@;      �Y4;^�4;��5;�7;ܫ9;<;ڟ>;�A;U@C;lE;��F;c�G;�}H;��H;�?I;]I;N`I;�UI;'GI;;9I;	-I;k"I;;I;^I;�
I;�I;) I;%�H;��H;%�H;��H;2�H;��H;��H;��H;��H;��H;��H;�H;��H;��H;3�H;��H;"�H;��H;%�H;' I;�I;�
I;\I;9I;j"I;-I;;9I;'GI;�UI;L`I;]I;�?I;��H;�}H;c�G;��F;kE;U@C;�A;ڟ>;<;�9;�7;��5;R�4;      k�;8�;��;0";�&;ֆ+;Ĺ0;��5;�:;y�>;� B;ߠD;�F;��G;1�H;I;8SI;-aI;�YI;\JI;P;I;+.I;�"I;;I;�I;:
I;iI;��H;��H;��H;��H;��H;6�H;�H;.�H;��H;��H;��H;-�H;�H;5�H;��H;��H;��H;��H;��H;gI;<
I;�I;9I;�"I;).I;K;I;]JI;�YI;0aI;8SI;I;3�H;��G;�F;ߠD;� B;v�>;�:;��5;Ĺ0;؆+;�&;0";��;(�;      $��:���:��:��:��;vN;�L;�, ;�f);Ɠ1;x8;�=;�&B;E;UG;JKH;��H;�GI;f`I;�[I;�KI;�;I;(.I;k"I;sI;QI;U	I;�I;��H;(�H;�H;��H;��H;X�H;{�H;��H;��H;��H;{�H;X�H;��H;��H;�H;#�H;��H;�I;S	I;SI;rI;i"I;$.I;�;I;�KI;�[I;f`I;�GI;��H;KKH;YG;E;�&B;�=;x8;Ǔ1;�f);�, ;�L;vN;��;��:��:���:      ���9غ:��":t�Q:�:���:�?�:���:�M
;$�;S�&;7'1;�`9;�m?;��C;lVF;[�G;��H;�=I;�_I;J\I;�KI;P;I;-I;!I;-I;�I;#I;�I;�H;q�H;��H;s�H;��H;��H;�H;��H;�H;��H;��H;s�H;��H;q�H;�H;�I;#I;�I;,I;!I;-I;N;I;�KI;H\I;�_I;�=I;��H;[�G;lVF;��C;�m?;�`9;9'1;V�&;#�;�M
;���:�?�:���:�:t�Q:�":��:      F�Ѻr�Ⱥ򈮺L��x��p%�P��9��Z:ܰ�:���:P0;>S;df);K�4;�<;LB;�E;V�G;��H;�:I;�_I;�[I;ZJI;@9I;�*I;�I;/I;;I;�I;JI;$�H;��H;L�H;i�H;4�H;n�H;"�H;n�H;3�H;h�H;I�H;��H;$�H;FI;�I;;I;-I;�I;�*I;99I;WJI;�[I;�_I;�:I;��H;W�G;�E;LB;�<;L�4;df);>S;N0;���:ܰ�:��Z:P��9p%�h��L��������Ⱥ      �5���R��P ��6��3�X�*�$��ۺpH[� Q�Xd,:�:p�:�>;v1";ָ0;��:;waA;dE;,�G;��H;�=I;f`I;�YI;)GI;6I;�'I;'I;�I;6I;�I; I;>�H;Z�H;0�H;��H;��H;y�H;��H;��H;0�H;X�H;?�H; I;�I;2I;�I;%I;�'I;6I;%GI;�YI;f`I;�=I;��H;,�G;dE;vaA;��:;ظ0;v1";�>;t�:�:Xd,:� Q�pH[��ۺ%�$�-�X�6��P ���R��      F",���(�5H�AG��.���jλR��{^e�;����� �W�(�Z:���:\�;��;��-;��9;�A;dE;Y�G;��H;�GI;/aI;�UI;{BI;�1I;%$I;I;'I;�I;-I;��H;��H;�H;D�H;N�H; �H;N�H;D�H;�H;��H;��H;-I;�I;#I;I;"$I;�1I;zBI;�UI;+aI;�GI;��H;Z�G;dE;�A;��9;��-;��;\�;���:4�Z: �W����;��~^e�R���jλ�.��AG�5H���(�      �d��A��������)���zl�RH��k"�n.���W��I�k�c� ��� �9���:���:9�;�-;��9;waA;�E;]�G;��H;;SI;N`I;"PI;�<I;�,I;�I;mI;II;�I;�I;��H;��H;�H;��H;��H;��H;�H;��H;��H;�I;�I;GI;iI;�I;�,I;�<I;!PI;I`I;4SI;��H;[�G;�E;xaA;��9;�-;9�;���:���:�9��c� �I�k��W��o.���k"�RH��zl��)������B���      ���i9�[5��;��Tb̼|֮�s�� d�",�����Q��+G5�.#����f9���:��:=�;��-;��:;LB;pVF;NKH;I;]I;Z\I;�HI;@6I;Y'I;UI;�I;R
I;yI;4 I;��H;��H;��H;$�H;��H;��H;��H;3 I;zI;R
I;�I;OI;W'I;=6I;�HI;Z\I;]I;I;LKH;mVF;LB;��:;��-;<�;��:���:жf9.#��+G5��Q�����",� d�s��|֮�Tb̼;��[5��j9�      �]��IY��ZN��`=���'�n����᷾������W��$�Z��R�X������9���:���:��;ո0;�<;��C;XG;3�H;�?I;baI;
UI;v@I;I/I;�!I;�I;HI;�I;�I;�H;��H;D�H;��H;D�H;��H;�H;�I;�I;HI;�I;�!I;I/I;u@I;
UI;caI;�?I;-�H;XG;��C;�<;ָ0;��;���:���:�9����R�X�Y���$��W�����᷾����n���'��`=��ZN��IY�      �A��!��e���*��轅�?�d��`=����_��c֮�K�y�x�(��һ|]e�����жf9 ��:_�;v1";Q�4;�m?;E;��G;��H;�WI;�^I;AKI;�7I;-(I;�I;_I;�
I;[I;UI;��H;�H;u�H;�H;��H;SI;XI;�
I;_I;�I;*(I;�7I;?KI;�^I;�WI;��H;��G;E;�m?;Q�4;v1";a�;���:жf9����z]e��һw�(�K�y�c֮�_�꼘���`=�?�d�轅��*��e��!��      ���HE	��������Wн�A�����h���3���� ¼�)��,x/��һP�X�*#���9���:�>;hf);�`9;�&B;�F;�}H;7I;�aI;�UI;�@I;/I;4!I;�I;]I;I;�I;� I;��H;3�H;��H;� I;�I;I;]I;I;2!I;/I;�@I;�UI;�aI;7I;�}H;�F;�&B;�`9;hf);�>;���:�9*#��P�X��һ,x/��)�� ¼�����3��h��󑽣A���Wн��콻��HE	�      �^Z�b
V��I��6�������ܽ!��۽���aG�[�	�ȼ�)��x�(�X��+G5���8�Z:r�:BS;9'1;�=;ݠD;a�G;$�H;�XI;N^I;�II;/6I;�&I;�I;�I;�
I;�I;�I;� I;��H;� I;�I;�I;�
I;�I;�I;�&I;,6I;�II;M^I;�XI;%�H;]�G;ڠD;�=;<'1;BS;r�:@�Z:��,G5�X��w�(��)��	�ȼ[��aG�۽��!���ܽ������6��I�c
V�      � �� f�����ݕ����q��I���"���������k���ZN�[� ¼L�y��$��Q��c� � �W��:P0;S�&;x8;� B;��F;�H;�@I;*bI;�RI;Q=I;H,I;I;I;�I;I;oI;QI;�I;QI;oI;I;�I;I;I;H,I;N=I;�RI;)bI;�@I;�H;��F;� B;x8;U�&;N0;�: �W�d� ��Q���$�L�y� ¼[��ZN�k������������"��I���q�ݕ����� f��      e5�������Y�Ҿ�a��|����l��6�EE	���Ƚk���aG����c֮��W����I�k����Xd,:���:$�;Ǔ1;y�>;lE;[�G;UI;Z_I;yZI;oDI;�1I;e#I;yI;.I;:
I;AI;I;UI;I;AI;9
I;-I;wI;g#I;�1I;lDI;yZI;X_I;SI;]�G;iE;w�>;Ǔ1;&�;���:Xd,:���I�k�����W�c֮�����aG�k����ȽEE	��6��l�|����a��Y�Ҿ������      }A��q<�ga/����:�~]׾� ��	w��>�EE	�����۽����3�`�꼘���",��W��;���Q�఩:�M
;�f);�:;S@C;'@G;��H;yTI;�_I;_KI;7I;�'I;�I;�I;sI;I;�I;�I;�I;I;rI;�I;�I;�'I;7I;\KI;�_I;vTI;��H;*@G;P@C;�:;�f);�M
;ް�:�Q�;���W��",�����`�꼙�3�۽������EE	�>�	w��� ��~]׾�:���ga/��q<�      w�������c�{�n$_��q<������~��	w���6�����!���h����᷾�~ d�n.��v^e�\H[���Z:���:�, ;��5;�A;WF;ۄH;AI;�bI;�QI; <I;u+I;�I;BI;pI;�	I;I;dI;!I;�	I;pI;@I;�I;u+I; <I;�QI;�bI;AI;لH;WF;�A;��5;�, ;���:��Z:hH[�t^e�p.��~ d�᷾�����h�!�������6�	w��~��������q<�n$_�c�{�����      >��������欿�������O��x����� ���l���"��ܽ���`=����t���k"�R���ۺ`��9�?�:�L;��0;؟>;�ME;�#H;&I;bI;<WI;�@I;)/I;v!I;rI;;I;DI;�I;�I;�I;DI;8I;oI;v!I;)/I;�@I;9WI;bI;�%I;�#H;�ME;՟>;��0;�L;�?�:P��9�ۺR���k"�t������`=����ܽ��"��l�� ����뾂x���O�������欿����      �������O��lȿl���������O���~]׾|����I�����A��@�d�n�|֮�RH��jλ-�$�`%����:nN;ц+;<;04D;�G;�I;�^I;�[I;EI;X2I;�#I;wI;�I;�I;�	I;�I;�	I;�I;�I;tI;�#I;X2I;EI;�[I;�^I;�I;�G;14D;<;ц+;nN;���:`%�/�$��jλRH�|֮�n�@�d��A������I�|���~]׾����O�����l���lȿO�Ῥ��      @�2i�������K�ѿl������q<��:��a����q����Wн轅���'�Tb̼�zl��.��-�X����"�:��;�&;�9;ZC;�MG;�H;kYI;�^I;�HI;5I;&I;I;>I;�I;�
I;�	I;�
I;�I;>I;I;&I;5I;�HI;�^I;kYI;�H;�MG;\C;�9;�&;��;$�:���-�X��.���zl�Tb̼��'�轅��Wн����q��a���:��q<���l���K�ѿ������2i�      H:�.5�/�'��������lȿ���n$_���Y�Ҿݕ���6�����*���`=�<�漬)��BG�6��H����Q:�:0";#�7;�&B;�F;��H;SI;�`I;�KI;U7I;�'I;rI;PI;�I;�I;�
I;�I;�I;OI;oI;�'I;U7I;�KI;�`I;SI;��H;�F;�&B;�7;0";�:��Q:J��6��BG��)��<���`=��*������6�ݕ��Y�Ҿ��n$_����lȿ�������/�'�.5�      ��U�\�O�J-?�/�'���O�῵欿d�{�ga/���뾟���I����e���ZN�]5������6H�T �� ���ث":��:��;��5;�`A;�F;i�H;KMI;+bI;�MI;�8I;)I;wI;I;uI;;I;=I;;I;uI;I;vI;)I;�8I;�MI;(bI;IMI;h�H;�F;�`A;��5;��;��:ܫ": ���T ��6H�����]5���ZN�e������I�������ga/�d�{��欿O����/�'�J-?�\�O�      ��i���b�\�O�.5�2i�������������q<���� f��b
V�HE	�!���IY�j9�B�����(��R����Ⱥ��:���:*�;S�4;w�@;vhF;͗H;CII;�bI;�NI;�9I;�)I;I;�I;�I;�I;�I;�I;�I;�I;I;�)I;�9I;�NI;�bI;CII;̗H;vhF;w�@;P�4;0�;���:��:��Ⱥ�R����(�B���j9��IY�!��HE	�b
V� f������q<������������2i�.5�\�O���b�      ᶕ�T���Ҭ��0�_���7�|�!}߿����,b��V�/l¾Kx�e.���Ž��t�)��c����?�N������x9���:��;��2;g@@;�fF;R�H;��I;��I;G|I;\I;�CI;<2I;�%I;�I;�I;eI;�I;�I;�%I;:2I;�CI;\I;F|I;��I;��I;R�H;�fF;g@@;��2;��;���:��x9��N����?�c��)����t���Že.�Kx�/l¾�V��,b����!}߿|���7�0�_�Ҭ��T���      T���E���%}��+Y��3�����$ڿ&��ƽ\����(���s��3�7����p�c�R���<<�*��@��� ��9���:�;d%3;|p@;zF;��H;/�I;(�I;�{I;�[I;�CI;�1I;�%I;ZI;�I;9I;�I;[I;�%I;�1I;�CI;�[I;�{I;%�I;/�I;��H;zF;|p@;a%3;�;���: ��9D���*���<<�R��c��p�7����3��s�(�����ƽ\�&���$ڿ����3��+Y�%}�F���      Ҭ��%}�?tf��lG�آ%��p�0�ʿ\����>M����V�����d�ʤ�̷�0�d��
��I����1�V������x��9���:_;�U4;��@;!�F;R�H;�I;�I;�yI;�YI;wBI;	1I;�$I;�I;I;�I;I;�I;�$I;1I;uBI;�YI;�yI;�I;�I;R�H;!�F;��@;�U4;b;���:x��9���V�����1��I���
�0�d�̷�ʤ���d�V�������>M�\���0�ʿ�p�آ%��lG�?tf�%}�      0�_��+Y��lG�!f.�|���꿳���O䂿��5���󾏰��P�N�W��S��"�Q����z����h!�xg����	:�
�:/�;v16;��A;�G;#I;j�I;��I;�vI;�WI;�@I;�/I;�#I;�I;@I;�I;@I;�I;�#I;�/I;�@I;�WI;�vI;��I;k�I;#I;�G;��A;r16;2�;�
�:�	:�xg���h!�z������"�Q�S��W��P�N���������5�O䂿�������|�!f.��lG��+Y�      ��7��3�آ%�|��<����ſ
���Ľ\�=����Ͼ����b�3��载z��}�9�^�἗���z�x7}��ct���^:�+�:ߣ#;ȍ8;��B;RsG;�%I;�I;$�I;5rI;HTI;>I;�-I;G"I;�I;I;�I;I;�I;G"I;�-I;>I;HTI;2rI;$�I;�I;�%I;RsG;��B;č8;�#;�+�:��^:�ct�w7}��z����^��~�9��z����b�3�������Ͼ=��Ľ\�
�����ſ�<��|�آ%��3�      |�����p������ſ&���Ps���1�4r���d���d�~I�ЈŽ��}�_*�JC���^��B�X�D�xE�� �:��;�);@7;;_D;w�G;~HI;�I;ߏI;�lI;&PI;;I;K+I;P I;�I;�I;aI;�I;�I;Q I;K+I;;I;&PI;�lI;ۏI;�I;|HI;v�G;^D;<7;;�);��;� �:�E�X�D��B��^�JC��_*���}�ЈŽ~I��d��d��4r����1��Ps�&����ſ��꿄p����      !}߿�$ڿ0�ʿ����
����Ps�SX:����'l¾�ǆ���7����95���Q�����t���75�\��w�� "�8)ʼ:��;��.;��=;�EE;�YH;�hI;X�I;��I;VfI;PKI;\7I;w(I;I;%I;�I;�I;�I;%I;I;w(I;]7I;PKI;UfI;�I;X�I;�hI;�YH;�EE;��=;��.;��;-ʼ:�!�8w��Z���75��t������Q�95�������7��ǆ�'l¾���SX:��Ps�
�������0�ʿ�$ڿ      ���&��\���O䂿Ľ\���1�����J˾Ꝓ�F�N�z��J������W�'�c�Ҽ��|��z��n���w����&:�P�:ڨ;�W4;��@;[gF;��H;A�I;R�I;j�I;L_I;FI;=3I;U%I;{I;�I;I;�I;I;�I;{I;T%I;=3I;FI;L_I;g�I;R�I;A�I;��H;ZgF;��@;�W4;ڨ;�P�:|�&:�w���n���z���|�c�ҼW�'����J���z��F�N�Ꝓ��J˾�����1�Ľ\�O䂿\���&��      �,b�ƽ\��>M���5�=��4r��'l¾Ꝓ�%&W��3�:Sؽ�z��[G����zI����?���̻i�-�X	��t��:��;��&;V|9;�C;�dG;�I;r�I;��I;�vI;�WI;`@I;�.I;�!I;�I;�I;
I;�I;	I;�I;�I;�!I;�.I;`@I;�WI;�vI;��I;q�I;�I;�dG;�C;V|9;��&;��;r��:X	��h�-���̻��?�zI�����[G��z��:Sؽ�3�%&W�Ꝓ�'l¾4r��=����5��>M�ƽ\�      �V������������Ͼ�d���ǆ�F�N��3��c�[����\�3��)C���o���	��눻����9v��:�h;�/;n�=;sE;/3H;�WI;�I;/�I;�kI;�OI;Y:I;*I;UI;�I;'I;�I;�I;�I;&I;�I;TI; *I;Y:I;�OI;�kI;/�I;�I;�WI;,3H;pE;n�=;�/;�h;r��:���9��눻��	��o�(C��3����\�[���cི3�F�N��ǆ��d����Ͼ���������      /l¾(��V������������d���7�z��:Sؽ[���d�D*�ckּ*\����'����R� }����:�Z;�#;j=7;`�A;G�F;��H;��I;�I;�I;!aI;�GI;'4I;Z%I;�I;�I;�I;
I;�	I;
I;�I;�I;�I;\%I;'4I;�GI;aI;�I;�I;��I;��H;C�F;]�A;j=7; �#;�Z;��:}���R�����'�*\��ckּD*��d�[��:Sؽz����7��d���������V���(��      Kx��s���d�P�N�b�3�~I����J����z����\�C*��ݼF���*<<���ڻ�V��ct���&:���:sC;�</;�D=;�D;��G;)9I; �I;ڔI;HtI;bVI;�?I;�-I;� I;�I;�I;�
I;,I;HI;,I;�
I;�I;�I;� I;�-I;�?I;bVI;JtI;ڔI; �I;'9I;��G;�D;�D=;�</;rC;���:��&:�ct��V���ڻ*<<�F����ݼC*���\��z��J������~I�b�3�P�N���d��s�      e.��3�ʤ�W����ЈŽ95�����[G�3��bkּF����xC��>�F6}�̬����x9���:8	;e�&;�;8;��A;՟F;�H;kyI;ƝI;*�I;ffI;�KI;�7I;�'I;�I;�I;�I;HI;�I;�I;�I;HI;�I;�I;�I;�'I;�7I;�KI;gfI;*�I;ɝI;iyI;�H;џF;��A;�;8;d�&;8	;���:p�x9ʬ��F6}��>��xC�F���bkּ3��[G����95��ЈŽ��W��ʤ��3�      ��Ž7���̷�S���z����}��Q�W�'����(C��*\��*<<��>�un�� �຀����:���:?�;�'3;��>;�E;�H;�<I;�I;ٕI;�vI;YI;�AI;�/I;�!I;I;%I;�	I;�I;WI;�I;WI;�I;�	I;%I;I;�!I;�/I;�AI;YI;�vI;ەI;�I;�<I;�H;�E;��>;�'3;?�;���:���:�����tn���>�*<<�*\��(C�����W�'��Q���}��z��S��̷�7���      ��t��p�/�d�"�Q�~�9�_*����d�ҼzI���o���'���ڻF6}� ��7� �:�m�:��;�.;L<;�oC;r7G;��H;�I;�I;�I;TfI;vLI;.8I;(I;I;�I;�I;~I;�I; I;� I; I;�I;�I;�I;�I;I;(I;-8I;wLI;RfI;�I;�I;�I;��H;r7G;�oC;M<;�.;��;�m�: �:07� ��G6}���ڻ��'��o�zI��d�Ҽ���_*�~�9�"�Q�/�d��p�      )��b��
����]��IC���t����|���?���	����V�Ь�� �
�:�: i;K�+;$�9;��A;�fF;��H;�_I;��I;͑I;9sI;�VI;�@I;/I;$!I;�I;AI;I;�I;� I;��H;?�H;��H;� I;�I;I;CI;�I;#!I;/I;�@I;�VI;<sI;ΑI;��I;�_I;��H;�fF;��A;$�9;K�+;�h;�:
�: �Ь���V�����	���?���|��t��IC��^������
�c�      b��P���I��y�������^��75��z���̻�눻�R��ct�p�x9���:�m�:�h;��*;�8;�@;�E;l(H;�8I;��I;M�I;�~I;�`I;�HI;�5I;�&I;�I;mI;2
I;�I;� I;(�H;��H;�H;��H;(�H;� I;�I;2
I;mI;�I;�&I;�5I;�HI;�`I;�~I;I�I;�I;�8I;k(H;�E;�@;
�8;��*;�h;�m�:���:`�x9�ct��R��눻��̻�z��75��^����y����I��R��      ��?��<<���1��h!��z��B�Z���n��h�-��}����&:���:��:��;G�+;�8;l�@;"^E;��G;{I; �I;��I;k�I;�iI;rPI;A<I;�+I;�I;�I;�I;cI;�I;�H;��H;��H;�H;��H;��H;�H;�I;cI;�I;�I;�I;�+I;?<I;sPI;�iI;g�I;��I; �I;xI;��G;"^E;m�@;�8;G�+;��;���:���:��&:}��
�h�-��n��Z���B黲z��h!���1��<<�      N��)��P���wg��{7}�Q�D�s��x��0	�����9��:���:8	;@�;�.;#�9;�@;"^E;��G;uI;�I;<�I;��I;�pI;�VI;�AI;�0I;�"I;�I;%I;)I;�I;��H;��H;��H;��H;�H;��H;��H;��H;��H;�I;)I;"I;�I;�"I;�0I;�AI;�VI;�pI;��I;>�I;�I;vI;��G;$^E;�@;"�9;�.;@�;8	;���:��:���90	�� x��s��M�D�w7}�wg��P���)��      ����������ct��E��!�8l�&:r��:v��:�Z;pC;b�&;�'3;I<;��A;�E;��G;sI;�|I;��I;ِI;�uI;�[I;DFI;�4I;g&I;�I;�I;
I;,I;q�H;��H;o�H;��H;��H;V�H;��H;��H;m�H;��H;q�H;,I;
I;�I;�I;d&I;�4I;FFI;�[I;�uI;ِI;��I;�|I;sI;��G;�E;��A;H<;�'3;a�&;oC;�Z;p��:n��:x�&:�!�8xE๘ct�����,���      P�x9���9���9�	:t�^:� �:/ʼ:�P�:��;�h;�#;�</;�;8;��>;�oC;�fF;n(H;{I;�I;��I;�I;5xI;�^I;sII;�7I;D)I;DI;�I;�I;�I;� I;��H;��H;q�H;��H;��H;��H;��H;��H;r�H;��H;��H;� I;�I;�I;�I;DI;F)I;�7I;oII;�^I;5xI;�I;��I;�I;|I;k(H;�fF;�oC;��>;�;8;�</; �#;�h;��;�P�:-ʼ:� �:x�^:�	:���9��9      ���:���:���:�
�:�+�:��;��;ި;��&;��/;n=7;�D=;��A;�E;r7G;��H;�8I; �I;<�I;ِI;4xI;�_I;KI;�9I;2+I;9I;sI;vI;�I;xI;<�H;��H;U�H;v�H;�H;H�H;"�H;H�H;�H;w�H;S�H;��H;<�H;tI;�I;vI;pI;:I;3+I;�9I;KI;�_I;1xI;ڐI;<�I;"�I;�8I;��H;s7G;�E;��A;�D=;l=7;�/;��&;�;��;��;�+�:�
�:���:���:      ��;�;_;(�;֣#;�);��.;�W4;Z|9;o�=;`�A;�D;՟F;�H;��H;�_I;��I;��I;��I;�uI;�^I;KI;_:I;Z,I;u I;�I;�I;�I;]I;��H;?�H;n�H;D�H;��H;��H;��H;��H;��H;��H;��H;C�H;n�H;?�H;��H;[I;�I;�I;�I;v I;W,I;]:I;KI;�^I;�uI;��I;��I;��I;�_I;��H;�H;ԟF;�D;a�A;n�=;X|9;�W4;��.;�);ߣ#;(�;a;	�;      ˼2;p%3;�U4;t16;Ǎ8;>7;;��=;��@;�C;sE;G�F;��G;�H;�<I;�I;��I;M�I;l�I;�pI;�[I;pII;�9I;X,I;� I;YI;]I;�I;I;��H;��H;��H;e�H;y�H;�H;&�H;��H;<�H;��H;'�H;�H;v�H;f�H;��H;��H;��H;I;�I;\I;ZI;� I;W,I;�9I;mII;�[I;�pI;o�I;L�I;��I;�I;�<I;�H;��G;F�F;pE;�C;��@;��=;@7;;ύ8;v16;�U4;e%3;      p@@;�p@;��@;��A;��B;aD;�EE;WgF;�dG;+3H;��H;,9I;kyI;�I;�I;ёI;�~I;�iI;�VI;JFI;�7I;6+I;z I;^I;�I;�I;{I;��H;�H;��H;[�H;\�H;��H;��H;��H;Y�H;7�H;Y�H;��H;��H;��H;]�H;[�H;��H;�H;��H;yI;�I;�I;\I;z I;6+I;�7I;KFI;�VI;�iI;�~I;БI;�I;�I;hyI;)9I;��H;+3H;�dG;WgF;�EE;bD;��B;��A;��@;�p@;      �fF;zF;�F;�G;RsG;o�G;�YH;��H;�I;�WI;��I;�I;ƝI;ڕI;�I;9sI;�`I;pPI;�AI;�4I;B)I;7I;�I;ZI;�I;�I;)�H;>�H;�H;��H;n�H;��H;Q�H;h�H;��H;H�H;N�H;H�H;��H;h�H;O�H;��H;m�H;��H;�H;=�H;(�H;�I;�I;ZI;�I;9I;=)I;�4I;�AI;sPI;�`I;8sI;�I;ڕI;ƝI;�I;��I;�WI;�I;��H;�YH;o�G;VsG;�G;�F;zF;      \�H;��H;N�H;%I;�%I;HI;�hI;=�I;q�I;�I;�I;ޔI;*�I;�vI;UfI;�VI;�HI;?<I;�0I;g&I;GI;tI;�I;�I;vI;,�H;D�H;&�H;��H;q�H;��H;0�H;!�H;F�H;��H;M�H;M�H;M�H;��H;F�H;�H;0�H;��H;o�H;��H;&�H;@�H;*�H;yI;�I;�I;tI;CI;g&I;�0I;A<I;�HI;�VI;UfI;�vI;*�I;ݔI;�I;�I;r�I;?�I;�hI;|HI;�%I;%I;N�H;��H;      ��I;4�I;�I;h�I;�I;�I;Y�I;W�I;��I;/�I;�I;OtI;ifI;YI;yLI;�@I;�5I;�+I;�"I;�I;�I;wI;�I;
I;��H;@�H;%�H;��H;��H;��H;%�H;��H;��H;<�H;��H;|�H;b�H;|�H;��H;<�H;��H;��H;#�H;��H;��H;��H;%�H;@�H;��H;
I;�I;wI;�I;�I;�"I;�+I;�5I;�@I;yLI;YI;dfI;MtI;�I;/�I;��I;Y�I;Y�I;�I;�I;g�I;�I;>�I;      ��I;&�I;�I;��I;!�I;ۏI;��I;i�I;�vI;�kI; aI;gVI;�KI;�AI;18I;/I;�&I;�I;�I;�I;�I;�I;]I;��H;�H;�H;��H;��H;��H;�H;��H;��H;��H;a�H;�H;��H;��H;��H;�H;a�H;��H;��H;��H;�H;��H;��H;��H;�H;�H;��H;\I;�I;�I;�I;�I;�I;�&I;/I;18I;�AI;�KI;dVI;aI;�kI;�vI;j�I;�I;ۏI;(�I;��I;�I;�I;      Q|I;�{I;�yI;�vI;CrI;�lI;[fI;O_I;�WI;�OI;�GI;�?I;�7I;�/I;(I;'!I;�I;�I;#I; 
I;�I;wI;��H;��H;��H;��H;o�H;��H;�H;��H;��H;��H;;�H;��H;H�H;�H;�H;�H;H�H;��H;7�H;��H;��H;��H;�H;��H;n�H;��H;��H;��H;��H;wI;�I; 
I;#I;�I;�I;'!I;(I;�/I;�7I;�?I;�GI;�OI;�WI;R_I;[fI;�lI;?rI;�vI;�yI;�{I;      \I;�[I;�YI;�WI;TTI;#PI;WKI;FI;h@I;]:I;.4I;�-I;�'I;�!I;I;�I;wI;�I;.I;3I;� I;=�H;@�H;��H;X�H;o�H;��H;%�H;��H;��H;��H;�H;��H;�H;��H;��H;��H;��H;��H;�H;��H;�H;��H;��H;��H;%�H;��H;n�H;Z�H;��H;=�H;=�H;� I;3I;-I;�I;vI;�I;I;�!I;�'I;�-I;.4I;_:I;h@I;FI;VKI;%PI;QTI;�WI;�YI;�[I;      �CI;�CI;{BI;�@I;>I; ;I;]7I;B3I;�.I; *I;^%I;� I;�I;I;�I;JI;=
I;fI;�I;{�H;��H;��H;q�H;i�H;Z�H;��H;0�H;��H;��H;��H;�H;��H;��H;��H;Q�H;�H;�H;�H;Q�H;��H;��H;��H;�H;��H;��H;��H;0�H;��H;]�H;i�H;o�H;��H;��H;{�H;�I;fI;<
I;JI;�I;I;�I;� I;^%I; *I;�.I;B3I;\7I;;I;>I;�@I;|BI;�CI;      ?2I;�1I;1I;�/I;�-I;H+I;v(I;W%I;�!I;TI;�I;�I;I;*I;�I;I;�I;�I;��H;�H;��H;V�H;G�H;}�H;��H;S�H;!�H;�H;��H;<�H;��H;��H;m�H;)�H;��H;��H;��H;��H;��H;(�H;j�H;��H;��H;>�H;��H;�H;�H;Q�H;��H;}�H;F�H;V�H;��H;�H;��H;�I;�I;I;�I;)I; I;�I;�I;UI;�!I;X%I;v(I;K+I;�-I;�/I;1I;�1I;      �%I;�%I;�$I;�#I;Q"I;I I;I;�I;�I;�I;�I;�I;�I;�	I;�I;�I;� I;�H;��H;v�H;|�H;z�H;��H;�H;��H;g�H;D�H;9�H;`�H;��H;�H;��H;"�H;��H;��H;z�H;_�H;z�H;��H;��H;!�H;��H;�H;��H;b�H;;�H;C�H;g�H;��H;�H;��H;z�H;y�H;v�H;��H;�H;� I;�I;�I;�	I;�I;�I;�I;�I;�I;�I;I;M I;F"I;�#I;�$I;�%I;      �I;mI;�I;�I;�I;�I;(I;�I;�I;)I;�I;�
I;MI;�I;�I;� I;2�H;��H;��H;��H;��H;�H;��H;(�H;��H;��H;��H;��H;�H;H�H;��H;R�H;��H;��H;P�H;D�H;M�H;D�H;P�H;��H;��H;U�H;��H;I�H;�H;��H;��H;��H;��H;*�H;��H;�H;��H;��H;��H;��H;0�H;� I;�I;�I;OI;�
I;�I;*I;�I;�I;(I;�I;�I;�I;�I;eI;      �I;�I;I;EI;+I;�I;�I; I;I;�I;�
I;8I;�I;cI;I;��H;��H;��H;��H;��H;��H;K�H;��H;��H;U�H;F�H;M�H;|�H;��H;�H;��H; �H;��H;}�H;D�H;+�H;&�H;+�H;C�H;z�H;��H;"�H;��H;�H;��H;|�H;J�H;D�H;V�H;��H;��H;K�H;��H;��H;��H;��H;��H;��H;I;`I;�I;8I;�
I;�I;I; I;�I;�I;!I;DI;I;�I;      cI;BI;�I;�I;�I;^I;�I;�I;�I;�I;�	I;SI;�I;�I;� I;F�H;#�H;�H;�H;_�H;��H;&�H;��H;>�H;3�H;J�H;J�H;g�H;��H;�H;��H;�H;��H;c�H;L�H;'�H;�H;'�H;L�H;e�H;��H;�H;��H;�H;��H;g�H;G�H;K�H;3�H;;�H;��H;&�H;��H;_�H;�H;�H;"�H;F�H;� I;�I;�I;SI;�	I;�I;�I;�I;�I;cI;�I;�I;�I;:I;      �I;�I;I;DI;+I;�I;�I; I;I;�I;�
I;8I;�I;aI;I;��H;��H;��H;��H;��H;��H;K�H;��H;��H;V�H;F�H;M�H;|�H;��H;�H;��H; �H;��H;}�H;C�H;+�H;&�H;+�H;D�H;z�H;��H;"�H;��H;�H;��H;|�H;J�H;D�H;U�H;��H;��H;K�H;��H;��H;��H;��H;��H;��H;I;aI;�I;8I;�
I;�I;I; I;�I;�I; I;EI;I;�I;      �I;mI;�I;�I;�I;�I;(I;�I;�I;)I;�I;�
I;OI;�I;�I;� I;2�H;��H;��H;��H;��H;�H;��H;+�H;��H;��H;��H;��H;�H;H�H;��H;R�H;��H;��H;P�H;D�H;M�H;D�H;P�H;��H;��H;V�H;��H;I�H;�H;��H;��H;��H;��H;&�H;��H;�H;��H;��H;��H;��H;0�H;� I;�I;�I;MI;�
I;�I;*I;�I;�I;(I;�I;�I;�I;�I;eI;      �%I;�%I;�$I;�#I;O"I;I I;I;�I;�I;�I;�I;�I;�I;�	I;�I;�I;� I;�H;��H;t�H;�H;z�H;��H;�H;��H;h�H;C�H;;�H;`�H;��H;�H;��H;"�H;��H;��H;z�H;_�H;z�H;��H;��H;!�H;��H;�H;��H;b�H;9�H;C�H;g�H;��H;�H;��H;z�H;y�H;w�H;��H;�H;� I;�I;�I;�	I;�I;�I;�I;�I;�I;�I;I;M I;F"I;�#I;�$I;�%I;      A2I;�1I;1I;�/I;�-I;G+I;u(I;U%I;�!I;TI;�I;�I; I;)I;�I;I;�I;�I;��H;�H;��H;V�H;G�H;}�H;��H;S�H;!�H;�H;��H;<�H;��H;��H;k�H;'�H;��H;��H;��H;��H;��H;(�H;j�H;��H;��H;>�H;��H;�H;�H;Q�H;��H;|�H;F�H;V�H;��H;�H;��H;�I;�I;I;�I;*I; I;�I;�I;UI;�!I;U%I;v(I;I+I;�-I;�/I;1I;�1I;      �CI;�CI;BI;�@I;>I;�:I;^7I;A3I;�.I; *I;^%I;� I;�I;I;�I;JI;=
I;fI;�I;|�H;��H;��H;q�H;i�H;]�H;��H;0�H;��H;��H;��H;�H;��H;��H;��H;Q�H;�H;�H;�H;Q�H;��H;��H;��H;�H;��H;��H;��H;0�H;��H;Z�H;i�H;o�H;��H;��H;{�H;�I;gI;<
I;JI;�I;I;�I;� I;^%I;!*I;�.I;A3I;^7I;;I;>I;�@I;BI;�CI;      \I;�[I;�YI;�WI;TTI;#PI;VKI;FI;h@I;]:I;.4I;�-I;�'I;�!I;I;�I;vI;�I;-I;3I;� I;=�H;@�H;��H;Z�H;o�H;��H;%�H;��H;��H;��H;�H;��H;�H;��H;��H;��H;��H;��H;�H;��H;
�H;��H;��H;��H;%�H;��H;n�H;X�H;��H;=�H;=�H;� I;3I;.I;�I;vI;�I;I;�!I;�'I;�-I;-4I;_:I;g@I;FI;WKI;%PI;QTI;�WI;�YI;�[I;      G|I;�{I;�yI;�vI;>rI;�lI;[fI;O_I;�WI;�OI;�GI;�?I;�7I;�/I;(I;'!I;�I;�I;#I;!
I;�I;wI;��H;��H;��H;��H;o�H;��H;�H;��H;��H;��H;8�H;��H;H�H;�H;�H;�H;H�H;��H;:�H;��H;��H;��H;�H;��H;n�H;��H;��H;��H;��H;wI;�I;!
I;#I;�I;�I;(!I;(I;�/I;�7I;�?I;�GI;�OI;�WI;P_I;[fI;�lI;?rI;�vI;�yI;�{I;      ��I;"�I;�I;��I;'�I;׏I;�I;j�I;�vI;�kI; aI;fVI;�KI;�AI;18I;/I;�&I;�I;�I;�I;�I;�I;]I;��H;�H;�H;��H;��H;��H;�H;��H;��H;��H;a�H;�H;��H;��H;��H;�H;a�H;��H;��H;��H;�H;��H;��H;��H;�H;�H;��H;\I;�I;�I;�I;�I;�I;�&I;/I;18I;�AI;�KI;gVI; aI;�kI;�vI;k�I;�I;ڏI;#�I;��I;�I;"�I;      ��I;2�I;�I;g�I;��I;�I;Y�I;X�I;��I;/�I;�I;MtI;dfI;YI;yLI;�@I;�5I;�+I;�"I;�I;�I;wI;�I;
I;��H;@�H;%�H;��H;��H;��H;#�H;��H;��H;;�H;��H;|�H;b�H;|�H;��H;<�H;��H;��H;%�H;��H;��H;��H;%�H;@�H;��H;
I;�I;wI;�I;�I;�"I;�+I;�5I;�@I;yLI;YI;ifI;OtI;�I;/�I;��I;Y�I;Y�I;ޝI;�I;h�I;�I;@�I;      W�H;��H;P�H;!I;�%I;{HI;�hI;=�I;r�I;�I; �I;ݔI;*�I;�vI;UfI;�VI;�HI;?<I;�0I;i&I;JI;tI;�I;�I;yI;,�H;B�H;&�H;��H;q�H;��H;0�H;�H;F�H;��H;M�H;M�H;L�H;��H;D�H;�H;1�H;��H;o�H;��H;&�H;@�H;,�H;vI;�I;�I;tI;CI;i&I;�0I;A<I;�HI;�VI;UfI;�vI;*�I;ޔI; �I;�I;q�I;=�I;�hI;{HI;�%I;!I;O�H;��H;      �fF;zF;�F;�G;TsG;p�G;�YH;��H;�I;�WI;��I;�I;ƝI;ڕI;�I;9sI;�`I;rPI;�AI;�4I;D)I;9I;�I;ZI;�I;�I;)�H;=�H;�H;��H;m�H;��H;P�H;h�H;��H;H�H;N�H;H�H;��H;h�H;O�H;��H;n�H;��H;�H;>�H;(�H;�I;�I;ZI;�I;7I;=)I;�4I;�AI;rPI;�`I;9sI;�I;ەI;ȝI;�I;��I;�WI;�I;��H;ZH;p�G;VsG;�G;�F;zF;      p@@;�p@;��@;��A;��B;aD;�EE;WgF;�dG;,3H;��H;)9I;hyI;�I;�I;ёI;�~I;�iI;�VI;KFI;�7I;6+I;| I;^I;�I;�I;{I;��H;�H;��H;[�H;\�H;��H;��H;��H;Y�H;7�H;Y�H;��H;��H;��H;^�H;[�H;��H;�H;��H;yI;�I;�I;]I;y I;6+I;�7I;KFI;�VI;�iI;�~I;ёI;�I;
�I;kyI;,9I;��H;)3H;�dG;WgF;�EE;aD;��B;��A;��@;�p@;      μ2;p%3;�U4;r16;��8;C7;;��=;��@; C;sE;F�F;��G;�H;�<I;�I;��I;M�I;l�I;�pI;�[I;qII;�9I;X,I;� I;ZI;\I;�I;I;��H;��H;��H;e�H;x�H;�H;$�H;��H;<�H;��H;'�H;�H;x�H;f�H;��H;��H;��H;I;�I;]I;YI;� I;W,I;�9I;lII;�[I;�pI;o�I;L�I;��I;�I;�<I;�H;��G;F�F;qE;�C;��@;��=;C7;;ύ8;r16;�U4;d%3;      ��;!�;p;)�;գ#;�);��.;�W4;Z|9;o�=;`�A;�D;ҟF;�H;��H;�_I;��I;��I;��I;�uI;�^I;KI;_:I;Z,I;v I;�I;�I;�I;]I;��H;?�H;n�H;D�H;��H;��H;��H;��H;��H;��H;��H;C�H;n�H;?�H;��H;[I;�I;�I;�I;u I;W,I;]:I;KI;�^I;�uI;��I;��I;��I;�_I;��H;�H;ԟF;�D;a�A;l�=;X|9;�W4;��.;�);ڣ#;)�;f;�;      ���:���:���:�
�:�+�:��;��;ި;��&;�/;n=7;�D=;��A;�E;r7G;��H;�8I; �I;<�I;ِI;5xI;�_I;KI;�9I;3+I;9I;qI;vI;�I;xI;<�H;��H;U�H;w�H;�H;H�H;"�H;H�H;�H;v�H;S�H;��H;<�H;tI;�I;vI;oI;:I;2+I;�9I;KI;�_I;1xI;ڐI;<�I;"�I;�8I;��H;s7G;�E;��A;�D=;l=7;��/;��&;�;��;��;�+�:�
�:���:���:      ��x9p��9ȭ�9�	:t�^:� �:1ʼ:�P�:��;�h;�#;�</;�;8;��>;�oC;�fF;l(H;{I;�I;��I;�I;5xI;�^I;sII;�7I;F)I;DI;�I;�I;�I;� I;��H;��H;q�H;��H;��H;��H;��H;��H;q�H;��H;��H;� I;�I;�I;�I;CI;F)I;�7I;oII;�^I;5xI;�I;��I;�I;|I;l(H;�fF;�oC;��>;�;8;�</;�#;�h;��;�P�:5ʼ:� �:��^:�	:ȭ�9��9      ��������񳺰ct��E��!�8p�&:r��:r��:�Z;oC;a�&;�'3;H<;��A;�E;��G;sI;�|I;��I;ِI;�uI;�[I;FFI;�4I;g&I;�I;�I;
I;,I;o�H;��H;m�H;��H;��H;V�H;��H;��H;o�H;��H;r�H;,I;
I;�I;�I;d&I;�4I;DFI;�[I;�uI;ِI;��I;�|I;sI;��G;�E;��A;I<;�'3;b�&;oC;�Z;p��:r��:x�&:�!�8xE๠ct�����0���      N��)��P���wg��|7}�S�D�s��x��8	�����9��:���:8	;@�;�.;"�9;�@;"^E;��G;uI;�I;>�I;��I;�pI;�VI;�AI;�0I;�"I;�I;%I;)I;�I;��H;��H;��H;��H;�H;��H;��H;��H;��H;�I;)I;"I;�I;�"I;�0I;�AI;�VI;�pI;��I;<�I;�I;vI;��G;$^E;�@;#�9;�.;@�;8	;���:��:���90	��x��s��M�D�w7}�wg��P���)��      ��?��<<���1��h!��z��B�Z���n��h�-�
�}����&:���:��:��;G�+;�8;l�@;"^E;��G;{I; �I;��I;k�I;�iI;rPI;A<I;�+I;�I;�I;�I;bI;�I;�H;��H;��H;�H;��H;��H;�H;�I;dI;�I;�I;�I;�+I;><I;sPI;�iI;g�I;��I; �I;wI;��G;"^E;m�@;�8;G�+;��;��:���:��&:}���h�-��n��Z���B黲z��h!���1��<<�      b��P���I��z�������^��75��z���̻�눻�R��ct�`�x9���:�m�:�h;��*;�8;�@;�E;l(H;�8I;��I;M�I;�~I;�`I;�HI;�5I;�&I;�I;mI;2
I;�I;� I;(�H;��H;�H;��H;(�H;� I;�I;3
I;mI;�I;�&I;�5I;�HI;�`I;�~I;I�I;�I;�8I;k(H;�E;�@;
�8;��*;�h;�m�:���:p�x9�ct��R��눻��̻�z��75��^����z����I��Q��      )��b��
����]��IC���t����|���?���	����V�Ь�� ��:�: i;J�+;$�9;��A;�fF;��H;�_I;��I;ΑI;<sI;�VI;�@I;/I;#!I;�I;AI;I;�I;� I;��H;?�H;��H;� I;�I;I;CI;�I;$!I;/I;�@I;�VI;;sI;͑I;��I;�_I;��H;�fF;��A;$�9;L�+;�h;�:�: �Ь���V�����	���?���|��t��IC��]������
�c�      ��t��p�/�d�"�Q�~�9�_*����d�ҼzI���o���'���ڻG6}� ��@7� �:�m�:��;�.;L<;�oC;r7G;��H;�I;�I;�I;TfI;wLI;18I;(I;I;�I;�I;�I;�I; I;� I; I;�I;I;�I;�I;I;(I;,8I;vLI;RfI;�I;�I;�I;��H;r7G;�oC;M<;�.;��;�m�: �:7� ��F6}���ڻ��'��o�zI��d�Ҽ���_*�~�9�!�Q�/�d��p�      ��Ž7���̷�S���z����}��Q�W�'����(C��*\��*<<��>�un����຀����:���:?�;�'3;��>;�E;�H;�<I;�I;ەI;�vI;YI;�AI;�/I;�!I;I;&I;�	I;�I;WI;�I;WI;�I;�	I;#I;I;�!I;�/I;�AI;YI;�vI;ڕI;�I;�<I;�H;�E;��>;�'3;?�;���:���:�� ��un���>�*<<�*\��(C�����W�'��Q���}��z��S��̷�7���      e.��3�ʤ�W����ЈŽ95�����[G�3��bkּF����xC��>�F6}�̬����x9���:8	;d�&;�;8;��A;՟F;�H;iyI;ɝI;*�I;gfI;�KI;�7I;�'I;�I;�I;�I;HI;�I;�I;�I;HI;�I;�I;�I;�'I;�7I;�KI;ffI;'�I;ɝI;kyI;߹H;џF;��A;�;8;d�&;8	;���:p�x9̬��F6}��>��xC�F���bkּ3��[G����95��ЈŽ��W��ʤ��3�      Kx��s���d�P�N�b�3�~I����J����z����\�C*��ݼF���+<<���ڻ�V��ct���&:���:rC;�</;�D=;�D;��G;'9I;�I;۔I;JtI;cVI;�?I;�-I;� I;�I;�I;�
I;-I;HI;-I;�
I;�I;�I;� I;�-I;�?I;`VI;HtI;ڔI; �I;)9I;��G;�D;�D=;�</;rC;���:��&:�ct��V���ڻ*<<�F����ݼC*���\��z��J������~I�b�3�P�N���d��s�      /l¾(��V������������d���7�z��:Sؽ[���d�D*�ckּ*\����'����R�}����:�Z;��#;j=7;`�A;G�F;��H;��I; �I;�I;!aI;�GI;'4I;Z%I;�I;�I;�I;
I;�	I;
I;�I;�I;�I;[%I;'4I;�GI;aI;�I;�I;��I;��H;B�F;]�A;j=7;��#;�Z;��:}���R�����'�*\��ckּD*��d�[��:Sؽz����7��d���������V���(��      �V������������Ͼ�d���ǆ�F�N��3��c�[����\�3��)C���o���	��눻����9v��:�h;�/;n�=;sE;,3H;�WI;�I;/�I;�kI;�OI;Y:I;*I;UI;�I;&I;�I;�I;�I;'I;�I;TI;*I;Y:I;�OI;�kI;/�I;�I;�WI;/3H;pE;l�=;�/;�h;r��:���9��눻��	��o�(C��3����\�[���cི3�F�N��ǆ��d����Ͼ���������      �,b�ƽ\��>M���5�=��4r��'l¾Ꝓ�%&W��3�:Sؽ�z��[G����zI����?���̻i�-�X	��t��:��;��&;V|9;�C;�dG;�I;r�I;��I;�vI;�WI;`@I;�.I;�!I;�I;�I;	I;�I;
I;�I;�I;�!I;�.I;`@I;�WI;�vI;��I;o�I;�I;�dG;�C;T|9;��&;��;r��:X	��h�-���̻��?�zI�����[G��z��:Sؽ�3�%&W�Ꝓ�'l¾4r��=����5��>M�ƽ\�      ���&��\���O䂿Ľ\���1�����J˾Ꝓ�F�N�z��J������W�'�c�Ҽ��|��z��n���w��|�&:�P�:ڨ;�W4;��@;ZgF;��H;C�I;R�I;k�I;L_I;FI;=3I;T%I;|I;�I;I;�I;I;�I;|I;T%I;;3I;FI;L_I;g�I;R�I;A�I;��H;[gF;��@;�W4;ڨ;�P�:x�&:�w���n���z���|�c�ҼW�'����J���z��F�N�Ꝓ��J˾�����1�Ľ\�O䂿\���&��      !}߿�$ڿ0�ʿ����
����Ps�SX:����'l¾�ǆ���7����95���Q�����t���75�\��w���!�8'ʼ:��;��.;��=;�EE;�YH;�hI;X�I;��I;VfI;PKI;\7I;y(I;	I;%I;�I;�I;�I;%I;I;v(I;\7I;PKI;UfI;�I;X�I;�hI;�YH;�EE;��=;��.;��;)ʼ:�!�8w��Z���75��t������Q�95�������7��ǆ�'l¾���SX:��Ps�
�������0�ʿ�$ڿ      |�����p������ſ&���Ps���1�4r���d���d�~I�ЈŽ��}�_*�JC���^��B�X�D�xE�� �:��;�);@7;;^D;w�G;~HI;�I;ߏI;�lI;&PI;;I;L+I;Q I;�I;�I;aI;�I;�I;P I;I+I;;I;&PI;�lI;ۏI;�I;|HI;v�G;_D;<7;;�);��;� �:�E�X�D��B��^�JC��_*���}�ЈŽ~I��d��d��4r����1��Ps�&����ſ��꿄p����      ��7��3�آ%�|��<����ſ
���Ľ\�=����Ͼ����b�3��轼z��}�9�^�἗���z�w7}��ct���^:�+�:ߣ#;ȍ8;��B;TsG;�%I;�I;'�I;5rI;HTI;>I;�-I;G"I;�I;I;�I;I;�I;G"I;�-I;>I;HTI;2rI;#�I;�I;�%I;QsG;��B;ō8;�#;�+�:��^:�ct�x7}��z����^��~�9��z����b�3�������Ͼ=��Ľ\�
�����ſ�<��|�آ%��3�      0�_��+Y��lG�!f.�|���꿳���O䂿��5���󾏰��P�N�W��S��"�Q����z����h!�xg����	:�
�:/�;v16;��A;�G;#I;k�I;��I;�vI;�WI;�@I;�/I;�#I;�I;@I;�I;@I;�I;�#I;�/I;�@I;�WI;�vI;��I;j�I;!I;�G;��A;r16;2�;�
�:�	:�xg���h!�z������"�Q�S��W��P�N���������5�O䂿�������|�!f.��lG��+Y�      Ҭ��%}�?tf��lG�آ%��p�0�ʿ\����>M����V�����d�ʤ�̷�/�d��
��I����1�V������p��9���:_;�U4;��@;!�F;R�H;�I;�I;�yI;�YI;wBI;	1I;�$I;�I;I;�I;I;�I;�$I;1I;uBI;�YI;�yI;�I;�I;R�H;!�F;��@;�U4;b;���:x��9���V�����1��I���
�0�d�̷�ʤ���d�V�������>M�\���0�ʿ�p�آ%��lG�?tf�%}�      T���E���%}��+Y��3�����$ڿ&��ƽ\����(���s��3�7����p�c�R���<<�*��>��� ��9���:�;d%3;|p@;zF;��H;/�I;(�I;�{I;�[I;�CI;�1I;�%I;ZI;�I;9I;�I;[I;�%I;�1I;�CI;�[I;�{I;%�I;/�I;��H;zF;|p@;b%3;�;���: ��9D���*���<<�R��c��p�7����3��s�(�����ƽ\�&���$ڿ����3��+Y�%}�E���      ����,������U���L�Q�Ǚ$�6�����>�}�I(�B�׾�T���L+���սk����L���iO���ͻ[���'m8�o�:��;l�1;��?; vF;� I;��I;��I;��I;�vI;�WI;BI;(2I;(I;"I;# I;"I;(I;(2I;BI;�WI;�vI;��I;��I;��I;� I; vF;��?;h�1;��;�o�:@(m8\����ͻ�iO�L����k����ս�L+��T��B�׾I(�>�}���6���Ǚ$�L�Q�U��������,��      �,��b��$P���{���K��x �����r�����w��$���Ҿh��� (���ѽҷ��'����۔K�4ɻ��� ��8���:��;��1;(@;��F;@I;�I;J�I;֞I;�uI;cWI;�AI;�1I;�'I;�!I; I;�!I;�'I;�1I;�AI;dWI;�uI;ԞI;H�I;�I;@I;��F;&@;��1;��;���: ��8���4ɻ۔K����'�ҷ����ѽ (�h�����Ҿ�$���w�r��������x ���K��{�$P��b��      ����$P�������d���;�$���㿴���#f�f�� ž��z���?�ƽ&0v�U5�.����o@�u���Hi��bu9�K�:U];�73;Y�@;/�F;jI;��I;��I;��I;tI;VI;w@I;1I;'I;B!I;dI;@!I;'I;1I;v@I;VI;tI;��I;��I;��I;jI;/�F;Y�@;�73;X];�K�:�bu9Ii�u����o@�/���U5�&0v�?�ƽ����z� žf��#f�������$����;���d����$P��      U����{���d��F�Ǚ$�;����ɿ0蒿��K�R���j��Zb�H�4���t�a����<�����.��d��
�غб�9Z�:mX;�25;Z�A;�!G;m7I;��I;��I;}�I;�pI;�SI;�>I;�/I;�%I;X I;fI;W I;�%I;�/I;�>I;�SI;�pI;|�I;��I;��I;m7I;�!G;Y�A;�25;pX;Z�:��9�غ�d����.�=������t�a�4���H�Zb��j��R����K�0蒿��ɿ;��Ǚ$��F���d��{�      L�Q���K���;�Ǚ$��;
��޿�����w�s,���澞���)�D������I��%�G�����N��~�������9:���: o!;��7;��B;��G;ZI;`�I;��I;�I;�lI;�PI;L<I;�-I;H$I;�I;�I;�I;F$I;�-I;J<I;�PI;�lI;�I;��I;`�I;ZI;��G;��B;��7;o!;���: �9:𓛺���}���N�����%�G��I������)�D��������s,���w�����޿�;
�Ǚ$���;���K�      Ǚ$��x �$��;���޿q���˅���F�~�
��~����z��$���ս���A2+���ϼPp�~���)�]�T�*�d��:D�;9';͌:;1�C;AH;�}I;R�I;��I;�I;�gI;�LI;Q9I;n+I;["I;*I;^I;*I;["I;n+I;Q9I;�LI;�gI;�I;��I;T�I;�}I;@H;/�C;Ɍ:;9';D�;j��:X�*�(�]�}���Pp���ϼA2+������ս�$���z��~��~�
��F�˅��q����޿;��$���x �      6��������㿌�ɿ���˅����P�e��>�׾�`��V�H����@��S�a���ʡ���D��ɻ� ��ѭ�#X�:�;�I-;^|=;[CE;܅H;;�I;�I;��I;�I;�aI;XHI;�5I;�(I; I;I;�I;I; I;�(I;�5I;XHI;�aI;�I;��I;�I;;�I;܅H;XCE;[|=;�I-;�;)X�:@ҭ�� ��ɻ�D�ʡ����S�a��@����V�H��`��>�׾e����P�˅�������ɿ�㿵���      ��r�������/蒿��w��F�e��Ͱ�"����Yb�+����ѽ�%��D4�ٟ�X������G��t潺p��9�r�: ;:3;RQ@;�vF;N�H;;�I;��I;��I;�zI;�ZI;ICI;�1I;�%I;xI;�I;YI;�I;xI;�%I;�1I;KCI;�ZI;�zI;��I;��I;:�I;N�H;�vF;NQ@;:3; ;�r�:`��9t潺�G�����X��ٟ�D4��%����ѽ+���Yb�"���Ͱ�e���F���w�/蒿����r���      >�}���w�#f���K�s,�~�
�>�׾"�����k���'�hz꽟I���;V�<M�����iO�ZG�IoE������:p� ;ֿ$;�8;��B;5�G;lKI;G�I;L�I;y�I;;qI;�SI;�=I;�-I;="I;�I;MI;�I;MI;�I;="I;�-I;�=I;�SI;;qI;v�I;L�I;E�I;lKI;2�G;��B;�8;ֿ$;p� ;���:��HoE�ZG໤iO����<M��;V��I��hz���'���k�"���>�׾~�
�s,���K�#f���w�      I(��$�f��R������~���`���Yb���'��U�J$��E�m�%����ϼ�/��6������L�غ�9�9���:G;H.;J|=;wE;�\H;X�I;��I;��I;0�I;6gI;7LI;8I;=)I;�I;�I;�I;_I;�I;�I;�I;<)I;8I;7LI;6gI;-�I;��I;��I;X�I;�\H;tE;I|=;H.;G;���:�9�9F�غ����6���/����ϼ%��E�m�J$���U���'��Yb��`���~�����R��f���$�      B�׾��Ҿ ž�j��������z�V�H�+��hz�I$���/v�2+�ܐ�����5��ɻ4��&�����:���:jo!;BP6;?lA;�F;��H;ȷI;��I;�I;�}I;�\I;�DI;<2I;�$I;�I;�I;�I;�I;�I;�I;�I;�$I;?2I;�DI;�\I;�}I;�I;��I;ʷI;��H;�F;=lA;BP6;jo!;���:���:�&��4��ɻ��5���ܐ�2+��/v�I$��hz�+��V�H���z������j�� ž��Ҿ      �T��h�����z�Zb�)�D��$�����ѽ�I��E�m�2+�������D�K���s�p�򖛺��9�T�:0;��-;��<;zD;�H;�mI;�I;��I;ƕI;�oI;�RI;�<I;7,I;�I;DI;iI;�I; I;�I;lI;EI;�I;:,I;�<I;�RI;�oI;ǕI;��I;�I;�mI;�H;}zD;��<;��-;0;�T�: ��9����s�p���D�K�������2+�E�m��I����ѽ���$�)�D�Zb���z�h���      �L+� (���H�������ս�@���%���;V�%��ܐ�����xMS�F����,D�@o8Vq�:�;��$;3_7;c�A;��F;/�H;��I;��I;��I;�I;�bI;�HI;D5I;[&I;eI;uI;%I;I;?
I;I;%I;uI;dI;\&I;D5I;�HI;�bI;�I;��I;��I;��I;+�H;��F;c�A;3_7;��$;�;^q�: o8*D���F��xMS�����ܐ�%���;V��%���@����ս����H��� (�      ��ս��ѽ>�ƽ3����I�����S�a�D4�<M���ϼ��D�K�F��<G��8f�@�o���:8C�:�Y;�1;�l>;E; 0H;SqI;9�I;!�I;�I;:sI;�UI;%?I;�-I;� I;�I;�I;�
I;JI;mI;JI;�
I;�I;�I;� I;�-I;&?I;�UI;:sI;�I;$�I;8�I;PqI;0H;E;�l>;�1;�Y;<C�:��:@�o�6f�:G��F��D�K�����ϼ<M�D4�S�a�����I��3���>�ƽ��ѽ      k��ҷ��&0v�s�a�%�G�@2+���ٟ�����/����5�����9f�p׬���g:��:7�;II-;Pg;;4OC;@SG;�I;��I;V�I;6�I;?�I;BcI;�II;�5I;�&I; I;nI;I;�I;�I;�I;�I;�I;I;nI;I;�&I;�5I;�II;DcI;>�I;9�I;V�I;��I;�I;@SG;3OC;Qg;;II-;:�;��:��g:p׬�9f�������5��/�����ٟ���@2+�%�G�s�a�&0v�ҷ��      
��'�T5���������ϼɡ��X���iO�6���ɻs�p�0D�`�o���g:K`�:vG;�*;�9;��A;�uF;S�H;��I;��I;�I;~�I;�pI;nTI;�>I;T-I;�I;�I;0I;�I;�I;�I;	I;�I;�I;�I;/I;�I;�I;T-I;�>I;nTI;�pI;��I;߻I;��I;��I;U�H;�uF;��A;�9;�*;rG;K`�:��g:@�o�0D�u�p��ɻ7���iO�X��ɡ����ϼ������T5�'�      L�����.���<����N��Pp��D����XG�����4�򖛺�o8��:��:rG;5�(;Ͷ7;��@;��E;�QH;NmI;��I;0�I;ԢI;_}I;�^I;�FI;4I;%I;�I;�I;)
I;FI;I; I;��H;  I;I;GI;(
I;�I;�I;%I;4I;�FI;�^I;a}I;ԢI;-�I;��I;NmI;�QH;��E;��@;ж7;5�(;rG;��:��:�o8����4�����XGເ���D�Pp��N��<���.������      �iO�ڔK��o@���.�~�������ɻ�G��EoE�F�غ�&����9Vq�:4C�:7�;�*;Ͷ7;�P@;�\E;'H;JI;��I;��I;D�I;��I;vhI;�NI;�:I;u*I;�I;�I;I;OI;FI;g�H;��H;�H;��H;g�H;GI;NI;I;�I;�I;r*I;�:I;�NI;yhI;��I;A�I;��I;��I;JI;)H;�\E;�P@;˶7;�*;7�;4C�:Tq�:��9�&��J�غEoE��G���ɻ���|����.��o@�ܔK�      ��ͻ2ɻo����d�����!�]�� �t潺����9�9���:�T�:�;�Y;KI-;�9;��@;�\E;��G;k5I;�I;~�I;�I;��I;�pI;�UI;�@I;n/I;�!I;�I;{I;�I;�I;W�H;��H;O�H;��H;O�H;��H;Y�H;�I;�I;{I;�I;�!I;n/I;�@I;�UI;�pI;��I;�I;~�I;�I;l5I;��G;�\E;��@;�9;LI-;�Y;�;�T�:���:�9�9 ��r潺� ��]�����d��o���2ɻ      X����Ei�
�غ�\�*� ҭ�@��9���:���:���:0;��$;�1;Mg;;��A;��E;$H;i5I;r�I;��I;��I;ϗI;�vI;�[I;�EI;�3I;o%I;�I;�I;�	I;�I;��H;��H;]�H;!�H;��H;#�H;]�H;��H;��H;�I;�	I;�I;�I;p%I;�3I;�EI;�[I;�vI;̗I;��I;��I;t�I;i5I;&H;��E;��A;Mg;;�1;��$;0;���:���:���:X��9 ҭ�T�*�ܓ���غCi���       *m8���8cu9���9�9:l��:-X�:�r�:r� ;G;jo!;��-;2_7;�l>;3OC;�uF;�QH;JI;�I;��I;�I;�I;�zI;�_I;II;�7I;�(I;�I;I;YI; I;b I;��H;��H;:�H;�H;��H;�H;:�H;��H;��H;b I; I;VI;I;�I;�(I;�7I;II;�_I;�zI;�I;�I;��I;�I;	JI;�QH;�uF;3OC;�l>;2_7;��-;ho!;G;r� ;�r�:)X�:r��:�9:���9�bu9���8      �o�:���:�K�:�Y�:���:M�;�;! ;ܿ$;H.;FP6;��<;`�A;E;@SG;R�H;NmI;��I;~�I;��I;�I;|I;�aI;�KI;�9I;+I;�I;�I;�I;cI;*I;-�H;	�H;��H;(�H;G�H;	�H;G�H;(�H;��H;�H;-�H;(I;`I;�I;�I;�I;+I;�9I;�KI;�aI;|I;�I;��I;~�I;��I;MmI;Q�H;@SG;E;`�A;��<;DP6;H.;ݿ$;$ ;�;O�;֨�:�Y�:�K�:��:      ��;��;X];gX;�n!;9';�I-;:3;�8;K|=;?lA;�zD;��F;#0H;�I;��I;��I;��I;�I;ЗI;�zI;�aI;�LI;Y;I;�,I;n I;`I;2I;vI;I;��H;7�H;��H;��H;B�H;��H;\�H;��H;B�H;��H;��H;6�H;��H;I;tI;3I;]I;p I;�,I;V;I;�LI;�aI;�zI;ӗI;�I;��I;��I;��I;�I;"0H;��F;�zD;@lA;J|=;�8;:3;�I-;9';o!;iX;Y];��;      ��1;��1;�73;�25;��7;ʌ:;e|=;MQ@;��B;xE;�F;�H;+�H;SqI;��I;��I;/�I;E�I;��I;�vI;�_I;�KI;W;I;-I;'!I;VI;I;SI;�I;5�H;��H;��H;a�H;��H;��H;�H;��H;�H;��H;��H;^�H;��H;��H;2�H;�I;SI;I;WI;(!I;-I;V;I;�KI;�_I;�vI;��I;F�I;-�I;��I;��I;SqI;*�H;�H;�F;vE;��B;OQ@;c|=;̌:;��7;�25;�73;��1;      ��?;0@;E�@;]�A;��B;1�C;WCE;�vF;3�G;�\H;��H;�mI;��I;;�I;X�I;�I;٢I;��I;�pI;�[I;�II;�9I;�,I;-!I;�I;�I;�I;3I;��H;��H;��H;e�H;��H;+�H;*�H;��H;k�H;��H;*�H;+�H;��H;h�H;��H;��H;��H;3I;�I;�I;�I;*!I;�,I;�9I;�II;�[I;�pI;��I;֢I;߻I;X�I;9�I;��I;�mI;��H;�\H;3�G;�vF;WCE;2�C;��B;]�A;D�@;/@;      ,vF;ʊF; �F;�!G;��G;9H;ۅH;I�H;oKI;X�I;ȷI;�I;��I;!�I;6�I;}�I;b}I;whI;�UI;�EI;�7I;+I;k I;SI;�I;	I;�I;��H;*�H;�H;c�H;x�H;��H;��H;��H;S�H;%�H;S�H;��H;��H;��H;y�H;c�H;�H;)�H;��H;�I;	I;�I;SI;k I;+I;�7I;�EI;�UI;yhI;a}I;}�I;6�I;"�I;��I;�I;ȷI;V�I;nKI;K�H;ۅH;9H;��G;�!G; �F;��F;      � I;@I;dI;q7I;ZI;�}I;>�I;7�I;I�I;��I;��I;��I;��I;�I;?�I;�pI;�^I;�NI;�@I;�3I;�(I;�I;_I;I;�I;�I;�H;`�H;�H;q�H;a�H;��H;T�H;V�H;��H;A�H;�H;A�H;��H;U�H;S�H;��H;a�H;p�H;�H;`�H;�H;�I;�I;I;]I;�I;�(I;�3I;�@I;�NI;�^I;�pI;?�I;�I;��I;��I;��I;��I;I�I;9�I;@�I;�}I; ZI;p7I;fI;BI;      ��I;�I;��I;��I;^�I;R�I;�I;��I;P�I;��I;�I;˕I;�I;=sI;EcI;oTI;�FI;�:I;o/I;q%I;�I;�I;5I;VI;0I;��H;^�H;5�H;~�H;a�H;��H;�H;�H;@�H;��H;<�H;+�H;=�H;��H;@�H;�H;�H;��H;^�H;}�H;7�H;^�H;��H;2I;VI;3I;�I;�I;q%I;n/I;�:I;�FI;oTI;DcI;;sI;�I;˕I;�I;��I;Q�I;��I;�I;T�I;h�I;��I;��I;$�I;      �I;G�I;��I;��I;��I;��I;��I;��I;x�I;/�I;�}I;�oI;�bI;�UI;�II;�>I;4I;t*I;�!I;�I;I;�I;uI;�I;��H;,�H;�H;~�H;h�H;��H;�H;��H;��H;8�H;��H;p�H;h�H;p�H;��H;8�H;��H;��H;
�H;��H;h�H;~�H;�H;*�H;��H;�I;tI;�I;I;�I;�!I;u*I;4I;�>I;�II;�UI;�bI;�oI;�}I;/�I;x�I;��I;��I;��I;��I;��I;��I;=�I;      ��I;۞I;��I;}�I;��I;�I;�I;�zI;CqI;=gI;�\I;�RI;�HI;-?I;6I;X-I;!%I;�I;�I;�I;ZI;bI;I;3�H;��H;�H;o�H;`�H;��H;�H;��H;��H;��H;[�H;��H;��H;��H;��H;��H;[�H;��H;��H;��H;�H;��H;`�H;m�H;�H;��H;5�H;I;bI;YI;�I;�I;�I; %I;X-I;�5I;,?I;�HI;�RI;�\I;=gI;CqI;�zI;�I;�I;��I;~�I;��I;۞I;      �vI;�uI;tI;�pI;�lI;�gI;�aI;[I;�SI;<LI;�DI;�<I;J5I;�-I;�&I;�I;�I;�I;�I;�	I;(I;+I;��H;��H;��H;e�H;^�H;��H;�H;��H;��H;��H;&�H;��H;H�H;�H;��H;�H;H�H;��H;#�H;��H;��H;��H;�H;��H;^�H;c�H;��H;��H;��H;+I;$I;�	I;�I;�I;�I;�I;�&I;�-I;J5I;�<I;�DI;>LI;�SI;[I;�aI;�gI;�lI;�pI;tI;�uI;      �WI;nWI;VI;�SI;�PI;�LI;XHI;OCI;�=I;8I;A2I;B,I;_&I;� I;
I;�I;�I;I;�I;�I;k I;2�H;:�H;��H;c�H;x�H;��H;�H;��H;��H;��H;"�H;��H;�H;��H;��H;��H;��H;��H;�H;}�H;#�H;��H;��H;��H;�H;��H;v�H;f�H;��H;7�H;2�H;h I;�I;�I;I;�I;�I;	I;� I;]&I;A,I;A2I;8I;�=I;OCI;WHI;�LI;�PI;�SI;VI;jWI;      BI;�AI;|@I;�>I;S<I;P9I;�5I;�1I;�-I;<)I;�$I; I;gI;�I;tI;5I;2
I;MI;�I;��H;��H;�H;��H;c�H;��H;��H;W�H;�H;��H;��H;'�H;��H;��H;��H;G�H;�H;%�H;�H;G�H;��H;��H;��H;'�H;��H;��H;�H;S�H;��H;��H;c�H;��H;�H;��H;��H;�I;NI;/
I;5I;qI;�I;eI;�I;�$I;=)I;�-I;�1I;�5I;Q9I;L<I;�>I;|@I;�AI;      32I;�1I;1I;�/I;�-I;h+I;�(I;�%I;C"I;�I;�I;LI;xI;�I;I;�I;QI;HI;`�H;��H;��H;��H;��H;��H;'�H;��H;R�H;?�H;5�H;X�H;��H;�H;��H;.�H;�H;��H;��H;��H;�H;.�H;��H;�H;��H;Z�H;8�H;?�H;R�H;��H;)�H;��H;��H;��H;��H;��H;`�H;JI;PI;�I;I;�I;xI;LI;�I;�I;D"I;�%I;�(I;m+I;�-I;�/I;1I;�1I;      (I;�'I;"'I;�%I;]$I;U"I; I;~I;�I;�I;�I;vI;+I; I;�I;�I;!I;g�H;��H;f�H;E�H;,�H;C�H;��H;#�H;��H;��H;��H;��H;��H;H�H;��H;G�H;�H;��H;��H;��H;��H;��H;�H;D�H;��H;H�H;��H;��H;��H;��H;��H;#�H;��H;B�H;,�H;B�H;f�H;��H;g�H; I;�I;�I; I;+I;vI;�I;�I;�I;~I; I;X"I;S$I;�%I;"'I;�'I;      "I;�!I;I!I;[ I;I;&I;I;�I;YI;�I;�I;�I;I;TI;�I;�I;, I;��H;V�H;*�H;(�H;J�H;��H;�H;��H;R�H;A�H;<�H;r�H;��H;�H;��H;�H;��H;��H;j�H;e�H;j�H;��H;��H;�H;��H;�H;��H;s�H;<�H;@�H;P�H;��H;�H;��H;J�H;&�H;+�H;V�H;��H;) I;�I;�I;SI;I;�I;�I;�I;YI;�I;I;*I;�I;Z I;I!I;�!I;        I;
 I;oI;jI;I;ZI;�I;]I;�I;\I;�I;I;A
I;tI;�I;I;��H;�H;��H;��H;��H;�H;]�H;��H;g�H;"�H;�H;/�H;i�H;��H;��H;��H;'�H;��H;��H;f�H;L�H;f�H;��H;��H;"�H;��H;��H;��H;l�H;/�H;�H;#�H;g�H;��H;]�H;�H;��H;��H;��H;�H;��H;I;�I;tI;A
I;I;�I;_I;�I;]I;�I;`I;�I;jI;oI; I;      "I;�!I;I!I;Z I;I;&I;I;�I;[I;�I;�I;�I;I;TI;�I;�I;, I;��H;V�H;*�H;)�H;J�H;��H;�H;��H;R�H;A�H;<�H;r�H;��H;�H;��H;�H;��H;��H;j�H;e�H;j�H;��H;��H;�H;��H;�H;��H;s�H;<�H;?�H;P�H;��H;�H;��H;J�H;&�H;+�H;V�H;��H;) I;�I;�I;SI;I;�I;�I;�I;YI;�I;I;*I;�I;[ I;F!I;�!I;      (I;�'I;!'I;�%I;]$I;U"I; I;~I;�I;�I;�I;vI;+I; I;�I;�I;!I;g�H;��H;f�H;F�H;,�H;C�H;��H;#�H;��H;��H;��H;��H;��H;H�H;��H;G�H;�H;��H;��H;��H;��H;��H;�H;D�H;��H;H�H;��H;��H;��H;��H;��H;#�H;��H;B�H;,�H;B�H;f�H;��H;g�H; I;�I;�I; I;+I;vI;�I;�I;�I;~I; I;X"I;S$I;�%I;!'I;�'I;      52I;�1I;1I;�/I;�-I;h+I;�(I;�%I;C"I;�I;�I;LI;xI;�I;I;�I;QI;HI;`�H;��H;��H;��H;��H;��H;)�H;��H;R�H;?�H;6�H;X�H;��H;�H;��H;.�H;�H;��H;��H;��H;�H;.�H;��H;�H;��H;Z�H;8�H;?�H;R�H;��H;'�H;��H;��H;��H;��H;��H;`�H;JI;PI;�I;I;�I;xI;LI;�I;�I;D"I;�%I;�(I;m+I;�-I;�/I;1I;�1I;      BI;�AI;}@I;�>I;Q<I;N9I;�5I;�1I;�-I;<)I;�$I;�I;eI;�I;qI;5I;2
I;MI;�I;��H;��H;�H;��H;c�H;��H;��H;V�H;�H;��H;��H;'�H;��H;��H;��H;G�H;�H;%�H;�H;G�H;��H;��H;��H;'�H;��H;��H;�H;S�H;��H;��H;b�H;��H;�H;��H;��H;�I;MI;/
I;5I;tI;�I;eI; I;�$I;=)I;�-I;�1I;�5I;Q9I;L<I;�>I;|@I;�AI;      �WI;nWI;	VI;�SI;�PI;�LI;ZHI;OCI;�=I;8I;A2I;A,I;]&I;� I;	I;�I;�I;I;�I;�I;n I;2�H;:�H;��H;f�H;x�H;��H;�H;��H;��H;��H;"�H;�H;�H;��H;��H;��H;��H;��H;�H;}�H;#�H;��H;��H;��H;�H;��H;v�H;c�H;��H;9�H;2�H;h I;�I;�I;I;�I;�I;
I;� I;_&I;B,I;A2I; 8I;�=I;OCI;ZHI;�LI;�PI;�SI;	VI;kWI;      �vI;�uI;tI;�pI;�lI;�gI;�aI; [I;�SI;<LI;�DI;�<I;J5I;�-I;�&I;�I;�I;�I;�I;�	I;*I;+I;��H;��H;��H;e�H;^�H;��H;�H;��H;��H;��H;%�H;��H;H�H;�H;��H;�H;H�H;��H;#�H;��H;��H;��H;�H;��H;^�H;c�H;��H;��H;��H;+I;$I;�	I;�I;�I;�I;�I;�&I;�-I;J5I;�<I;�DI;>LI;�SI;[I;�aI;�gI;�lI;�pI;tI;�uI;      ��I;۞I;��I;}�I;�I;�I;�I;�zI;DqI;;gI;�\I;�RI;�HI;-?I;�5I;X-I;!%I;�I;�I;�I;]I;bI;I;3�H;��H;�H;o�H;`�H;��H;�H;��H;��H;��H;Z�H;��H;��H;��H;��H;��H;[�H;��H;��H;��H;�H;��H;`�H;m�H;�H;��H;5�H;I;bI;YI;�I;�I;�I; %I;Z-I;6I;-?I;�HI;�RI;�\I;;gI;DqI;�zI;�I;�I;��I;}�I;��I;ޞI;      ��I;C�I;��I;��I;��I;��I;��I;��I;x�I;/�I;�}I;�oI;�bI;�UI;�II;�>I;4I;u*I;�!I;�I;I;�I;vI;�I;��H;,�H;�H;~�H;h�H;��H;
�H;��H;��H;8�H;��H;p�H;h�H;p�H;��H;8�H;��H;��H;�H;��H;h�H;~�H;�H;*�H;��H;�I;tI;�I;I;�I;�!I;u*I;4I;�>I;�II;�UI;�bI;�oI;�}I;-�I;y�I;ĤI;��I;��I;��I;��I;��I;D�I;      ��I;�I;��I;��I;\�I;T�I;�I;��I;P�I;��I;�I;˕I;�I;=sI;EcI;oTI;�FI;�:I;n/I;q%I;�I;�I;5I;VI;2I;��H;^�H;7�H;~�H;a�H;��H;�H;�H;?�H;��H;<�H;+�H;=�H;��H;@�H;�H;�H;��H;^�H;}�H;5�H;^�H;��H;0I;VI;3I;�I;�I;q%I;o/I;�:I;�FI;pTI;EcI;;sI;�I;͕I;�I;��I;P�I;��I;�I;O�I;j�I;��I;��I;$�I;      � I;?I;gI;k7I;ZI;�}I;>�I;7�I;I�I;��I;��I;��I;��I;�I;?�I;�pI;�^I;�NI;�@I;�3I;�(I;�I;_I;I;�I;�I;�H;`�H;�H;q�H;a�H;��H;T�H;U�H;��H;A�H;�H;@�H;��H;U�H;S�H;��H;a�H;p�H;�H;`�H;�H;�I;�I;I;]I;�I;�(I;�3I;�@I;�NI;�^I;�pI;?�I;�I;��I;��I;��I;��I;H�I;7�I;=�I;�}I;ZI;k7I;fI;6I;      0vF;ƊF;+�F;�!G;��G;:H;ۅH;J�H;nKI;X�I;ȷI;�I;��I;"�I;5�I;}�I;b}I;yhI;�UI;�EI;�7I;+I;k I;SI;�I;	I;�I;��H;*�H;�H;c�H;x�H;��H;��H;��H;S�H;%�H;S�H;��H;��H;��H;y�H;c�H;�H;)�H;��H;�I;	I;�I;SI;k I;+I;�7I;�EI;�UI;yhI;a}I;}�I;6�I;"�I;��I;�I;ȷI;U�I;lKI;I�H;ޅH;9H;��G;�!G;+�F;��F;      ��?;0@;E�@;]�A;��B;1�C;WCE;�vF;3�G;�\H;��H;�mI;��I;9�I;X�I;�I;آI;��I;�pI;�[I;�II;�9I;�,I;-!I;�I;�I;�I;3I;��H;��H;��H;f�H;��H;+�H;(�H;��H;k�H;��H;*�H;)�H;��H;h�H;��H;��H;��H;3I;�I;�I;�I;+!I;�,I;�9I;II;�[I;�pI;��I;֢I;�I;X�I;9�I;��I;�mI;��H;�\H;2�G;�vF;WCE;1�C;�B;]�A;D�@;0@;      ��1;��1;83;�25;��7;Ќ:;a|=;NQ@;��B;xE;�F;�H;-�H;SqI;��I;��I;/�I;E�I;��I;�vI;�_I;�KI;Y;I;-I;(!I;WI;I;SI;�I;5�H;��H;��H;_�H;��H;��H;�H;��H;�H;��H;��H;_�H;��H;��H;2�H;�I;SI;I;VI;'!I;-I;V;I;�KI;�_I;�vI;��I;F�I;-�I;��I;��I;TqI;+�H;�H;�F;vE;��B;NQ@;a|=;Ќ:;��7;�25;83;��1;      ��;��;i];iX;�n!;9';�I-;:3;�8;K|=;@lA;�zD;��F;"0H;�I;��I;��I;��I;�I;ЗI;�zI;�aI;�LI;Y;I;�,I;o I;_I;3I;vI;I;��H;6�H;��H;��H;B�H;��H;\�H;��H;B�H;��H;��H;7�H;��H;I;tI;2I;\I;o I;�,I;V;I;�LI;�aI;�zI;ӗI;�I;��I;��I;��I;�I;#0H;��F;�zD;@lA;J|=;�8;:3;�I-;9';�n!;iX;]];��;      �o�:���:�K�:�Y�:���:M�;�;! ;ܿ$;H.;FP6;��<;`�A;E;>SG;R�H;MmI;��I;~�I;��I;�I;|I;�aI;�KI;�9I;+I;�I;�I;�I;dI;(I;-�H;�H;��H;(�H;G�H;	�H;G�H;(�H;��H;�H;-�H;*I;`I;�I;�I;�I;+I;�9I;�KI;�aI;|I;�I;��I;~�I;��I;MmI;R�H;ASG;E;`�A;��<;DP6;H.;ܿ$;# ;�;M�;Ԩ�:�Y�:�K�:��:      @(m8 ��8Pcu9���9�9:^��:/X�:�r�:r� ;G;jo!;��-;2_7;�l>;3OC;�uF;�QH;JI;�I;��I;�I;�I;�zI;�_I;II;�7I;�(I;�I;I;WI; I;a I;��H;��H;:�H;�H;��H;�H;:�H;��H;��H;d I; I;VI;I;�I;�(I;�7I;II;�_I;�zI;�I;�I;��I;�I;	JI;�QH;�uF;3OC;�l>;2_7;��-;jo!;G;t� ;�r�:/X�:r��: �9:���9Pcu9���8      Y����Ai��غ擛�X�*� ҭ�H��9���:���:���:0;��$;�1;Kg;;��A;��E;$H;i5I;r�I;��I;��I;ЗI;�vI;�[I;�EI;�3I;p%I;�I;�I;�	I;�I;��H;��H;]�H;#�H;��H;#�H;]�H;��H;��H;�I;�	I;�I;�I;o%I;�3I;�EI;�[I;�vI;̗I;��I;��I;t�I;i5I;&H;��E;��A;Mg;;�1;��$;0;���:���:���:`��9 ҭ�T�*�ܓ���غCi���      ��ͻ2ɻo����d�����"�]�� �t潺 ���9�9���:�T�:�;�Y;KI-;�9;��@;�\E;��G;k5I;�I;~�I;�I;��I;�pI;�UI;�@I;n/I;�!I;�I;{I;�I;�I;Y�H;��H;O�H;��H;O�H;��H;W�H;�I;�I;{I;�I;�!I;n/I;�@I;�UI;�pI;��I;�I;~�I;�I;l5I;��G;�\E;��@;�9;LI-;�Y;�;�T�:���:�9�9���t潺� ��]�����d��o���2ɻ      �iO�ٔK��o@���.�~�������ɻ�G��EoE�L�غ�&����9Tq�:2C�:7�;�*;Ͷ7;�P@;�\E;'H;JI;��I;��I;E�I;��I;whI;�NI;�:I;u*I;�I;�I;I;OI;GI;g�H;��H;�H;��H;g�H;FI;NI;I;�I;�I;r*I;�:I;�NI;yhI;��I;>�I;��I;��I;JI;)H;�\E;�P@;̶7;�*;7�;4C�:Vq�:��9�&��F�غFoE��G���ɻ~���|����.��o@�۔K�      L�����.���<����N��Pp��D����XG�����4������o8��:��:rG;7�(;Ͷ7;��@;��E;�QH;NmI;��I;1�I;ԢI;_}I;�^I;�FI;4I;%I;�I;�I;)
I;GI;I; I;��H; I;I;GI;(
I;�I;�I;%I;4I;�FI;�^I;a}I;ԢI;,�I;��I;NmI;�QH;��E;��@;ж7;5�(;rG;��:��:�o8򖛺4�����XGເ���D�Pp��N��<���.������      ��&�T5���������ϼɡ��X���iO�6���ɻu�p�0D�`�o���g:K`�:uG;�*;�9;��A;�uF;U�H;��I;��I;߻I;��I;�pI;nTI;�>I;T-I;�I;�I;0I;�I;�I;�I;	I;�I;�I;�I;/I;�I;�I;T-I;�>I;nTI;�pI;��I;�I;��I;��I;S�H;�uF;��A;�9;�*;uG;K`�:��g:@�o�0D�s�p��ɻ6���iO�X��ɡ����ϼ������T5�'�      k��ҷ��&0v�s�a�%�G�@2+���ٟ�����/����5�����9f�p׬���g:��:7�;II-;Pg;;3OC;@SG;�I;�I;V�I;8�I;?�I;DcI;�II;�5I;�&I; I;pI;I;�I;�I;�I;�I;�I;I;nI;I;�&I;�5I;�II;BcI;>�I;8�I;V�I;��I;�I;@SG;3OC;Qg;;II-;:�;��:��g:p׬�8f�������5��/�����ٟ���@2+�%�G�s�a�&0v�ҷ��      ��ս��ѽ>�ƽ3����I�����S�a�D4�<M���ϼ��D�K�F��<G��6f�@�o���::C�:�Y;�1;�l>;E; 0H;TqI;8�I;"�I;�I;:sI;�UI;%?I;�-I;� I;�I;�I;�
I;JI;mI;JI;�
I;�I;�I;� I;�-I;%?I;�UI;:sI;�I;"�I;9�I;PqI;0H;E;�l>;�1;�Y;<C�:��:@�o�8f�:G��F��D�K�����ϼ<M�D4�S�a�����I��3���>�ƽ��ѽ      �L+� (���H�������ս�@���%���;V�%��ܐ�����xMS�F����,D⺀o8\q�:�;��$;2_7;c�A;��F;/�H;��I;��I;��I;�I;�bI;�HI;D5I;[&I;dI;uI;%I;I;?
I;I;%I;uI;dI;[&I;D5I;�HI;�bI;�I;��I;��I;��I;(�H;��F;c�A;2_7;��$;�;^q�:@o8,D���E��xMS�����ܐ�%���;V��%���@����ս����H��� (�      �T��h�����z�Zb�)�D��$�����ѽ�I��E�m�2+�������D�K���s�p�򖛺��9�T�:0;��-;��<;zD;�H;�mI;�I;��I;ǕI;�oI;�RI;�<I;7,I;�I;GI;lI;�I; I;�I;iI;DI;�I;8,I;�<I;�RI;�oI;ƕI;��I;�I;�mI;�H;}zD;��<;��-;0;�T�: ��9����v�p���D�K�������2+�E�m��I����ѽ���$�)�D�Zb���z�h���      B�׾��Ҿ ž�j��������z�V�H�+��hz�J$���/v�2+�ܐ�����5��ɻ4��&�����:���:ho!;BP6;@lA;�F;��H;ʷI;��I;�I;�}I;�\I;�DI;<2I;�$I;�I;�I;�I;�I;�I;�I;�I;�$I;=2I;�DI;�\I;�}I;�I;��I;ȷI;��H;�F;=lA;BP6;jo!;���:���:�&��4��ɻ��5���ܐ�2+��/v�I$��hz�+��V�H���z������j�� ž��Ҿ      I(��$�f��R������~���`���Yb���'��U�J$��E�m�%����ϼ�/��6������J�غ�9�9���:G;H.;J|=;xE;�\H;Y�I;��I;��I;0�I;6gI;7LI;8I;=)I;�I;�I;�I;_I;�I;�I;�I;<)I;8I;7LI;6gI;-�I;��I;��I;X�I;�\H;tE;I|=;H.;G;���:�9�9F�غ����6���/����ϼ%��E�m�J$���U���'��Yb��`���~�����R��f���$�      >�}���w�#f���K�s,�~�
�=�׾"�����k���'�hz꽟I���;V�<M�����iO�YG�HoE������:n� ;ֿ$;�8;��B;2�G;nKI;H�I;L�I;y�I;9qI;�SI;�=I;�-I;="I;�I;MI;�I;MI;�I;="I;�-I;�=I;�SI;9qI;v�I;L�I;E�I;lKI;5�G;��B;�8;ֿ$;p� ;���:��FoE�ZG໤iO����<M��;V��I��hz���'���k�"���=�׾~�
�s,���K�#f���w�      ��r�������/蒿��w��F�e��Ͱ�"����Yb�+����ѽ�%��D4�ٟ�X������G��t潺p��9�r�: ;:3;QQ@;�vF;P�H;;�I;��I;¤I;�zI;�ZI;ICI;�1I;�%I;zI;�I;YI;�I;xI;�%I;�1I;HCI;�ZI;�zI;��I;��I;:�I;M�H;�vF;NQ@;:3; ;�r�:X��9t潺�G�����X��ٟ�D4��%����ѽ+���Yb�"���Ͱ�e���F���w�/蒿����r���      6��������㿌�ɿ���˅����P�e��>�׾�`��V�H����@��S�a���ʡ���D��ɻ� � ҭ�#X�:�;�I-;_|=;XCE;ޅH;;�I;�I;��I;�I;�aI;XHI;�5I;�(I; I;I;�I;I; I;�(I;�5I;WHI;�aI;�I;��I;�I;:�I;܅H;[CE;[|=;�I-;�;'X�:@ҭ�� ��ɻ�D�ʡ����S�a��@����V�H��`��>�׾e����P�˅�������ɿ�㿵���      Ǚ$��x �$��;���޿q���˅���F�~�
��~����z��$���ս���A2+���ϼPp�~���(�]�X�*�`��:D�;9';͌:;/�C;AH;�}I;T�I;��I;�I;�gI;�LI;Q9I;n+I;["I;*I;^I;+I;["I;n+I;P9I;�LI;�gI;�I;��I;R�I;�}I;@H;1�C;Ɍ:;9';D�;f��:X�*�)�]�}���Pp���ϼA2+������ս�$���z��~��~�
��F�˅��q����޿;��$���x �      L�Q���K���;�Ǚ$��;
��޿�����w�s,���澞���)�D������I��%�G�����N��~�����𓛺�9:���: o!;��7;��B;��G;ZI;`�I;��I;�I;�lI;�PI;J<I;�-I;H$I;�I;�I;�I;F$I;�-I;J<I;�PI;�lI;�I;��I;`�I;ZI;��G;��B;��7;o!;���: �9:𓛺���}���N�����%�G��I������)�D��������s,���w�����޿�;
�Ǚ$���;���K�      U����{���d��F�Ǚ$�;����ɿ0蒿��K�R���j��Zb�H�4���t�a����<�����.��d��
�غȱ�9Z�:mX;�25;Y�A;�!G;m7I;��I;��I;~�I;�pI;�SI;�>I;�/I;�%I;W I;fI;X I;�%I;�/I;�>I;�SI;�pI;|�I;��I;��I;m7I;�!G;Z�A;�25;pX;Z�:��9�غ�d����.�=������t�a�3���H�Zb��j��R����K�0蒿��ɿ;��Ǚ$��F���d��{�      ����$P�������d���;�$���㿴���#f�f�� ž��z���?�ƽ&0v�U5�.����o@�u���Ii��bu9�K�:U];�73;Y�@;/�F;kI;��I;��I;��I;tI;VI;w@I;1I;'I;@!I;dI;B!I;'I;1I;v@I;VI;tI;��I;��I;��I;hI;/�F;Y�@;�73;X];�K�:�bu9Ii�u����o@�/���U5�&0v�?�ƽ����z� žf��#f�������$����;���d����$P��      �,��b��$P���{���K��x �����r�����w��$���Ҿh��� (���ѽҷ��'����۔K�4ɻ��� ��8���:��;��1;&@;��F;@I;�I;J�I;מI;�uI;cWI;�AI;�1I;�'I;�!I; I;�!I;�'I;�1I;�AI;dWI;�uI;ԞI;H�I;�I;?I;��F;(@;��1;��;���: ��8���4ɻ۔K����'�ҷ����ѽ (�h�����Ҿ�$���w�r��������x ���K��{�$P��b��      E(��r'���o��O�d��X1�x�Ŀ����3�y���x����4�m��Z+���'���ü2yY��kٻ�o&���p����:{;��0;��?;
�F;� I;2�I;��I;X�I;��I;�dI;�KI;:I;�.I;�'I;�%I;�'I;�.I;:I;�KI;�dI;��I;W�I;��I;2�I;� I;
�F;��?;��0;};���: �p��o&��kٻ2yY���ü�'�Z+��m�ཿ�4��x��y���3����Ŀx��X1�d�O��o��r'��      r'���X��g^�������]]���,�Q9�7g��U�����/����o��i1��hܽ���-$�^l���|U�V�ԻM!� �,���:;�51;��?;��F;a'I;��I;N�I;k�I;ՆI;dI;tKI;�9I;[.I;�'I;�%I;�'I;\.I;�9I;rKI;dI;ՆI;i�I;K�I;��I;a'I;��F;��?;�51;";��: �,�O!�V�Ի�|U�^l���-$����hܽi1��o���ྜ�/�U���7g��Q9���,��]]�����g^���X��      �o��g^���ē��4z�6K�i��T��(ﱿV�v��X#���Ѿń�	�&�r�нd̀�`��s���D�I�{ǻ�4�P$9-�:s�;;�2;��@;�F;;I;&�I;2�I;ʲI;��I;�bI;2JI;�8I;�-I;�&I;%I;�&I;�-I;�8I;0JI;�bI;��I;ȲI;1�I;&�I;;I;�F;��@;7�2;x�;-�:`$9�4�|ǻC�I�t���`��d̀�r�н�&�ń���Ѿ�X#�V�v�(ﱿT��i��6K��4z��ē�g^��      O������4z���V��X1��<�uؿ����RZ��	�*���LUo����_y��/l�Z��R��;�7� �������Ƴ9H��:�;x�4;�tA;�2G;�XI;��I;��I;9�I;+�I;�_I;0HI;W7I;3,I;�%I;�#I;�%I;3,I;Y7I;.HI;�_I;+�I;7�I;��I;��I;�XI;�2G;�tA;s�4;�;H��: ǳ9��� ���:�7��R��Z�/l�_y�����LUo�*����	��RZ����uؿ�<��X1���V��4z�����      d��]]�6K��X1�[f��pQ��U���]58��A���נ���O���a什�Q����<ߓ��� ��V��氺��":'��:@ ;17;<�B;w�G;|I;�I;��I;�I;p|I;o\I;EI;Q5I;m*I;d$I;`"I;d$I;k*I;S5I;~EI;o\I;p|I;�I;��I;�I;|I;u�G;<�B;17;D ;'��:��":氺�V���� �<ߓ�����Q�a什����O��נ��A��]58�U���pQ���[f��X1�6K��]]�      �X1���,�i���<��7g��f_���U�ς�،Ⱦ
ń�,�-�k��R ��&�2�	?ټ\�{��!��n�T�O�8�u:Q ;&;R#:;x�C;8&H;E�I;Y�I; �I;�I;�vI;
XI;$BI;�2I;I(I;w"I;� I;w"I;I(I;�2I;$BI;XI;�vI;�I;��I;Y�I;D�I;7&H;u�C;K#:;&;Q ;<�u:X�O��n��!�]�{�	?ټ&�2�R ��k��,�-�
ń�،Ⱦς��U�f_��7g��<�i����,�      x�Q9�T��uؿpQ��f_��8�_��X#�s���f��<�S�{�����l�B�w���M���Ի��+��9T���:�e;�\,;#0=;�BE;��H;��I;�I;��I;�I;�oI;�RI;H>I;�/I;�%I;' I;{I;' I;�%I;�/I;H>I;�RI;�oI;�I;��I;�I;��I;��H;�BE;0=;�\,;�e;��: :T���+���Ի�M�w��B�l�����{�<�S��f��s���X#�8�_�f_��pQ��uؿT��Q9�      Ŀ7g��(ﱿ���U����U��X#�v��f���KUo�	�#��hܽ����n<����9����� ��᝻�Ժ0v�9���:�V;�2;� @;��F;I;.�I;v�I;b�I;��I;7hI;DMI;�9I;%,I;�"I;�I;�I;�I;�"I;%,I;�9I;FMI;7hI;��I;_�I;v�I;-�I;I;��F;� @;�2;�V;���:0v�9�Ժ�᝻�� �9�������n<�����hܽ	�#�KUo�f���v���X#��U�U������(ﱿ7g��      ���U���V�v��RZ�]58�ς�s��f���ioy�_1�bO��]什�`�N�����iyY���m�T�`�1�X�u:\��:v#;H98;8�B;��G;*mI;D�I;3�I;d�I;��I;`I;9GI;*5I;[(I;�I;�I;CI;�I;�I;](I;*5I;9GI;`I;��I;a�I;5�I;A�I;*mI;��G;6�B;H98;x#;^��:P�u:`�1�k�T���iyY����N���`�]什bO��_1�ioy�f���s��ς�]58��RZ�V�v�U���      �3���/��X#��	��A��،Ⱦ�f��KUo�_1�Ͱ��}n��ռx��'��>ټ�@���k�����Ĵ��39$�:\R;=e-;�/=;
E;�xH;��I;D�I;��I;9�I;GvI;�WI;�@I;*0I;Z$I;vI;�I;nI;�I;vI;[$I;*0I;�@I;�WI;HvI;6�I;��I;D�I;��I;�xH;�	E;�/=;=e-;\R;	$�:��39��𺼼���k��@���>ټ�'�ռx�}n��Ͱ��_1�KUo��f��،Ⱦ�A���	��X#���/�      y���྅�Ѿ*����נ�
ń�<�S�	�#�bO��}n��J̀���2����|�>��Իd�B�#��m::H�:� ;̼5;�FA;��F;�I;��I;��I;پI;��I;�jI;�NI;D:I;+I;1 I;	I;�I;�I;�I;	I;3 I;+I;G:I;�NI;�jI;��I;ھI;��I;��I;�I;��F;�FA;ͼ5;� ;8H�:�m:#�e�B��Ի|�>�������2�J̀�}n��bO��	�#�<�S�
ń��נ�*�����Ѿ��      �x���o��ń�LUo���O�,�-�{��hܽ]什ռx���2�rb��SR��P|U�K2��(���鰺�v�9�:CD;��,;�h<;�rD;�%H; �I;��I;�I;=�I;A�I;_I;?FI;�3I;�%I;I;�I;�I;nI;�I;�I;
I;�%I;�3I;@FI;_I;?�I;=�I;�I;��I;��I;~%H;�rD;�h<;��,;BD;�:w�9�鰺(��K2��P|U�SR��sb����2�ռx�]什�hܽ{�,�-���O�LUo�ń��o��      ��4�h1��&������k�ཆ�������`��'���SR��>�]�x��V���X���<o����:��;\#;L�6;�tA;��F;�	I;��I;�I;��I;O�I;qI;�SI;�=I;�,I;� I;�I;�I;zI;tI;{I;�I;�I;� I; -I;�=I;�SI;qI;P�I;��I;�I;��I;�	I;��F;�tA;L�6;^#;��;��:@=o��X��V��x��>�]�SR����'��`��������k��������&�h1�      m�ཹhܽq�н_y��`什Q ��l��n<�N���>ټ��O|U�x������a1�X�����u:�l�:8�;�71;�)>;�	E;DJH;��I;��I;��I;�I;�I;�bI;�HI;_5I;�&I;�I;�I;uI;YI;V
I;YI;uI;�I;�I;�&I;a5I;�HI;�bI;�I;�I;��I;��I;��I;AJH;�	E;�)>;�71;8�;�l�:��u:X���_1�����x��O|U��𛼿>ټN���n<�l�Q ��`什_y��q�н�hܽ      Z+����c̀�.l��Q�&�2�B��������@��|�>�K2��V��c1�P��$R:��:;�\,;p;; <C;�eG;�9I;��I;n�I;�I;x�I;�qI;�TI;�>I;p-I;d I;�I;�I;I;II;HI;II;I;�I;�I;h I;q-I;�>I;�TI;�qI;w�I;�I;l�I;��I;�9I;�eG;<C;q;;�\,;;��:�$R:P��c1�V��K2��|�>��@��������B�&�2��Q�.l�c̀���      �'��-$�_��Y����?ټw��9���hyY��k��Ի(���X��`����$R:��:�R;�);�8;��A;��F;k�H;a�I;��I;��I;�I;@�I;aI;,HI;�4I;�%I;~I;I;�I;�I;II;�I;JI;�I;�I;I;I;�%I;�4I;'HI;aI;=�I;�I;��I;��I;]�I;k�H;��F;��A;�8;�);�R;��:�$R:X����X��(���Ի�k�hyY�9���w��?ټ���Y�_���-$�      ��ü[l��s����R��<ߓ�[�{��M��� ��컹���`�B��鰺�<o���u:��:�R;a�';E17;�@;4�E;�lH;g�I;��I;��I;C�I;��I;mI;�QI;b<I;�+I;�I;�I;�I;I;|I;bI;�I;bI;|I;I;�I;�I;�I;�+I;`<I;�QI;�lI;��I;C�I;��I;��I;g�I;�lH;5�E;�@;H17;a�';�R;��:��u:@=o��鰺a�B������컄� ��M�Z�{�<ߓ��R��s���]l��      2yY��|U�B�I�9�7��� ��!���Ի�᝻h�T����#� w�9���:�l�:;�);E17;^ @;p]E;�$H;�kI;A�I;��I;0�I;g�I;�wI;�ZI;�CI;�1I;�#I;aI;�I;h	I;�I;oI;��H;7�H;��H;oI;�I;h	I;�I;aI;�#I;�1I;�CI;�ZI;�wI;g�I;,�I;��I;A�I;�kI;�$H;p]E;a @;B17;�);;�l�:���:�v�9#�Ĵ�j�T��᝻��Ի�!��� �9�7�B�I��|U�      �kٻS�Իtǻ�����V���n���+��ԺD�1���39�m:�:��;;�;�\,;�8;�@;p]E;�
H;�VI;��I;%�I;*�I;��I;=�I;�bI;�JI;^7I;(I;�I;iI;I;sI;pI;��H;�H;��H;�H;��H;pI;qI;I;iI;�I;(I;^7I;�JI;�bI;=�I;��I;$�I;%�I;��I;�VI;�
H;q]E;�@;�8;�\,;;�;��;�:m:��39D�1��Ժ��+��n��V������tǻS�Ի      �o&�:!��4����氺X�O��9T�v�9X�u:$�::H�:@D;\#;�71;l;;��A;1�E;�$H;�VI;G�I;��I;N�I;��I;5�I;IiI;ePI;Z<I;1,I;YI;�I;�I;�I;�I;i�H;
�H;��H;@�H;��H;
�H;j�H;�I;�I; I;�I;UI;1,I;W<I;dPI;JiI;1�I;��I;N�I;��I;I�I;�VI;�$H;1�E;��A;l;;�71;\#;@D;:H�:	$�:L�u:(v�9�9T�P�O�
氺���4�B!�      ��p� �,��$9�Ƴ9|�":H�u:��:���:`��:^R;� ;��,;J�6;�)>;<C;��F;�lH;�kI;��I;��I;��I;S�I;��I;�mI;�TI;d@I;�/I;]"I;�I;�I;I;�I;��H;��H;��H;��H;�H;��H;��H;��H;��H;�I;I;�I;�I;]"I;�/I;d@I;�TI;�mI;��I;S�I;��I;��I;��I;�kI;�lH;��F;<C;�)>;J�6;��,;� ;\R;`��:���:��:X�u:��":�Ƴ9�$9 �,�      ���:��:O�:@��:%��:$Q ;�e;�V;~#;>e-;м5;�h<;�tA;�	E;�eG;h�H;g�I;@�I;&�I;O�I;P�I;0�I;BpI;�WI;*CI;|2I;�$I;�I;�I;	I;�I;2�H;��H;;�H;��H;g�H;	�H;g�H;��H;;�H;��H;3�H;�I;{	I;�I;�I;�$I;~2I;,CI;�WI;>pI;0�I;O�I;P�I;%�I;C�I;d�I;f�H;�eG;�	E;�tA;�h<;ϼ5;=e-;~#;�V;�e;&Q ;O��:@��:O�:��:      �; ;y�;�;: ;&;�\,;�2;O98; 0=;�FA;�rD;��F;EJH;�9I;^�I;��I;��I;*�I;��I;��I;CpI;�XI;�DI;%4I;�&I;`I;$I;�
I;�I;��H;��H;$�H;�H;q�H;~�H;F�H;~�H;s�H;�H;#�H;��H;��H;�I;�
I;"I;\I;�&I;'4I;�DI;�XI;CpI;��I;��I;*�I;��I;��I;]�I;�9I;EJH;��F;�rD;�FA;�/=;N98;�2;�\,;&;@ ;�;{�;;      �0;�51;D�2;y�4;17;Q#:;*0=;� @;;�B;
E;��F;�%H;�	I;��I;��I;��I;��I;1�I;��I;3�I;�mI;�WI;�DI;�4I;|'I;oI;>I;�I;sI;l I;k�H;�H;��H;��H;��H;��H;��H;��H;��H;��H;��H;�H;k�H;i I;pI;�I;=I;nI;|'I;�4I;�DI;�WI;�mI;4�I;��I;4�I;��I;��I;��I;��I;�	I;�%H;��F;�	E;;�B;� @;'0=;Q#:;17;y�4;A�2;�51;      Ƕ?;��?;��@;�tA;:�B;y�C;�BE;��F;��G;�xH;�I;��I;��I;��I;n�I;��I;H�I;g�I;C�I;MiI;�TI;0CI;,4I;�'I;�I;�I;QI;I;� I;��H;Q�H;��H;��H;�H;��H;a�H;.�H;b�H;�H;�H;��H;��H;S�H;��H;� I;I;OI;�I;�I;}'I;)4I;/CI;�TI;PiI;C�I;j�I;F�I;��I;n�I;��I;��I;��I;�I;�xH;��G;��F;�BE;y�C;:�B;�tA;��@;��?;      �F;��F;�F;�2G;u�G;1&H;��H;I;*mI;��I;��I;��I;�I;��I;�I;�I;��I;�wI;�bI;bPI;a@I;|2I;�&I;nI;�I;}I;]I;<I;�H;��H;��H;��H;��H;c�H;��H;�H;��H;�H;��H;b�H;��H;��H;��H;��H;�H;=I;\I;}I;�I;lI;�&I;{2I;[@I;bPI;�bI;�wI;��I;�I;�I;��I;�I;��I;��I;��I;*mI;I;��H;1&H;x�G;�2G;	�F;��F;      � I;c'I;;I;�XI;|I;H�I;��I;)�I;D�I;C�I;��I;�I;��I;�I;x�I;?�I;mI;�ZI;�JI;[<I;�/I;�$I;`I;@I;MI;`I;DI;(�H;��H;��H;��H;��H;�H;��H;R�H;��H;��H;��H;P�H;��H;�H;��H;��H;��H;��H;*�H;CI;_I;QI;>I;]I;�$I;�/I;Z<I;�JI;�ZI;mI;=�I;x�I;�I;��I;�I;��I;B�I;E�I;*�I;��I;E�I;|I;�XI;;I;a'I;      '�I;��I;*�I;��I;�I;W�I;�I;y�I;8�I;��I;޾I;A�I;P�I;�I;�qI;aI;�QI;�CI;^7I;4,I;_"I;�I;'I;�I;I;?I;(�H;��H;��H;��H;��H;��H;��H;��H;�H;��H;��H;��H;�H;��H;��H;��H;��H;��H;��H;��H;(�H;?I;I;�I;%I;�I;\"I;5,I;^7I;�CI;�QI;aI;�qI;�I;O�I;A�I;ݾI;��I;8�I;}�I;�I;W�I;!�I;��I;)�I;��I;      �I;J�I;+�I;��I;��I;��I;��I;_�I;d�I;8�I;��I;C�I;qI;�bI;�TI;*HI;g<I;�1I;(I;ZI;�I;�I;�
I;vI;� I;�H;��H;��H;��H;��H;��H;��H;~�H;��H;$�H;��H;��H;��H;$�H;��H;{�H;��H;��H;��H;��H;��H;��H;�H;� I;wI;�
I;�I;�I;ZI;(I;�1I;e<I;*HI;�TI;�bI;qI;C�I;��I;6�I;f�I;_�I;��I;��I;��I;��I;+�I;>�I;      _�I;q�I;ϲI;:�I;�I;�I;�I;��I;��I;MvI;�jI;_I;�SI;�HI;�>I;�4I;�+I;�#I;�I;I;�I;~	I;�I;l I;��H;��H;��H;��H;��H;��H;j�H;Q�H;t�H;��H;M�H;
�H;��H;
�H;M�H;��H;q�H;R�H;k�H;��H;��H;��H;��H;��H;��H;l I;�I;~	I;�I;I;�I;�#I;�+I;�4I;�>I;�HI;�SI;_I;�jI;NvI;��I;��I;�I;�I;�I;;�I;ʲI;n�I;      ��I;�I;��I;4�I;z|I;�vI;�oI;8hI;`I;�WI;�NI;JFI;�=I;f5I;v-I;�%I;�I;bI;nI;I;I;�I;��H;n�H;N�H;��H;��H;��H;��H;m�H;J�H;M�H;��H;�H;��H;n�H;0�H;n�H;��H;�H;��H;N�H;J�H;k�H;��H;��H;��H;��H;Q�H;o�H;��H;�I;I;I;nI;bI;�I;�%I;v-I;e5I;�=I;HFI;�NI;�WI;`I;:hI;�oI;�vI;w|I;4�I;��I;�I;      �dI;dI;�bI;`I;r\I;
XI;�RI;JMI;=GI;�@I;J:I;�3I;-I;�&I;l I;�I;	I;�I;I;�I;�I;9�H;��H; �H;��H;��H;��H;��H;��H;Q�H;J�H;��H;��H;d�H;�H;��H;��H;��H;�H;d�H;��H;��H;L�H;R�H;��H;��H;��H;��H;��H; �H;��H;9�H;�I;�I;I;�I;I;�I;l I;�&I;-I;�3I;J:I;�@I;=GI;JMI;�RI;XI;p\I;`I;�bI;dI;      �KI;�KI;7JI;:HI;�EI;$BI;D>I;�9I;/5I;)0I;+I;�%I;� I;�I;�I;I;�I;e	I;xI;�I;��H;��H;&�H;��H;��H;��H;�H;��H;�H;w�H;��H;��H;N�H;��H;��H;Y�H;g�H;Y�H;��H;��H;K�H;��H;��H;x�H;��H;��H;�H;��H;��H;��H;$�H;��H;��H;�I;xI;f	I;�I;I;�I;�I;� I;�%I;+I;*0I;.5I;�9I;D>I;%BI;EI;:HI;7JI;yKI;      :I;�9I;�8I;a7I;X5I;�2I;�/I;*,I;a(I;[$I;8 I;I;�I;�I;�I;�I;&I;�I;xI;q�H;��H;=�H;	�H;��H;�H;b�H;��H;��H;��H;��H;�H;c�H;��H;w�H;5�H;�H;��H;�H;5�H;w�H;��H;e�H;�H;��H;��H;��H;��H;a�H;�H;��H;�H;=�H;��H;r�H;xI;�I;%I;�I;�I;�I;�I;I;7 I;[$I;b(I;-,I;�/I;�2I;N5I;a7I;�8I;�9I;      �.I;k.I;�-I;<,I;�*I;E(I;�%I;�"I;�I;yI;I;�I;�I;{I;I;�I;�I;mI;��H;�H;��H;��H;t�H;��H;��H;��H;O�H;�H;$�H;M�H;��H;�H;��H;6�H;��H;��H;��H;��H;��H;7�H;��H;�H;��H;O�H;'�H;�H;N�H;��H;��H;��H;s�H;��H;��H;�H;��H;oI;�I;�I;I;{I;�I;�I;I;zI;�I;�"I;�%I;H(I;x*I;<,I;�-I;c.I;      �'I;�'I;�&I;�%I;s$I;r"I;- I;�I;�I;�I;�I;�I;I;cI;OI;PI;kI;��H;&�H;��H;��H;j�H;��H;��H;_�H;�H;��H;��H;��H;�H;n�H;��H;V�H;�H;��H;��H;��H;��H;��H;�H;U�H;��H;n�H;
�H;��H;��H;��H;�H;a�H;��H;��H;j�H;��H;��H;&�H;��H;jI;PI;OI;aI;I;�I;�I;�I;�I;�I;- I;w"I;i$I;�%I;�&I;�'I;      �%I;�%I;%I;�#I;j"I;� I;zI;�I;GI;kI;�I;vI;wI;]
I;KI;�I;�I;0�H;��H;G�H;�H;�H;H�H;��H;+�H;��H;��H;��H;��H;��H;4�H;��H;i�H;��H;��H;��H;��H;��H;��H;��H;f�H;��H;4�H;��H;��H;��H;��H;��H;+�H;��H;H�H;�H;�H;G�H;��H;2�H;�I;�I;KI;]
I;wI;vI;�I;nI;GI;�I;zI;� I;_"I;�#I;%I;�%I;      �'I;�'I;�&I;�%I;s$I;q"I;- I;�I;�I;�I;�I;�I;I;cI;OI;PI;kI;��H;&�H;��H;��H;j�H;��H;��H;a�H;
�H;��H;��H;��H;�H;n�H;��H;V�H;�H;��H;��H;��H;��H;��H;�H;U�H;��H;n�H;
�H;��H;��H;��H;�H;_�H;��H;��H;j�H;��H;��H;&�H;��H;jI;PI;OI;aI;I;�I;�I;�I;�I;�I;- I;w"I;h$I;�%I;�&I;�'I;      �.I;m.I;�-I;;,I;�*I;E(I;�%I;�"I;�I;yI;I;�I;�I;{I;I;�I;�I;mI;��H;�H;��H;��H;t�H;��H;��H;��H;O�H;�H;&�H;M�H;��H;�H;��H;7�H;��H;��H;��H;��H;��H;6�H;��H;�H;��H;O�H;'�H;�H;N�H;��H;��H;��H;t�H;��H;��H;�H;��H;oI;�I;�I;I;{I;�I;�I;I;zI;�I;�"I;�%I;H(I;x*I;<,I;�-I;c.I;      :I;�9I;�8I;a7I;X5I;�2I;�/I;*,I;a(I;[$I;8 I;I;�I;�I;�I;�I;&I;�I;xI;q�H;��H;=�H;	�H;��H;�H;b�H;��H;��H;��H;��H;�H;c�H;��H;w�H;5�H;�H;��H;�H;5�H;w�H;��H;e�H;�H;��H;��H;��H;��H;b�H;�H;��H;�H;=�H;��H;q�H;xI;�I;%I;�I;�I;�I;�I;I;8 I;[$I;b(I;-,I;�/I;�2I;M5I;a7I;�8I;�9I;      �KI;�KI;9JI;;HI;�EI;"BI;D>I;�9I;/5I;)0I;+I;�%I;� I;�I;�I;I;�I;e	I;xI;�I;��H;��H;&�H;��H;��H;��H;�H;��H;�H;w�H;��H;��H;L�H;��H;��H;X�H;g�H;Y�H;��H;��H;K�H;��H;��H;x�H;��H;��H;�H;��H;��H;��H;$�H;��H;��H;�I;xI;e	I;�I;I;�I;�I;� I;�%I;+I;*0I;/5I;�9I;D>I;$BI;EI;;HI;6JI;KI;      �dI;dI;�bI;`I;r\I;
XI;�RI;JMI;=GI;�@I;J:I;�3I;-I;�&I;l I;�I;I;�I;I;�I;�I;9�H;��H; �H;��H;��H;��H;��H;��H;Q�H;L�H;��H;��H;d�H;�H;��H;��H;��H;�H;d�H;��H;��H;J�H;R�H;��H;��H;��H;��H;��H; �H;��H;9�H;�I;�I;I;�I;I;�I;l I;�&I;-I;�3I;J:I;�@I;>GI;JMI;�RI;XI;o\I;`I;�bI;dI;      ��I;�I;��I;4�I;y|I;�vI;�oI;8hI;`I;�WI;�NI;HFI;�=I;f5I;v-I;�%I;�I;bI;nI;I;I;�I;��H;o�H;Q�H;��H;��H;��H;��H;m�H;J�H;M�H;��H;�H;��H;n�H;0�H;n�H;��H;�H;��H;N�H;J�H;k�H;��H;��H;��H;��H;N�H;o�H;��H;�I;I;I;nI;bI;�I;�%I;v-I;h5I;�=I;JFI;�NI;�WI;`I;:hI;�oI;�vI;w|I;4�I;��I;�I;      W�I;q�I;ͲI;:�I;�I;�I;�I;��I;��I;MvI;�jI;_I;�SI;�HI;�>I;�4I;�+I;�#I;�I;I;�I;~	I;�I;l I;��H;��H;��H;��H;��H;��H;k�H;Q�H;s�H;��H;M�H;
�H;��H;
�H;M�H;��H;s�H;R�H;j�H;��H;��H;��H;��H;��H;��H;l I;�I;~	I;�I;I;�I;�#I;�+I;�4I;�>I;�HI;�SI;_I;�jI;KvI;��I;��I;�I;�I;�I;:�I;ͲI;r�I;      
�I;E�I;2�I;��I;��I;��I;��I;_�I;d�I;8�I;��I;C�I;qI;�bI;�TI;*HI;g<I;�1I;(I;\I;�I;�I;�
I;vI;� I;�H;��H;��H;��H;��H;��H;��H;|�H;��H;#�H;��H;��H;��H;$�H;��H;|�H;��H;��H;��H;��H;��H;��H;�H;� I;wI;�
I;�I;�I;ZI;(I;�1I;e<I;,HI;�TI;�bI;qI;C�I;��I;8�I;d�I;a�I;��I;��I;��I;��I;1�I;E�I;      '�I;��I;*�I;��I;�I;W�I;�I;z�I;8�I;��I;޾I;A�I;O�I;�I;�qI;aI;�QI;�CI;^7I;5,I;b"I;�I;'I;�I;I;?I;(�H;��H;��H;��H;��H;��H;��H;��H;�H;��H;��H;��H;�H;��H;��H;��H;��H;��H;��H;��H;(�H;?I;I;�I;%I;�I;\"I;5,I;^7I;�CI;�QI;aI;�qI;�I;P�I;B�I;ݾI;��I;8�I;|�I;�I;T�I;"�I;��I;)�I;��I;      � I;a'I;;I;�XI;|I;D�I;��I;)�I;E�I;C�I;��I;�I;��I;�I;x�I;?�I;mI;�ZI;�JI;[<I;�/I;�$I;`I;@I;QI;`I;DI;*�H;��H;��H;��H;��H;�H;��H;P�H;��H;��H;��H;R�H;��H;�H;��H;��H;��H;��H;(�H;CI;`I;MI;>I;]I;�$I;�/I;[<I;�JI;�ZI;mI;=�I;x�I; �I;��I;�I;��I;C�I;D�I;)�I;��I;B�I;|I;�XI;;I;X'I;      �F;��F;�F;�2G;u�G;3&H;��H;I;)mI;��I;��I;��I;�I;��I;�I;�I;��I;�wI;�bI;bPI;a@I;{2I;�&I;lI;�I;~I;]I;=I;�H;��H;��H;��H;��H;b�H;��H;�H;��H;�H;��H;c�H;��H;��H;��H;��H;�H;<I;\I;}I;�I;lI;�&I;|2I;]@I;bPI;�bI;�wI;��I;�I;�I;��I;�I;��I;��I;��I;)mI;I;��H;1&H;z�G;�2G;�F;��F;      Ƕ?;��?;��@;�tA;:�B;y�C;�BE;��F;��G;�xH;�I;��I;��I;��I;n�I;��I;G�I;i�I;C�I;NiI;�TI;/CI;*4I;�'I;�I;�I;PI;I;� I;��H;S�H;��H;��H;�H;��H;a�H;.�H;b�H;��H;�H;��H;��H;Q�H;��H;� I;I;PI;�I;�I;�'I;*4I;0CI;�TI;NiI;C�I;j�I;F�I;��I;n�I;��I;��I;��I;�I;�xH;��G;��F;�BE;x�C;8�B;�tA;��@;��?;      �0;�51;H�2;v�4;17;V#:;%0=;� @;=�B;
E;��F;�%H;�	I;��I;��I;��I;��I;1�I;��I;4�I;�mI;�WI;�DI;�4I;|'I;oI;>I;�I;sI;k I;k�H;�H;��H;��H;��H;��H;��H;��H;��H;��H;��H;�H;k�H;i I;qI;�I;=I;oI;|'I;�4I;�DI;�WI;�mI;4�I;��I;3�I;��I;��I;��I;��I;�	I;�%H;��F;�	E;=�B;� @;%0=;U#:;17;v�4;E�2;�51;      �;*;��;�;8 ;
&;�\,;�2;O98; 0=;�FA;�rD;��F;EJH;�9I;^�I;��I;��I;*�I;��I;��I;CpI;�XI;�DI;'4I;�&I;^I;"I;�
I;�I;��H;��H;$�H;�H;s�H;~�H;F�H;~�H;q�H;�H;#�H;��H;��H;�I;�
I;$I;]I;�&I;%4I;�DI;�XI;CpI;��I;��I;*�I;��I;��I;^�I;�9I;GJH;��F;�rD;�FA;�/=;N98;�2;�\,;&;> ;�;�;;      ���:��:O�:@��:%��:$Q ;�e;�V;~#;=e-;м5;�h<;�tA;�	E;�eG;h�H;e�I;A�I;%�I;O�I;R�I;0�I;BpI;�WI;,CI;~2I;�$I;�I;�I;	I;�I;3�H;��H;;�H;��H;g�H;	�H;g�H;��H;;�H;��H;2�H;�I;{	I;�I;�I;�$I;~2I;*CI;�WI;>pI;0�I;O�I;P�I;&�I;C�I;e�I;h�H;�eG;�	E;�tA;�h<;м5;>e-;~#;�V;�e;$Q ;Q��:@��:M�:��:      ��p� �,�0%9�Ƴ9|�":4�u:��:���:`��:\R;� ;��,;J�6;�)>;<C;��F;�lH;�kI;��I;��I;��I;S�I;��I;�mI;�TI;d@I;�/I;]"I;�I;�I;I;�I;��H;��H;��H;��H;�H;��H;��H;��H;��H;�I;I;�I;�I;]"I;�/I;d@I;�TI;�mI;��I;S�I;��I;��I;��I;�kI;�lH;��F;<C;�)>;J�6;��,;� ;\R;d��:���:��:P�u:��":�Ƴ9%9 �,�      �o&�8!��4����氺X�O��9T� v�9X�u:$�::H�:@D;\#;�71;l;;��A;1�E;�$H;�VI;G�I;��I;N�I;��I;5�I;JiI;ePI;X<I;1,I;YI; I; I;�I;�I;j�H;
�H;��H;@�H;��H;
�H;i�H;�I;�I;�I;�I;SI;1,I;V<I;dPI;IiI;1�I;��I;N�I;��I;I�I;�VI;�$H;1�E;��A;l;;�71;\#;?D;8H�:	$�:X�u:0v�9�9T�P�O�氺���4�C!�      �kٻS�Իtǻ�����V���n���+��ԺD�1���39m:�:��;;�;�\,;�8;�@;p]E;�
H;�VI;��I;%�I;*�I;��I;=�I;�bI;�JI;^7I;(I;�I;iI;I;sI;pI;��H;�H;��H;�H;��H;pI;qI;I;iI;�I;(I;^7I;�JI;�bI;=�I;��I;$�I;%�I;��I;�VI;�
H;q]E;�@;�8;�\,;;�;��;�:�m:��39D�1��Ժ��+��n��V������tǻS�Ի      2yY��|U�B�I�9�7��� ��!���Ի�᝻h�T�Ĵ�#��v�9���:�l�:;�);E17;` @;p]E;�$H;�kI;A�I;��I;0�I;g�I;�wI;�ZI;�CI;�1I;�#I;aI;�I;h	I;�I;oI;��H;7�H;��H;oI;�I;f	I;�I;aI;�#I;�1I;�CI;�ZI;�wI;g�I;,�I;��I;A�I;�kI;�$H;p]E;a @;D17;�);;�l�:���: w�9#����h�T��᝻��Ի�!��� �9�7�B�I��|U�      ��ü[l��s����R��<ߓ�[�{��M��� ��컺���`�B��鰺@=o���u:��:�R;d�';E17;�@;4�E;�lH;g�I;��I;��I;C�I;��I;mI;�QI;b<I;�+I;�I;�I;�I;I;|I;bI;�I;bI;|I;I;�I;�I;�I;�+I;`<I;�QI;�lI;��I;C�I;��I;��I;g�I;�lH;5�E;�@;H17;b�';�R;��:��u:�<o��鰺`�B������컄� ��M�Z�{�<ߓ��R��s���]l��      �'��-$�_��Y����?ټw��9���hyY��k��Ի(���X��`����$R:��:�R;�);�8;��A;��F;k�H;_�I;��I;��I;�I;@�I;aI;,HI;�4I;�%I;~I;I;�I;�I;II;�I;II;�I;�I;I;I;�%I;�4I;'HI;aI;=�I;�I;��I;��I;]�I;k�H;��F;��A;�8;�);�R;��:�$R:X����X��(���Ի�k�gyY�9���w��?ټ���Y�_���-$�      Z+����c̀�.l��Q�&�2�B��������@��|�>�K2��V��c1�P��$R:��:;�\,;p;;<C;�eG;�9I;��I;l�I;�I;x�I;�qI;�TI;�>I;q-I;e I;�I;�I;I;II;HI;II;I;�I;�I;g I;p-I;�>I;�TI;�qI;w�I;�I;n�I;��I;�9I;�eG;<C;q;;�\,;;��:�$R:P��c1�V��K2��|�>��@��������B�&�2��Q�.l�c̀���      m�ཹhܽq�н_y��`什Q ��l��n<�N���>ټ��P|U�x������`1�X�����u:�l�:8�;�71;�)>;�	E;EJH;��I;��I;��I;�I;�I;�bI;�HI;a5I;�&I;�I;�I;uI;YI;V
I;YI;uI;�I;�I;�&I;_5I;�HI;�bI;�I;�I;��I;��I;��I;@JH;�	E;�)>;�71;8�;�l�:��u:X���c1�����x��O|U��𛼿>ټN���n<�l�Q ��`什_y��q�н�hܽ      ��4�h1��&������k�ཆ�������`��'���SR��>�]�x��V���X���<o���:��;\#;J�6;�tA;��F;�	I;��I;�I;��I;P�I;qI;�SI;�=I;�,I;� I;�I;�I;zI;tI;zI;�I;�I;� I;�,I;�=I;�SI;qI;O�I;��I;�I;��I;�	I;��F;�tA;L�6;^#;��;��:@=o��X��V��x��>�]�SR����'��`��������k��������&�h1�      �x���o��ń�LUo���O�,�-�{��hܽ]什ռx���2�sb��SR��P|U�K2��(���鰺 w�9�:BD;��,;�h<;�rD;�%H;��I;��I;�I;=�I;A�I;_I;@FI;�3I;�%I;I;�I;�I;nI;�I;�I;I;�%I;�3I;?FI;_I;?�I;=�I;�I;��I; �I;~%H;�rD;�h<;��,;BD;�:w�9�鰺(��K2��P|U�SR��sb����2�ռx�]什�hܽ{�,�-���O�LUo�ń��o��      y���྅�Ѿ*����נ�
ń�<�S�	�#�bO��}n��J̀���2����|�>��Իd�B�#��m::H�:� ;ͼ5;�FA;��F;�I;��I;��I;ھI;��I;�jI;�NI;D:I;+I;3 I;	I;�I;�I;�I;	I;1 I;+I;D:I;�NI;�jI;��I;پI;��I;��I;�I;��F;�FA;̼5;� ;8H�:�m:#�e�B��Ի|�>�������2�J̀�}n��bO��	�#�<�S�
ń��נ�*�����Ѿ��      �3���/��X#��	��A��،Ⱦ�f��KUo�_1�Ͱ��}n��ռx��'��>ټ�@���k�����Ĵ��39$�:[R;=e-;�/=;
E;�xH;��I;F�I;��I;9�I;GvI;�WI;�@I;*0I;[$I;vI;�I;nI;�I;vI;Z$I;)0I;�@I;�WI;GvI;6�I;��I;C�I;��I;�xH;�	E;�/=;=e-;\R;	$�:��39��𺼼���k��@���>ټ�'�ռx�}n��Ͱ��_1�KUo��f��،Ⱦ�A���	��X#���/�      ���U���V�v��RZ�]58�ς�s��f���ioy�_1�bO��]什�`�N�����iyY���m�T�`�1�X�u:X��:x#;J98;8�B;��G;,mI;D�I;5�I;d�I;��I;`I;7GI;+5I;](I;�I;�I;CI;�I;�I;[(I;(5I;7GI;`I;��I;a�I;3�I;A�I;*mI;��G;4�B;G98;v#;^��:P�u:`�1�k�T���iyY����N���`�]什bO��_1�ioy�f���s��ς�]58��RZ�V�v�U���      Ŀ7g��(ﱿ���U����U��X#�v��f���KUo�	�#��hܽ����n<����9����� ��᝻�Ժ@v�9���:�V;�2;� @;��F;I;.�I;v�I;b�I;��I;7hI;DMI;�9I;&,I;�"I;�I;�I;�I;�"I;&,I;�9I;DMI;7hI;��I;_�I;v�I;-�I;I;��F;� @;�2;�V;���:(v�9�Ժ�᝻�� �9�������n<�����hܽ	�#�KUo�f���v���X#��U�U������(ﱿ7g��      x�Q9�T��uؿpQ��f_��8�_��X#�s���f��<�S�{�����l�B�w���M���Ի��+��9T���:�e;�\,;#0=;�BE;��H;��I;�I;��I;�I;�oI;�RI;H>I;�/I;�%I;' I;{I;' I;�%I;�/I;G>I;�RI;�oI;�I;��I;�I;��I;��H;�BE;0=;�\,;�e;��: :T���+���Ի�M�w��B�l�����{�<�S��f��s���X#�8�_�f_��pQ��uؿT��Q9�      �X1���,�i���<��7g��f_���U�ς�،Ⱦ
ń�,�-�k��R ��&�2�?ټ\�{��!��n�X�O�,�u:Q ;&;O#:;u�C;8&H;E�I;Y�I;�I;�I;�vI;
XI;%BI;�2I;I(I;w"I;� I;x"I;I(I;�2I;"BI;XI;�vI;�I;��I;Y�I;D�I;7&H;x�C;M#:;&;Q ;<�u:X�O��n��!�]�{�	?ټ&�2�R ��k��,�-�
ń�،Ⱦς��U�f_��7g��<�i����,�      d��]]�6K��X1�[f��pQ��U���]58��A���נ���O���a什�Q����<ߓ��� ��V��氺��":'��:@ ;17;<�B;w�G;|I;�I;��I;�I;p|I;o\I;EI;S5I;m*I;d$I;`"I;d$I;k*I;Q5I;~EI;o\I;p|I;�I;��I;�I;|I;u�G;<�B;17;D ;'��:��":氺�V���� �=ߓ�����Q�a什����O��נ��A��]58�U���pQ���[f��X1�6K��]]�      O������4z���V��X1��<�uؿ����RZ��	�*���LUo����_y��/l�Z��R��;�7� �������Ƴ9H��:�;x�4;�tA;�2G;�XI;��I;��I;:�I;+�I;�_I;0HI;Y7I;3,I;�%I;�#I;�%I;3,I;W7I;.HI;�_I;+�I;7�I;��I;��I;�XI;�2G;�tA;u�4;�;H��:�Ƴ9��� ���:�7��R��Z�/l�_y�����LUo�*����	��RZ����uؿ�<��X1���V��4z�����      �o��g^���ē��4z�6K�i��T��(ﱿV�v��X#���Ѿń�	�&�r�нd̀�`��s���D�I�{ǻ�4�0$9-�:u�;;�2;��@;�F;;I;&�I;2�I;ʲI;��I;�bI;2JI;�8I;�-I;�&I;%I;�&I;�-I;�8I;0JI;�bI;��I;ȲI;1�I;&�I;;I;�F;��@;7�2;v�;-�:`$9�4�{ǻC�I�t���`��d̀�r�н	�&�ń���Ѿ�X#�V�v�(ﱿT��i��6K��4z��ē�g^��      r'���X��g^�������]]���,�Q9�7g��U�����/����o��i1��hܽ���-$�^l���|U�V�ԻM!� �,���:;�51;��?;��F;a'I;��I;N�I;k�I;ՆI;dI;tKI;�9I;[.I;�'I;�%I;�'I;\.I;�9I;rKI;dI;ՆI;i�I;K�I;��I;`'I;��F;��?;�51;";��: �,�O!�V�Ի�|U�^l���-$����hܽi1��o���ྜ�/�U���7g��Q9���,��]]�����g^���X��      m����������Ѣ��1�j��5���	��ȿ(8����7�G�꾄S���7�3�L���)���Ƽ��\��ݻW+� Rɸ��:\x;��0;ؤ?;��F;,I;��I;�I; �I;Z�I;	iI;/OI;�<I;1I;�)I;�'I;�)I;1I;�<I;-OI;	iI;Z�I;��I;�I;��I;,I;��F;ؤ?;��0;_x;��:�QɸY+��ݻ��\���Ƽ�)�L��3��7��S��G�꾪�7�(8���ȿ��	��5�1�j�Ѣ����������      ��������B��^�����c�821�&X��ÿjڇ�t�3��s��7��~74�c�?ى���&�Nü$�X���ػZ�%���J���:�b;��0;��?;M�F;�2I;�I;z�I;�I;~�I;�hI;�NI;g<I;�0I;�)I;�'I;�)I;�0I;g<I;�NI;�hI;~�I;�I;w�I;�I;�2I;M�F;��?;��0;�b;��:��J�\�%���ػ#�X�Nü��&�?ى�c�~74��7���s�t�3�jڇ��ÿ&X�821���c�^����B�����      �����B����F��y�P���#�P�������x|��'�[D־�X��q�)� Խ�Ă�I<�7_��w-M���ʻ&��`*�8	��:�;:K2;Jv@;��F;�FI;��I;C�I;Y�I;6�I;gI;sMI;y;I;�/I;�(I;�&I;�(I;�/I;y;I;qMI;gI;6�I;U�I;A�I;��I;�FI;��F;Jv@;4K2;�;	��:`*�8)����ʻv-M�8_��J<��Ă� Խq�)��X��[D־�'��x|����P�����#�y�P�F�����B��      Ѣ��^���F���/]��5�O���,ݿ-8��sm_��K��t��Z�s�%>����:�o��3��۩���:�]T������)�9�f�:�<;�_4;ChA;P8G;�dI;9�I;i�I;��I;��I;adI;PKI;�9I;�.I;�'I;�%I;�'I;�.I;�9I;OKI;`dI;��I;��I;f�I;9�I;�dI;M8G;AhA;�_4;�<;�f�:()�9����]T����:��۩��3�:�o����%>�Z�s��t���K�sm_�-8���,ݿO���5��/]�F��^���      1�j���c�y�P��5���u��J���jڇ�Iv<�*���r���_S��������+T��� �)$���G#�����1����:��:o�;P7;��B;��G;�I;J�I;��I;��I;��I;�`I;~HI;�7I;�,I;=&I;5$I;=&I;�,I;�7I;}HI;�`I;��I;��I;��I;K�I;�I;��G;��B;L7;p�;��:��:
1�������G#�)$���� �+T���������_S�r��*���Iv<�jڇ�J���u�����5�y�P���c�      �5�821���#�O��u���ÿ�ҕ�Z������̾�X����0�3�1W����5��zܼ9��Q��9�s��T\� �n:/��:�%;��9;��C;!/H;F�I;G�I;?�I;��I;�{I;B\I;EI;�4I;b*I;L$I;N"I;L$I;b*I;�4I;EI;C\I;�{I;��I;;�I;H�I;E�I; /H;��C;��9;�%;1��:�n:�T\�9�s�Q��:���zܼ��5�1W��3佁�0��X����̾���Z��ҕ��ÿu��O����#�821�      ��	�&X�P����,ݿJ����ҕ��d��'�B��%���{�W����m���3�o��G��*���Q���ػڮ0�@�~�8�:��;i,;�=;tBE;ȬH;��I;��I;�I;�I;�tI;�VI;AI;�1I;�'I;�!I; I;�!I;�'I;�1I;AI;�VI;�tI;�I;}�I;��I;��I;ȬH;qBE;�=;i,;��;:�:@�~�ڮ0���ػ�Q��*���G�3�o�m������{�W�%���B�꾎'��d��ҕ�J����,ݿP���&X�      �ȿ�ÿ���-8��jڇ�Z��'�����n8��Z�s�.�&�Z�1j??��V�琼PG#�N7��(Tܺ�9dW�:��;RL2;|@;�F;4I;��I;��I;��I;u�I;�lI;QI;�<I;2.I;�$I;YI;~I;YI;�$I;2.I;�<I;QI;�lI;u�I;��I;��I;��I;4I;�F;z@;TL2;��;fW�:�9(TܺN7��PG#�琼�V�j??�1Z�.�&�Z�s�n8�������'�Z�jڇ�-8������ÿ      '8��jڇ��x|�sm_�Iv<����B��n8��'6~�q74��l��|���8nc�4���^����\��9�Z�8�=���n:���:&#;�8;��B;��G;�xI;��I;��I;��I;�I;ldI;�JI;�7I;O*I;o!I;�I;�I;�I;o!I;O*I;�7I;�JI;ldI;�I;��I;��I;��I;�xI;��G;��B;�8;&#;���:��n:8�=�Z��9���\��^��4��8nc�|����l��q74�'6~�n8��B�꾐��Iv<�sm_��x|�jڇ�      ��7�t�3��'��K�*�����̾%���Z�s�q74����#N��Ї|��)�9zܼ�Y��8 �y�������V9;��:N�;2-;A=;�E;:�H;��I;d�I;��I;ߥI;L{I;�[I;�CI;�2I;K&I;I;aI;�I;aI;I;K&I;�2I;�CI;�[I;N{I;ߥI;��I;b�I;��I;7�H;�E;?=;2-;R�;9��:�V9����z��8 ��Y��9zܼ�)�Ї|�#N�����q74�Z�s�%�����̾*����K��'�t�3�      G���s�[D־�t��r���X��{�W�.�&��l��#N���Ă�j�5�����{Q����A�4�ػ��G�h!/��f:fb�:�;��5;�9A;w�F;+I;
�I;�I;?�I;��I;coI;�RI;�<I;P-I;�!I;{I;6I;�I;7I;|I;�!I;N-I;�<I;�RI;coI;��I;@�I;
�I;�I;+I;s�F;�9A;��5;�;fb�:�f:\!/���G�4�ػ��A�{Q������j�5��Ă�#N���l��.�&�{�W��X��r���t��[D־�s�      �S���7���X��Z�s��_S���0����Z�|���χ|�j�5�j���ک�2�X�c �g􃻄3�� �9g��:�;0�,;�L<;�oD;?.H;��I;��I;��I;��I;��I;kcI;�II;6I; (I;I;�I;�I;�I;�I;�I;�I; (I;6I;�II;mcI;��I;��I;��I;��I;��I;<.H;�oD;�L<;2�,;�;g��:H�9�3��f�c �2�X��ک�j��j�5�χ|�|���Zཤ����0��_S�Z�s��X���7��      �7�~74�q�)�%>����3�m���08nc��)������ک�pa��Q�A����M���ȸv��:�;�#;��6;5hA;��F;�I;q�I;��I;H�I;��I;�uI;�WI;�@I;=/I;�"I;MI;6I;�I;�I;�I;6I;MI;�"I;>/I;�@I;�WI;�uI;��I;E�I;��I;o�I;�I;��F;6hA;��6;�#;�;z��: �ȸ�M�A����Q�pa��ک������)�8nc�0m���3����%>�q�)�~74�      3�c�Խ�������0W��2�o�i??�4��9zܼzQ��1�X��Q��6�������Ϲ<�n:�m�:@>;��0;�>;dE;�SH;}�I;�I;��I;u�I;��I;gI;XLI;�7I;�(I;BI;*I;�I;SI;vI;SI;�I;(I;BI;�(I;�7I;ZLI;gI;��I;t�I;��I; �I;z�I;�SH;dE;�>;��0;B>;�m�:8�n:��Ϲ����6���Q�1�X�zQ��8zܼ4��i??�3�o�0W���������Խc�      ~L��>ى��Ă�:�o�+T���5��G��V��^���Y����A�c �A����������J:�l�:f;P,;��:;=5C;DlG;EI;3�I;��I;��I;ƝI;�vI;�XI;zAI;�/I;D"I;I;�I;�I;1	I;�I;1	I;�I;�I;I;G"I;�/I;zAI;�XI;�vI;ŝI;��I;��I;/�I;EI;ElG;<5C;�:;P,;f;�l�:��J:�����B���c ���A��Y���^���V��G���5�+T�:�o��Ă�?ى�      �)���&�I<��3��� ��zܼ�*��琼��\�8 �2�ػf��M���Ϲ��J:�j�:��;��(;�e8;ΕA;D�F;�H;V�I;��I;9�I;1�I;��I;�eI;�KI;N7I;�'I;I;EI; I;�I;I;aI;I;�I; I;DI;I;�'I;O7I;�KI;�eI;��I;2�I;9�I;��I;R�I;�H;C�F;ΕA;�e8;��(;��;�j�:��J:��Ϲ�M�f�2�ػ8 ���\�琼�*���zܼ�� ��3�H<���&�      ��ƼNü6_���۩�)$��8���Q�NG#��9�w����G��3����ȸ8�n:�l�:��;H�';�7;�v@;W�E;GvH;*�I;��I;
�I;u�I;��I;�qI;�UI;g?I;.I;� I;HI;�I;	I;xI;!I;YI;!I;xI;	I;�I;HI;� I;.I;d?I;�UI;�qI;��I;u�I;�I;��I;*�I;GvH;Y�E;�v@;�7;H�';��;�l�:<�n:��ȸ�3����G�w���9�NG#��Q�8��)$���۩�6_��Nü      ��\�"�X�u-M���:��G#�R����ػN7��Z�����X!/� �9v��:�m�:f;��(;�7;�@;U]E;�-H;iwI;��I;��I; �I;��I;}I;
_I;GI;&4I;�%I;�I;I;
I;sI;XI;a I;��H;a I;VI;sI;|
I;I;�I;�%I;#4I;GI;_I;}I;��I;��I;��I;��I;fwI;�-H;U]E;�@;�7;��(;f;�m�:v��:0�9X!/�����Z�N7����ػQ���G#���:�v-M�$�X�      �ݻ��ػ��ʻ[T������1�s�Ѯ0�"Tܺ�=��V9�f:q��:�;C>;Q,;�e8;�v@;U]E;bH;8bI;F�I;��I;t�I;ʭI;��I;9gI;9NI;:I;"*I;�I;�I;1I;mI;=I;}�H;��H;��H;��H;}�H;<I;kI;3I;�I;�I; *I;:I;5NI;:gI;��I;ȭI;p�I;��I;C�I;9bI;bH;W]E;�v@;�e8;T,;C>;�;q��:�f:�V9�=�$TܺѮ0�-�s�����[T����ʻ��ػ      T+�E�%�%������
1���T\�@�~���9��n:;��:hb�:�;�#;��0;��:;ɕA;U�E;�-H;5bI;��I;��I;��I;<�I;�I;nI;7TI;A?I;k.I;#!I;�I;6I;�I;�I;2�H;��H;A�H;��H;B�H;��H;2�H;�I;�I;6I;�I;!I;m.I;>?I;7TI;nI;�I;9�I;��I;��I;��I;5bI;�-H;U�E;ɕA;��:;��0;�#;�;fb�:9��:��n:�90�~��T\��0������%��O�%�      �Pɸ �J�@+�8�(�9|�:�n:@�:dW�:���:R�;�;0�,;��6;�>;=5C;A�F;GvH;iwI;F�I;��I;l�I;��I;��I;�rI;�XI;oCI;$2I;a$I;I;&I;	I;yI;x�H;d�H;�H;��H;��H;��H;�H;d�H;v�H;yI;	I;%I;	I;b$I;"2I;oCI;�XI;�rI;��I;��I;i�I;��I;F�I;jwI;FvH;A�F;=5C;�>;��6;/�,;�;R�;���:dW�:>�: �n:��:�(�9 +�8@�J�      
�:E��:/��:�f�:���:E��:��;��;-#;2-;��5;�L<;5hA;cE;ElG;�H;*�I;��I;��I;��I;��I;'�I;(uI;�[I;�FI;�4I;�&I;jI;�I;�
I;�I;��H;F�H;��H;��H;��H;��H;��H;��H;��H;C�H;��H;�I;�
I;�I;kI;�&I;�4I;�FI;�[I;$uI;&�I;��I;��I;��I;��I;'�I;�H;GlG;cE;5hA;�L<;��5;2-;-#;��;��;K��:'��:�f�:/��:7��:      cx;�b;�;�<;f�;�%;m,;RL2;�8;B=;�9A;�oD;��F;�SH;EI;S�I;��I;��I;t�I;?�I;��I;+uI;�\I;�GI;�6I;�(I;I;xI;�I;�I;} I;��H;��H;:�H;��H;�H;��H;�H;��H;;�H;��H;��H;} I;�I;�I;yI;I;�(I;�6I;�GI;�\I;+uI;��I;@�I;t�I;��I;��I;R�I;EI;�SH;��F;�oD;�9A;A=;�8;RL2;m,;�%;o�;�<;�;�b;      ��0;��0;BK2;�_4;R7;��9;�=;z@;��B;�E;w�F;?.H;�I;}�I;3�I;��I;
�I;�I;̭I;�I;�rI;�[I;�GI;Y7I;�)I;7I;�I;�I;iI;&I;��H;��H;3�H;(�H;��H;=�H;��H;=�H;��H;*�H;2�H;��H;��H;$I;gI;�I;�I;7I;�)I;V7I;�GI;�[I;�rI;�I;̭I;�I;�I;��I;3�I;}�I;�I;?.H;v�F;�E;��B;|@;�=;��9;X7;�_4;@K2;��0;      �?;��?;8v@;GhA;��B;��C;pBE;�F;��G;6�H;+I;��I;n�I;�I;��I;9�I;z�I;��I;��I;nI;�XI;�FI;�6I;�)I;�I;I;pI;�I;�I;q�H;��H;�H;��H;c�H;M�H;��H;i�H;��H;M�H;a�H;��H;�H;��H;q�H;�I;�I;oI;I;�I;�)I;�6I;�FI;�XI;nI;��I;��I;v�I;7�I;��I;�I;m�I;��I;+I;5�H;��G;�F;pBE;��C;��B;FhA;6v@;��?;      ��F;a�F;��F;S8G;��G;/H;ƬH;-I;�xI;��I;	�I;��I;��I;��I;��I;1�I;��I;}I;6gI;5TI;mCI;�4I;�(I;5I;I;�I;nI;�I;��H;�H;4�H;��H;�H;��H;��H;0�H;'�H;0�H;��H;��H;�H;��H;4�H;�H;��H;�I;mI;�I;I;3I;�(I;�4I;hCI;5TI;7gI;}I;��I;/�I;��I;��I;��I;��I;	�I;��I;�xI;/I;ȬH;/H;��G;Q8G;��F;V�F;      #,I;�2I;�FI;�dI;�I;I�I;��I;��I;��I;d�I;�I;��I;E�I;u�I;ƝI;��I;�qI;_I;9NI;B?I;%2I;�&I;I;�I;lI;oI;'I;��H;K�H;9�H;��H;��H;q�H;Z�H;e�H;��H;��H;��H;d�H;X�H;p�H;��H;��H;9�H;K�H;��H;%I;oI;oI;�I;I;�&I;"2I;B?I;9NI;
_I;�qI;��I;ɝI;u�I;F�I;��I;�I;b�I;��I;��I;��I;E�I;�I;�dI;�FI;�2I;      ��I;�I;��I;6�I;I�I;E�I;��I;��I;��I;��I;E�I;��I;��I;��I;�vI;�eI;�UI;GI;:I;n.I;b$I;kI;{I;�I;�I;�I;��H;k�H;W�H;��H;��H;9�H;��H;��H;[�H;��H;��H;��H;[�H;��H;��H;9�H;��H;��H;V�H;m�H;��H;�I;�I;�I;yI;kI;`$I;n.I;:I;GI;�UI;�eI;�vI;��I;��I;��I;C�I;��I;��I;��I;��I;E�I;S�I;5�I;��I;(�I;      +�I;v�I;<�I;m�I;��I;9�I;~�I;��I;µI;ߥI;��I;��I;�uI;gI;�XI;�KI;k?I;#4I;$*I;!!I;I;�I;�I;mI;�I;��H;K�H;W�H;��H;��H;�H;��H;��H;��H;v�H;�H;��H;�H;t�H;��H;��H;��H;�H;��H;��H;V�H;M�H;��H;�I;kI;�I;�I;I;#!I;$*I;%4I;j?I;�KI;�XI;gI;�uI;��I;��I;ޥI;µI;��I;~�I;;�I;��I;m�I;<�I;i�I;      �I;!�I;\�I;��I;�I;��I;�I;w�I;�I;S{I;joI;vcI;�WI;bLI;~AI;R7I; .I;%I;�I;�I;)I;�
I;�I;'I;m�H;�H;:�H;��H;��H;$�H;��H;��H;��H;��H;]�H;0�H;0�H;0�H;]�H;��H;��H;��H;��H;#�H;��H;��H;7�H;�H;o�H;'I;�I;�
I;&I;�I;�I;�%I;.I;R7I;AI;aLI;�WI;xcI;hoI;S{I;�I;{�I; �I;��I;�I;��I;X�I;�I;      Z�I;��I;:�I;��I;ɁI;�{I;�tI;�lI;sdI;�[I;�RI;�II;�@I;8I;�/I;(I;� I;�I;�I;=I;#	I;�I;� I;��H;��H;7�H;��H;��H;�H;��H;x�H;t�H;��H; �H;��H;��H;h�H;��H;��H; �H;��H;v�H;x�H;��H;�H;��H;��H;6�H;��H;��H;| I;�I;	I;<I;�I;�I;� I;(I;�/I;8I;�@I;�II;�RI;�[I;rdI;�lI;�tI;�{I;ǁI;��I;:�I;��I;      iI;�hI;gI;hdI;�`I;A\I;�VI;	QI;�JI;�CI;�<I;6I;A/I;�(I;M"I;"I;TI;I;:I;�I;�I;��H;��H;��H;�H;��H;��H;;�H;��H;��H;q�H;��H;��H;q�H;%�H;��H;��H;��H;%�H;q�H;��H;��H;s�H;��H;��H;;�H;��H;��H;�H;��H;��H;��H;�I;�I;8I;I;RI;"I;M"I;�(I;A/I;6I;�<I;�CI;�JI;	QI;�VI;C\I;�`I;hdI;gI;�hI;      0OI;�NI;wMI;WKI;�HI;EI;AI;�<I;�7I;�2I;S-I;(I;�"I;FI; I;II;�I;z
I;qI;�I;��H;H�H;��H;7�H;��H;�H;t�H;��H;��H;��H;��H; �H;P�H; �H;��H;r�H;g�H;r�H;��H; �H;N�H;�H;��H;��H;��H;��H;q�H;�H;��H;9�H;��H;H�H;}�H;�I;qI;{
I;�I;II;I;FI;�"I;(I;S-I;�2I;�7I;�<I;AI;EI;|HI;WKI;wMI;�NI;      �<I;o<I;o;I;�9I;�7I;�4I;�1I;6.I;T*I;K&I;�!I;�I;PI;/I;�I;I;$	I;tI;DI;:�H;n�H;��H;=�H;.�H;`�H;��H;W�H;��H;��H;��H;�H;o�H;��H;��H;G�H;.�H;�H;.�H;H�H;��H;��H;r�H;�H;��H;��H;��H;W�H;��H;a�H;-�H;;�H;��H;k�H;9�H;DI;vI;!	I;I;�I;1I;PI;�I;�!I;K&I;U*I;9.I;�1I;�4I;�7I;�9I;q;I;h<I;      	1I;�0I;�/I;�.I;�,I;]*I;�'I;�$I;v!I;I;�I;�I;;I;�I;�I;�I;�I;UI;��H;��H;�H;��H;��H;�H;H�H;��H;c�H;[�H;v�H;]�H;��H;&�H;��H;K�H;��H;��H;��H;��H;��H;K�H;��H;)�H;��H;`�H;x�H;[�H;a�H;��H;H�H; �H;��H;��H;�H;��H;��H;VI;�I;�I;�I;�I;;I;�I;I;I;t!I;�$I;�'I;`*I;�,I;�.I;�/I;�0I;      �)I;�)I;�(I;�'I;M&I;H$I;�!I;aI;�I;cI;=I;�I;�I;^I;8	I;I;,I;] I;��H;H�H;��H;��H;�H;@�H;��H;.�H;��H;��H;�H;0�H;��H;��H;q�H;2�H;��H;��H;��H;��H;��H;/�H;p�H;��H;��H;0�H;�H;��H;��H;-�H;��H;@�H;�H;��H;��H;I�H;��H;^ I;*I;I;8	I;]I;�I;�I;<I;eI;�I;aI;�!I;L$I;C&I;�'I;�(I;�)I;      �'I;�'I;'I;�%I;>$I;M"I; I;�I;�I;�I;�I;�I;�I;I;�I;fI;bI;��H;��H;��H;��H;��H;��H;��H;h�H;%�H;��H;��H;��H;5�H;m�H;��H;i�H;	�H;��H;��H;��H;��H;��H;	�H;f�H;��H;m�H;7�H;��H;��H;��H;&�H;h�H;��H;��H;��H;��H;��H;��H;��H;`I;fI;�I;I;�I;�I;�I;�I;�I;�I; I;Q"I;3$I;�%I;'I;�'I;      �)I;�)I;�(I;�'I;M&I;H$I;�!I;aI;�I;bI;=I;�I;�I;^I;8	I;I;,I;] I;��H;H�H;��H;��H;�H;@�H;��H;.�H;��H;��H;�H;.�H;��H;��H;q�H;2�H;��H;��H;��H;��H;��H;/�H;p�H;��H;��H;1�H;�H;��H;��H;-�H;��H;@�H;�H;��H;��H;I�H;��H;^ I;*I;I;8	I;]I;�I;�I;=I;cI;�I;aI;�!I;L$I;C&I;�'I;�(I;�)I;      1I;�0I;�/I;�.I;�,I;\*I;�'I;�$I;t!I;I;I;�I;;I;�I;�I;�I;�I;UI;��H;��H;�H;��H;��H;�H;H�H;��H;c�H;[�H;w�H;]�H;��H;(�H;��H;K�H;��H;��H;��H;��H;��H;K�H;��H;*�H;��H;`�H;x�H;[�H;a�H;��H;H�H; �H;��H;��H;�H;��H;��H;VI;�I;�I;�I;�I;;I;�I;�I;I;v!I;�$I;�'I;b*I;�,I;�.I;�/I;�0I;      �<I;o<I;o;I;�9I;�7I;�4I;�1I;6.I;T*I;K&I;�!I;�I;PI;/I;�I;I;$	I;tI;DI;9�H;o�H;��H;;�H;.�H;a�H;��H;W�H;��H;��H;��H;�H;o�H;��H;��H;H�H;.�H;�H;.�H;G�H;��H;��H;r�H;�H;��H;��H;��H;W�H;��H;`�H;-�H;=�H;��H;l�H;:�H;DI;vI;!	I;I;�I;1I;PI;�I;�!I;K&I;U*I;9.I;�1I;�4I;�7I;�9I;q;I;h<I;      3OI;�NI;xMI;YKI;�HI;EI;AI;�<I;�7I;�2I;S-I;(I;�"I;FI;I;II;�I;z
I;qI;�I;��H;H�H;��H;9�H;��H;	�H;t�H;��H;��H;��H;��H; �H;O�H;��H;��H;r�H;g�H;r�H;��H;��H;N�H;�H;��H;��H;��H;��H;q�H;�H;��H;7�H;��H;H�H;�H;�I;qI;z
I;�I;II; I;GI;�"I;(I;Q-I;�2I;�7I;�<I;AI;EI;|HI;ZKI;vMI;�NI;      iI;�hI;gI;hdI;�`I;A\I;�VI;	QI;�JI;�CI;�<I;6I;A/I;�(I;M"I;"I;TI;I;8I;�I;�I;��H;��H;��H;�H;��H;��H;;�H;��H;��H;s�H;��H;��H;q�H;%�H;��H;��H;��H;%�H;q�H;��H;��H;q�H;��H;��H;;�H;��H;��H;�H;��H;��H;��H;�I;�I;:I;I;RI;"I;M"I;�(I;A/I;6I;�<I;�CI;�JI;	QI;�VI;B\I;�`I;hdI;gI;�hI;      Z�I;��I;:�I;��I;ɁI;�{I;�tI;�lI;sdI;�[I;�RI;�II;�@I;8I;�/I;(I;� I;�I;�I;:I;#	I;�I;~ I;��H;��H;7�H;��H;��H;�H;��H;x�H;t�H;��H; �H;��H;��H;h�H;��H;��H; �H;��H;v�H;x�H;��H;�H;��H;��H;6�H;��H;��H;} I;�I;	I;=I;�I;�I;� I;(I;�/I;8I;�@I;�II;�RI;�[I;rdI;�lI;�tI;�{I;ǁI;��I;:�I;��I;      �I;!�I;Z�I;��I;��I;��I;�I;w�I;�I;R{I;joI;vcI;�WI;bLI;~AI;R7I; .I;%I;�I;�I;*I;�
I;�I;&I;o�H;�H;9�H;��H;��H;$�H;��H;��H;��H;��H;]�H;0�H;0�H;0�H;]�H;��H;��H;��H;��H;#�H;��H;��H;9�H;�H;m�H;(I;�I;�
I;'I;�I;�I;�%I;.I;S7I;~AI;aLI;�WI;vcI;joI;S{I;�I;z�I; �I;��I;�I;��I;Z�I;"�I;      &�I;r�I;C�I;k�I;��I;7�I;�I;��I;��I;ޥI;��I;��I;�uI;gI;�XI;�KI;k?I;#4I;$*I;#!I;I;�I;�I;kI;�I;��H;J�H;V�H;��H;��H;�H;��H;��H;��H;s�H;�H;��H;�H;v�H;��H;��H;��H;�H;��H;��H;W�H;M�H;��H;�I;mI;�I;�I;I;#!I;$*I;%4I;j?I;�KI;�XI;gI;�uI;��I;��I;ޥI;µI;��I;��I;8�I;��I;i�I;A�I;r�I;      ��I;�I;��I;5�I;I�I;E�I;��I;��I;��I;��I;E�I;��I;��I;��I;�vI;�eI;�UI;GI;:I;n.I;e$I;kI;{I;�I;�I;�I;��H;m�H;V�H;��H;��H;9�H;��H;��H;Y�H;��H;��H;��H;[�H;��H;��H;;�H;��H;��H;V�H;k�H;��H;�I;�I;�I;yI;kI;`$I;n.I;:I;GI;�UI;�eI;�vI;��I;��I;��I;C�I;��I;��I;��I;��I;B�I;T�I;6�I;��I;(�I;      ,I;�2I;�FI;�dI;�I;D�I;��I;��I;��I;d�I;�I;��I;F�I;u�I;ȝI;��I;�qI;	_I;9NI;D?I;(2I;�&I;I;�I;oI;rI;'I;��H;M�H;:�H;��H;��H;p�H;X�H;d�H;��H;��H;��H;e�H;X�H;q�H;��H;��H;9�H;K�H;��H;%I;oI;lI;�I;I;�&I;!2I;B?I;9NI;	_I;�qI;��I;ƝI;u�I;E�I;��I;�I;d�I;��I;��I;��I;B�I;�I;�dI;�FI;�2I;      ��F;Z�F;��F;S8G;��G;/H;ȬH;/I;�xI;��I;	�I;��I;��I;��I;��I;1�I;��I;}I;7gI;5TI;nCI;�4I;�(I;5I;I;�I;mI;�I;��H;�H;4�H;��H;�H;��H;��H;0�H;'�H;0�H;��H;��H;�H;��H;4�H;�H;��H;�I;kI;�I;I;3I;�(I;�4I;gCI;5TI;6gI;}I;��I;1�I;��I;��I;��I;��I;	�I;��I;�xI;/I;ȬH;/H;��G;S8G;��F;Q�F;      �?;��?;8v@;FhA;��B;��C;pBE;�F;��G;6�H;+I;��I;m�I;�I;��I;9�I;w�I;��I;��I;nI;�XI;�FI;�6I;�)I;�I;I;pI;�I;�I;q�H;��H;�H;��H;a�H;K�H;��H;i�H;��H;M�H;a�H;��H;�H;��H;p�H;�I;�I;oI;I;�I;�)I;�6I;�FI;�XI;nI;��I;��I;w�I;9�I;��I;�I;n�I;��I;+I;5�H;��G;�F;pBE;��C;��B;GhA;6v@;��?;      ��0;��0;DK2;�_4;L7;��9;�=;{@;��B;�E;w�F;?.H;�I;}�I;3�I;��I;
�I;�I;̭I;�I;�rI;�[I;�GI;Y7I;�)I;7I;�I;�I;iI;&I;��H;��H;2�H;(�H;��H;=�H;��H;=�H;��H;(�H;2�H;��H;��H;#I;fI;�I;�I;7I;�)I;W7I;�GI;�[I;�rI;�I;̭I;�I;�I;��I;2�I;}�I;�I;?.H;v�F;�E;��B;{@;�=;��9;\7;�_4;DK2;��0;      ax;�b;�;�<;f�;�%;r,;RL2;�8;B=;�9A;�oD;��F;�SH;EI;S�I;��I;��I;t�I;?�I;��I;+uI;�\I;�GI;�6I;�(I;I;yI;�I;�I;} I;��H;��H;;�H;��H;�H;��H;�H;��H;:�H;��H;��H;} I;�I;�I;xI;I;�(I;�6I;�GI;�\I;+uI;��I;A�I;t�I;��I;��I;S�I;EI;�SH;��F;�oD;�9A;?=;�8;TL2;p,;�%;l�;�<;�;�b;      
�:C��:/��:�f�:���:G��:��;��;-#;2-;��5;�L<;5hA;cE;ElG;�H;)�I;��I;��I;��I;��I;&�I;(uI;�[I;�FI;�4I;�&I;kI;�I;�
I;�I;��H;E�H;��H;��H;��H;��H;��H;��H;��H;E�H;��H;�I;�
I;�I;jI;�&I;�4I;�FI;�[I;&uI;'�I;��I;��I;��I;��I;)�I;�H;GlG;cE;5hA;�L<;��5;2-;-#;��;��;E��:+��:�f�:+��:;��:      �Qɸ��J��+�8�(�9��:��n:B�:jW�:���:R�;�;/�,;��6;�>;<5C;A�F;GvH;iwI;F�I;��I;l�I;��I;��I;�rI;�XI;oCI;"2I;b$I;I;&I;	I;xI;v�H;b�H;�H;��H;��H;��H;�H;d�H;x�H;{I;	I;#I;	I;a$I;!2I;oCI;�XI;�rI;��I;��I;h�I;��I;F�I;jwI;FvH;A�F;<5C;�>;��6;/�,;�;N�;���:lW�:F�:�n:��:)�9�+�8@�J�      V+�D�%�������1���T\��~� �9��n:;��:hb�:�;�#;��0;��:;ɕA;U�E;�-H;5bI;��I;��I;��I;=�I;�I;nI;7TI;A?I;m.I;#!I;�I;6I;�I;�I;2�H;��H;B�H;��H;B�H;��H;2�H;�I;�I;6I;�I;!I;k.I;>?I;7TI;nI;�I;9�I;��I;��I;��I;5bI;�-H;U�E;ɕA;��:;��0;�#;�;fb�:9��:��n:�90�~��T\��0������#��O�%�      �ݻ��ػ��ʻ[T������1�s�Ѯ0�$Tܺ�=��V9�f:q��:�;C>;S,;�e8;�v@;W]E;bH;8bI;F�I;��I;t�I;ʭI;��I;9gI;7NI;:I;"*I;�I;�I;1I;kI;<I;}�H;��H;��H;��H;}�H;=I;kI;3I;�I;�I; *I;:I;5NI;:gI;��I;ƭI;p�I;��I;B�I;9bI;bH;X]E;�v@;�e8;S,;C>;�;q��:�f:�V9�=�$TܺѮ0�-�s�����[T����ʻ��ػ      ��\�!�X�u-M���:��G#�R����ػN7��Z�����X!/�0�9v��:�m�:f;��(;�7;�@;U]E;�-H;gwI;��I;��I; �I;��I;}I;
_I;GI;&4I;�%I;�I;I;|
I;sI;VI;a I;��H;a I;XI;sI;|
I;I;�I;�%I;#4I;GI;_I;}I;��I;��I;��I;��I;dwI;�-H;U]E;�@;�7;��(;f;�m�:v��: �9X!/�����Z�P7����ػQ���G#���:�u-M�#�X�      ��ƼNü6_���۩�)$��8���Q�NG#��9�w����G��3����ȸ<�n:�l�:��;J�';�7;�v@;W�E;GvH;*�I;��I;
�I;u�I;��I;�qI;�UI;g?I;.I;� I;HI;�I;	I;xI;!I;YI;!I;xI;	I;�I;JI;� I;.I;d?I;�UI;�qI;��I;u�I;�I;��I;*�I;FvH;Y�E;�v@;�7;H�';��;�l�:8�n:��ȸ�3����G�x���9�NG#��Q�8��)$���۩�6_��Nü      �)���&�I<��3��� ��zܼ�*��琼��\�8 �4�ػg��M���Ϲ��J:�j�:��;��(;�e8;ΕA;C�F;�H;U�I;��I;9�I;1�I;��I;�eI;�KI;N7I;�'I;I;EI; I;�I;I;aI;I;�I; I;DI;I;�'I;N7I;�KI;�eI;��I;2�I;:�I;��I;R�I;�H;A�F;ΕA;�e8;��(;��;�j�:��J:��Ϲ�M�f�2�ػ8 ���\�琼�*���zܼ�� ��3�H<���&�      ~L��>ى��Ă�:�o�+T���5��G��V��^���Y����A�c �A����������J:�l�:f;P,;��:;<5C;ElG;EI;3�I;��I;��I;ȝI;�vI;�XI;zAI;�/I;D"I;I;�I;�I;1	I;�I;1	I;�I;�I;I;F"I;�/I;xAI;�XI;�vI;ŝI;��I;��I;/�I;EI;DlG;<5C;�:;P,;f;�l�:��J:�����A���c ���A��Y���^���V��G���5�+T�:�o��Ă�?ى�      3�c�Խ�������0W��3�o�i??�4��9zܼzQ��1�X��Q��6�������Ϲ<�n:�m�:B>;��0;�>;dE;�SH;}�I; �I;��I;u�I;��I;gI;XLI;�7I;�(I;CI;*I;�I;SI;vI;SI;�I;(I;@I;�(I;�7I;XLI;gI;��I;t�I;��I;�I;y�I;�SH;dE;�>;��0;@>;�m�:8�n:��Ϲ����6���Q�1�X�zQ��8zܼ4��i??�2�o�0W���������Խc�      �7�~74�q�)�%>����3�m���08nc��)������ک�pa��Q�A����M���ȸx��:�;�#;��6;6hA;��F;�I;o�I;��I;H�I;��I;�uI;�WI;�@I;=/I;�"I;MI;6I;�I;�I;�I;6I;MI;�"I;;/I;�@I;�WI;�uI;��I;E�I;��I;q�I;�I;��F;5hA;��6;�#;�;z��: �ȸ�M�A����Q�pa��ک������)�8nc�0m���3����%>�q�)�~74�      �S���7���X��Z�s��_S���0����Z�|���χ|�j�5�j���ک�2�X�c �f􃻄3��8�9g��:�;.�,;�L<;�oD;?.H;��I;��I;��I;��I;��I;mcI;�II;6I;(I;�I;�I;�I;�I;�I;�I;I;�'I;6I;�II;kcI;��I;��I;��I;��I;��I;<.H;�oD;�L<;0�,;�;g��:H�9�3��h�c �2�X��ک�j��j�5�χ|�|���Zཤ����0��_S�Z�s��X���7��      G���s�[D־�t��r���X��{�W�.�&��l��#N���Ă�j�5�����{Q����A�4�ػ��G�\!/��f:hb�:�;��5;�9A;w�F;+I;�I;�I;@�I;��I;coI;�RI;�<I;P-I;�!I;|I;7I;�I;6I;{I;�!I;N-I;�<I;�RI;coI;��I;?�I;
�I;
�I;+I;s�F;�9A;��5;�;fb�:�f:X!/���G�6�ػ��A�{Q������j�5��Ă�#N���l��.�&�{�W��X��r���t��[D־�s�      ��7�t�3��'��K�*�����̾%���Z�s�q74����#N��Ї|��)�9zܼ�Y��8 �x�������V9;��:N�;2-;A=;�E;7�H;��I;d�I;��I;�I;L{I;�[I;�CI;�2I;K&I;I;bI;�I;aI;I;K&I;�2I;�CI;�[I;L{I;ܥI;��I;b�I;��I;:�H;�E;?=;2-;N�;9��:�V9����y��8 ��Y��9zܼ�)�Ї|�#N�����q74�Z�s�%�����̾*����K��'�t�3�      (8��jڇ��x|�sm_�Iv<����B��n8��'6~�q74��l��|���8nc�4���^����\��9�Z�8�=���n:���:&#;�8;��B;��G;�xI;��I;��I;ĵI;�I;ldI;�JI;�7I;O*I;o!I;�I;�I;�I;o!I;O*I;�7I;�JI;ldI;�I;��I;��I;��I;�xI;��G;��B;�8;&#;���:��n:8�=�Z��9���\��^��4��8nc�|����l��q74�'6~�n8��B�꾐��Iv<�sm_��x|�jڇ�      �ȿ�ÿ���-8��jڇ�Z��'�����n8��Z�s�.�&�Z�1j??��V�琼PG#�N7��(Tܺ�9bW�:��;TL2;|@;�F;4I;��I;��I;��I;u�I;�lI;QI;�<I;3.I;�$I;YI;~I;ZI;�$I;3.I;�<I;QI;�lI;u�I;��I;��I;��I;3I;�F;x@;RL2;��;fW�:�9(TܺN7��PG#�琼�V�j??�1Z�.�&�Z�s�n8�������'�Z�jڇ�-8������ÿ      ��	�&X�P����,ݿJ����ҕ��d��'�B��%���{�W����m���3�o��G��*���Q���ػڮ0�0�~�4�:��;k,;�=;qBE;ȬH;��I;��I;�I;�I;�tI;�VI;AI;�1I;�'I;�!I; I;�!I;�'I;�1I;AI;�VI;�tI;�I;~�I;��I;��I;ȬH;tBE;�=;h,;��;:�:P�~�ڮ0���ػ�Q��*���G�3�o�m������{�W�%���B�꾎'��d��ҕ�J����,ݿP���&X�      �5�821���#�O��u���ÿ�ҕ�Z������̾�X����0�3�1W����5��zܼ9��Q��9�s��T\���n:1��:�%;��9;��C;!/H;F�I;H�I;?�I;��I;�{I;B\I;	EI;�4I;b*I;L$I;N"I;M$I;b*I;�4I;EI;C\I;�{I;��I;;�I;G�I;E�I; /H;��C;��9;�%;/��:�n:�T\�9�s�P��:���zܼ��5�1W��3佁�0��X����̾���Z��ҕ��ÿu��O����#�821�      1�j���c�y�P��5���u��J���jڇ�Iv<�*���r���_S��������+T��� �)$���G#�����
1����:��:o�;P7;��B;��G;�I;K�I;��I;��I;��I;�`I;~HI;�7I;�,I;?&I;5$I;=&I;�,I;�7I;}HI;�`I;��I;��I;��I;J�I;�I;��G;��B;N7;p�;��:��:
1�������G#�*$���� �+T���������_S�r��*���Iv<�jڇ�J���u�����5�y�P���c�      Ѣ��^���F���/]��5�O���,ݿ-8��sm_��K��t��Z�s�%>����:�o��3��۩���:�]T������)�9�f�:�<;�_4;AhA;M8G;�dI;9�I;i�I;��I;��I;adI;PKI;�9I;�.I;�'I;�%I;�'I;�.I;�9I;OKI;^dI;��I;��I;f�I;9�I;�dI;P8G;ChA;�_4;�<;�f�:()�9����]T����:��۩��3�:�o����%>�Z�s��t���K�sm_�-8���,ݿO���5��/]�F��^���      �����B����F��y�P���#�P�������x|��'�[D־�X��q�)� Խ�Ă�J<�7_��v-M���ʻ)��@*�8	��:�;:K2;Jv@;��F;�FI;��I;C�I;X�I;6�I;gI;sMI;y;I;�/I;�(I;�&I;�(I;�/I;y;I;qMI;gI;6�I;V�I;A�I;��I;�FI;��F;Jv@;4K2;�;	��:`*�8(����ʻw-M�8_��J<��Ă� Խq�)��X��[D־�'��x|����P�����#�y�P�F�����B��      ��������B��^�����c�821�&X��ÿjڇ�t�3��s��7��~74�c�?ى���&�Nü$�X���ػZ�%���J���:�b;��0;��?;M�F;�2I;�I;z�I;�I;~�I;�hI;�NI;g<I;�0I;�)I;�'I;�)I;�0I;g<I;�NI;�hI;~�I;�I;w�I;�I;�2I;M�F;��?;��0;�b;��:��J�\�%���ػ#�X�Nü��&�?ى�c�~74��7���s�t�3�jڇ��ÿ&X�821���c�^����B�����      E(��s'���o��O�d��X1��x�Ŀ����3�z���x����4�o��[+���'���ü4yY��kٻ�o&���p����:y;��0;��?;	�F;� I;2�I;��I;W�I;��I;�dI;�KI;�9I;�.I;�'I;�%I;�'I;�.I;�9I;�KI;�dI;��I;W�I;��I;2�I;� I;	�F;��?;��0;|;���:@�p��o&��kٻ3yY���ü�'�[+��o�ཿ�4��x��z���3����Ŀ�x��X1�d�O��o��s'��      s'���X��f^�������]]���,�Q9�8g��V�����/����o��i1��hܽ���-$�^l���|U�X�ԻQ!� �,���:;�51;��?;��F;`'I;��I;K�I;i�I;ӆI;dI;rKI;�9I;X.I;�'I;�%I;�'I;Y.I;�9I;qKI;dI;ӆI;f�I;H�I;��I;`'I;��F;��?;�51;;��: �,�Q!�X�Ի�|U�_l���-$����hܽi1��o���ྛ�/�V���8g��Q9���,��]]�����f^���X��      �o��f^���ē��4z�6K�j��T��(ﱿX�v��X#���Ѿń��&�q�нd̀�`��u���H�I�~ǻ�4� $9+�:q�;:�2;��@;�F;;I;%�I;2�I;ɲI;��I;�bI;0JI;�8I;�-I;�&I;%I;�&I;�-I;�8I;0JI;�bI;��I;ƲI;/�I;%�I;;I;�F;��@;4�2;s�;+�:0$9�4�~ǻG�I�u���`��d̀�q�н�&�ń���Ѿ�X#�X�v�(ﱿT��j��6K��4z��ē�f^��      O������4z���V��X1��<�wؿ����RZ��	�*���LUo����`y��/l�Z��R��<�7��������Ƴ9F��:�;v�4;�tA;�2G;�XI;��I;��I;7�I;*�I;�_I;0HI;V7I;0,I;�%I;�#I;�%I;0,I;W7I;.HI;�_I;*�I;6�I;��I;��I;�XI;�2G;�tA;q�4;�;F��:�Ƴ9������<�7��R��Z�/l�`y�����LUo�*����	��RZ����wؿ�<��X1���V��4z�����      d��]]�6K��X1�[f��pQ��V���]58��A���נ���O���b什�Q�	���=ߓ��� ��V��"氺��":!��:< ;17;:�B;t�G;|I;�I;��I;�I;o|I;n\I;~EI;P5I;k*I;b$I;_"I;b$I;j*I;P5I;}EI;n\I;o|I;�I;��I;�I;|I;t�G;9�B;17;> ;%��:��":$氺�V���� �=ߓ�	����Q�b什����O��נ��A��]58�V���pQ���[f��X1�6K��]]�      �X1���,�i���<��7g��g_���U�ς�،Ⱦ
ń�,�-�l��Q ��'�2�	?ټ\�{��!��n�`�O�(�u:Q ;&;N#:;u�C;6&H;D�I;W�I; �I;�I;�vI;XI;"BI;�2I;H(I;w"I;� I;w"I;H(I;�2I;"BI;
XI;�vI;�I;��I;W�I;B�I;6&H;s�C;J#:;&;Q ;,�u:`�O��n��!�\�{�	?ټ'�2�Q ��l��,�-�
ń�،Ⱦς��U�g_��7g��<�i����,�      �x�Q9�T��wؿpQ��g_��8�_��X#�t���f��<�S�{�����l�C�w���M���Ի��+��9T���:�e;�\,; 0=;�BE;��H;��I;�I;��I;�I;�oI;�RI;F>I;�/I;�%I;) I;zI;) I;�%I;�/I;F>I;�RI;�oI;�I;��I;�I;��I;��H;�BE;0=;�\,;�e;��: :T���+���Ի�M�w��C�l�����{�<�S��f��t���X#�8�_�g_��pQ��wؿT��Q9�      Ŀ8g��(ﱿ���V����U��X#�v��f���KUo�	�#��hܽ����n<����:����� ��᝻��Ժ v�9���:�V;�2;� @;��F;I;-�I;u�I;a�I;��I;5hI;CMI;�9I;#,I;�"I;�I;�I;�I;�"I;#,I;�9I;DMI;5hI;��I;^�I;u�I;*�I;I;��F;� @;�2;�V;���:v�9��Ժ�᝻�� �:�������n<�����hܽ	�#�KUo�f���w���X#��U�V������(ﱿ8g��      ���V���W�v��RZ�]58�ς�t��f���ioy�`1�bO��^什�`�N�����jyY���q�T�p�1�H�u:V��:t#;H98;7�B;��G;*mI;B�I;3�I;c�I;��I;`I;7GI;(5I;[(I;�I;�I;BI;�I;�I;[(I;(5I;9GI;`I;��I;a�I;3�I;>�I;,mI;��G;3�B;H98;t#;\��:@�u:p�1�o�T���jyY����N���`�^什bO��`1�ioy�f���t��ς�]58��RZ�W�v�V���      �3���/��X#��	��A��،Ⱦ�f��KUo�`1�ΰ��~n��ռx��'��>ټ�@���k�����̴�`�39	$�:[R;:e-;�/=;�	E;�xH;��I;C�I;��I;8�I;FvI;�WI;�@I;)0I;Z$I;uI;�I;mI;�I;uI;Z$I;)0I;�@I;�WI;GvI;5�I;��I;B�I;��I;�xH;�	E;�/=;:e-;[R;$�:��39ʴ𺼼���k��@���>ټ�'�ռx�~n��Ͱ��`1�KUo��f��،Ⱦ�A���	��X#���/�      z���྅�Ѿ*����נ�
ń�<�S�	�#�bO��~n��K̀���2����}�>��Իh�B� #��m:2H�:� ;ɼ5;�FA;��F;�I;��I;��I;پI;��I;�jI;�NI;C:I;+I;1 I;I;�I;�I;�I;I;1 I;+I;F:I;�NI;�jI;��I;پI;��I;��I;�I;��F;�FA;˼5;� ;2H�:�m:#�h�B��Ի}�>�������2�K̀�~n��bO��	�#�<�S�
ń��נ�*�����Ѿ��      �x���o��ń�LUo���O�,�-�{��hܽ^什ռx���2�tb��TR��Q|U�N2��)���鰺�v�9�:BD;��,;�h<;�rD;%H;��I;��I;�I;;�I;?�I;_I;?FI;�3I;�%I;I;�I;�I;lI;�I;�I;I;�%I;�3I;?FI;_I;>�I;;�I;�I;��I;��I;|%H;�rD;�h<;��,;@D;�: w�9�鰺)��M2��Q|U�TR��sb����2�ռx�^什�hܽ{�,�-���O�LUo�ń��o��      ��4�i1��&������l�཈�������`��'���TR��?�]�y��V���X���=o����:��;\#;H�6;�tA;��F;�	I;��I;�I;��I;N�I;qI;�SI;�=I;�,I;� I;�I;�I;xI;tI;zI;�I;�I;� I;�,I;�=I;�SI;qI;N�I;��I;�I;��I;�	I;��F;�tA;H�6;\#;��;���:�=o��X��V��x��?�]�TR����'��`��������l��������&�i1�      n�ླྀhܽq�н_y��b什Q ��l��n<�N���>ټ��P|U�y������f1�x�����u:�l�:5�;�71;�)>;�	E;CJH;��I;��I;��I;�I;�I;�bI;�HI;^5I;�&I;�I;�I;tI;WI;U
I;WI;tI;�I;�I;�&I;a5I;�HI;�bI;�I;�I;��I;��I;��I;>JH;�	E;�)>;�71;7�;�l�:��u:p���c1�����x��P|U����>ټN���n<�l�P ��b什_y��p�н�hܽ      Z+����d̀�/l��Q�&�2�C��������@��}�>�M2��V��g1�`��$R:���:;�\,;l;;<C;�eG;�9I;��I;k�I;�I;w�I;�qI;�TI;�>I;o-I;b I;�I;�I;I;HI;GI;HI;I;�I;�I;e I;p-I;�>I;�TI;�qI;u�I;�I;k�I;��I;�9I;�eG;<C;n;;�\,;;���:�$R:`��f1�V��N2��|�>��@��������C�&�2��Q�/l�d̀���      �'��-$�_��Z����	?ټw��:���hyY��k��Ի)���X��x����$R:��:�R;�);�8;��A;��F;h�H;_�I;��I;��I;�I;?�I;aI;*HI;�4I;�%I;|I;I;�I;�I;II;|I;II;�I;�I;I;~I;�%I;�4I;&HI;aI;<�I;�I;��I;��I;[�I;i�H;��F;��A;�8;�);�R;��:�$R:p����X��(���Ի�k�hyY�:���w��?ټ���Z�_���-$�      ��ü\l��t����R��=ߓ�Z�{��M��� ��컹���c�B��鰺�=o���u:��:�R;`�';D17;�@;4�E;�lH;e�I;��I;��I;A�I;��I;mI;�QI;a<I;�+I;�I;�I;�I;I;zI;`I;�I;`I;zI;I;�I;�I;�I;�+I;^<I;�QI;�lI;��I;A�I;��I;��I;e�I;�lH;5�E;�@;F17;`�';�R;��:��u:�=o��鰺e�B������컅� ��M�Z�{�=ߓ��R��t���^l��      3yY��|U�E�I�:�7��� ��!���Ի�᝻m�T�ʴ�#��v�9���:�l�:;�);B17;] @;m]E;�$H;�kI;@�I;��I;/�I;f�I;�wI;�ZI;�CI;�1I;�#I;`I;�I;f	I;�I;mI;��H;7�H;��H;mI;�I;e	I;�I;`I;�#I;�1I;�CI;�ZI;�wI;f�I;*�I;��I;@�I;�kI;�$H;m]E;^ @;A17;�);;�l�:���:�v�9#�ʴ�m�T��᝻��Ի�!��� �:�7�E�I��|U�      �kٻU�Իvǻ ����V���n���+��ԺH�1���39�m:�:��;9�;�\,;�8;�@;p]E;�
H;�VI;��I;#�I;)�I;��I;<�I;�bI;�JI;]7I;(I;�I;fI;I;qI;oI;��H;�H;��H;�H;��H;oI;pI;I;gI;�I;
(I;]7I;�JI;�bI;<�I;��I;#�I;#�I;��I;�VI;�
H;q]E;�@;�8;�\,;9�;��;�:�m:��39H�1��Ժ��+��n��V�� ���vǻV�Ի      �o&�<!��4����$氺`�O� :T�v�9H�u:	$�:6H�:@D;Z#;�71;l;;��A;1�E;�$H;�VI;F�I;��I;K�I;��I;4�I;FiI;dPI;W<I;0,I;WI;�I;�I;�I;�I;g�H;
�H;��H;?�H;��H;
�H;g�H;�I;�I;�I;�I;SI;0,I;T<I;bPI;FiI;.�I;��I;K�I;��I;G�I;�VI;�$H;1�E;��A;l;;�71;Z#;?D;6H�:$�:@�u:v�9 :T�X�O�氺���4�F!�      ��p� �,��$9�Ƴ9p�":<�u:��:���:\��:\R;� ;��,;H�6;�)>;<C;��F;�lH;�kI;��I;��I;��I;R�I;��I;�mI;�TI;a@I;�/I;]"I;�I;�I;
I;�I;��H;��H;��H;��H;�H;��H;��H;��H;��H;�I;
I;�I;�I;\"I;�/I;a@I;�TI;�mI;��I;R�I;��I;��I;��I;�kI;�lH;��F;<C;�)>;H�6;��,;� ;[R;^��:���:��:H�u:t�":�Ƴ9�$9 �,�      ���:��:I�::��:��:"Q ;�e;�V;z#;:e-;ͼ5;�h<;�tA;�	E;�eG;f�H;e�I;A�I;#�I;K�I;O�I;/�I;?pI;�WI;)CI;|2I;�$I;�I;�I;~	I;�I;2�H;��H;9�H;��H;f�H;�H;f�H;��H;9�H;��H;0�H;�I;z	I;�I;�I;�$I;|2I;*CI;WI;<pI;/�I;N�I;N�I;#�I;C�I;d�I;e�H;�eG;�	E;�tA;�h<;̼5;:e-;z#;�V;�e;&Q ;E��::��:I�:��:      �;;v�;�;6 ;&;�\,;�2;N98;�/=;�FA;�rD;��F;DJH;�9I;^�I;��I;��I;)�I;��I;��I;BpI;�XI;�DI;%4I;�&I;^I;"I;�
I;�I;��H;��H;&�H;�H;q�H;~�H;E�H;}�H;q�H;�H;#�H;��H;��H;�I;�
I;!I;ZI;�&I;%4I;�DI;�XI;BpI;��I;��I;)�I;��I;��I;[�I;�9I;DJH;��F;�rD;�FA;�/=;M98;�2;�\,;&;@ ;�;x�;;      �0;�51;A�2;{�4;17;N#:;'0=;� @;;�B;�	E;��F;%H;�	I;��I;��I;��I;��I;0�I;��I;1�I;�mI;�WI;�DI;�4I;{'I;nI;=I;�I;qI;k I;i�H;�H;��H;��H;��H;��H;��H;��H;��H;��H;��H;�H;k�H;h I;pI;�I;;I;lI;|'I;�4I;�DI;�WI;�mI;3�I;��I;1�I;��I;��I;��I;��I;�	I;%H;��F;�	E;:�B;� @;&0=;O#:;17;y�4;@�2;�51;      ƶ?;��?;��@;�tA;9�B;v�C;�BE;��F;��G;�xH;�I;��I;��I;��I;l�I;��I;G�I;f�I;C�I;LiI;�TI;-CI;*4I;�'I;�I;�I;PI;I;� I;��H;Q�H;��H;��H;�H;�H;a�H;.�H;a�H;�H;�H;��H;��H;S�H;��H;� I;I;OI;�I;�I;}'I;'4I;-CI;�TI;LiI;B�I;i�I;D�I;��I;l�I;��I;��I;��I;�I;�xH;��G;��F;�BE;u�C;:�B;�tA;��@;��?;      �F;��F;�F;�2G;q�G;0&H;��H;
I;,mI;��I;��I;��I;�I;��I;��I;�I;��I;�wI;�bI;bPI;`@I;{2I;�&I;lI;�I;|I;\I;;I;�H;��H;��H;��H;��H;a�H;��H;�H;��H;�H;��H;b�H;��H;��H;��H;��H;�H;<I;[I;|I;�I;kI;�&I;{2I;[@I;aPI;�bI;�wI;��I;ߩI;��I;��I;�I;��I;��I;��I;*mI;I;��H;0&H;w�G;�2G;�F;��F;      � I;a'I;;I;�XI;|I;H�I;��I;'�I;D�I;C�I;��I;�I;��I;�I;w�I;=�I;mI;�ZI;�JI;Z<I;�/I;�$I;^I;@I;LI;]I;CI;'�H;��H;��H;��H;��H;�H;��H;P�H;��H;��H;��H;O�H;��H;�H;��H;��H;��H;��H;(�H;BI;\I;PI;>I;\I;�$I;�/I;Z<I;�JI;�ZI;mI;<�I;w�I;�I;��I;�I;��I;B�I;E�I;)�I;��I;E�I;|I;�XI;;I;_'I;      $�I;��I;*�I;��I;�I;V�I;�I;y�I;6�I;��I;ݾI;?�I;O�I;�I;�qI;aI;�QI;�CI;^7I;3,I;]"I;�I;%I;�I;I;=I;'�H;��H;��H;��H;��H;��H;��H;��H;�H;��H;��H;��H;�H;��H;��H;��H;��H;��H;��H;��H;'�H;=I;I;�I;"I;�I;["I;4,I;^7I;�CI;�QI;aI;�qI;�I;N�I;?�I;۾I;��I;6�I;|�I;�I;V�I;�I;��I;)�I;��I;      �I;J�I;+�I;��I;��I;��I;��I;^�I;d�I;8�I;��I;B�I;qI;�bI;�TI;*HI;e<I;�1I;(I;YI;�I;�I;�
I;tI;� I;�H;��H;��H;��H;��H;��H;��H;{�H;��H;#�H;��H;��H;��H;#�H;��H;z�H;��H;��H;��H;��H;��H;��H;�H;� I;vI;�
I;�I;�I;YI;(I;�1I;d<I;*HI;�TI;�bI;qI;A�I;��I;6�I;d�I;^�I;��I;��I;��I;��I;*�I;<�I;      a�I;p�I;ϲI;:�I;�I;�I;�I;��I;��I;MvI;�jI;_I;�SI;�HI;�>I;�4I;�+I;�#I;�I;I;�I;}	I;�I;k I;��H;��H;��H;��H;��H;��H;h�H;N�H;q�H;��H;L�H;�H;��H;�H;L�H;��H;p�H;O�H;h�H;��H;��H;��H;��H;�H;��H;k I;�I;}	I;�I;I;�I;�#I;�+I;�4I;�>I;�HI;�SI;_I;�jI;MvI;��I;��I;�I;�I;�I;9�I;ɲI;m�I;      ��I;�I;��I;5�I;y|I;�vI;�oI;8hI;`I;�WI;�NI;HFI;�=I;h5I;v-I;�%I;�I;aI;mI;I;I;�I;��H;l�H;M�H;��H;��H;��H;��H;m�H;J�H;M�H;��H;�H;��H;m�H;/�H;m�H;��H;�H;��H;M�H;H�H;j�H;��H;��H;��H;��H;P�H;l�H;��H;�I;I;I;mI;bI;�I;�%I;v-I;e5I;�=I;GFI;�NI;�WI;`I;:hI;�oI;�vI;v|I;4�I;��I;�I;      �dI;dI;�bI; `I;o\I;XI;�RI;IMI;;GI;�@I;H:I;�3I;-I;�&I;l I;�I;I;�I;I;�I;�I;6�H;��H;�H;��H;��H;��H;��H;��H;Q�H;J�H;��H;��H;d�H;�H;��H;��H;��H;�H;c�H;��H;��H;J�H;R�H;��H;��H;��H;��H;��H;�H;��H;7�H;�I;�I;I;�I;I;�I;k I;�&I;-I;�3I;H:I;�@I;;GI;IMI;�RI;XI;n\I; `I;�bI;dI;      �KI;�KI;7JI;8HI;�EI;!BI;C>I;�9I;.5I;'0I;+I;�%I;� I;�I;�I;I;�I;b	I;vI;�I;��H;��H;$�H;��H;��H;��H;�H;��H;�H;w�H;��H;��H;O�H;��H;��H;Y�H;i�H;X�H;��H;��H;L�H;��H;��H;x�H;��H;��H;�H;��H;��H;��H;#�H;��H;��H;�I;vI;c	I;�I;I;�I;�I;� I;�%I;+I;)0I;-5I;�9I;C>I;$BI;~EI;8HI;7JI;xKI;      :I;�9I;�8I;`7I;W5I;�2I;�/I;*,I;`(I;[$I;7 I;I;�I;�I;�I;�I;&I;�I;wI;p�H;��H;<�H;�H;��H;
�H;a�H;��H;��H;��H;��H;�H;c�H;��H;w�H;2�H;�H;��H;�H;2�H;w�H;��H;e�H;�H;��H;��H;��H;��H;^�H;�H;��H;�H;<�H;��H;p�H;wI;�I;%I;�I;�I;�I;�I;I;5 I;[$I;b(I;,,I;�/I;�2I;M5I;`7I;�8I;�9I;      �.I;j.I;�-I;:,I;*I;C(I;�%I;�"I;�I;wI;I;�I;�I;{I;I;�I;�I;lI;��H;�H;��H;��H;s�H;��H;��H;��H;O�H;�H;$�H;M�H;��H;�H;��H;7�H;��H;��H;��H;��H;��H;6�H;��H;�H;��H;P�H;'�H;�H;N�H;��H;��H;��H;q�H;��H;��H;�H;��H;mI;�I;�I;I;|I;�I;�I;I;yI;�I;�"I;�%I;F(I;w*I;:,I;�-I;b.I;      �'I;�'I;�&I;�%I;r$I;q"I;, I;�I;�I;�I;�I;�I;~I;cI;OI;PI;kI;��H;#�H;��H;��H;i�H;��H;��H;^�H;�H;��H;��H;��H;�H;n�H;��H;V�H;�H;��H;��H;��H;��H;��H;�H;V�H;��H;n�H;
�H;��H;��H;��H;�H;_�H;��H;��H;i�H;��H;��H;#�H;��H;jI;PI;OI;aI;~I;�I;�I;�I;�I;�I;, I;u"I;h$I;�%I;�&I;�'I;      �%I;�%I;%I;�#I;g"I;� I;xI;�I;FI;jI;�I;sI;vI;\
I;II;�I;�I;0�H;��H;F�H;�H;�H;F�H;��H;*�H;��H;��H;��H;��H;��H;4�H;��H;i�H;��H;��H;��H;��H;��H;��H;��H;g�H;��H;4�H;��H;��H;��H;��H;��H;*�H;��H;F�H;�H;
�H;F�H;��H;2�H;�I;�I;II;\
I;vI;sI;�I;mI;GI;�I;xI;� I;]"I;�#I;%I;�%I;      �'I;�'I;�&I;�%I;r$I;q"I;, I;�I;�I;�I;�I;�I;~I;cI;OI;PI;kI;��H;#�H;��H;��H;i�H;��H;��H;_�H;�H;��H;��H;��H;�H;n�H;��H;V�H;�H;��H;��H;��H;��H;��H;�H;V�H;��H;n�H;
�H;��H;��H;��H;�H;^�H;��H;��H;i�H;��H;��H;#�H;��H;jI;PI;OI;aI;~I;�I;�I;�I;�I;�I;, I;u"I;h$I;�%I;�&I;�'I;      �.I;j.I;�-I;:,I;*I;C(I;�%I;�"I;�I;wI;I;�I;�I;{I;I;�I;�I;lI;��H;�H;��H;��H;s�H;��H;��H;��H;O�H;�H;&�H;M�H;��H;�H;��H;6�H;��H;��H;��H;��H;��H;7�H;��H;�H;��H;O�H;'�H;�H;N�H;��H;��H;��H;q�H;��H;��H;�H;��H;mI;�I;�I;I;|I;�I;�I;I;yI;�I;�"I;�%I;H(I;w*I;:,I;�-I;b.I;      :I;�9I;�8I;`7I;U5I;�2I;�/I;*,I;a(I;[$I;7 I;I;�I;�I;�I;�I;&I;�I;wI;p�H;��H;<�H;�H;��H;�H;a�H;��H;��H;��H;��H;�H;c�H;��H;w�H;2�H;�H;��H;�H;2�H;w�H;��H;e�H;�H;��H;��H;��H;��H;a�H;
�H;��H;�H;<�H;��H;p�H;wI;�I;%I;�I;�I;�I;�I;I;7 I;[$I;b(I;,,I;�/I;�2I;L5I;`7I;�8I;�9I;      �KI;�KI;9JI;;HI;�EI;!BI;C>I;�9I;.5I;'0I;+I;�%I;� I;�I;�I;I;�I;c	I;vI;�I;��H;��H;$�H;��H;��H;��H;�H;��H;�H;w�H;��H;��H;N�H;��H;��H;X�H;i�H;Y�H;��H;��H;L�H;��H;��H;x�H;��H;��H;�H;��H;��H;��H;#�H;��H;��H;�I;vI;b	I;�I;I;�I;�I;� I;�%I;+I;)0I;.5I;�9I;C>I;"BI;~EI;:HI;6JI;}KI;      �dI;dI;�bI;�_I;p\I;XI;�RI;IMI;;GI;�@I;H:I;�3I;-I;�&I;k I;�I;I;�I;I;�I;�I;7�H;��H;�H;��H;��H;��H;��H;��H;Q�H;J�H;��H;��H;c�H;�H;��H;��H;��H;�H;d�H;��H;��H;J�H;R�H;��H;��H;��H;��H;��H;�H;��H;6�H;�I;�I;I;�I;I;�I;l I;�&I;-I;�3I;H:I;�@I;=GI;IMI;�RI;
XI;n\I;�_I;�bI;dI;      ��I;�I;��I;4�I;y|I;�vI;�oI;8hI;`I;�WI;�NI;GFI;�=I;f5I;v-I;�%I;�I;aI;mI;I;I;�I;��H;n�H;P�H;��H;��H;��H;��H;k�H;H�H;L�H;��H;�H;��H;m�H;/�H;m�H;��H;�H;��H;M�H;J�H;k�H;��H;��H;��H;��H;M�H;n�H;��H;�I;I;I;mI;bI;�I;�%I;v-I;i5I;�=I;HFI;�NI;�WI;`I;:hI;�oI;�vI;w|I;5�I;��I;�I;      Z�I;n�I;ͲI;9�I;�I;�I;�I;��I;��I;KvI;�jI;_I;�SI;�HI;�>I;�4I;�+I;�#I;�I;I;�I;}	I;�I;k I;��H;��H;��H;��H;��H;��H;h�H;N�H;q�H;��H;L�H;�H;��H;�H;L�H;��H;q�H;O�H;h�H;��H;��H;��H;��H;�H;��H;k I;�I;}	I;�I;I;�I;�#I;�+I;�4I;�>I;�HI;�SI;_I;�jI;MvI;��I;��I;�I;�I;�I;9�I;ͲI;q�I;      �I;E�I;/�I;��I;��I;��I;��I;^�I;d�I;6�I;��I;B�I;qI;�bI;�TI;*HI;e<I;�1I;(I;ZI;�I;�I;�
I;tI;� I;�H;��H;��H;��H;��H;��H;��H;z�H;��H;!�H;��H;��H;��H;#�H;��H;z�H;��H;��H;��H;��H;��H;��H;�H;� I;vI;�
I;�I;�I;YI;(I;�1I;d<I;,HI;�TI;�bI;qI;B�I;��I;8�I;d�I;a�I;��I;��I;��I;��I;/�I;E�I;      $�I;��I;*�I;��I;�I;V�I;�I;y�I;8�I;��I;ݾI;?�I;N�I;�I;�qI;aI;�QI;�CI;^7I;4,I;`"I;�I;%I;�I;I;=I;'�H;��H;��H;��H;��H;��H;��H;��H;�H;��H;��H;��H;�H;��H;��H;��H;��H;��H;��H;��H;'�H;=I;I;�I;"I;�I;["I;4,I;^7I;�CI;�QI;aI;�qI;�I;O�I;?�I;۾I;��I;8�I;|�I;�I;S�I;"�I;��I;)�I;��I;      � I;`'I;;I;�XI;|I;D�I;��I;'�I;D�I;C�I;��I;�I;��I;�I;w�I;=�I;mI;�ZI;�JI;[<I;�/I;�$I;^I;>I;PI;_I;CI;(�H;��H;��H;��H;��H;�H;��H;O�H;��H;��H;��H;P�H;��H;�H;��H;��H;��H;��H;'�H;BI;]I;LI;=I;\I;�$I;�/I;Z<I;�JI;�ZI;mI;<�I;w�I;�I;��I;�I;��I;B�I;D�I;)�I;��I;B�I;|I;�XI;;I;U'I;      �F;��F;�F;�2G;s�G;1&H;��H;I;*mI;��I;��I;��I;�I;��I;��I;�I;��I;�wI;�bI;aPI;a@I;{2I;�&I;lI;�I;|I;\I;<I;�H;��H;��H;��H;��H;b�H;��H;�H;��H;�H;��H;a�H;��H;��H;��H;��H;�H;;I;[I;|I;�I;iI;�&I;{2I;[@I;bPI;�bI;�wI;��I;�I;��I;��I;�I;��I;��I;��I;)mI;I;��H;0&H;w�G;�2G;�F;��F;      ƶ?;��?;��@;�tA;9�B;v�C;�BE;��F;��G;�xH;�I;��I;��I;��I;l�I;��I;F�I;g�I;B�I;LiI;�TI;-CI;*4I;�'I;�I;�I;PI;I;� I;��H;S�H;��H;��H;�H;��H;a�H;.�H;a�H;�H;�H;��H;��H;Q�H;��H;� I;I;OI;�I;�I;'I;'4I;-CI;�TI;MiI;C�I;i�I;D�I;��I;l�I;��I;��I;��I;�I;�xH;��G;��F;�BE;v�C;8�B;�tA;��@;��?;      �0;�51;E�2;v�4;17;T#:;"0=;� @;=�B;�	E;��F;%H;�	I;��I;��I;��I;��I;0�I;��I;3�I;�mI;�WI;�DI;�4I;|'I;nI;=I;�I;sI;k I;k�H;�H;��H;��H;��H;��H;��H;��H;��H;��H;��H;�H;i�H;h I;pI;�I;;I;nI;{'I;�4I;�DI;�WI;�mI;3�I;��I;1�I;��I;��I;��I;��I;�	I;%H;��F;�	E;;�B;� @;"0=;T#:;17;x�4;D�2;�51;      };(;��;�;6 ;&;�\,;�2;N98;�/=;�FA;�rD;��F;DJH;�9I;]�I;��I;��I;)�I;��I;��I;BpI;�XI;�DI;%4I;�&I;]I;!I;�
I;�I;��H;��H;$�H;�H;q�H;}�H;E�H;~�H;q�H;�H;$�H;��H;��H;�I;�
I;"I;\I;�&I;%4I;�DI;�XI;BpI;��I;��I;)�I;��I;��I;^�I;�9I;DJH;��F;�rD;�FA;�/=;M98;�2;�\,;
&;< ;�;{�;;      ���:��:I�::��:��:$Q ;�e;�V;z#;:e-;ͼ5;�h<;�tA;�	E;�eG;f�H;d�I;A�I;#�I;L�I;P�I;/�I;ApI;�WI;*CI;|2I;�$I;�I;�I;}	I;�I;0�H;��H;9�H;��H;f�H;�H;f�H;��H;9�H;��H;2�H;�I;z	I;�I;�I;�$I;~2I;)CI;�WI;<pI;/�I;N�I;N�I;#�I;C�I;d�I;f�H;�eG;�	E;�tA;�h<;̼5;:e-;z#;�V;�e;"Q ;K��::��:I�:��:      ��p� �,� %9�Ƴ9p�":(�u:��:���:^��:[R;� ;��,;H�6;�)>;<C;��F;�lH;�kI;��I;��I;��I;R�I;��I;�mI;�TI;b@I;�/I;\"I;�I;�I;
I;�I;��H;��H;��H;��H;�H;��H;��H;��H;��H;�I;
I;�I;�I;]"I;�/I;a@I;�TI;�mI;��I;R�I;��I;��I;��I;�kI;�lH;��F;<C;�)>;H�6;��,;� ;YR;\��:���:��:H�u:��":�Ƴ9�$9 �,�      �o&�<!��4����氺`�O��9T�v�9L�u:	$�:6H�:?D;Z#;�71;l;;��A;1�E;�$H;�VI;F�I;��I;K�I;��I;3�I;FiI;dPI;W<I;0,I;WI;�I;�I;�I;�I;g�H;
�H;��H;?�H;��H;
�H;g�H;�I;�I;�I;�I;RI;0,I;T<I;bPI;FiI;.�I;��I;K�I;��I;G�I;�VI;�$H;1�E;��A;l;;�71;Z#;=D;2H�:$�:L�u:(v�9�9T�T�O�氺���4�H!�      �kٻU�Իwǻ ����V���n���+��ԺP�1���39�m:�:��;9�;�\,;�8;�@;p]E;�
H;�VI;��I;#�I;)�I;��I;<�I;�bI;�JI;]7I;(I;�I;gI;I;qI;oI;��H;�H;��H;�H;��H;oI;pI;I;fI;�I;
(I;]7I;�JI;�bI;<�I;��I;#�I;#�I;��I;�VI;�
H;q]E;�@;�8;�\,;9�;��;�:�m:��39H�1��Ժ��+��n��V�� ���vǻV�Ի      2yY��|U�E�I�:�7��� ��!���Ի�᝻m�T�̴�#��v�9���:�l�:;�);D17;] @;m]E;�$H;�kI;@�I;��I;-�I;f�I;�wI;�ZI;�CI;�1I;�#I;`I;�I;f	I;�I;mI;��H;7�H;��H;mI;�I;e	I;�I;`I;�#I;�1I;�CI;�ZI;�wI;f�I;)�I;��I;@�I;�kI;�$H;m]E;^ @;B17;�);;�l�:���:�v�9#�ʴ�m�T��᝻��Ի�!��� �:�7�E�I��|U�      ��ü\l��t����R��=ߓ�Z�{��M��� ��컹���d�B��鰺�=o���u:��:�R;a�';D17;�@;4�E;�lH;e�I;��I;��I;A�I;��I;mI;�QI;a<I;�+I;�I;�I;�I;I;zI;`I;�I;`I;zI;I;�I;�I;�I;�+I;^<I;�QI;�lI;��I;A�I;��I;��I;e�I;�lH;5�E;�@;F17;`�';�R;��:��u:�=o��鰺c�B������컅� ��M�Z�{�<ߓ��R��t���]l��      �'��-$�_��Z����	?ټw��:���hyY��k��Ի(���X��x����$R:��:�R;�);�8;��A;��F;i�H;^�I;��I;��I;�I;?�I;aI;*HI;�4I;�%I;|I;I;�I;�I;II;|I;II;�I;�I;I;~I;�%I;�4I;&HI;aI;;�I;�I;��I;��I;[�I;h�H;��F;��A;�8;�);�R;��:�$R:x����X��)���Ի�k�hyY�:���w��?ټ���Z�_���-$�      Z+����d̀�/l��Q�&�2�C��������@��}�>�N2��V��f1�`��$R:���:;�\,;m;;<C;�eG;�9I;��I;k�I;�I;w�I;�qI;�TI;�>I;p-I;b I;�I;�I;I;HI;GI;HI;I;�I;�I;e I;o-I;�>I;�TI;�qI;u�I;�I;k�I;��I;�9I;�eG;<C;m;;�\,;;���:�$R:`��g1�V��N2��}�>��@��������C�&�2��Q�/l�d̀���      n�ླྀhܽq�н_y��b什Q ��l��n<�N���>ټ��P|U�x������c1�p�����u:�l�:7�;�71;�)>;�	E;CJH;��I;��I;��I;�I;�I;�bI;�HI;a5I;�&I;�I;�I;tI;WI;U
I;WI;tI;�I;�I;�&I;^5I;�HI;�bI;�I;�I;��I;��I;��I;>JH;�	E;�)>;�71;5�;�l�:��u:x���f1�����y��P|U����>ټN���n<�l�P ��b什_y��q�н�hܽ      ��4�i1��&������l�཈�������`��'���TR��?�]�x��V���X��@=o����:��;\#;H�6;�tA;��F;�	I;��I;�I;��I;N�I;qI;�SI;�=I;�,I;� I;�I;�I;zI;tI;xI;�I;�I;� I;�,I;�=I;�SI;qI;N�I;��I;�I;��I;�	I;��F;�tA;H�6;\#;��;���:@>o��X��V��y��?�]�TR����'��`��������l��������&�i1�      �x���o��ń�LUo���O�,�-�{��hܽ^什ռx���2�sb��TR��Q|U�M2��)���鰺�v�9�:@D;��,;�h<;�rD;%H;��I;��I;�I;;�I;?�I;_I;?FI;�3I;�%I;
I;�I;�I;lI;�I;�I;I;�%I;�3I;?FI;_I;>�I;;�I;�I;��I;��I;|%H;�rD;�h<;��,;@D;�:�v�9�鰺*��N2��Q|U�TR��tb����2�ռx�^什�hܽ{�,�-���O�LUo�ń��o��      z���྅�Ѿ*����נ�
ń�<�S�	�#�bO��~n��K̀���2����}�>��Իe�B�#��m:8H�:� ;˼5;�FA;��F;�I;��I;��I;پI;��I;�jI;�NI;C:I;+I;1 I;I;�I;�I;�I;I;1 I;+I;D:I;�NI;�jI;��I;پI;��I;��I;�I;��F;�FA;ɼ5;� ;2H�:�m:#�j�B��Ի}�>�������2�K̀�~n��bO��	�#�<�S�
ń��נ�*�����Ѿ��      �3���/��X#��	��A��،Ⱦ�f��KUo�`1�Ͱ��~n��ռx��'��>ټ�@���k�����̴��39	$�:YR;:e-;�/=;�	E;�xH;��I;C�I;��I;8�I;FvI;�WI;�@I;)0I;Z$I;uI;�I;mI;�I;uI;Z$I;'0I;�@I;�WI;FvI;5�I;��I;B�I;��I;�xH;�	E;�/=;:e-;[R;$�:`�39ƴ𺻼���k��@���>ټ�'�ռx�~n��ΰ��`1�KUo��f��،Ⱦ�A���	��X#���/�      ���V���W�v��RZ�]58�ς�t��f���ioy�`1�bO��^什�`�N�����jyY���q�T�p�1�H�u:V��:t#;J98;6�B;��G;*mI;B�I;3�I;d�I;��I;`I;7GI;*5I;[(I;�I;�I;BI;�I;�I;[(I;'5I;6GI;`I;��I;a�I;3�I;>�I;*mI;��G;3�B;G98;t#;X��:H�u:p�1�o�T���jyY����N���`�^什bO��`1�ioy�f���t��ς�]58��RZ�W�v�V���      Ŀ8g��(ﱿ���V����U��X#�v��f���KUo�	�#��hܽ����n<����:����� ��᝻��Ժ v�9���:�V;�2;� @;��F;I;-�I;u�I;a�I;��I;5hI;CMI;�9I;%,I;�"I;�I;�I;�I;�"I;%,I;�9I;CMI;5hI;��I;^�I;u�I;*�I;I;��F;� @;�2;�V;���:v�9��Ժ�᝻�� �:�������n<�����hܽ	�#�KUo�f���w���X#��U�V������(ﱿ8g��      �x�Q9�T��wؿpQ��g_��8�_��X#�t���f��<�S�{�����l�C�w���M���Ի��+� :T���:�e;�\,; 0=;�BE;��H;��I;�I;��I;�I;�oI;�RI;G>I;�/I;�%I;) I;zI;) I;�%I;�/I;D>I;�RI;�oI;�I;��I;�I;��I;��H;�BE;0=;�\,;�e;��: :T���+���Ի�M�w��C�l�����{�<�S��f��t���X#�8�_�g_��pQ��wؿT��Q9�      �X1���,�i���<��7g��g_���U�ς�،Ⱦ
ń�,�-�l��Q ��'�2�	?ټ\�{��!��n�`�O��u:Q ;&;N#:;s�C;7&H;D�I;W�I; �I;�I;�vI;XI;$BI;�2I;H(I;w"I;� I;x"I;H(I;�2I;!BI;
XI;�vI;�I;��I;W�I;B�I;4&H;u�C;J#:;&;Q ;,�u:d�O��n��!�\�{�
?ټ'�2�Q ��l��,�-�
ń�،Ⱦς��U�g_��7g��<�i����,�      d��]]�6K��X1�[f��pQ��V���]58��A���נ���O���b什�Q�	���=ߓ��� ��V��$氺|�":%��:< ;17;9�B;u�G;|I;�I;��I;�I;o|I;l\I;~EI;P5I;k*I;b$I;_"I;b$I;j*I;P5I;}EI;n\I;o|I;�I;��I;�I;|I;s�G;:�B;17;> ;!��:��":$氺�V���� �>ߓ�	����Q�b什����O��נ��A��]58�V���pQ���[f��X1�6K��]]�      O������4z���V��X1��<�wؿ����RZ��	�*���LUo����`y��/l�Z��R��<�7��������Ƴ9F��:�;v�4;�tA;�2G;�XI;��I;��I;9�I;*�I;�_I;0HI;W7I;0,I;�%I;�#I;�%I;0,I;V7I;.HI;�_I;*�I;6�I;��I;��I;�XI;�2G;�tA;q�4;�;F��:�Ƴ9������;�7��R��Z�/l�`y�����LUo�*����	��RZ����wؿ�<��X1���V��4z�����      �o��f^���ē��4z�6K�i��T��(ﱿX�v��X#���Ѿń��&�q�нd̀�`��u���G�I�~ǻ�4� $9+�:q�;:�2;��@;�F;;I;%�I;2�I;ɲI;��I;�bI;0JI;�8I;�-I;�&I;%I;�&I;�-I;�8I;0JI;�bI;��I;ƲI;/�I;%�I;;I;�F;��@;4�2;u�;+�: $9�4�~ǻG�I�u���`��d̀�q�н�&�ń���Ѿ�X#�X�v�(ﱿT��i��6K��4z��ē�f^��      s'���X��f^�������]]���,�Q9�8g��V�����/����o��i1��hܽ���-$�^l���|U�X�ԻQ!� �,���:;�51;��?;��F;`'I;��I;K�I;i�I;ӆI;dI;rKI;�9I;X.I;�'I;�%I;�'I;Y.I;�9I;qKI;dI;ӆI;f�I;H�I;��I;_'I;��F;��?;�51;;��: �,�Q!�X�Ի�|U�_l���-$����hܽi1��o���ྛ�/�V���8g��Q9���,��]]�����f^���X��      ����,������U���L�Q�ș$�5�����>�}�J(�C�׾�T���L+���սl����L���iO���ͻ`�� &m8�o�:��;f�1;��?;vF;� I;��I;��I;��I;�vI;�WI;�AI;%2I;(I;"I;  I;"I;(I;%2I;�AI;�WI;�vI;��I;��I;��I;� I;vF;��?;d�1;��;�o�:�&m8a����ͻ�iO� L����l����ս�L+��T��C�׾J(�>�}���5���ș$�L�Q�U��������,��      �,��b��$P���{���K��x �����s�����w��$���Ҿh��� (���ѽӷ��(������K�<ɻ�����8���:��;��1;#@;��F;<I;�I;H�I;ԞI;�uI;`WI;�AI;�1I;�'I;�!I;�I;�!I;�'I;�1I;�AI;aWI;�uI;ҞI;E�I;�I;<I;��F;#@;��1;��;���:��8���<ɻߔK����(�ӷ����ѽ (�h�����Ҿ�$���w�s��������x ���K��{�$P��b��      ����$P�������d���;�$���㿴���#f�f�� ž��z���?�ƽ(0v�V5�0����o@�z���Oi�@bu9|K�:Q];�73;S�@;,�F;fI;��I;��I;��I;tI;�UI;s@I;1I;'I;?!I;cI;?!I;'I;1I;r@I;�UI;tI;}�I;��I;��I;fI;,�F;S�@;�73;U];~K�:@bu9Pi�z����o@�0���V5�(0v�?�ƽ����z� žf��#f�������$����;���d����$P��      U����{���d��F�ș$�;����ɿ0蒿��K�R���j��Zb�G�4���u�a����?�����.��d���غ���9�Y�:iX;�25;U�A;�!G;i7I;��I;��I;z�I;�pI;�SI;�>I;�/I;�%I;T I;cI;T I;�%I;�/I;�>I;�SI;�pI;y�I;~�I;��I;i7I;�!G;S�A;�25;kX;�Y�:���9�غ�d����.�?������u�a�4���G�Zb��j��R����K�0蒿��ɿ;��ș$��F���d��{�      L�Q���K���;�ș$��;
��޿�����w�s,���澟���)�D������I��&�G�����N�������������9:���:�n!;��7;�B;��G;ZI;\�I;��I;�I;�lI;�PI;I<I;�-I;F$I;�I;�I;�I;E$I;�-I;H<I;�PI;�lI;�I;��I;]�I;ZI;��G;�B;��7;�n!;���:�9:����������N�����&�G��I������)�D��������s,���w�����޿�;
�ș$���;���K�      ș$��x �$��;���޿r���˅���F��
��~����z��$���ս���B2+���ϼPp�����0�]�`�*�V��:>�;9';Ȍ:;+�C;?H;�}I;Q�I;��I;�I;�gI;�LI;N9I;k+I;X"I;*I;]I;(I;X"I;m+I;N9I;�LI;�gI;�I;��I;Q�I;�}I;=H;+�C;Ì:;9';>�;X��:h�*�0�]�����Pp���ϼB2+������ս�$���z��~���
��F�˅��r����޿;��$���x �      5��������㿌�ɿ���˅����P�e��?�׾�`��W�H����@��T�a���̡���D��ɻ� ��ҭ�X�:�;�I-;Y|=;WCE;ۅH;9�I;�I;��I;�I;�aI;WHI;�5I;�(I; I;I;�I;I; I;�(I;�5I;XHI;�aI;�I;��I;�I;6�I;ۅH;UCE;U|=;�I-;�;X�:�ҭ�� ��ɻ�D�̡����T�a��@����W�H��`��?�׾e����P�˅�������ɿ�㿵���      ��s�������0蒿��w��F�e��Ͱ�"����Yb�+����ѽ�%��D4�ڟ�X������G��~潺@��9�r�: ;:3;MQ@;�vF;M�H;7�I;��I;��I;�zI;�ZI;GCI;�1I;�%I;wI;�I;WI;�I;wI;�%I;�1I;HCI;�ZI;�zI;��I;��I;4�I;M�H;�vF;HQ@;:3; ;�r�:8��9~潺�G�����X��ڟ�D4��%����ѽ+���Yb�"���Ͱ�e���F���w�0蒿����s���      =�}���w�#f���K�s,��
�?�׾"�����k���'�iz꽟I���;V�=M�����iO�\G�NoE�4�����:l� ;ҿ$;ߴ8;��B;2�G;kKI;D�I;I�I;s�I;;qI;�SI;�=I;�-I;<"I;�I;MI;�I;MI;�I;<"I;�-I;�=I;�SI;9qI;r�I;J�I;A�I;kKI;/�G;��B;ݴ8;ӿ$;n� ;���:0��MoE�\G໦iO����=M��;V��I��iz���'���k�"���?�׾�
�s,���K�#f���w�      J(��$�f��R������~���`���Yb���'��U�J$��G�m�&����ϼ�/��8������X�غ�9�9���:G;	H.;G|=;qE;�\H;X�I;��I;��I;-�I;4gI;7LI;8I;<)I;�I;�I;�I;]I;�I;�I;�I;;)I;8I;7LI;6gI;,�I;��I;��I;V�I;�\H;qE;D|=;	H.;G;���:�9�9T�غ����8���/����ϼ&��G�m�J$���U���'��Yb��`���~�����R��f���$�      C�׾��Ҿ ž�j��������z�W�H�+��iz�J$���/v�2+�ސ�����5��ɻ4�0'�����:���:fo!;>P6;<lA;�F;��H;ŷI;��I;�I;�}I;�\I;�DI;92I;�$I;�I;�I;�I;�I;�I;�I;�I;�$I;<2I;�DI;�\I;}I;�I;��I;ǷI;��H;�F;8lA;>P6;fo!;���:���:'��4��ɻ��5���ސ�2+��/v�J$��iz�+��W�H���z������j�� ž��Ҿ      �T��h�����z�Zb�)�D��$�����ѽ�I��G�m�2+�������H�K���}�p����ؓ�9xT�:0;��-;��<;{zD;�H;�mI;�I;��I;ĕI;�oI;�RI;�<I;5,I;�I;DI;hI;�I;�I;�I;iI;DI;�I;8,I;�<I;�RI;�oI;ĕI;��I;�I;�mI;�H;xzD;��<;��-;0;|T�:��9���y�p���H�K�������2+�G�m��I����ѽ���$�)�D�Zb���z�h���      �L+� (���G�������ս�@���%���;V�&��ސ�����zMS�H����:D�@o8Lq�:�;��$;-_7;_�A;��F;+�H;��I;��I;��I;�I;�bI;�HI;D5I;Y&I;cI;uI;$I;I;=
I;I;$I;uI;cI;[&I;D5I;�HI;�bI;�I;��I;��I;��I;'�H;��F;`�A;-_7;��$;�;Pq�:@o88D���G��zMS�����ސ�&���;V��%���@����ս����G��� (�      ��ս��ѽ?�ƽ4����I�����T�a�D4�<M���ϼ��H�K�H��?G��=f���o���:,C�:�Y;�1;�l>;E; 0H;NqI;5�I; �I;�I;6sI;�UI;#?I;�-I;� I;�I;�I;�
I;II;jI;II;�
I;�I;�I;� I;�-I;%?I;�UI;7sI;�I;"�I;5�I;LqI;0H;E;�l>;�1;�Y;4C�:��:��o�<f�>G��H��H�K�����ϼ<M�D4�T�a�����I��4���>�ƽ��ѽ      l��ӷ��'0v�t�a�&�G�A2+���ڟ�����/����5�����?f��׬�|�g:��:2�;DI-;Kg;;0OC;;SG;�I;��I;U�I;6�I;;�I;AcI;�II;�5I;�&I; I;mI;I;�I;�I;�I;�I;�I;I;mI;I;�&I;�5I;�II;AcI;:�I;8�I;S�I;��I;�I;=SG;0OC;Ng;;DI-;5�;��:|�g:�׬�?f�������5��/�����ڟ���A2+�&�G�t�a�'0v�ӷ��      ��'�U5���������ϼʡ��X���iO�8���ɻz�p�:D���o���g:?`�:pG;�*;�9;��A;�uF;Q�H;��I;��I;ݻI;~�I;�pI;lTI;�>I;S-I;�I;�I;/I;�I;�I;�I;I;�I;�I;�I;.I;�I;�I;S-I;�>I;lTI;�pI;~�I;ܻI;��I;��I;R�H;�uF;��A;�9;�*;oG;?`�:��g:��o�:D�z�p��ɻ8���iO�X��ʡ����ϼ������U5�(�      L�����0���>����N��Pp��D����YG�����4������o8��:��:nG;1�(;ɶ7;��@;��E;�QH;JmI;��I;-�I;ҢI;^}I;�^I;�FI;4I;%I;�I;�I;(
I;DI;I; I;��H; I;I;FI;'
I;�I;�I;%I;4I;�FI;�^I;_}I;ҢI;'�I;��I;LmI;�QH;��E;��@;˶7;1�(;nG;��:��:�o8����4�����YGໂ���D�Pp��N��>���0������      �iO�ޔK��o@���.���������ɻ�G��KoE�X�غ'����9Hq�:,C�:5�;�*;ȶ7;�P@;�\E;$H;JI;��I;��I;B�I;��I;vhI;�NI;�:I;t*I;�I;�I;I;NI;FI;e�H;��H;�H;��H;e�H;FI;MI;I;�I;�I;q*I;�:I;�NI;vhI;��I;=�I;��I;��I; JI;&H;�\E;�P@;ƶ7;�*;5�;.C�:Lq�:��9'��T�غJoE��G���ɻ����~����.��o@���K�      ��ͻ9ɻr����d�����(�]�� �|潺���9�9���:�T�:�;�Y;HI-;�9;��@;�\E;��G;h5I;�I;{�I;�I;��I;�pI;�UI;�@I;k/I;�!I;�I;xI;�I;�I;V�H;��H;N�H;��H;N�H;��H;V�H;�I;�I;zI;�I;�!I;m/I;�@I;�UI;�pI;��I;�I;{�I;�I;i5I;��G;�\E;��@;�9;II-;�Y;�;�T�:���:�9�9��x潺� �$�]�����d��r���9ɻ      ]����Li��غ����h�*��ҭ� ��9���:���:���: 0;��$;�1;Jg;;��A;��E;#H;e5I;o�I;��I;��I;ϗI;�vI;�[I;�EI;�3I;l%I;�I;�I;�	I;�I;��H;��H;\�H;�H;��H; �H;\�H;��H;��H;�I;�	I;�I;�I;l%I;�3I;�EI;�[I;�vI;ɗI;��I;��I;q�I;e5I;#H;��E;��A;Jg;;�1;��$; 0;���:���:���:(��9�ҭ�\�*�쓛��غJi����      �(m8 ��8�bu9x��9��9:`��:!X�:�r�:p� ;G;fo!;��-;,_7;~l>;0OC;�uF;�QH;JI;�I;��I;�I;�I;�zI;�_I;}II;�7I;�(I;�I;
I;VI;I;^ I;��H;��H;8�H;�H;��H;�H;8�H;��H;��H;` I;I;SI;	I;�I;�(I;�7I;}II;�_I;�zI;�I;�I;��I;�I;JI;�QH;�uF;0OC;~l>;,_7;��-;fo!;G;p� ;�r�:X�:f��:��9:���9�bu9���8      �o�:��:�K�:�Y�:���:I�;�;  ;ؿ$;H.;BP6;��<;]�A;E;>SG;N�H;LmI;��I;{�I;��I;�I;|I;�aI;�KI;�9I;+I;�I;�I;�I;`I;'I;+�H;�H;��H;'�H;D�H;�H;D�H;'�H;��H;�H;+�H;'I;\I;�I;�I;�I;+I;�9I;�KI;�aI;|I;�I;��I;{�I;��I;ImI;L�H;@SG;E;]�A;��<;@P6;H.;ٿ$;  ;�;K�;Ȩ�:�Y�:�K�:��:      ��;��;V];dX;�n!;9';�I-;:3;�8;G|=;<lA;}zD;��F; 0H;�I;��I;��I;��I;�I;ϗI;�zI;�aI;�LI;V;I;�,I;k I;\I;0I;uI;I;��H;5�H;��H;��H;?�H;��H;Z�H;��H;?�H;��H;��H;5�H;��H;I;qI;0I;YI;l I;�,I;S;I;�LI;�aI;�zI;їI;�I;��I;��I;��I;�I; 0H;��F;}zD;;lA;F|=;�8;:3;�I-;9';�n!;dX;X];��;      |�1;��1;�73;�25;��7;Ȍ:;b|=;KQ@;��B;sE;�F;�H;'�H;PqI;��I;��I;/�I;D�I;��I;�vI;�_I;�KI;U;I;-I;&!I;SI;I;QI;�I;2�H;��H;��H;_�H;��H;��H;	�H;��H;�H;��H;��H;[�H;��H;��H;.�H;�I;PI;I;SI;&!I;-I;S;I;�KI;�_I;�vI;��I;E�I;,�I;��I;��I;PqI;'�H;�H;�F;pE;��B;MQ@;a|=;Ɍ:;��7;�25;�73;��1;      ��?;-@;A�@;Z�A;�B;/�C;TCE;�vF;1�G;�\H;��H;�mI;��I;8�I;X�I;߻I;آI;��I;�pI;�[I;II;�9I;�,I;-!I;�I;�I;�I;0I;��H;��H;��H;c�H;��H;)�H;'�H;��H;i�H;��H;(�H;'�H;��H;c�H;��H;��H;��H;0I;�I;�I;�I;'!I;�,I;�9I;~II;�[I;�pI;��I;բI;ݻI;V�I;6�I;��I;�mI;��H;�\H;/�G;�vF;TCE;.�C;�B;Z�A;A�@;-@;      )vF;ʊF; �F;�!G;��G;9H;مH;F�H;kKI;U�I;ķI;�I;��I; �I;5�I;|�I;^}I;uhI;�UI;�EI;�7I;+I;i I;SI;�I;	I;�I;��H;)�H;�H;b�H;u�H;��H;��H;��H;R�H;#�H;R�H;��H;��H;��H;v�H;a�H;�H;&�H;��H;�I;	I;�I;PI;h I;+I;�7I;�EI;�UI;vhI;\}I;z�I;6�I; �I;��I;�I;÷I;R�I;iKI;G�H;مH;8H;��G;�!G;�F;��F;      � I;=I;dI;p7I;ZI;�}I;=�I;4�I;G�I;��I;��I;��I;��I;�I;<�I;�pI;�^I;�NI;�@I;�3I;�(I;�I;]I;I;�I;�I;�H;]�H;�H;p�H;^�H;��H;S�H;S�H;��H;@�H;�H;@�H;��H;R�H;P�H;��H;`�H;m�H;�H;]�H;�H;�I;�I;I;[I;�I;�(I;�3I;�@I;�NI;�^I;�pI;<�I;�I;��I;��I;��I;��I;G�I;4�I;=�I;�}I; ZI;p7I;cI;;I;      ��I;�I;��I;��I;\�I;Q�I;�I;��I;N�I;��I;�I;ȕI;�I;;sI;BcI;lTI;�FI;�:I;m/I;p%I;�I;�I;3I;TI;-I;��H;]�H;4�H;}�H;^�H;��H;�H;�H;?�H;��H;;�H;(�H;;�H;��H;?�H;�H;�H;��H;]�H;z�H;4�H;]�H;��H;/I;TI;2I;�I;�I;o%I;k/I;�:I;�FI;lTI;BcI;;sI;�I;ʕI;�I;��I;N�I;��I;�I;Q�I;e�I;��I;��I;"�I;      �I;G�I;��I;��I;��I;��I;��I;��I;u�I;-�I;}I;�oI;�bI;�UI;�II;�>I;4I;r*I;�!I;�I;I;�I;tI;�I;��H;*�H;�H;{�H;g�H;��H;�H;��H;��H;5�H;��H;p�H;g�H;p�H;��H;5�H;��H;��H;�H;��H;g�H;}�H;�H;)�H;��H;�I;rI;�I;I;�I;�!I;r*I;4I;�>I;�II;�UI;�bI;�oI;~}I;*�I;u�I;��I;��I;��I;��I;��I;��I;:�I;      ��I;ڞI;��I;|�I;�I;
�I;�I;�zI;@qI;=gI;�\I;�RI;�HI;,?I;�5I;U-I; %I;�I;�I;�I;YI;_I;I;3�H;��H;�H;m�H;]�H;��H; �H;��H;��H;��H;X�H;��H;��H;��H;��H;��H;X�H;��H;��H;��H;��H;��H;^�H;m�H;��H;��H;2�H;I;`I;WI;�I;�I;�I;%I;T-I;�5I;,?I;�HI;�RI;�\I;=gI;BqI;�zI;�I;
�I;�I;z�I;��I;מI;      �vI;�uI;tI;�pI;�lI;�gI;�aI;�ZI;�SI;<LI;�DI;�<I;I5I;�-I;�&I;�I;�I;�I;I;�	I;&I;(I;��H;��H;��H;c�H;]�H;��H;�H;��H;��H;��H;%�H;��H;G�H;�H;��H;�H;G�H;��H;"�H;��H;��H;��H;�H;��H;]�H;a�H;��H;��H;��H;(I;#I;�	I;I;�I;�I;�I;�&I;�-I;I5I;�<I;�DI;<LI;�SI; [I;�aI;�gI;�lI;�pI;tI;�uI;      �WI;oWI;VI;�SI;�PI;�LI;VHI;NCI;�=I;8I;@2I;?,I;]&I;� I;	I;�I;�I;I;�I;�I;h I;1�H;7�H;��H;b�H;u�H;��H;�H;��H;��H;��H;�H;}�H;�H;��H;�H;��H;�H;��H;�H;|�H; �H;��H;��H;��H;�H;��H;t�H;f�H;��H;6�H;1�H;g I;�I;�I;I;�I;�I;I;� I;]&I;?,I;@2I;8I;�=I;NCI;VHI;�LI;�PI;�SI;VI;jWI;      BI;�AI;z@I;�>I;P<I;N9I;�5I;�1I;�-I;<)I;�$I;�I;eI;�I;qI;3I;/
I;KI;�I;��H;��H;�H;��H;b�H;��H;��H;T�H;�H;��H;��H;'�H;��H;��H;��H;G�H;�H;$�H;�H;G�H;��H;��H;��H;&�H;��H;��H;�H;Q�H;��H;��H;b�H;��H;�H;��H;��H;�I;MI;.
I;2I;pI;�I;eI;�I;�$I;=)I;�-I;�1I;�5I;P9I;J<I;�>I;z@I;�AI;      32I;�1I;1I;�/I;�-I;g+I;�(I;�%I;A"I;�I;�I;II;vI;�I;I;�I;PI;FI;]�H;��H;��H;��H;��H;��H;$�H;��H;P�H;?�H;4�H;X�H;��H;�H;��H;,�H;��H;��H;��H;��H;��H;,�H;��H;�H;��H;X�H;8�H;=�H;P�H;��H;%�H;��H;��H;��H;��H;��H;]�H;GI;NI;�I;I;�I;vI;II;�I;�I;C"I;�%I;�(I;k+I;�-I;�/I;1I;�1I;      (I;�'I;'I;�%I;[$I;R"I; I;}I;�I;�I;�I;sI;)I;�
I;�I;�I; I;d�H;��H;c�H;B�H;)�H;A�H;��H;!�H;��H;��H;��H;��H;��H;E�H;��H;F�H;�H;��H;��H;��H;��H;��H;�H;C�H;��H;G�H;��H;��H;��H;��H;��H;!�H;��H;A�H;)�H;A�H;c�H;��H;e�H;I;�I;�I; I;+I;sI;�I;�I;�I;}I; I;V"I;S$I;�%I;'I;�'I;      "I;�!I;G!I;X I;I;$I;I;�I;YI;�I;�I;�I;I;SI;�I;�I;) I;��H;U�H;(�H;%�H;I�H;��H;�H;��H;N�H;?�H;<�H;s�H;��H;�H;��H;�H;��H;��H;j�H;e�H;j�H;��H;��H;�H;��H;�H;��H;v�H;;�H;=�H;L�H;��H;�H;��H;I�H;#�H;(�H;U�H;��H;' I;�I;�I;SI;I;�I;�I;�I;YI;�I;I;*I;�I;X I;G!I;�!I;        I; I;oI;gI;I;ZI;�I;\I;�I;[I;�I;I;?
I;rI;�I;I;��H;�H;��H;��H;��H;�H;\�H;��H;e�H;�H;�H;.�H;i�H;��H;��H;��H;$�H;��H;��H;f�H;J�H;f�H;��H;��H;"�H;��H;��H;��H;l�H;.�H;�H;�H;e�H;��H;\�H;�H;��H;��H;��H;�H;��H;I;�I;rI;?
I;I;�I;]I;�I;\I;�I;^I;�I;gI;oI;  I;      "I;�!I;G!I;X I;I;&I;I;�I;YI;�I;�I;�I;I;TI;�I;�I;) I;��H;U�H;(�H;&�H;I�H;��H;�H;��H;N�H;?�H;;�H;s�H;��H;�H;��H;�H;��H;��H;j�H;e�H;j�H;��H;��H;�H;��H;�H;��H;v�H;<�H;=�H;L�H;��H;�H;��H;I�H;#�H;(�H;U�H;��H;' I;�I;�I;QI;I;�I;�I;�I;YI;�I;I;(I;�I;X I;D!I;�!I;      (I;�'I;'I;�%I;[$I;R"I; I;}I;�I;�I;�I;sI;+I;�
I;�I;�I; I;d�H;��H;c�H;C�H;)�H;A�H;��H;!�H;��H;��H;��H;��H;��H;G�H;��H;F�H;�H;��H;��H;��H;��H;��H;�H;C�H;��H;E�H;��H;��H;��H;��H;��H;!�H;��H;A�H;)�H;A�H;c�H;��H;e�H;I;�I;�I; I;)I;sI;�I;�I;�I;}I; I;V"I;S$I;�%I;'I;�'I;      52I;�1I;1I;�/I;�-I;g+I;�(I;�%I;A"I;�I;�I;II;vI;�I;I;�I;PI;FI;]�H;��H;��H;��H;��H;��H;%�H;��H;P�H;=�H;4�H;W�H;��H;�H;��H;,�H;�H;��H;��H;��H;��H;,�H;��H;�H;��H;Z�H;6�H;?�H;P�H;��H;$�H;��H;��H;��H;��H;��H;]�H;GI;NI;�I;I;�I;vI;II;�I;�I;C"I;�%I;�(I;k+I;�-I;�/I;1I;�1I;      BI;�AI;|@I;�>I;P<I;N9I;�5I;�1I;�-I;<)I;�$I;�I;eI;�I;pI;2I;/
I;KI;�I;��H;��H;�H;��H;b�H;��H;��H;T�H;�H;��H;��H;&�H;��H;��H;��H;G�H;�H;$�H;�H;F�H;��H;��H;��H;'�H;��H;��H;�H;Q�H;��H;��H;a�H;��H;�H;��H;��H;�I;KI;.
I;3I;qI;�I;dI;�I;�$I;=)I;�-I;�1I;�5I;P9I;I<I;�>I;y@I;�AI;      �WI;oWI;VI;�SI;�PI;�LI;XHI;NCI;�=I;8I;@2I;?,I;]&I;� I;I;�I;�I;I;�I;�I;k I;1�H;7�H;��H;f�H;u�H;��H;�H;��H;��H;��H;�H;|�H;�H;��H;�H;��H;�H;��H;�H;{�H;�H;��H;��H;��H;�H;��H;t�H;b�H;��H;6�H;1�H;g I;�I;�I;I;�I;�I;I;� I;]&I;?,I;@2I; 8I;�=I;NCI;XHI;�LI;�PI;�SI;VI;kWI;      �vI;�uI;tI;�pI;�lI;�gI;�aI;�ZI;�SI;;LI;�DI;�<I;I5I;�-I;�&I;�I;�I;�I;I;�	I;'I;(I;��H;��H;��H;c�H;]�H;��H;�H;��H;��H;��H;#�H;��H;G�H;�H;��H;�H;G�H;��H;"�H;��H;��H;��H;�H;��H;]�H;a�H;��H;��H;��H;(I;#I;�	I;I;�I;�I;�I;�&I;�-I;I5I;�<I;�DI;>LI;�SI; [I;�aI;�gI;�lI;�pI;tI;�uI;      ��I;ٞI;��I;z�I;�I;�I;�I;�zI;CqI;;gI;�\I;�RI;�HI;,?I;�5I;T-I; %I;�I;�I;�I;ZI;`I;I;3�H;��H;�H;o�H;^�H;��H; �H;��H;��H;��H;W�H;��H;��H;��H;��H;��H;X�H;��H;��H;��H;��H;��H;]�H;l�H;��H;��H;5�H;I;_I;WI;�I;�I;�I;%I;W-I;�5I;,?I;�HI;�RI;�\I;;gI;CqI;�zI;�I;�I;�I;z�I;��I;ڞI;      ��I;C�I;��I;��I;��I;��I;��I;��I;u�I;,�I;}I;�oI;�bI;�UI;�II;�>I;4I;q*I;�!I;�I;I;�I;tI;�I;��H;*�H;�H;}�H;g�H;��H;�H;��H;��H;5�H;��H;p�H;g�H;p�H;��H;5�H;��H;��H;�H;��H;g�H;{�H;�H;)�H;��H;�I;rI;�I;I;�I;�!I;t*I;4I;�>I;�II;�UI;�bI;�oI;}I;-�I;v�I;��I;��I;��I;��I;�I;��I;C�I;      ��I;�I;��I;��I;\�I;Q�I;�I;��I;N�I;��I;�I;ʕI;�I;;sI;BcI;lTI;�FI;�:I;k/I;o%I;�I;�I;3I;TI;/I;��H;]�H;4�H;{�H;`�H;��H;�H;�H;=�H;��H;;�H;(�H;;�H;��H;?�H;�H;�H;��H;]�H;{�H;4�H;]�H;��H;-I;TI;2I;�I;�I;p%I;m/I;�:I;�FI;nTI;BcI;;sI;�I;ȕI;�I;��I;P�I;��I;�I;N�I;h�I;��I;��I;!�I;      � I;=I;cI;j7I;ZI;�}I;;�I;4�I;G�I;��I;��I;��I;��I;�I;;�I;�pI;�^I;�NI;�@I;�3I;�(I;�I;\I;I;�I;�I;�H;]�H;�H;o�H;`�H;��H;Q�H;R�H;��H;@�H;�H;?�H;��H;R�H;Q�H;��H;^�H;o�H;�H;]�H;�H;�I;�I;I;\I;�I;�(I;�3I;�@I;�NI;�^I;�pI;;�I;�I;��I;��I;��I;��I;G�I;6�I;;�I;�}I;ZI;j7I;`I;2I;      /vF;F;*�F;�!G;��G;:H;مH;I�H;iKI;S�I;ķI;�I;��I; �I;4�I;|�I;^}I;uhI;�UI;�EI;�7I;+I;h I;RI;�I;	I;�I;��H;(�H;�H;a�H;t�H;��H;��H;��H;R�H;#�H;R�H;��H;��H;��H;v�H;b�H; �H;(�H;��H;�I;	I;�I;PI;i I;+I;�7I;�EI;�UI;vhI;\}I;|�I;5�I; �I;��I;�I;ķI;S�I;iKI;I�H;ۅH;9H;��G;�!G;'�F;��F;      ��?;-@;A�@;Z�A;�B;/�C;TCE;�vF;/�G;�\H;��H;�mI;��I;6�I;V�I;߻I;֢I;��I;�pI;�[I;II;�9I;�,I;+!I;�I;�I;�I;0I;��H;��H;��H;b�H;��H;'�H;'�H;��H;i�H;��H;'�H;(�H;��H;f�H;��H;��H;��H;0I;�I;�I;�I;*!I;�,I;�9I;}II;�[I;�pI;��I;բI;߻I;X�I;6�I;��I;�mI;��H;�\H;/�G;�vF;TCE;/�C;�B;Z�A;A�@;,@;      ��1;��1;�73;�25;��7;͌:;\|=;MQ@;��B;sE;�F;�H;*�H;PqI;��I;��I;-�I;D�I;��I;�vI;�_I;�KI;U;I;-I;&!I;SI;I;PI;�I;0�H;��H;��H;[�H;��H;��H;�H;��H;	�H;��H;��H;^�H;��H;��H;/�H;�I;QI;I;SI;&!I;	-I;S;I;�KI;�_I;�vI;��I;E�I;-�I;��I;��I;PqI;(�H;�H;�F;pE;��B;NQ@;\|=;͌:;��7;�25;�73;��1;      ��;��;d];dX;�n!;9';�I-;:3;�8;G|=;;lA;}zD;��F; 0H;�I;��I;��I;��I;�I;ЗI;�zI;�aI;�LI;V;I;�,I;k I;\I;0I;tI;I;��H;5�H;��H;��H;?�H;��H;Z�H;��H;?�H;��H;��H;5�H;��H;I;rI;0I;[I;l I;�,I;S;I;�LI;�aI;�zI;їI;�I;��I;��I;��I;�I; 0H;��F;}zD;<lA;F|=;�8;:3;�I-;9';�n!;dX;[];��;      �o�:��:�K�:�Y�:���:I�;�; ;ؿ$;H.;BP6;��<;]�A;E;>SG;N�H;JmI;��I;{�I;��I;�I;|I;�aI;�KI;�9I;+I;�I;�I;�I;`I;'I;+�H;�H;��H;'�H;F�H;�H;D�H;'�H;��H;�H;*�H;'I;\I;�I;�I;�I;+I;�9I;�KI;�aI;|I;�I;��I;{�I;��I;JmI;N�H;@SG;E;]�A;��<;BP6;H.;ٿ$;  ;�;I�;Ψ�:�Y�:�K�:��:       'm8@��8cu9���9��9:V��:#X�:�r�:p� ;G;fo!;��-;,_7;~l>;0OC;�uF;�QH;JI;�I;��I;�I;�I;�zI;�_I;}II;�7I;�(I;�I;
I;VI;I;^ I;��H;��H;8�H;�H;��H;�H;8�H;��H;��H;` I;I;SI;I;�I;�(I;�7I;}II;�_I;�zI;�I;�I;��I;�I;JI;�QH;�uF;0OC;~l>;,_7;��-;fo!;G;p� ;�r�:#X�:f��:�9:���9�bu9��8      ]����Fi��غ𓛺h�*��ҭ�(��9���:���:���: 0;��$;�1;Jg;;��A;��E;"H;e5I;o�I;��I;��I;͗I;�vI;�[I;�EI;�3I;l%I;�I;�I;�	I;�I;��H;��H;\�H;!�H;��H; �H;\�H;��H;��H;�I;�	I;�I;�I;l%I;�3I;�EI;�[I;�vI;ʗI;��I;��I;q�I;e5I;$H;��E;��A;Jg;;�1;��$; 0;���:���:���:@��9�ҭ�\�*�擛��غIi����      ��ͻ9ɻs����d�����(�]�� �x潺���9�9���:�T�:�;�Y;HI-;�9;��@;�\E;��G;i5I;�I;{�I;�I;��I;�pI;�UI;�@I;m/I;�!I;�I;zI;�I;�I;V�H;��H;N�H;��H;N�H;��H;V�H;�I;�I;xI;�I;�!I;k/I;�@I;�UI;�pI;��I;�I;{�I;�I;k5I;��G;�\E;��@;�9;II-;�Y;�;�T�:���:�9�9��x潺� �$�]�����d��r���9ɻ      �iO�ݔK��o@���.���������ɻ�G��KoE�X�غ'����9Lq�:,C�:5�;�*;ȶ7;�P@;�\E;$H;JI;��I;��I;A�I;��I;uhI;�NI;�:I;t*I;�I;�I;I;NI;FI;e�H;��H;�H;��H;e�H;FI;MI;I;�I;�I;q*I;�:I;�NI;vhI;��I;>�I;��I;��I; JI;&H;�\E;�P@;ȶ7;�*;5�;,C�:Hq�:��9'��X�غJoE��G���ɻ����~����.��o@���K�      L�����0���>����N��Pp��D����YG�����4������o8��:��:nG;3�(;ɶ7;��@;��E;�QH;LmI;��I;,�I;ҢI;^}I;�^I;�FI;4I;%I;�I;�I;(
I;FI;I; I;��H; I;I;FI;'
I;�I;�I;%I;4I;�FI;�^I;_}I;ҢI;'�I;��I;JmI;�QH;��E;��@;̶7;1�(;nG;��:��:�o8����4�����YGໂ���D�Pp��N��>���0������      ��'�U5���������ϼʡ��X���iO�8���ɻz�p�:D���o���g:?`�:pG;�*;�9;��A;�uF;R�H;��I;��I;ܻI;~�I;�pI;lTI;�>I;S-I;�I;�I;/I;�I;�I;�I;I;�I;�I;�I;.I;�I;�I;S-I;�>I;lTI;�pI;��I;ݻI;��I;��I;Q�H;�uF;��A;�9;�*;oG;?`�:��g:��o�:D�z�p��ɻ8���iO�X��ʡ����ϼ������U5�(�      l��ӷ��'0v�t�a�%�G�A2+���ڟ�����/����5�����?f��׬�|�g:��:2�;DI-;Mg;;.OC;=SG;�I;��I;S�I;6�I;<�I;AcI;�II;�5I;�&I; I;mI;I;�I;�I;�I;�I;�I;I;mI;I;�&I;�5I;�II;AcI;:�I;8�I;U�I;��I;�I;;SG;.OC;Ng;;DI-;5�;��:|�g:�׬�?f�������5��/�����ڟ���A2+�%�G�t�a�'0v�ӷ��      ��ս��ѽ?�ƽ4����I�����T�a�D4�<M���ϼ��H�K�H��?G��<f���o���:2C�:�Y;�1;~l>;E; 0H;NqI;5�I;!�I;�I;7sI;�UI;#?I;�-I;� I;�I;�I;�
I;II;jI;II;�
I;�I;�I;� I;�-I;%?I;�UI;6sI;�I;!�I;5�I;LqI;0H;E;~l>;�1;�Y;2C�:��:��o�=f�?G��H��H�K�����ϼ<M�D4�T�a�����I��4���?�ƽ��ѽ      �L+� (���G�������ս�@���%���;V�&��ސ�����zMS�G����:D⺀o8Nq�:�;��$;,_7;`�A;��F;+�H;��I;��I;��I;�I;�bI;�HI;D5I;Y&I;cI;uI;$I;I;=
I;I;$I;uI;aI;X&I;D5I;�HI;�bI;�I;��I;��I;��I;&�H;��F;_�A;-_7;��$;�;Pq�:�o8:D���H��zMS�����ސ�&���;V��%���@����ս����G��� (�      �T��h�����z�Zb�)�D��$�����ѽ�I��G�m�2+�������H�K���y�p� �����9|T�:0;��-;��<;}zD;�H;�mI;�I;��I;ĕI;�oI;�RI;�<I;5,I;�I;EI;jI;�I;�I;�I;iI;DI;�I;7,I;�<I;�RI;�oI;ĕI;��I;�I;�mI;�H;xzD;��<;��-;0;xT�: ��9���~�p���H�K�������2+�G�m��I����ѽ���$�)�D�Zb���z�h���      C�׾��Ҿ ž�j��������z�W�H�+��iz�J$���/v�2+�ސ�����5��ɻ4� '�����:���:do!;>P6;<lA;�F;��H;ŷI;��I;�I;�}I;�\I;�DI;92I;�$I;�I;�I;�I;�I;�I;�I;�I;�$I;:2I;�DI;�\I;~}I;�I;��I;ǷI;��H;�F;8lA;>P6;fo!;���:���: '��4��ɻ��5���ސ�2+��/v�J$��iz�+��W�H���z������j�� ž��Ҿ      J(��$�f��R������~���`���Yb���'��U�J$��G�m�&����ϼ�/��8������X�غ�9�9���:G;	H.;G|=;sE;�\H;V�I;��I;��I;/�I;4gI;7LI;8I;<)I;�I;�I;�I;]I;�I;�I;�I;;)I;8I;7LI;6gI;*�I;��I;��I;X�I;�\H;oE;D|=;	H.;G;���:�9�9T�غ����8���/����ϼ&��G�m�J$���U���'��Yb��`���~�����R��f���$�      >�}���w�#f���K�s,��
�?�׾"�����k���'�iz꽟I���;V�=M�����iO�ZG�NoE�0�����:l� ;ӿ$;ߴ8;��B;/�G;iKI;D�I;J�I;u�I;8qI;�SI;�=I;�-I;<"I;�I;MI;�I;MI;�I;<"I;�-I;�=I;�SI;9qI;r�I;I�I;A�I;kKI;2�G;��B;ݴ8;ҿ$;n� ;���:4��MoE�\G໦iO����=M��;V��I��iz���'���k�"���?�׾�
�s,���K�#f���w�      ��s�������0蒿��w��F�e��Ͱ�"����Yb�+����ѽ�%��D4�ڟ�X������G��~潺@��9�r�: ;:3;KQ@;�vF;M�H;7�I;��I;��I;�zI;�ZI;GCI;�1I;�%I;xI;�I;WI;�I;wI;�%I;�1I;GCI;�ZI;�zI;��I;��I;6�I;K�H;�vF;HQ@;:3; ;�r�:8��9~潺�G�����X��ڟ�D4��%����ѽ+���Yb�"���Ͱ�e���F���w�0蒿����s���      5��������㿌�ɿ���˅����P�e��?�׾�`��W�H����@��T�a���̡���D��ɻ� ��ҭ�X�:�;�I-;Y|=;UCE;ۅH;9�I;�I;��I;�I;�aI;WHI;�5I;�(I; I;I;�I;I; I;�(I;�5I;WHI;�aI;�I;��I;�I;7�I;ۅH;WCE;W|=;�I-;�;X�:�ҭ�� ��ɻ�D�̡����T�a��@����W�H��`��?�׾e����P�˅�������ɿ�㿵���      ș$��x �$��;���޿r���˅���F��
��~����z��$���ս���B2+���ϼPp�����0�]�h�*�P��:>�;9';Ȍ:;+�C;?H;�}I;Q�I;��I;�I;�gI;�LI;P9I;m+I;X"I;*I;]I;*I;X"I;k+I;M9I;�LI;�gI;�I;��I;Q�I;�}I;=H;+�C;Ì:;9';>�;X��:h�*�0�]�����Pp���ϼB2+������ս�$���z��~���
��F�˅��r����޿;��$���x �      L�Q���K���;�ș$��;
��޿�����w�s,���澟���)�D������I��&�G�����N��������������9:���:�n!;��7;�B;��G;ZI;]�I;��I;�I;�lI;�PI;I<I;�-I;F$I;�I;�I;�I;E$I;�-I;H<I;�PI;�lI;�I;��I;\�I;ZI;��G;�B;��7;�n!;���:�9:����������N�����&�G��I������)�D��������s,���w�����޿�;
�ș$���;���K�      U����{���d��F�ș$�;����ɿ0蒿��K�R���j��Zb�G�4���t�a����?�����.��d���غ���9�Y�:iX;�25;S�A;�!G;i7I;��I;��I;|�I;�pI;�SI;�>I;�/I;�%I;T I;cI;T I;�%I;�/I;�>I;�SI;�pI;y�I;~�I;��I;i7I;�!G;U�A;�25;kX;�Y�:���9�غ�d����.�?������u�a�4���G�Zb��j��R����K�0蒿��ɿ;��ș$��F���d��{�      ����$P�������d���;�$���㿴���#f�f�� ž��z���?�ƽ(0v�V5�0����o@�z���Pi�0bu9~K�:R];�73;S�@;,�F;fI;��I;��I;��I;tI;�UI;s@I;1I;'I;?!I;cI;?!I;'I;1I;r@I;�UI;tI;}�I;��I;��I;fI;,�F;S�@;�73;S];|K�:@bu9Pi�z����o@�0���V5�(0v�?�ƽ����z� žf��#f�������$����;���d����$P��      �,��b��$P���{���K��x �����s�����w��$���Ҿh��� (���ѽӷ��(������K�<ɻ�����8���:��;��1;#@;��F;<I;�I;H�I;ԞI;�uI;`WI;�AI;�1I;�'I;�!I;�I;�!I;�'I;�1I;�AI;aWI;�uI;ҞI;E�I;�I;;I;��F;#@;��1;��;���:��8���<ɻߔK����(�ӷ����ѽ (�h�����Ҿ�$���w�s��������x ���K��{�$P��b��      ᶕ�T���Ҭ��/�_���7�|�!}߿����,b��V�0l¾Lx�f.���Ž��t�+��e����?�N�����P�x9���:��;��2;b@@;�fF;M�H;��I;��I;E|I;�[I;�CI;72I;�%I;�I;�I;aI;�I;�I;�%I;62I;�CI;�[I;E|I;��I;��I;M�H;�fF;b@@;��2;��;���:`�x9���N����?�e��+����t���Žf.�Lx�0l¾�V��,b����!}߿|���7�/�_�Ҭ��T���      T���G���&}��+Y��3�����$ڿ'��ƽ\����(���s��3�8����p�d�T���<<�1��T���ؗ�9|��:�;_%3;up@;zF;��H;,�I;%�I;�{I;[I;�CI;�1I;�%I;UI;�I;6I;�I;XI;�%I;�1I;�CI;[I;�{I;"�I;,�I;��H;zF;up@;[%3;�;|��:ؗ�9T���1���<<�T��d��p�8����3��s�(�����ƽ\�'���$ڿ����3��+Y�&}�G���      Ҭ��&}�@tf��lG�آ%��p�1�ʿ\����>M����X�����d�ʤ�̷�1�d��
��I���1�\����� ��9���:W;�U4;��@;�F;L�H;�I;�I;�yI;�YI;rBI;1I;�$I;�I;I;�I;I;�I;�$I;1I;rBI;�YI;�yI;�I;�I;L�H;�F;��@;�U4;Z;���: ��9��\����1��I���
�1�d�̷�ʤ���d�X�������>M�\���1�ʿ�p�آ%��lG�@tf�&}�      /�_��+Y��lG� f.�|���꿳���O䂿��5���󾎰��R�N�X��U��#�Q����|����h!�~g��񳺰	:�
�:(�;r16;��A;�G;I;h�I;��I;�vI;}WI;�@I;�/I;�#I;�I;;I;�I;;I;�I;�#I;�/I;�@I;WI;�vI;��I;h�I;I;�G;��A;n16;+�;�
�:�	:�~g���h!�|������#�Q�U��X��R�N���������5�O䂿�������|� f.��lG��+Y�      ��7��3�آ%�|��<����ſ���Ž\�>����Ͼ����c�3��载z���9�`�Ἑ���z��7}��ct�h�^:�+�:أ#;8;��B;NsG;�%I;��I; �I;0rI;CTI;>I;�-I;C"I;�I;I;�I;I;I;D"I;�-I;>I;ETI;.rI;�I;��I;�%I;NsG;��B;��8;ڣ#;�+�:t�^:�ct��7}��z����`���9��z����c�3�������Ͼ>��Ž\������ſ�<��|�آ%��3�      |�����p������ſ'���Ps���1�4r���d���d�I�шŽ��}�a*�LC���^��B�d�D��E�� �:��;�);<7;;ZD;t�G;xHI;ޝI;ۏI;�lI;"PI;�:I;G+I;O I;�I;�I;^I;�I;�I;O I;G+I;�:I;"PI;�lI;׏I;ܝI;wHI;s�G;XD;77;;�);��;� �:�E�d�D��B��^�LC��a*���}�шŽI��d��d��4r����1��Ps�'����ſ��꿄p����       }߿�$ڿ0�ʿ��������Ps�RX:����)l¾�ǆ���7����:5���Q�����t���75�b������ �8ʼ:��;��.;��=;�EE;�YH;�hI;U�I;�I;TfI;NKI;W7I;u(I;I;"I;�I;�I;�I;"I;I;u(I;Y7I;NKI;RfI;�I;U�I;�hI;�YH;�EE;��=;��.;��;ʼ:� �8���`���75��t������Q�:5�������7��ǆ�)l¾���RX:��Ps��������0�ʿ�$ڿ      ���'��\���O䂿Ž\���1�����J˾띒�H�N�z��K������X�'�e�Ҽ��|��z��n��x��\�&:�P�:ը;�W4;��@;WgF;��H;=�I;P�I;f�I;H_I;FI;93I;S%I;vI;�I;I;�I;I;�I;vI;P%I;:3I;FI;H_I;c�I;P�I;:�I;��H;TgF;�@;�W4;ը;�P�:X�&:x���n���z���|�e�ҼW�'����K���z��H�N�띒��J˾�����1�Ž\�O䂿\���'��      �,b�ƽ\��>M���5�>��4r��)l¾띒�%&W��3�;Sؽ�z��\G����}I����?���̻t�-��	��d��:��;��&;P|9;�C;�dG;�I;l�I;�I;�vI;�WI;]@I;�.I;�!I;�I;�I;I;�I;I;�I;�I;�!I;�.I;]@I;�WI;�vI;�I;j�I;�I;�dG;�C;M|9;��&;��;d��:�	��s�-���̻��?�}I�����\G��z��;Sؽ�3�%&W�띒�)l¾4r��>����5��>M�ƽ\�      �V������������Ͼ�d���ǆ�H�N��3��c�[����\�4��*C���o���	��눻𳺘��9d��:�h;x�/;i�=;mE;)3H;�WI;�I;)�I;�kI;�OI;U:I;*I;RI;�I;%I;�I;�I;�I;%I;�I;QI;*I;V:I;�OI;�kI;)�I;�I;�WI;&3H;jE;h�=;x�/;�h;b��:���9��눻��	��o�*C��4����\�[���cཱི3�H�N��ǆ��d����Ͼ���������      0l¾(��X������������d���7�z��;Sؽ[���d�E*�ekּ,\����'�"���R�`}����:�Z;��#;d=7;]�A;@�F;��H;��I;�I;�I;aI;�GI;%4I;U%I;�I;�I;�I;
I;�	I;~
I;�I;�I;�I;Z%I;&4I;�GI;aI;�I;�I;��I;��H;>�F;Y�A;d=7;��#;�Z;��:H}���R�"����'�,\��dkּD*��d�[��;Sؽz����7��d���������X���(��      Kx��s���d�R�N�c�3�~I����K����z����\�D*��ݼH���.<<���ڻ�V��ct���&:���:lC;�</;{D=;	�D;��G;%9I;��I;֔I;DtI;_VI;�?I;�-I;� I;�I;�I;�
I;,I;HI;,I;�
I;�I;�I;� I;�-I;�?I;]VI;DtI;ӔI;��I;$9I;��G;�D;{D=;�</;kC;���:��&:�ct��V���ڻ-<<�H����ݼD*���\��z��K������~I�c�3�R�N���d��s�      e.��3�ʤ�X����ЈŽ:5�����\G�4��dkּH����xC��>�P6}�଼��x9���:0	;^�&;�;8;��A;џF;߹H;iyI;ŝI;&�I;bfI;�KI;7I;�'I;�I;�I;�I;FI;�I;�I;�I;FI;�I;�I;�I;�'I;7I;�KI;cfI;!�I;ƝI;gyI;۹H;͟F;��A;�;8;]�&;0	;���: �x9ެ��N6}��>��xC�H���dkּ4��\G����:5��ЈŽ��X��ʤ��3�      ��Ž7���̷�T���z����}��Q�W�'����*C��+\��,<<��>�zn��
�� �z��:u��:7�;�'3;��>;�E;�H;�<I;�I;וI;�vI; YI;�AI;�/I;�!I;I;"I;�	I;�I;VI;�I;VI;�I;�	I;#I;I;�!I;�/I;�AI; YI;�vI;ٕI;�I;�<I;�H;�E;��>;�'3;7�;w��:x��:����zn���>�,<<�+\��*C�����W�'��Q���}��z��T��̷�7���      ��t��p�0�d�#�Q��9�`*����e�Ҽ|I���o���'� �ڻP6}��ະ7���:�m�:��;�.;H<;�oC;n7G;��H;�I;�I;
�I;QfI;sLI;,8I;(I;I;�I;�I;~I;�I;� I;� I;� I;�I;I;�I;�I;I;(I;*8I;sLI;OfI;�I;�I; �I;��H;n7G;�oC;H<;�.;��;�m�:��:�7���P6}� �ڻ��'��o�|I��e�Ҽ���`*��9�#�Q�0�d��p�      *��d��
����_��KC���t����|���?���	�!���V�ެ�� ���:�:�h;E�+;�9;��A;�fF;��H;�_I;��I;ˑI;8sI;�VI;�@I;/I; !I;�I;@I;I;�I;� I;��H;<�H;��H;� I;�I;I;AI;�I;!!I;/I;�@I;�VI;8sI;ʑI;��I;�_I;��H;�fF;��A;�9;H�+;�h;�:��:��ڬ���V� ����	���?���|��t��JC��_������
�d�      d��R���I��{�������^��75��z���̻�눻�R��ct� �x9x��:�m�:�h;��*;�8;�@;�E;i(H;�8I;��I;I�I;�~I;�`I;�HI;�5I;�&I;�I;lI;/
I;�I;� I;%�H;��H;�H;��H;%�H;� I;�I;0
I;lI;�I;�&I;�5I;�HI;�`I;�~I;D�I;�I;�8I;h(H;�E;�@;�8;��*;�h;�m�:x��: �x9�ct��R��눻��̻�z��75��^����{����I��S��      ��?��<<���1��h!��z��B�`���n��r�-��@}����&:���:q��:��;D�+;�8;e�@;^E;��G;wI;�I;��I;g�I;�iI;pPI;<<I;�+I;�I;�I;�I;`I;�I;�H;��H;��H;�H;��H;��H;�H;�I;bI;�I;�I;�I;�+I;:<I;pPI;�iI;c�I;��I;�I;tI;��G;^E;f�@; �8;D�+;��;u��:���:��&:@}���p�-��n��`���B黶z��h!� �1��<<�      N��.��U���|g���7}�^�D�{��x��p	�����9��:���:0	;9�;�.;�9;�@;^E;��G;qI;�I;8�I;��I;�pI;�VI;�AI;�0I;�"I;�I;"I;%I;�I;��H;��H;��H;��H;�H;��H;��H;��H;��H;�I;%I;I;�I;�"I;�0I;�AI;�VI;�pI;|�I;9�I;
�I;rI;��G;^E;�@;�9;�.;9�;0	;���:��:���9p	��x��~��Y�D��7}�|g��U���.��      ���*��������ct��Eเ �8L�&:d��:d��:�Z;iC;[�&;�'3;E<;��A;�E;��G;oI;�|I;��I;ԐI;�uI;�[I;AFI;�4I;d&I;�I;�I;
I;)I;n�H;��H;l�H;��H;��H;U�H;��H;��H;l�H;��H;o�H;)I;
I;I;�I;`&I;�4I;AFI;�[I;�uI;ԐI;�I;�|I;nI;��G;�E;��A;C<;�'3;[�&;iC;�Z;b��:d��:P�&:� �8�E��ct�����D���      ��x9X��9H��9�	:X�^:� �:ʼ:�P�:��;�h;��#;�</;�;8;��>;�oC;�fF;i(H;xI;�I;��I;�I;0xI;�^I;qII;�7I;B)I;CI;�I;�I;�I;� I;}�H;��H;o�H;��H;��H;��H;��H;��H;n�H;��H;~�H;� I;I;�I;�I;@I;@)I;�7I;lII;�^I;1xI;ߑI;��I;�I;xI;h(H;�fF;�oC;��>;�;8;�</;��#;�h;��;�P�:ʼ:� �:X�^:�	:X��9ؗ�9      ���:���:���:�
�:�+�:��;��;ܨ;��&;x�/;h=7;|D=;��A;�E;o7G;��H;�8I;�I;8�I;֐I;0xI;�_I;KI;�9I;-+I;6I;pI;qI;�I;tI;8�H;��H;R�H;s�H;�H;D�H;�H;D�H;�H;s�H;O�H;��H;9�H;pI;�I;sI;lI;6I;0+I;�9I;KI;�_I;-xI;אI;8�I;�I;�8I;��H;q7G;�E;��A;|D=;g=7;x�/;��&;ܨ;��;��;�+�:�
�:���:���:      ��;�;Z;$�;ң#;�);��.;�W4;T|9;i�=;]�A;	�D;ϟF;�H;��H;�_I;�I;��I;��I;�uI;�^I;KI;\:I;W,I;r I;�I;�I;�I;[I;��H;:�H;j�H;C�H;��H;��H;��H;��H;��H;��H;��H;@�H;j�H;:�H;��H;YI;�I;�I;�I;s I;Q,I;Y:I;KI;�^I;�uI;��I;��I;�I;�_I;��H;�H;ϟF;	�D;Z�A;h�=;S|9;�W4;��.;�);ڣ#;!�;[;�;      Ǽ2;s%3;�U4;v16;č8;:7;;��=;�@;�C;mE;C�F;��G;ܹH;�<I;�I;��I;H�I;j�I;�pI;�[I;mII;�9I;T,I;� I;UI;YI;�I;I;��H;��H;��H;_�H;u�H;�H;#�H;��H;8�H;��H;$�H;�H;r�H;b�H;��H;��H;�H;I;�I;WI;VI;� I;Q,I;�9I;iII;�[I;�pI;j�I;F�I;��I;�I;�<I;ܹH;��G;@�F;lE;�C;�@;��=;<7;;ɍ8;r16;�U4;e%3;      k@@;�p@;��@;��A;��B;]D;�EE;SgF;�dG;(3H;��H;%9I;gyI;�I;�I;͑I;�~I;�iI;�VI;GFI;�7I;2+I;v I;ZI;�I;�I;xI;��H;�H;��H;X�H;W�H;��H;��H;��H;V�H;3�H;V�H;��H;��H;��H;Y�H;X�H;��H;�H;��H;vI;�I;�I;WI;v I;2+I;�7I;GFI;�VI;�iI;�~I;ˑI;�I;�I;eyI;'9I;��H;%3H;�dG;SgF;�EE;]D;��B;��A;��@;�p@;      �fF;zF;�F;�G;LsG;o�G;�YH;��H;�I;�WI;��I; �I;I;וI;	�I;6sI;�`I;oPI;�AI;�4I;?)I;4I;�I;YI;�I;�I;&�H;;�H;�H;��H;j�H;��H;P�H;e�H;��H;G�H;K�H;F�H;��H;d�H;L�H;��H;j�H;��H;�H;:�H;#�H;�I;�I;VI;�I;4I;;)I;�4I;�AI;oPI;�`I;5sI;	�I;וI;I;��I;��I;�WI;�I;��H;�YH;m�G;RsG;�G;�F;zF;      ^�H;��H;L�H;#I;�%I;|HI;�hI;:�I;q�I;�I;�I;ؔI;$�I;�vI;RfI;�VI;�HI;;<I;�0I;d&I;CI;pI;�I;�I;tI;)�H;@�H; �H;��H;n�H;��H;.�H;�H;C�H;��H;L�H;L�H;L�H;��H;@�H;�H;-�H;��H;m�H;��H;"�H;=�H;%�H;uI;�I;�I;pI;BI;d&I;�0I;;<I;�HI;�VI;QfI;�vI;$�I;ؔI;�I;�I;q�I;:�I;�hI;xHI;�%I;#I;K�H;��H;      ��I;/�I;�I;d�I;ߙI;ޝI;X�I;U�I;��I;0�I;�I;JtI;cfI;YI;vLI;�@I;�5I;�+I;�"I;�I;�I;tI;�I;	I;��H;=�H;"�H;��H;��H;��H; �H;��H;��H;9�H;��H;z�H;a�H;z�H;��H;9�H;��H;��H;�H;��H;}�H;��H; �H;;�H;��H;I;�I;sI;�I;�I;�"I;�+I;�5I;�@I;vLI;YI;cfI;JtI;�I;/�I;��I;X�I;X�I;ܝI;�I;e�I;�I;<�I;      ��I;%�I;�I;��I;�I;؏I;�I;g�I;�vI;�kI;aI;bVI;�KI;�AI;-8I;/I;�&I;�I;�I;�I;�I;�I;[I;��H;�H;�H;��H;��H;��H;�H;��H;��H;��H;`�H;�H;��H;��H;��H;�H;`�H;��H;��H;��H;�H;��H;�H;��H;�H;�H;��H;XI;�I;�I;�I;�I;�I;�&I;/I;-8I;�AI;�KI;`VI;aI;�kI;�vI;g�I;�I;؏I;$�I;��I;�I;�I;      P|I;�{I;�yI;�vI;>rI;�lI;XfI;N_I;�WI;�OI;�GI;�?I;�7I;�/I;(I;$!I;�I;�I;"I;
I;�I;sI;��H;��H;��H;��H;m�H;��H;�H;��H;��H;��H;7�H;��H;G�H;�H; �H;�H;G�H;��H;5�H;��H;��H;��H;�H;��H;k�H;��H;��H;��H;��H;sI;�I;
I;!I;�I;�I;#!I;(I;�/I;�7I;�?I;�GI;�OI;�WI;P_I;XfI;�lI;;rI;�vI;�yI;�{I;       \I;�[I;�YI;�WI;PTI;"PI;UKI;FI;e@I;]:I;-4I;�-I;�'I;�!I;I;�I;tI;�I;*I;.I;� I;;�H;=�H;��H;T�H;m�H;��H;#�H;��H;��H;��H;�H;��H;�H;��H;��H;��H;��H;��H;�H;��H;�H;��H;��H;��H;#�H;��H;k�H;W�H;��H;:�H;9�H;� I;-I;)I;�I;qI;�I;I;�!I;�'I;�-I;,4I;]:I;g@I;FI;UKI;"PI;MTI;�WI;�YI;�[I;      �CI;�CI;zBI;�@I;>I;�:I;Z7I;@3I;�.I;*I;^%I;� I;�I;I;�I;GI;9
I;cI;�I;v�H;��H;��H;n�H;f�H;W�H;��H;-�H;��H;��H;��H;�H;�H;��H;��H;N�H;�H;�H;�H;N�H;��H;��H;��H;�H;��H;��H;��H;-�H;��H;Z�H;f�H;m�H;��H;��H;v�H;�I;cI;7
I;GI;�I;I;�I;� I;^%I;*I;�.I;@3I;Y7I; ;I;>I;�@I;xBI;�CI;      :2I;�1I;1I;�/I;�-I;E+I;u(I;U%I;�!I;TI;�I;�I; I;)I;�I;I;�I;�I;��H;��H;��H;S�H;D�H;{�H;��H;O�H;�H;��H;��H;;�H;��H;��H;m�H;'�H;��H;��H;��H;��H;��H;'�H;j�H;��H;��H;<�H;��H;��H;�H;M�H;��H;{�H;C�H;S�H;��H;��H;��H;�I;�I;I;�I;)I;�I;�I;�I;UI;�!I;U%I;u(I;G+I;�-I;�/I;1I;�1I;      �%I;�%I;�$I;�#I;N"I;I I;I;�I;�I;�I;�I;�I;�I;�	I;�I;�I;� I;�H;��H;s�H;x�H;v�H;��H;�H;��H;d�H;@�H;9�H;^�H;��H;�H;��H;!�H;��H;��H;x�H;\�H;x�H;��H;��H; �H;��H;�H;��H;a�H;9�H;@�H;c�H;��H;	�H;��H;v�H;v�H;s�H;��H;�H;� I;�I;�I;�	I;�I;�I;�I;�I;�I;�I;I;L I;D"I;�#I;�$I;�%I;      �I;iI;�I;�I;�I;�I;&I;�I;�I;)I;�I;�
I;LI;�I;�I;� I;0�H;��H;��H;��H;��H;�H;��H;(�H;��H;��H;��H;��H;�H;G�H;��H;Q�H;��H;��H;M�H;B�H;J�H;B�H;M�H;��H;��H;T�H;��H;H�H;�H;��H;��H;��H;��H;'�H;��H;�H;��H;��H;��H;��H;/�H;� I;�I;�I;LI;�
I;�I;*I;�I;�I;&I;�I;�I;�I;�I;aI;      �I;�I;I;>I;(I;�I;�I;I;I;�I;�
I;5I;�I;aI;I;��H;��H;��H;��H;��H;��H;G�H;��H;��H;R�H;C�H;J�H;|�H;��H;�H;��H;�H;��H;}�H;B�H;*�H;&�H;+�H;B�H;z�H;��H;!�H;��H;�H;��H;|�H;I�H;A�H;S�H;��H;��H;G�H;��H;��H;��H;��H;��H;��H;I;`I;�I;7I;�
I;�I;I;I;�I;�I;I;=I;I;�I;      ^I;>I;�I;�I;�I;\I;�I;�I;�I;�I;�	I;PI;�I;�I;� I;D�H; �H;�H;�H;[�H;��H;!�H;��H;<�H;2�H;F�H;I�H;e�H;��H;�H;��H;�H;��H;b�H;J�H;'�H;�H;'�H;J�H;b�H;��H;�H;��H;�H;��H;e�H;G�H;G�H;2�H;:�H;��H;!�H;��H;[�H;�H;�H;�H;D�H;� I;�I;�I;PI;�	I;�I;�I;�I;�I;`I;�I;�I;�I;6I;      �I;�I;I;=I;(I;�I;�I;I;I;�I;�
I;7I;�I;`I;I;��H;��H;��H;��H;��H;��H;G�H;��H;��H;S�H;C�H;J�H;|�H;��H;�H;��H;�H;��H;}�H;B�H;*�H;&�H;+�H;B�H;z�H;��H;!�H;��H;�H;��H;|�H;I�H;A�H;R�H;��H;��H;G�H;��H;��H;��H;��H;��H;��H;I;`I;�I;7I;�
I;�I;I;I;�I;�I;I;>I;I;�I;      �I;iI;�I;�I;�I;�I;&I;�I;�I;)I;�I;�
I;MI;�I;�I;� I;/�H;��H;��H;��H;��H;�H;��H;(�H;��H;��H;��H;��H;�H;G�H;��H;Q�H;��H;��H;M�H;B�H;J�H;B�H;M�H;��H;��H;U�H;��H;H�H;�H;��H;��H;��H;��H;&�H;��H;�H;��H;��H;��H;��H;/�H;� I;�I;�I;MI;�
I;�I;*I;�I;�I;&I;�I;�I;�I;�I;aI;      �%I;�%I;�$I;�#I;M"I;I I;I;�I;�I;�I;�I;�I;�I;�	I;�I;�I;� I;�H;��H;s�H;y�H;v�H;��H;�H;��H;d�H;@�H;9�H;^�H;��H;�H;��H;!�H;��H;��H;x�H;\�H;x�H;��H;��H; �H;��H;�H;��H;a�H;9�H;@�H;d�H;��H;	�H;��H;v�H;v�H;s�H;��H;�H;� I;�I;�I;�	I;�I;�I;�I;�I;�I;�I;I;M I;A"I;�#I;�$I;�%I;      =2I;�1I;1I;�/I;�-I;E+I;u(I;T%I;�!I;TI;�I;�I;�I;(I;�I;I;�I;�I;��H;��H;��H;S�H;D�H;{�H;��H;O�H;�H;��H;��H;;�H;��H;��H;k�H;%�H;��H;��H;��H;��H;��H;%�H;j�H;��H;��H;<�H;��H;��H;�H;M�H;��H;y�H;C�H;S�H;��H; �H;��H;�I;�I;I;�I;)I;�I;�I;�I;UI;�!I;T%I;u(I;G+I;�-I;�/I;1I;�1I;      �CI;�CI;xBI;�@I;>I;�:I;]7I;A3I;�.I;*I;^%I;� I;�I;I;�I;GI;9
I;bI;�I;x�H;��H;��H;n�H;f�H;Z�H;��H;-�H;��H;��H;��H;�H;�H;��H;��H;N�H;�H;�H;�H;N�H;��H;��H;��H;�H;��H;��H;��H;-�H;��H;W�H;f�H;m�H;��H;��H;v�H;�I;dI;7
I;GI;�I;I;�I;� I;^%I; *I;�.I;A3I;]7I;�:I;>I;�@I;xBI;�CI;       \I;�[I;�YI;�WI;QTI;"PI;UKI;FI;g@I;\:I;-4I;�-I;�'I;�!I;I;�I;qI;�I;)I;-I;� I;9�H;=�H;��H;W�H;m�H;��H;#�H;��H;��H;��H;�H;��H;�H;��H;��H;��H;��H;��H;�H;��H;�H;��H;��H;��H;#�H;��H;j�H;T�H;��H;:�H;;�H;� I;.I;*I;�I;sI;�I;I;�!I;�'I;�-I;,4I;_:I;e@I;FI;UKI;"PI;OTI;�WI;�YI;�[I;      J|I;�{I;�yI;�vI;:rI;�lI;XfI;N_I;�WI;�OI;�GI;�?I;�7I;�/I;(I;#!I;�I;�I;!I;
I;�I;sI;��H;��H;��H;��H;m�H;��H;�H;��H;��H;��H;7�H;��H;G�H;�H; �H;�H;G�H;��H;7�H;��H;��H;��H;�H;��H;k�H;��H;��H;��H;��H;sI;�I;
I;"I;�I;�I;&!I;(I;�/I;�7I;�?I;�GI;�OI;�WI;R_I;YfI;�lI;;rI;�vI;�yI;�{I;      ��I;!�I;�I;��I;#�I;ՏI;��I;g�I;�vI;�kI;aI;bVI;�KI;�AI;-8I;/I;�&I;�I;�I;�I;�I;�I;YI;��H;�H;�H;��H;�H;��H;�H;��H;��H;��H;`�H;�H;��H;��H;��H;�H;`�H;��H;��H;��H;�H;��H;��H;��H;�H;�H;��H;YI;�I;�I;�I;�I;�I;�&I;/I;-8I;�AI;�KI;bVI;aI;�kI;�vI;i�I;�I;؏I;!�I;��I;�I;"�I;      ��I;2�I;�I;e�I;��I;ޝI;X�I;W�I;��I;/�I;�I;JtI;cfI;YI;vLI;�@I;�5I;�+I;�"I;�I;�I;sI;�I;I;��H;;�H; �H;��H;�H;��H;�H;��H;��H;8�H;��H;z�H;a�H;z�H;��H;9�H;��H;��H; �H;��H;�H;��H;"�H;=�H;��H;I;�I;tI;�I;�I;�"I;�+I;�5I;�@I;vLI;YI;cfI;HtI;�I;0�I;��I;Y�I;X�I;۝I;�I;d�I;�I;:�I;      X�H;��H;I�H;I;�%I;xHI;�hI;:�I;q�I;�I;�I;ؔI;$�I;�vI;QfI;�VI;�HI;;<I;�0I;f&I;FI;pI;�I;�I;uI;(�H;@�H;"�H;��H;n�H;��H;-�H;�H;@�H;��H;L�H;L�H;J�H;��H;A�H;�H;.�H;��H;m�H;��H; �H;>�H;(�H;tI;�I;�I;pI;@I;d&I;�0I;<<I;�HI;�VI;RfI;�vI;$�I;ؔI;�I;�I;q�I;<�I;�hI;wHI;�%I;I;G�H;��H;      �fF;zF;�F;�G;NsG;o�G;�YH;��H;�I;�WI;��I;��I;I;וI;�I;6sI;�`I;nPI;�AI;�4I;?)I;4I;�I;WI;�I;�I;%�H;:�H;�H;��H;j�H;��H;M�H;d�H;��H;G�H;K�H;G�H;��H;e�H;M�H;��H;j�H;��H;�H;;�H;%�H;�I;�I;VI;�I;4I;;)I;�4I;�AI;pPI;�`I;6sI;	�I;וI;I; �I;��I;�WI;�I;��H;�YH;m�G;RsG;�G;�F;zF;      k@@;�p@;��@;��A;��B;]D;�EE;SgF;�dG;&3H;��H;'9I;eyI;�I;�I;͑I;�~I;�iI;�VI;GFI;�7I;2+I;v I;ZI;�I;�I;xI;��H;�H;��H;X�H;W�H;��H;��H;��H;V�H;3�H;V�H;��H;��H;��H;Z�H;X�H;��H;�H;��H;vI;�I;�I;YI;u I;2+I;�7I;HFI;�VI;�iI;�~I;͑I;�I;�I;gyI;%9I;��H;&3H;�dG;TgF;�EE;^D;��B;��A;��@;p@;      ͼ2;o%3;�U4;p16;��8;@7;;��=;�@;�C;oE;B�F;��G;޹H;�<I;�I;��I;H�I;g�I;�pI;�[I;lII;�9I;S,I;� I;VI;YI;�I;I;��H;��H;��H;a�H;t�H;�H;!�H;��H;8�H;��H;$�H;�H;t�H;a�H;��H;��H;~�H;I;�I;YI;UI;� I;S,I;�9I;jII;�[I;�pI;k�I;F�I;��I;�I;�<I;ܹH;��G;B�F;lE;�C;�@;��=;>7;;΍8;r16;�U4;d%3;      ��;�;h;!�;ѣ#;�);��.;�W4;T|9;i�=;Z�A;	�D;ΟF;�H;��H;�_I;�I;��I;��I;�uI;�^I;KI;[:I;V,I;s I;�I;�I;�I;[I;��H;:�H;j�H;@�H;��H;��H;��H;��H;��H;��H;��H;B�H;j�H;:�H;��H;YI;�I;�I;�I;r I;S,I;\:I;KI;�^I;�uI;��I;��I;��I;�_I;��H;�H;ΟF;	�D;]�A;g�=;T|9;�W4;��.;�);֣#;"�;^;�;      ���:���:���:�
�:�+�:��;��;ܨ;��&;x�/;h=7;|D=;��A;�E;o7G;��H;�8I;�I;8�I;֐I;0xI;�_I;KI;�9I;0+I;6I;pI;sI;�I;tI;9�H;��H;P�H;s�H;�H;E�H;�H;D�H;�H;s�H;P�H;��H;8�H;pI;�I;qI;lI;6I;-+I;�9I;KI;�_I;.xI;אI;8�I;�I;�8I;��H;q7G;�E;��A;~D=;h=7;x�/;��&;ݨ;��;��;�+�:�
�:���:���:      ��x9 ��9x��9�	:T�^:� �:!ʼ:�P�:��;�h;��#;�</;�;8;��>;�oC;�fF;i(H;wI;�I;��I;�I;1xI;�^I;pII;�7I;B)I;BI;�I;�I;�I;� I;}�H;��H;m�H;��H;��H;��H;��H;��H;o�H;��H;}�H;� I;I;�I;�I;@I;B)I;�7I;lII;�^I;0xI;ߑI;��I;�I;yI;i(H;�fF;�oC;��>;�;8;�</;��#;�h;��;�P�:#ʼ:� �:p�^:�	:p��9ؗ�9      ���0��������ct��E�� �8P�&:f��:d��:�Z;iC;[�&;�'3;C<;��A;�E;��G;nI;�|I;��I;ԐI;�uI;�[I;AFI;�4I;d&I;�I;�I;
I;)I;n�H;��H;l�H;��H;��H;U�H;��H;��H;l�H;��H;o�H;)I;
I;I;�I;`&I;�4I;AFI;�[I;�uI;ԐI;�I;�|I;oI;��G;�E;��A;C<;�'3;[�&;hC;�Z;b��:f��:\�&:� �8�E��ct�����D���      N��.��U���|g���7}�^�D�~��x��x	�����9��:���:0	;9�;�.;�9;�@;^E;��G;qI;�I;9�I;��I;�pI;�VI;�AI;�0I;�"I;�I;"I;%I;�I;��H;��H;��H;��H;�H;��H;��H;��H;��H;�I;%I;I;�I;�"I;�0I;�AI;�VI;�pI;|�I;8�I;
�I;rI;��G;^E;�@;�9;�.;9�;0	;���:��:���9p	��x��{��Z�D�~7}�|g��T���.��      ��?��<<� �1��h!��z��B�`���n��r�-��@}����&:���:q��:��;D�+;�8;e�@;^E;��G;wI;�I;��I;g�I;�iI;oPI;<<I;�+I;�I;�I;�I;`I;�I;�H;��H;��H;�H;��H;��H;�H;�I;bI;�I;�I;�I;�+I;:<I;rPI;�iI;c�I;��I;�I;tI;��G;^E;f�@; �8;D�+;��;q��:���:��&:@}���p�-��n��`���B黶z��h!� �1��<<�      d��R���I��{�������^��75��z���̻�눻�R��ct� �x9x��:�m�:�h;��*;�8;�@;�E;i(H;�8I;��I;H�I;�~I;�`I;�HI;�5I;�&I;�I;lI;0
I;�I;� I;%�H;��H;�H;��H;'�H;� I;�I;/
I;lI;�I;�&I;�5I;�HI;�`I;�~I;D�I;�I;�8I;h(H;�E;�@;�8;��*;�h;�m�:x��: �x9�ct��R��눻��̻�z��75��^����{����I��S��      *��c��
����_��KC���t����|���?���	� ���V�ڬ�� ���:�:�h;G�+;�9;��A;�fF;��H;�_I;��I;ʑI;6sI;�VI;�@I;/I;!!I;�I;@I;I;�I;� I;��H;<�H;��H;� I;�I;I;@I;�I; !I;/I;�@I;�VI;8sI;ˑI;��I;�_I;��H;�fF;��A;�9;G�+;�h;�:��: �ެ���V�!����	���?���|��t��JC��_������
�d�      ��t��p�0�d�#�Q��9�`*����e�Ҽ|I���o���'� �ڻP6}��ະ7���:�m�:��;�.;F<;�oC;n7G;��H;�I;�I;�I;QfI;sLI;.8I;(I;I;�I;�I;I;�I;� I;� I;� I;�I;I;�I;�I;I;(I;)8I;sLI;OfI;�I;�I; �I;��H;n7G;�oC;I<;�.;��;�m�:��:�7���P6}� �ڻ��'��o�|I��e�Ҽ���`*��9�#�Q�0�d��p�      ��Ž7���̷�T���z����}��Q�W�'����*C��+\��-<<��>�zn������z��:w��:7�;�'3;��>;�E;�H;�<I;�I;֕I;�vI; YI;�AI;�/I;�!I;I;#I;�	I;�I;VI;�I;VI;�I;�	I;!I;I;�!I;�/I;�AI; YI;�vI;ٕI;�I;�<I;�H;�E;��>;�'3;7�;y��:x��: �
��zn���>�,<<�+\��*C�����W�'��Q���}��z��T��̷�7���      e.��3�ʤ�X����ЈŽ:5�����\G�4��dkּH����xC��>�N6}�଼��x9���:0	;]�&;�;8;��A;џF;߹H;gyI;ŝI;&�I;cfI;�KI;7I;�'I;�I;�I;�I;FI;�I;�I;�I;FI;�I;�I;�I;�'I;7I;�KI;bfI;!�I;ȝI;iyI;ڹH;͟F;��A;�;8;]�&;0	;���: �x9଼�P6}��>��xC�H���dkּ4��\G����:5��ЈŽ��X��ʤ��3�      Kx��s���d�R�N�b�3�~I����K����z����\�D*��ݼH���.<<���ڻ�V��ct���&:���:kC;�</;{D=;	�D;��G;$9I; �I;֔I;DtI;_VI;�?I;�-I;� I;�I;�I;�
I;-I;HI;-I;�
I;�I;�I;� I;�-I;�?I;]VI;DtI;ӔI;��I;%9I;��G;�D;{D=;�</;kC;���:��&:�ct���V���ڻ.<<�H����ݼD*���\��z��K������~I�b�3�R�N���d��s�      0l¾(��X������������d���7�z��;Sؽ[���d�E*�ekּ,\����'�"���R�X}����:�Z;��#;d=7;]�A;@�F;��H;��I;�I;�I;aI;�GI;&4I;U%I;�I;�I;�I;
I;�	I;
I;�I;�I;�I;W%I;%4I;�GI;aI;�I;�I;��I;��H;>�F;Y�A;d=7;��#;�Z;��:H}���R�#����'�,\��ekּE*��d�[��;Sؽz����7��d���������X���(��      �V������������Ͼ�d���ǆ�H�N��3��c�[����\�4��*C���o���	��눻𳺘��9d��:�h;x�/;k�=;mE;&3H;�WI;�I;)�I;�kI;�OI;V:I;*I;RI;�I;%I;�I;�I;�I;%I;�I;QI;*I;U:I;�OI;�kI;)�I;�I;�WI;)3H;jE;h�=;x�/;�h;b��:���9��눻��	��o�*C��4����\�[���cཱི3�H�N��ǆ��d����Ͼ���������      �,b�ƽ\��>M���5�>��4r��)l¾띒�%&W��3�;Sؽ�z��\G����}I����?���̻t�-��	��f��:��;��&;P|9;�C;�dG;�I;l�I;�I;�vI;�WI;]@I;�.I;�!I;�I;�I;I;�I;I;�I;�I;�!I;�.I;]@I;�WI;�vI;�I;j�I;�I;�dG;�C;M|9;��&;��;`��:�	��r�-���̻��?�}I�����\G��z��;Sؽ�3�%&W�띒�)l¾4r��>����5��>M�ƽ\�      ���'��\���O䂿Ž\���1�����J˾띒�H�N�z��K������W�'�e�Ҽ��|��z��n��x��\�&:�P�:ը;�W4;�@;TgF;��H;<�I;P�I;f�I;H_I;FI;:3I;Q%I;xI;�I;I;�I;I;�I;xI;Q%I;93I;FI;H_I;c�I;P�I;:�I;��H;WgF;�@;�W4;ը;�P�:X�&:x���n���z���|�f�ҼX�'����K���z��H�N�띒��J˾�����1�Ž\�O䂿\���'��       }߿�$ڿ0�ʿ��������Ps�RX:����)l¾�ǆ���7����:5���Q�����t���75�a������ �8ʼ:��;��.;��=;�EE;�YH;�hI;U�I;�I;RfI;NKI;W7I;v(I;I;"I;�I;�I;�I;"I;I;s(I;W7I;NKI;RfI;�I;U�I;�hI;�YH;�EE;��=;��.;��;ʼ:� �8���`���75��t������Q�:5�������7��ǆ�)l¾���RX:��Ps��������0�ʿ�$ڿ      |�����p������ſ'���Ps���1�4r���d���d�I�шŽ��}�a*�LC���^��B�d�D��E๼ �:��;�);<7;;XD;t�G;xHI;ܝI;ۏI;�lI;"PI;�:I;H+I;O I;�I;�I;^I;�I;�I;O I;E+I;�:I;"PI;�lI;׏I;ޝI;wHI;s�G;ZD;77;;�);��;� �:�E�d�D��B��^�LC��a*���}�шŽI��d��d��4r����1��Ps�'����ſ��꿄p����      ��7��3�آ%�|��<����ſ���Ž\�>����Ͼ����c�3��载z���9�`�Ἑ���z��7}��ct�h�^:�+�:أ#;č8;��B;OsG;�%I;��I;!�I;1rI;ETI;>I;�-I;D"I;�I;I;�I;I;I;C"I;�-I;>I;CTI;.rI;�I;��I;�%I;LsG;��B;��8;ڣ#;�+�:p�^:�ct��7}��z����`���9��z����c�3�������Ͼ>��Ž\������ſ�<��|�آ%��3�      /�_��+Y��lG� f.�|���꿳���O䂿��5���󾎰��R�N�X��U��#�Q����|����h!�~g��񳺨	:�
�:(�;r16;��A;�G;I;h�I;��I;�vI;WI;�@I;�/I;�#I;�I;;I;�I;;I;�I;�#I;�/I;�@I;}WI;�vI;��I;h�I;I;�G;��A;l16;+�;�
�:�	:�~g���h!�|������#�Q�U��X��R�N���������5�O䂿�������|� f.��lG��+Y�      Ҭ��&}�@tf��lG�آ%��p�1�ʿ\����>M����X�����d�ʤ�̷�1�d��
��I���1�\�������9���:W;�U4;��@;�F;L�H;�I;�I;�yI;�YI;rBI;1I;�$I;�I;I;�I;I;�I;�$I;1I;rBI;�YI;�yI;�I;�I;L�H;�F;��@;�U4;Z;���: ��9��\����1��I��	�
�1�d�̷�ʤ���d�X�������>M�\���1�ʿ�p�آ%��lG�@tf�&}�      T���G���&}��+Y��3�����$ڿ'��ƽ\����(���s��3�8����p�d�T���<<�1��R���ؗ�9|��:�;a%3;up@;zF;��H;,�I;%�I;�{I;[I;�CI;�1I;�%I;UI;�I;6I;�I;XI;�%I;�1I;�CI;[I;�{I;"�I;,�I;��H;zF;up@;]%3;�;|��:ؗ�9T���1���<<�T��d��p�8����3��s�(�����ƽ\�'���$ڿ����3��+Y�&}�G���      �Aq���i���U�I:�@�����=���x���}A�f5�� ���^Z�����A���]�����d��J",��5��b�Ѻx��9��:_�;dY4;s�@;�VF;��H;�GI;�bI;=OI;M:I;	*I;OI;�I;�I;�I;�I;�I;�I;�I;NI;*I;M:I;<OI;�bI;�GI;��H;�VF;s�@;bY4;b�;��:���9d�Ѻ�5��J",��d������]��A������^Z�� ��f5�}A�x���=�������@�I:���U���i�      ��i���b�\�O�.5�4i�������������q<����f��c
V�IE	�!���IY�k9�D�����(��R����Ⱥ|�:{��:"�;K�4;m�@;ohF;ŗH;@II;�bI;�NI;�9I;�)I;I;�I;�I;�I;�I;�I;�I;�I;I;�)I;�9I;�NI;�bI;@II;ŗH;ohF;m�@;F�4;(�;{��:|�:��Ⱥ�R����(�E���k9��IY�!��IE	�c
V�f������q<������������4i�.5�\�O���b�      ��U�\�O�J-?�0�'���O�ῶ欿c�{�ha/���뾟���I����f���ZN�`5������;H�\ �������":��:��;��5;�`A;��F;a�H;FMI;&bI;�MI;�8I;)I;qI;I;rI;8I;7I;8I;qI;I;pI;)I;�8I;�MI;$bI;FMI;a�H;��F;�`A;��5;��;��:��":���\ ��;H�����`5���ZN�f������I�������ha/�c�{��欿O����0�'�J-?�\�O�      I:�.5�0�'� ������lȿ���m$_���Z�Ҿޕ���6�����*���`=�?�漮)��HG�6��`��X�Q:��:0";�7;�&B;�F;��H;SI;�`I;�KI;O7I;�'I;lI;LI;�I;�I;�
I;�I;�I;LI;kI;�'I;O7I;�KI;�`I;SI;��H;�F;�&B;�7;0";��:d�Q:d��6��GG��)��?���`=��*������6�ޕ��Z�Ҿ��m$_����lȿ���� ��0�'�.5�      @�4i�������K�ѿm������q<��:��a����q����Wн齅���'�Wb̼�zl��.��;�X�����:��;�&;ܫ9;TC;MG;�H;hYI;�^I;�HI;5I;&I;I;;I;�I;�
I;�	I;�
I;�I;;I;I;&I;5I;�HI;�^I;hYI;	�H;}MG;RC;٫9;
�&;��;�:���;�X��.���zl�Wb̼��'�齅��Wн����q��a���:��q<���m���K�ѿ������4i�      �������O��lȿm���������O���}]׾}����I�����A��A�d�o�֮�
RH��jλ;�$�&����:dN;ʆ+;�<;*4D;�G;�I;�^I;�[I;EI;T2I;�#I;qI;�I;�I;�	I;�I;�	I;�I;�I;qI;�#I;T2I;EI;�[I;�^I;�I;�G;)4D;�<;ʆ+;dN;���:0&�;�$��jλRH�֮�o�A�d��A������I�}���}]׾����O�����m���lȿO�Ῥ��      =��������欿�������O��x����� ���l���"��ܽ���`=����v���k"�%R��ۺ ��9�?�:|L;��0;П>;�ME;�#H;�%I;bI;6WI;�@I;%/I;q!I;mI;7I;@I;~I;�I;~I;@I;5I;nI;s!I;%/I;�@I;3WI;bI;�%I;�#H;�ME;̟>;��0;|L;�?�:�9ۺ$R���k"�v������`=����ܽ��"��l�� ����뾃x���O�������欿����      x�������c�{�m$_��q<������~��
w���6�����!���h����䷾�� d�w.���^e��H[�x�Z:���:�, ;��5;�A;WF;ׄH;AI;�bI;�QI;<I;r+I;�I;=I;kI;�	I;I;bI;I;�	I;kI;<I;�I;q+I;<I;�QI;�bI;AI;քH;�VF;�A;��5;�, ;���:x�Z:�H[��^e�x.��� d�䷾�����h�!�������6�
w��~��������q<�m$_�c�{�����      }A��q<�ha/����:�}]׾� ��
w��>�FE	�����ܽ����3�`�꼙���",��W��I���Q�ϰ�:�M
;�f);�:;L@C;#@G;��H;sTI;�_I;[KI;7I;�'I;�I;�I;oI;I;�I;�I;�I;I;pI;�I;�I;'I;7I;XKI;�_I;oTI;��H; @G;I@C;��:;�f);�M
;˰�:�Q�H���W��",�����`�꼜�3�ܽ������FE	�>�
w��� ��}]׾�:���ha/��q<�      f5�������Z�Ҿ�a��}����l��6�FE	���Ƚk���aG����f֮��W����U�k���$d,:���:�;��1;r�>;dE;V�G;QI;T_I;uZI;kDI;�1I;d#I;uI;*I;6
I;=I;I;SI;I;?I;7
I;)I;vI;c#I;�1I;hDI;uZI;S_I;QI;T�G;aE;p�>;��1;�;���:,d,:���V�k�����W�f֮�����aG�k����ȽFE	��6��l�}����a��Z�Ҿ������      � ��f�����ݕ����q��I���"���������k���ZN�\�#¼N�y��$��Q��q� � �W��:G0;L�&;x8;� B;��F;	�H;�@I;$bI;�RI;M=I;C,I;
I;I;�I;I;kI;OI;�I;OI;lI;I;�I;I;
I;C,I;J=I;�RI;#bI;�@I;�H;��F;� B;x8;K�&;F0;�: �W�r� ��Q���$�N�y�#¼\��ZN�k������������"��I���q�ݕ�����f��      �^Z�c
V��I��6�������ܽ!��ܽ���aG�\��ȼ�)��|�(�`��7G5�@�� �Z:^�::S;2'1;��=;ؠD;Z�G; �H;�XI;J^I;�II;)6I;�&I;�I;�I;�
I;�I;�I;� I;��H;� I;�I;�I;�
I;�I;�I;�&I;(6I;�II;G^I;�XI;�H;W�G;ӠD;��=;2'1;8S;^�:�Z:D��7G5�`��{�(��)���ȼ\��aG�ܽ��!���ܽ������6��I�c
V�      ���IE	��������Wн�A�����h���3����#¼�)��.x/�
�һ\�X�D#����9���:�>;`f);�`9;�&B;�F;�}H;
7I;�aI;�UI;�@I;
/I;.!I;|I;XI;I;�I;� I;��H;0�H;��H;� I;�I;I;YI;|I;.!I;	/I;�@I;�UI;�aI;7I;�}H;ߊF;�&B;�`9;^f);�>;���:��9>#��]�X�
�һ.x/��)��#¼�����3��h��󑽤A���Wн��콼��IE	�      �A��!��f���*��轅�@�d��`=����`��f֮�N�y�{�(�
�һ�]e����� �f9鱩:U�;l1";H�4;�m?;E;��G;��H;�WI;�^I;<KI;�7I;'(I;�I;[I;�
I;UI;QI;��H;	�H;r�H;	�H;��H;PI;WI;�
I;[I;�I;&(I;�7I;;KI;�^I;�WI;��H;��G;E;�m?;H�4;l1";W�;鱩: �f9�����]e�
�һ{�(�N�y�e֮�_�꼚���`=�@�d�齅��*��e��!��      �]��IY��ZN��`=���'�o����䷾������W��$�`��^�X������9���:���:��;̸0;�<;��C;QG;-�H;�?I;_aI;UI;p@I;D/I;�!I;�I;DI;�I;�I;�H;��H;A�H;��H;A�H;��H;�H;�I;�I;DI;�I;�!I;D/I;o@I;UI;^aI;�?I;(�H;QG;��C;�<;̸0;��;���:���:�9����^�X�`���$��W�����䷾����o���'��`=��ZN��IY�      ���k9�^5��>��Vb̼~֮�u��� d�
",�����Q��7G5�D#���f9���:��:4�;��-;��:;LB;iVF;GKH;I;]I;X\I;�HI;:6I;S'I;PI;�I;N
I;uI;0 I;��H;��H;��H;!�H;��H;��H;��H;0 I;vI;N
I;�I;LI;S'I;76I;�HI;V\I;]I;
I;GKH;fVF;LB;��:;��-;2�;��:���: �f9D#��7G5��Q�����
",�� d�u��~֮�Vb̼>��^5��k9�      �d��C��������)���zl�	RH��k"�t.���W��T�k�n� �@����9鱩:���:1�;�-;�9;qaA;�E;V�G;��H;6SI;I`I;PI;�<I;�,I;�I;hI;CI;�I;�I;��H;��H;�H;��H;��H;��H;�H;��H;��H;�I;�I;CI;eI;�I;�,I;�<I;PI;D`I;0SI;��H;T�G;�E;qaA;�9;�-;1�;���:鱩:��9@��p� �T�k��W��v.���k"�RH��zl��)������D���      J",���(�8H�FG��.���jλ$R���^e�F����� �W��Z:���:T�;��;��-;�9;�A;dE;S�G;��H;�GI;+aI;�UI;uBI;�1I; $I;�I;"I;�I;)I;��H;��H;�H;@�H;K�H;�H;K�H;@�H;�H;��H;��H;*I;�I;I;�I;$I;�1I;uBI;�UI;(aI;�GI;��H;T�G;dE;�A;�9;��-;��;U�;���:�Z: �W����E���^e�$R���jλ�.��FG�8H���(�      �5���R��V ��6��<�X�4�$�ۺ�H[�@Q�,d,:
�:b�:�>;n1";ϸ0;��:;qaA;dE;%�G;��H;�=I;``I;�YI;%GI;6I;�'I;#I;�I;2I;�I; I;:�H;W�H;-�H;��H;��H;v�H;��H;��H;,�H;U�H;;�H; I;�I;/I;�I; I;�'I;6I; GI;�YI;b`I;�=I;��H;%�G;dE;paA;��:;Ѹ0;n1";�>;b�:
�:,d,:�Q��H[�ۺ0�$�8�X�6��V ���R��      Z�Ѻ��Ⱥ���`�����&����9l�Z:˰�:���:F0;6S;[f);C�4;	�<;LB;�E;P�G;��H;�:I;�_I;�[I;WJI;99I;�*I;�I;-I;6I;�I;FI; �H;��H;H�H;e�H;0�H;h�H;�H;j�H;0�H;e�H;G�H;��H;!�H;CI;�I;5I;(I;�I;�*I;59I;UJI;�[I;�_I;�:I;��H;R�G;�E;LB;	�<;D�4;[f);6S;G0;���:ɰ�:l�Z:���9&����`��
�����Ⱥ      ���9ĺ:��":@�Q:��:���:�?�:���:�M
;�;L�&;/'1;�`9;�m?;��C;gVF;W�G;��H;�=I;�_I;F\I;�KI;K;I;-I;!I;)I;�I;I;�I;�H;m�H;��H;o�H;��H;��H;�H;��H;�H;��H;��H;m�H;��H;m�H;�H;~I;I;�I;&I;!I;-I;I;I;�KI;C\I;�_I;�=I;��H;V�G;fVF;��C;�m?;�`9;0'1;I�&;�;�M
;���:�?�:���:��:L�Q:ī":��:      ��:���:��:��:��;pN;�L;�, ;�f);��1;x8;��=;�&B;E;RG;EKH;��H;�GI;``I;�[I;�KI;�;I;!.I;g"I;lI;MI;S	I;�I;��H;%�H;�H;��H;��H;T�H;w�H;��H;��H;��H;w�H;T�H;��H;��H;�H;!�H;��H;�I;M	I;LI;nI;b"I; .I;�;I;�KI;�[I;_`I;�GI;��H;DKH;TG;E;�&B;��=;x8;��1;�f);�, ;�L;pN;��;��:��:���:      d�;&�;��;0"; �&;ˆ+;��0;��5;�:;r�>;� B;ؠD;�F;��G;,�H;I;4SI;)aI;�YI;WJI;I;I;$.I;�"I;8I;�I;5
I;eI;��H;��H;��H;��H;��H;2�H;�H;*�H;��H;��H;��H;*�H;�H;0�H;��H;��H;��H;��H;�H;aI;5
I;�I;4I;�"I;$.I;G;I;YJI;�YI;)aI;1SI;
I;,�H;��G;�F;ؠD;� B;p�>;�:;��5;��0;ˆ+;
�&;0";��;�;      zY4;^�4;��5;�7;ݫ9;�<;ן>;�A;L@C;bE;��F;[�G;�}H;��H;�?I;
]I;H`I;�UI;#GI;69I;-I;f"I;5I;[I;�
I;�I;% I; �H;��H; �H;��H;.�H;��H;��H;��H;��H;��H;��H;��H;��H;��H;/�H;��H;�H;��H; �H;" I;�I;�
I;UI;4I;d"I;�,I;69I;#GI;�UI;G`I;
]I;�?I;��H;�}H;[�G;��F;aE;K@C;�A;ן>;�<;�9;�7;��5;O�4;      ~�@;x�@;�`A;�&B;VC;,4D;�ME;�VF;%@G;T�G;	�H;!�H;7I;�WI;`aI;Y\I;$PI;wBI;6I;�*I;	!I;pI;�I;�
I;&I;V I;k�H;�H;[�H;�H;9�H;��H;��H;��H;�H;��H;��H;��H;�H;��H;��H;��H;9�H;�H;X�H;�H;g�H;T I;&I;�
I;�I;oI;!I;�*I;6I;zBI;!PI;V\I;`aI;�WI;7I;!�H;	�H;Q�G;#@G;�VF;�ME;,4D;XC;�&B;�`A;x�@;      �VF;hF;қF;�F;~MG;�G;�#H;ЄH;��H;OI;�@I;�XI;�aI;�^I;UI;�HI;�<I;�1I;�'I;�I;&I;LI;2
I;�I;O I;��H;N�H;��H;&�H;3�H;��H;�H;z�H;��H;?�H;��H;��H;��H;@�H;��H;u�H;��H;��H;2�H;%�H;��H;M�H;}�H;O I;�I;0
I;JI;!I;�I;�'I;�1I;�<I;�HI;UI;�^I;�aI;�XI;�@I;LI;��H;ЄH;�#H;�G;�MG;�F;қF;rhF;      ��H;ŗH;a�H;��H;�H;�I;�%I;AI;tTI;U_I;&bI;M^I;�UI;>KI;r@I;<6I;�,I;$I;%I;.I;�I;S	I;dI;' I;d�H;Q�H;��H;I�H;c�H;��H;c�H;G�H;t�H;��H;s�H;�H;�H;�H;r�H;��H;p�H;F�H;c�H;��H;b�H;J�H;��H;P�H;e�H;# I;aI;Q	I;�I;-I;#I; $I;�,I;96I;r@I;>KI;�UI;M^I;&bI;T_I;vTI;AI;�%I;�I;�H;��H;_�H;ƗH;      �GI;?II;LMI;SI;gYI;�^I;bI;�bI;`I;zZI;�RI;�II;�@I;�7I;E/I;U'I;�I;�I;�I;9I;I;�I;��H;#�H;�H;��H;I�H;?�H;��H;c�H;:�H;C�H;��H;�H;��H;y�H;o�H;y�H;��H;�H;��H;C�H;<�H;`�H;��H;?�H;I�H;��H;�H;#�H;��H;�I;I;8I;�I;�I;�I;U'I;E/I;�7I;�@I;�II;�RI;zZI;`I;�bI;bI;�^I;rYI;SI;LMI;KII;       cI;�bI;bI;�`I;�^I;�[I;9WI;�QI;]KI;nDI;N=I;.6I;
/I;'(I;�!I;PI;jI; I;2I;�I;�I;��H;��H;��H;T�H;'�H;`�H;��H;V�H;:�H;1�H;s�H;��H;d�H;�H;��H;��H;��H;�H;d�H;��H;s�H;/�H;7�H;V�H;��H;b�H;&�H;V�H;��H;��H;��H;�I;�I;3I;"I;iI;OI;�!I;)(I;
/I;,6I;M=I;kDI;]KI;�QI;9WI;�[I;�^I;�`I;!bI;�bI;      HOI;�NI;�MI;�KI;�HI;EI;�@I;"<I;7I;�1I;M,I;�&I;4!I;�I;�I;�I;II;�I;�I;II;�H;"�H;��H;!�H;�H;2�H;��H;a�H;9�H;9�H;b�H;��H;0�H;��H;|�H;\�H;X�H;\�H;|�H;��H;-�H;��H;a�H;6�H;6�H;c�H;��H;/�H;�H; �H;��H;"�H;�H;GI;�I;�I;GI;�I;�I;�I;5!I;�&I;L,I;�1I;7I;&<I;�@I;EI;�HI;�KI;�MI;�NI;      Q:I;�9I;�8I;\7I;!5I;T2I;//I;x+I;�'I;k#I;I;�I;�I;dI;JI;V
I;�I;*I; I;&�H;r�H;�H;��H;��H;6�H;��H;a�H;?�H;/�H;e�H;��H;)�H;��H;J�H;�H;��H;��H;��H;�H;K�H;��H;*�H;��H;d�H;1�H;?�H;`�H;��H;6�H;��H;��H;�H;p�H;&�H; I;*I;�I;U
I;JI;cI;�I;�I;I;k#I;�'I;x+I;//I;T2I; 5I;\7I;�8I;�9I;      *I;�)I;)I;�'I;&I;�#I;t!I;�I;�I;yI;!I;�I;]I;�
I;�I;~I;�I;��H;A�H;��H;��H;��H;��H;3�H;��H;��H;F�H;D�H;r�H;��H;&�H;��H;)�H;��H;��H;��H;q�H;��H;��H;��H;'�H;��H;)�H;��H;u�H;D�H;F�H;�H;��H;2�H;��H;��H;��H;��H;A�H;��H;�I;|I;�I;�
I;_I;�I; I;yI;�I;�I;t!I;�#I;&I;�'I;)I;�)I;      TI;+I;}I;yI;I;qI;nI;FI;�I;.I;�I;�
I;I;^I;�I;5 I;��H;}�H;Z�H;K�H;t�H;��H;2�H;��H;��H;x�H;s�H;��H;��H;3�H;��H;,�H;��H;��H;G�H;?�H;L�H;?�H;G�H;��H;��H;.�H;��H;4�H;��H;��H;q�H;w�H;��H;��H;0�H;��H;s�H;L�H;Z�H;�H;��H;7 I;�I;^I;I;�
I;�I;0I;�I;FI;nI;tI;I;yI;zI;$I;      �I;�I;I;TI;DI;�I;:I;uI;vI;<
I;I;�I;�I;XI;�H; �H;��H;�H;3�H;j�H;��H;U�H;�H;��H;��H;��H;��H;�H;c�H;��H;H�H;��H;��H;X�H;�H;�H;��H;�H;�H;X�H;��H;��H;H�H;��H;e�H;�H;��H;��H;��H;��H;�H;U�H;��H;j�H;2�H;�H;��H; �H;�H;XI;�I;�I;I;:
I;yI;uI;8I;�I;:I;TI;I;�I;      �I;�I;{I;�I;�I;�I;GI;�	I;I;DI;vI;�I;� I;��H;��H;��H;�H;>�H;��H;5�H;��H;z�H;)�H;�H;�H;<�H;n�H;��H;�H;|�H;�H;��H;G�H; �H;	�H;��H;��H;��H;	�H; �H;D�H;��H;�H;�H;
�H;��H;n�H;<�H;�H;��H;)�H;z�H;��H;5�H;��H;A�H;�H;��H;��H;��H;� I;�I;uI;FI;I;�	I;EI;�I;�I;�I;{I;�I;      �I;�I;AI;�I;�
I;�	I;�I;)I;�I;
I;XI;� I;��H;�H;H�H;��H;��H;H�H;��H;o�H;�H;��H;��H;��H;��H;��H;�H;y�H;��H;\�H;��H;��H;?�H;�H;��H;��H;��H;��H;��H;�H;=�H;��H;��H;]�H;��H;y�H;�H;��H;��H;��H;��H;��H;�H;o�H;��H;J�H;��H;��H;H�H;�H;��H;� I;VI;I;�I;(I;�I;�	I;�
I;�I;?I;�I;      �I;�I;HI;�
I;�	I;�I;�I;iI;�I;SI;�I;��H;6�H;|�H;��H;*�H;��H;�H;y�H;#�H;��H;��H;��H;��H;��H;��H; �H;u�H;��H;[�H;��H;x�H;L�H;��H;��H;��H;��H;��H;��H;��H;J�H;z�H;��H;\�H;��H;u�H; �H;��H;��H;��H;��H;��H;��H;#�H;y�H;�H;��H;*�H;��H;|�H;6�H;��H;�I;VI;�I;gI;�I;�I;�	I;�
I;GI;�I;      �I;�I;AI;�I;�
I;�	I;�I;)I;�I;I;XI;� I;��H;�H;H�H;��H;��H;H�H;��H;o�H;�H;��H;��H;��H;��H;��H;�H;y�H;��H;\�H;��H;��H;=�H;�H;��H;��H;��H;��H;��H;�H;=�H;��H;��H;]�H;��H;y�H;�H;��H;��H;��H;��H;��H;�H;o�H;��H;J�H;��H;��H;I�H;�H;��H;� I;XI;
I;�I;(I;�I;�	I;�
I;�I;<I;�I;      �I;�I;yI;�I;�I;�I;EI;�	I;I;DI;uI;�I;� I;��H;��H;��H;�H;@�H;��H;5�H;��H;z�H;)�H; �H;�H;<�H;n�H;��H;	�H;|�H;�H;��H;G�H; �H;	�H;��H;��H;��H;	�H; �H;D�H;��H;�H;~�H;
�H;��H;n�H;<�H;�H;��H;)�H;z�H;��H;5�H;��H;A�H;�H;��H;��H;��H;� I;�I;uI;FI;I;�	I;GI;�I;�I;�I;xI;�I;      �I;�I;I;TI;BI;�I;8I;uI;wI;:
I;I;�I;�I;XI;�H; �H;��H;�H;2�H;j�H;��H;U�H;�H;��H;��H;��H;��H;�H;c�H;��H;H�H;��H;��H;X�H;�H;�H;��H;�H;�H;X�H;��H;��H;H�H;��H;e�H;�H;��H;��H;��H;��H;�H;U�H;��H;j�H;3�H;�H;��H; �H;�H;XI;�I;�I;I;<
I;yI;wI;:I;�I;7I;TI;I;�I;      VI;+I;{I;zI;I;qI;nI;DI;�I;.I;�I;�
I;I;^I;�I;7 I;��H;}�H;Z�H;K�H;t�H;��H;2�H;��H;��H;x�H;t�H;��H;��H;3�H;��H;,�H;��H;��H;G�H;?�H;L�H;?�H;G�H;��H;��H;/�H;��H;4�H;��H;��H;q�H;w�H;��H;��H;0�H;��H;t�H;L�H;Z�H;}�H;��H;5 I;�I;^I;I;�
I;�I;0I;�I;CI;nI;sI;I;zI;xI;(I;      *I;�)I;)I;�'I;&I;�#I;w!I;�I;�I;yI;!I;�I;_I;�
I;�I;}I;�I;��H;A�H;��H;��H;��H;��H;2�H;��H;��H;F�H;D�H;r�H;��H;)�H;��H;(�H;��H;��H;��H;q�H;��H;��H;��H;'�H;��H;&�H;��H;u�H;D�H;F�H;��H;��H;3�H;��H;��H;��H;��H;A�H;��H;�I;~I;�I;�
I;_I;�I;!I;zI;�I;�I;w!I;�#I;&I;�'I;)I;�)I;      Q:I;�9I;�8I;\7I;#5I;T2I;//I;x+I;�'I;j#I;I;�I;�I;dI;JI;V
I;�I;)I; I;&�H;t�H;�H;��H;��H;6�H;��H;`�H;=�H;/�H;e�H;��H;)�H;��H;K�H;�H;��H;��H;��H;�H;J�H;��H;*�H;��H;b�H;1�H;?�H;a�H;��H;6�H;��H;��H;�H;p�H;&�H; I;*I;�I;V
I;JI;dI;�I;�I;I;m#I;�'I;y+I;//I;T2I; 5I;\7I;�8I;�9I;      AOI;�NI;�MI;�KI;�HI;EI;�@I;#<I;7I;�1I;L,I;�&I;6!I;�I;�I;�I;II;�I;�I;JI;�H;"�H;��H; �H;�H;0�H;��H;c�H;7�H;9�H;a�H;��H;/�H;��H;|�H;\�H;X�H;\�H;|�H;��H;/�H;��H;b�H;8�H;9�H;a�H;��H;0�H;�H; �H;��H;"�H;�H;II;�I;�I;GI;�I;�I;�I;5!I;�&I;M,I;�1I;7I;&<I;�@I;EI;�HI;�KI;�MI;�NI;      �bI;�bI;$bI;�`I;�^I;�[I;<WI;�QI;\KI;kDI;N=I;.6I;
/I;'(I;�!I;OI;jI; I;3I;�I;�I;��H;��H;��H;V�H;'�H;`�H;��H;V�H;9�H;/�H;p�H;��H;d�H;�H;��H;��H;��H;�H;d�H;��H;u�H;1�H;9�H;V�H;��H;b�H;&�H;T�H;��H;��H;��H;�I;�I;2I;"I;iI;RI;�!I;'(I;
/I;.6I;N=I;lDI;_KI;�QI;=WI;�[I;�^I;�`I;%bI;�bI;      �GI;AII;LMI;SI;hYI;�^I;bI;�bI;`I;zZI;�RI;�II;�@I;�7I;E/I;U'I;�I;�I;�I;9I; I;�I;��H;#�H;�H;��H;I�H;?�H;��H;d�H;<�H;B�H;��H;�H;��H;y�H;o�H;y�H;��H;�H;��H;D�H;:�H;`�H;��H;?�H;I�H;��H;�H;#�H;�H;�I;I;9I;�I;�I;�I;V'I;E/I;�7I;�@I;�II;�RI;zZI;`I;�bI;bI;�^I;uYI;SI;LMI;KII;      ��H;ƗH;_�H;��H;	�H;�I;�%I;AI;tTI;U_I;&bI;M^I;�UI;>KI;r@I;:6I;�,I;$I;#I;.I;�I;Q	I;bI;& I;e�H;Q�H;��H;J�H;c�H;��H;c�H;F�H;q�H;��H;r�H;�H;�H;�H;s�H;��H;s�H;H�H;c�H;��H;b�H;I�H;��H;Q�H;d�H;% I;bI;S	I;�I;.I;%I; $I;�,I;:6I;r@I;>KI;�UI;M^I;'bI;T_I;tTI;AI;�%I;�I;
�H;��H;[�H;��H;      �VF;xhF;ܛF;�F;~MG;�G;�#H;҄H;��H;NI;�@I;�XI;�aI;�^I;UI;�HI;�<I;�1I;�'I;�I;%I;JI;0
I;�I;O I;~�H;N�H;��H;&�H;3�H;��H;�H;w�H;��H;=�H;��H;��H;��H;@�H;��H;w�H;��H;��H;0�H;%�H;��H;M�H;��H;O I;�I;2
I;LI;"I;�I;�'I;�1I;�<I;�HI;UI;�^I;�aI;�XI;�@I;NI;��H;҄H;�#H;�G;�MG;�F;ڛF;nhF;      ~�@;z�@;�`A;�&B;XC;,4D;�ME;�VF;#@G;S�G;�H;!�H;7I;�WI;`aI;X\I;"PI;wBI;6I;�*I;	!I;oI;�I;�
I;&I;T I;h�H;�H;[�H;�H;9�H;��H;��H;��H;�H;��H;��H;��H;�H;��H;��H;��H;9�H;�H;X�H;�H;h�H;V I;&I;�
I;�I;pI;!I;�*I;6I;zBI;!PI;Y\I;`aI;�WI;7I;!�H;	�H;S�G;#@G;�VF;�ME;,4D;TC;�&B;�`A;x�@;      ~Y4;Y�4;��5;�7;٫9;<;ӟ>;�A;N@C;dE;��F;[�G;�}H;��H;�?I;
]I;H`I;�UI;#GI;69I;-I;d"I;5I;XI;�
I;�I;# I; �H;��H; �H;��H;.�H;��H;��H;��H;��H;��H;��H;��H;��H;��H;/�H;��H;�H;��H; �H;# I;�I;�
I;XI;4I;f"I; -I;69I;#GI;�UI;G`I;
]I;�?I;��H;�}H;[�G;��F;aE;N@C;�A;ӟ>;<;�9;�7;��5;O�4;      a�;4�;��;0"; �&;φ+;��0;��5;�:;r�>;� B;ؠD;��F;��G;,�H;I;3SI;&aI;�YI;WJI;K;I;$.I;�"I;6I;�I;3
I;dI;�H;��H;��H;��H;��H;2�H;�H;*�H;��H;��H;��H;*�H;�H;0�H;��H;��H;��H;��H;��H;bI;6
I;�I;4I;�"I;$.I;E;I;YJI;�YI;+aI;4SI;I;-�H;��G;��F;ؠD;� B;o�>;�:;��5;��0;҆+;�&;0";��;$�;      ��:���:��:��:��;pN;�L;�, ;�f);��1;x8;��=;�&B;E;RG;EKH;��H;�GI;_`I;�[I;�KI;�;I;".I;f"I;nI;JI;Q	I;�I;��H;%�H;�H;��H;��H;T�H;w�H;��H;��H;��H;w�H;T�H;��H;��H;�H;!�H;��H;�I;N	I;MI;lI;d"I; .I;�;I;�KI;�[I;``I;�GI;��H;EKH;TG;E;�&B; �=;x8;��1;�f);�, ;�L;pN;��;��:��:���:      ���9��:Ы":H�Q:��:���:�?�:���:�M
;�;K�&;0'1;�`9;�m?;��C;fVF;W�G;��H;�=I;�_I;E\I;�KI;K;I;-I;!I;(I;�I;I;�I;�H;m�H;��H;o�H;��H;��H;�H;��H;�H;��H;��H;o�H;��H;m�H;�H;I;I;�I;)I;!I;-I;I;I;�KI;C\I;�_I;�=I;��H;V�G;gVF;��C;�m?;�`9;0'1;K�&;�;�M
;���:�?�:���:�:H�Q:Ы":|�:      V�Ѻ��Ⱥ���d�����@&� ��9l�Z:ϰ�:���:G0;6S;[f);D�4;	�<;LB;�E;P�G;��H;�:I;�_I;�[I;WJI;99I;�*I;�I;+I;5I;�I;FI;!�H;��H;H�H;e�H;0�H;k�H;�H;j�H;0�H;e�H;G�H;��H; �H;CI;�I;6I;*I;�I;�*I;59I;UJI;�[I;�_I;�:I;��H;R�G;�E;LB;	�<;C�4;[f);6S;D0;���:˰�:x�Z: ��9 &����d�������Ⱥ      �5���R��V ��6��<�X�4�$�ۺ�H[��Q�,d,:
�:b�:�>;n1";ϸ0;��:;qaA;dE;%�G;��H;�=I;b`I;�YI;%GI;6I;�'I;#I;�I;2I;�I; I;:�H;W�H;,�H;��H;��H;v�H;��H;��H;-�H;U�H;;�H; I;�I;/I;�I; I;�'I;6I; GI;�YI;``I;�=I;��H;%�G;dE;paA;��:;Ѹ0;n1";�>;b�:
�:,d,:�Q��H[�ۺ0�$�5�X�6��V ���R��      J",���(�9H�FG��.���jλ$R���^e�F����� �W��Z:���:T�;��;��-;�9;�A;dE;S�G;��H;�GI;+aI;�UI;uBI;�1I; $I;�I; I;�I;*I;��H;��H;�H;@�H;K�H;�H;K�H;A�H;�H;��H;��H;)I;�I;I;�I;$I;�1I;uBI;�UI;(aI;�GI;��H;T�G;dE;�A;�9;��-;��;T�;���:�Z: �W����E���^e�$R���jλ�.��FG�8H���(�      �d��C��������)���zl�	RH��k"�v.���W��T�k�n� �@����9鱩:���:1�;�-;�9;qaA;�E;V�G;��H;6SI;H`I;PI;�<I;�,I;�I;hI;CI;�I;�I;��H;��H;�H;��H;��H;��H;�H;��H;��H;�I;�I;CI;eI;�I;�,I;�<I;PI;D`I;0SI;��H;T�G;�E;qaA;��9;�-;1�;���:鱩:��9@��n� �U�k��W��t.���k"�RH��zl��)������D���      ���k9�^5��>��Vb̼~֮�u��� d�
",�����Q��7G5�D#���f9���:��:4�;��-;��:;LB;gVF;GKH;I;]I;V\I;�HI;:6I;S'I;PI;�I;N
I;uI;1 I;��H;��H;��H;!�H;��H;��H;��H;. I;uI;N
I;�I;LI;S'I;76I;�HI;X\I;]I;I;GKH;fVF;LB;��:;��-;2�;��:���:�f9D#��6G5��Q�����
",�� d�u��~֮�Vb̼>��^5��k9�      �]��IY��ZN��`=���'�o����䷾������W��$�`��^�X������9���:���:��;̸0;�<;�C;QG;-�H;�?I;^aI;UI;p@I;D/I;�!I;�I;DI;�I;�I;�H;��H;A�H;��H;A�H;��H;�H;�I;�I;DI;�I;�!I;D/I;o@I;UI;_aI;�?I;(�H;QG;�C;�<;̸0;��;���:���:�9����^�X�`���$��W�����䷾����o���'��`=��ZN��IY�      �A��!��f���*��轅�@�d��`=����_��f֮�N�y�{�(�
�һ�]e����� �f9�:U�;l1";G�4;�m?;E;��G;��H;�WI;�^I;<KI;�7I;'(I;�I;[I;�
I;XI;QI;��H;	�H;r�H;	�H;��H;PI;TI;�
I;[I;�I;&(I;�7I;;KI;�^I;�WI;��H;��G;E;�m?;G�4;l1";X�;籩: �f9�����]e�
�һ{�(�N�y�f֮�_�꼚���`=�@�d�轅��*��f��!��      ���IE	��������Wн�A�����h���3����#¼�)��.x/�
�һ]�X�B#����9���:�>;^f);�`9;�&B;�F;�}H;7I;�aI;�UI;�@I;
/I;.!I;|I;XI;I;�I;� I;��H;0�H;��H;� I;�I;I;XI;|I;.!I;/I;�@I;�UI;�aI;
7I;�}H;ފF;�&B;�`9;^f);�>;���:��9D#��\�X�
�һ.x/��)��#¼�����3��h��󑽤A���Wн��콼��IE	�      �^Z�c
V��I��6�������ܽ!��ܽ���aG�\��ȼ�)��|�(�`��7G5�@���Z:^�:8S;/'1;��=;ؠD;Y�G;�H;�XI;J^I;�II;)6I;�&I;�I;�I;�
I;�I;�I;� I;��H;� I;�I;�I;�
I;�I;�I;�&I;(6I;�II;G^I;�XI; �H;W�G;ӠD;��=;2'1;:S;^�:�Z:D��9G5�`��|�(��)���ȼ\��aG�ܽ��!���ܽ������6��I�c
V�      � ��f�����ݕ����q��I���"���������k���ZN�\�#¼O�y��$��Q��q� � �W��:G0;I�&;x8;� B;��F;�H;�@I;$bI;�RI;M=I;C,I;
I;I;�I;I;lI;OI;�I;OI;kI;I;�I;I;
I;C,I;J=I;�RI;#bI;�@I;	�H;��F;� B;x8;K�&;F0;�: �W�r� ��Q���$�O�y�#¼\��ZN�k������������"��I���q�ݕ�����f��      f5�������Z�Ҿ�a��}����l��6�FE	���Ƚk���aG����f֮��W����U�k����,d,:���:�;��1;r�>;dE;T�G;QI;T_I;uZI;kDI;�1I;c#I;uI;*I;7
I;?I;I;SI;I;=I;6
I;)I;uI;d#I;�1I;hDI;uZI;S_I;QI;V�G;bE;p�>;��1;�;���:$d,:���V�k�����W�f֮�����aG�k����ȽFE	��6��l�}����a��Z�Ҿ������      }A��q<�ha/����:�}]׾� ��
w��>�FE	�����ܽ����3�`�꼙���",��W��I���Q�ϰ�:�M
;�f);�:;L@C; @G;��H;rTI;�_I;[KI;7I;'I;�I;�I;pI;I;�I;�I;�I;I;oI;�I;�I;�'I;7I;XKI;�_I;oTI;��H;#@G;I@C;��:;�f);�M
;˰�:�Q�H���W��",�����`�꼜�3�ܽ������FE	�>�
w��� ��}]׾�:���ha/��q<�      x�������c�{�m$_��q<������~��
w���6�����!���h����䷾�� d�v.���^e��H[���Z:���:�, ;��5;�A;�VF;քH;AI;�bI;�QI;<I;q+I;�I;=I;mI;�	I;I;bI;I;�	I;mI;<I;�I;r+I;<I;�QI;�bI;AI;ԄH;WF;�A;��5;�, ;���:x�Z:�H[��^e�x.��� d�䷾�����h�!�������6�
w��~��������q<�m$_�c�{�����      =��������欿�������O��x����� ���l���"��ܽ���`=����v���k"�$R��ۺ���9�?�:|L;��0;П>;�ME;�#H;�%I;bI;6WI;�@I;%/I;q!I;oI;7I;@I;~I;�I;~I;@I;7I;kI;q!I;%/I;�@I;6WI;bI;�%I;�#H;�ME;͟>;��0;|L;�?�:�9ۺ$R���k"�w������`=����ܽ��"��l�� ����뾃x���O�������欿����      �������O��lȿm���������O���}]׾}����I�����A��A�d�o�֮�
RH��jλ;�$�0&����:dN;ʆ+;�<;)4D;�G;�I;�^I;�[I;EI;T2I;�#I;sI;�I;�I;�	I;�I;�	I;�I;�I;pI;�#I;T2I;EI;�[I;�^I;�I;�G;*4D;�<;ʆ+;dN;���:0&�;�$��jλRH�֮�o�A�d��A������I�}���}]׾����O�����m���lȿO�Ῥ��      @�4i�������K�ѿm������q<��:��a����q����Wн齅���'�Wb̼�zl��.��;�X�����:��;�&;ܫ9;RC;MG;�H;hYI;�^I;�HI;5I;&I;I;;I;�I;�
I;�	I;�
I;�I;;I;I;&I;5I;�HI;�^I;hYI;�H;~MG;TC;٫9;
�&;��;�:���;�X��.���zl�Wb̼��'�齅��Wн����q��a���:��q<���m���K�ѿ������4i�      I:�.5�0�'� ������lȿ���m$_���Z�Ҿޕ���6�����*���`=�?�漮)��GG�6��`��X�Q:��:0";�7;�&B;�F;��H;SI;�`I;�KI;O7I;�'I;lI;LI;�I;�I;�
I;�I;�I;LI;kI;�'I;O7I;�KI;�`I;SI;��H;�F;�&B;�7;0";��:\�Q:d��6��GG��)��?���`=��*������6�ޕ��Z�Ҿ��m$_����lȿ���� ��0�'�.5�      ��U�\�O�J-?�0�'���O�ῶ欿c�{�ha/���뾟���I����f���ZN�`5������;H�\ �������":��:��;��5;�`A;��F;a�H;FMI;%bI;�MI;�8I;)I;qI;I;rI;8I;7I;8I;rI;I;pI;)I;�8I;�MI;$bI;FMI;a�H;ޛF;�`A;��5;��;��:��":���\ ��;H�����`5���ZN�f������I�������ha/�c�{��欿O����0�'�J-?�\�O�      ��i���b�\�O�.5�4i�������������q<����f��c
V�IE	�!���IY�k9�D�����(��R����Ⱥ|�:{��:"�;K�4;m�@;ohF;ŗH;@II;�bI;�NI;�9I;�)I;I;�I;�I;�I;�I;�I;�I;�I;I;�)I;�9I;�NI;�bI;@II;×H;ohF;m�@;H�4;(�;{��:|�:��Ⱥ�R����(�E���k9��IY�!��IE	�c
V�f������q<������������4i�.5�\�O���b�      �>���8���*�O������˿p��H�b�E\�7m־^��T�:��J�+��J�B�A��������,/�������>:�t�:Pp ;�J6;EA;�IF;�NH;�H;"I;�I; I;�I;}I;I;� I;��H;9�H;��H;� I;I;|I;�I; I;�I;
"I;�H;�NH;�IF;EA;�J6;Sp ;�t�:�>: ���,/���������A��J�B�+���J�T�:�^��7m־E\�H�b�p���˿����O���*���8�      ��8��4��g&�7��>����<ƿ򲗿�>]�î�S�Ѿ�p���*7����(W��PR?�}�r8�������������G:� �:�!;�6;#lA;�YF;�TH;x�H;("I;�I;�I;�I;VI; I;r I;��H;!�H;��H;s I; I;UI;�I;�I;�I;%"I;x�H;�TH;�YF;#lA;�6;�!;� �:��G:���������r8��}�PR?�(W�����*7��p��S�Ѿî��>]�򲗿�<ƿ>���7���g&��4�      ��*��g&��#�v�X[�rL�������M�t5��>ľ����,��D�쒐��5�6�ݼ���q
��x�|tk���b:Sl�:#;ϗ7;��A;�F;�dH;�I;h"I;I;xI;OI; I;�I;0 I;��H;��H;��H;. I;�I;�I;OI;xI;I;e"I;�I;�dH;�F;��A;˗7;#;Sl�:��b:�tk��x��q
���6�ݼ�5�쒐��DὬ�,����>ľt5���M����rL��X[�v��#��g&�      O�7��v����˿B1��9�y�Ǝ6��z �����5�l�+��ͽ&�����&���˼B�k�#�����X�`� ����:O�;&;�9;��B;�F;�}H;�	I;s"I;=I;�I;�I;�I;XI;��H;5�H;��H;6�H;��H;XI;I;�I;�I;;I;q"I;�	I;�}H;�F;��B;�9;&;O�;���:d� ���X�"���B�k���˼��&�&����ͽ+�5�l������z �Ǝ6�9�y�B1���˿���v�7��      ����>���X[忸˿�T���~�R�î��E۾՗����M���	� �����j��3�d����O�9�׻��/���V��:� 
;*;b;;�jC;�'G;�H; I;"I;I;�I;�
I;�I;�I;V�H;��H;�H;��H;U�H;�I;�I;�
I;�I;�I;"I; I;�H;�'G;�jC;_;;*;� 
;X��:����/�8�׻��O�d���3���j� �����	���M�՗���E۾î�~�R���T���˿X[�>���      �˿�<ƿrL��B1����>]���)�%��	ֳ���{���,�u��*��U`I��J���,���3/��+��� �`/69�4�:�;p.;*.=;naD;��G;p�H;�I;N!I;iI;]I;�	I;�I;� I;��H;$�H;u�H;$�H;��H;� I;�I;�	I;]I;gI;J!I;�I;n�H;��G;laD;%.=;p.;�;�4�:`/69� ��+���3/��,���J��U`I�*��u�齧�,���{�	ֳ�%����)��>]��B1��rL���<ƿ      p��򲗿���9�y�~�R���)�ov��>ľ^���I�Zl����������&�خҼ�}�0B�Ȯ������ �!:	+�:?z;�3;ej?;�\E;��G;��H;zI;�I;�I;�I;�I;�I;, I;��H;s�H;��H;s�H;��H;, I;�I;�I;�I;�I;�I;{I;��H;��G;�\E;`j?;�3;?z;+�:�!:����Ʈ��0B��}�خҼ��&��������[l��I�^���>ľov���)�~�R�9�y����򲗿      H�b��>]���M�Ŏ6�î�%���>ľ$q��|�Z�+�U9ݽ#W����L����$F���G��׻�;��n��Ȋ:�i;#P$;ޘ7;t�A;JF;@CH;��H;� I;yI;�I;(I;=I;�I;)�H;��H;��H;!�H;��H;��H;)�H;�I;>I;(I;�I;vI;� I;��H;>CH;JF;p�A;ݘ7;"P$;�i;�Ȋ:�n��;�	�׻�G�$F�������L�#W��U9ݽ+�|�Z�$q���>ľ%��î�Ŏ6���M��>]�      E\�î�s5��z ��E۾ֳ�^��|�Z�N?#����A����j�(��Hϼ�����ĵ���lۺ :�9�4�:[�;h�,;��;;@�C;�G;[�H;�I;�!I;�I;OI;9I;�I;PI;.�H;�H;��H;3�H;��H;�H;.�H;PI;�I;7I;NI;�I;�!I;�I;Y�H;�G;>�C;��;;g�,;\�;�4�:0:�9�lۺĵ�������Hϼ(����j��A�����N?#�|�Z�^��ֳ��E۾�z �s5�î�      7m־S�Ѿ�>ľ����՗����{��I�+�����V���{�A�/�)���,��@=�B�һZ�@��� ��k:�:b;��3;:j?;t2E;��G;x�H;?I;� I;�I;�I;1	I;I;��H;�H;��H;��H;i�H;��H;��H;�H;��H;I;1	I;�I;�I;� I;?I;x�H;��G;q2E;:j?;��3;b;�:�k:� �\�@�B�һ@=��,��)��A�/��{��V�����+��I���{�՗�������>ľS�Ѿ      ^���p����4�l���M���,�Zl�U9ݽ�A���{��5��J��;���T[�!?�����,P���P�9��:��;/*;*�9;gkB;݇F;�NH;��H;+ I;�I;�I;-I;I;QI;r�H;��H;��H;��H;}�H;��H;��H;��H;q�H;TI;I;-I;�I;�I;) I;��H;�NH;؇F;dkB;*�9;.*;��;��:�P�9.P������!?��T[�;���J���5��{��A��U9ݽZl���,���M�5�l����p��      T�:��*7���,�+���	�u�齅���#W����j�A�/��J���I���k�l�.��W��p ���Ȋ:io�:;er3;*�>;7�D;w�G;Y�H;I;:!I;�I;�I;�
I;	I;r I;��H;��H;��H;��H;u�H;��H;��H;��H;��H;u I;	I;�
I;�I;�I;:!I;I;V�H;r�G;4�D;)�>;er3;;io�:�Ȋ:x ��W��.��l��k��I���J��A�/���j�#W������u�齄�	�+���,��*7�      �J�����D��ͽ ���)�������L�'��)��;���k����hI����/�T/���>:I��:�B;l�,;��:;:�B;�xF;�<H; �H;I;�I;�I;TI;�I;�I;��H;��H;J�H;��H;��H;��H;��H;��H;J�H;��H;��H;�I;�I;RI;�I;�I;I;��H;�<H;�xF;8�B;��:;l�,;�B;O��:��>:L/���/�hI������k�;��(��'����L����)�� ����ͽ�D����      +��'W��뒐�&�����j�T`I���&����Gϼ�,���T[�k�hI��V;�dnk��:,5�:�;&;�6;�!@;B2E;�G;��H;�I;!I;_I;!I;I;JI;� I;��H;�H;��H;u�H;��H;\�H;��H;u�H;��H;�H;��H;� I;LI;I;!I;]I;!I;�I;��H;�G;B2E;�!@;�6;&;�;(5�:�:\nk�T;�hI��k��T[��,��Gϼ�����&�T`I���j�&���뒐�'W��      I�B�PR?��5���&��3��J��׮Ҽ$F����@=�!?�
.����/�pnk����9P׳:��;;!;b3;��=;��C;,�F;#dH;�H;�I;!I;�I;6I;�I;�I;X�H;�H;��H;��H;X�H;��H;P�H;��H;Z�H;��H;��H;�H;X�H;�I;�I;6I;�I;!I;�I;�H;dH;+�F;��C;��=;b3;=!;��;P׳:���9pnk���/�
.��!?�?=���$F��׮Ҽ�J���3���&��5�PR?�      @��}�4�ݼ��˼d���,���}��G����B�һ����U��T/��:Z׳:
�;tb;��0;�<;��B;�IF;{H;8�H;�I;� I;+I;LI;n
I;�I;4 I;C�H;h�H;!�H;<�H;8�H;��H;R�H;��H;8�H;<�H;�H;i�H;C�H;5 I;�I;n
I;II;+I;� I;�I;2�H;{H;�IF;��B;�<;��0;tb;
�;Z׳:�:T/�U������B�һ����G��}��,��d����˼4�ݼ}�      ����p8����@�k���O��3/�.B��׻µ��X�@�,P��p ����>:(5�:��;pb;��/;7;;H�A;��E;οG;�H;�
I;y I;I;I;�I;�I;�I;��H;R�H;��H;��H;�H;,�H;��H;J�H;��H;,�H;�H;��H;��H;R�H;��H;�I;�I;�I;I;I;s I;�
I;�H;ͿG;��E;H�A;9;;��/;pb;��;(5�:��>:p ��.P��X�@�µ���׻.B��3/���O�@�k���q8��      ������q
� ���9�׻ ,��Ʈ���;��lۺ�� ��P�9�Ȋ:I��:�;<!;��0;8;;ʓA;�pE;��G;ގH;��H;�I;KI;kI;7I;�I;�I;�H;Y�H;��H;�H;7�H;�H;�H;z�H;T�H;z�H;�H;�H;5�H;�H;��H;W�H;�H;�I;�I;7I;jI;EI;�I;��H;ێH;��G;�pE;˓A;7;;��0;<!;�;I��:�Ȋ:�P�9�� ��lۺ�;�Ʈ���+��6�׻ ����q
���      &/������x���X���/�� ������n�H:�9�k:��:ko�:�B;&;d3;�<;H�A;�pE;otG;
}H;=�H;;I;�I;XI;I;�
I;I;h I;g�H;;�H;��H;��H;��H;��H;�H;��H;~�H;��H;�H;��H;��H;��H;��H;8�H;b�H;h I;	I;�
I;I;SI;�I;;I;9�H;}H;otG;�pE;G�A;�<;f3;&;�B;ko�:��:�k:P:�9�n������� ���/���X��x����      ����^���ltk�\� ���`/69�!:�Ȋ:�4�:�:��;;k�,;ۡ6;��=;��B;��E;��G;	}H;��H;�I;' I;�I;pI;�I;@I;�I;_�H;�H;V�H;��H;*�H;��H;��H;�H;��H;��H;��H;�H;��H;��H;*�H;��H;R�H;��H;_�H;�I;?I;�I;kI;�I;& I;�I;��H;}H;��G;��E;��B;��=;ݡ6;k�,;;��;�:�4�:�Ȋ:�!:�/69���`� �htk�r���      �>:��G:��b:���:J��:�4�:+�:�i;[�;b;/*;br3;��:;�!@;��C;�IF;пG;ގH;<�H;�I;1 I;XI;PI;�I;*I;uI;7�H;��H;��H;��H;d�H;��H;��H;��H;-�H;��H;��H;��H;-�H;��H;��H;��H;c�H;��H;��H;��H;5�H;uI;*I;�I;OI;WI;- I;�I;=�H;ގH;οG;�IF;��C;�!@;��:;dr3;,*;b;\�;�i;+�:�4�:L��:���:�b:��G:      �t�:� �:ql�:F�;� 
;��;Gz;*P$;l�,;��3;/�9;+�>;:�B;D2E;.�F;{H;�H;��H;;I;) I;WI;�I;PI;�I;I;��H;;�H;g�H;��H;��H;��H;��H;��H;��H;Q�H;�H;��H;�H;Q�H;��H;��H;��H;��H;��H;��H;g�H;9�H;��H;I;�I;MI;�I;TI;) I;;I;��H;�H;yH;/�F;D2E;:�B;+�>;-�9;��3;n�,;)P$;Iz;��;� 
;F�;ul�:� �:      Tp ;�!;#;&;*;p.;�3;ݘ7;��;;<j?;ikB;8�D;�xF;�G;"dH;3�H;�
I;�I;�I;�I;PI;QI;�I;oI;N�H;��H;��H;C�H;�H;/�H;��H;��H;��H;�H;p�H;6�H;!�H;6�H;p�H;�H;��H;��H;��H;+�H;��H;A�H;��H;��H;N�H;mI;�I;QI;KI;�I;�I;�I;�
I;2�H;"dH;�G;�xF;8�D;gkB;:j?;��;;ۘ7;�3;	p.;*;&;#;�!;      �J6;)�6;֗7;�9;e;;'.=;mj?;q�A;C�C;t2E;އF;y�G;�<H;��H;�H;�I;w I;LI;WI;nI;�I;�I;nI;e�H;��H;��H;|�H;I�H;X�H;��H;��H;��H;��H;C�H;��H;��H;e�H;��H;��H;C�H;��H;��H;��H;��H;T�H;H�H;z�H;��H;��H;a�H;mI;�I;�I;mI;VI;LI;v I;�I;�H;��H;�<H;y�G;݇F;r2E;C�C;s�A;lj?;(.=;j;;�9;ח7;�6;      EA;0lA;m�A;��B;�jC;qaD;�\E;JF;�G;��G;�NH;Z�H; �H; I;�I;� I;I;mI;I;�I;-I;I;R�H;��H;�H;��H;Q�H;f�H;��H;��H;��H;��H;��H;|�H;�H;��H;��H;��H;�H;z�H;��H;��H;��H;��H;��H;d�H;M�H;��H;�H;��H;P�H;I;,I;�I;I;pI;I;� I;�I; I;��H;[�H;�NH;��G;�G;JF;�\E;qaD; kC;��B;n�A;0lA;      �IF;�YF;�F;�F;�'G;�G;��G;9CH;X�H;w�H;��H;I;I;!I;!I;+I;I;4I;�
I;?I;tI;��H;��H;��H;��H;|�H;��H;��H;��H;��H;��H;��H;Q�H;��H;n�H;P�H;A�H;P�H;o�H;��H;O�H;��H;��H;��H;��H;��H;~�H;z�H;��H;��H;��H;��H;nI;=I;�
I;6I;
I;(I;!I;!I;I;I;��H;u�H;X�H;9CH;��G;�G;�'G;�F;�F;�YF;      �NH;�TH;�dH;�}H;��H;u�H;��H;��H;�I;BI;, I;@!I;�I;aI;�I;LI;�I;�I;I;�I;9�H;=�H;��H;�H;M�H;��H;��H;��H;��H;��H;��H;�H;��H;&�H;��H;��H;��H;��H;��H;%�H;��H;�H;��H;��H;��H;��H;��H;��H;M�H;|�H;��H;=�H;6�H;�I;I;�I;�I;JI;�I;aI;�I;@!I;, I;?I;�I;��H;��H;q�H;��H;�}H;�dH;�TH;      �H;y�H;�I;�	I; I;�I;~I;� I;�!I;� I;�I;�I;�I;%I;7I;p
I;�I;�I;h I;c�H;��H;h�H;C�H;L�H;b�H;��H;��H;��H;}�H;��H;�H;j�H;�H;��H;k�H;<�H;3�H;:�H;j�H;��H;�H;j�H;�H;��H;{�H;��H;��H;��H;b�H;J�H;A�H;g�H;��H;b�H;g I;�I;�I;n
I;7I;$I;�I;�I;�I;� I;�!I;� I;�I;�I;I;�	I;�I;��H;      "I;+"I;a"I;v"I;"I;J!I;�I;|I;�I;�I;�I;�I;UI;I;�I;�I;�I;�H;g�H;�H;��H;��H; �H;[�H;��H;��H;��H;}�H;��H;�H;`�H;��H;{�H;,�H;��H;��H;��H;��H;��H;+�H;x�H;��H;^�H;�H;��H;}�H;��H;��H;��H;Y�H;��H;��H;��H;�H;e�H;�H;�I;�I;�I;I;TI;�I;�I;�I;�I;zI;�I;J!I;"I;v"I;c"I;""I;      �I;�I;I;>I;I;oI;�I;�I;YI;�I;6I;�
I;�I;TI;�I;: I;��H;V�H;9�H;W�H;��H;��H;+�H;��H;��H;��H;��H;��H;�H;R�H;��H;u�H;��H;��H;��H;}�H;i�H;}�H;��H;��H;��H;w�H;��H;O�H;�H;��H;��H;��H;��H;��H;)�H;��H;��H;W�H;9�H;W�H;��H;8 I;�I;TI;�I;�
I;5I;�I;[I;�I;�I;lI;I;=I;I;�I;      #I;I;�I;�I;�I;]I;�I;1I;BI;8	I;(I;I;�I;� I;_�H;M�H;[�H;��H;��H;�H;j�H;��H;��H;��H;��H;��H;��H;�H;^�H;��H;Y�H;��H;��H;p�H;=�H; �H;�H; �H;=�H;o�H;��H;��H;X�H;��H;^�H;�H;��H;��H;��H;��H;��H;��H;g�H;�H;��H;��H;Y�H;L�H;_�H;� I;�I;I;&I;9	I;BI;1I;�I;^I;�I;�I;�I;I;      �I;�I;WI;�I;�
I;�	I;�I;EI;�I;I;XI;| I;��H;��H;�H;s�H;��H;�H;��H;3�H;��H;��H;��H;��H;��H;��H;�H;m�H;��H;w�H;��H;��H;U�H;.�H;��H;��H;��H;��H;��H;-�H;S�H;��H;��H;x�H;��H;m�H;�H;��H;��H;��H;��H;��H;��H;3�H;��H; �H;��H;s�H;�H;��H;��H;} I;YI;I;�I;DI;�I;�	I;�
I;�I;VI;�I;      �I;jI;
I;�I;�I;�I;�I;�I;XI;��H;x�H;��H;��H; �H;��H;(�H;��H;5�H;��H;��H;��H;��H;��H;��H;��H;P�H;��H;	�H;~�H;�H;��H;W�H;�H;��H;��H;��H;��H;��H;��H;��H;�H;Z�H;��H;�H;�H;	�H;��H;O�H;��H;��H;��H;��H;��H;��H;��H;7�H;��H;(�H;��H;!�H;��H;��H;x�H;��H;XI;�I;�I;�I;�I;�I;
I;dI;      I;I;�I;bI;�I;� I;1 I;3�H;3�H;�H;��H;��H;P�H;��H;��H;G�H;�H;�H;��H;��H;��H;��H;�H;G�H;u�H;��H;#�H;��H;,�H;��H;o�H;.�H;��H;��H;��H;��H;n�H;��H;��H;��H;��H;2�H;o�H;��H;/�H;��H;#�H;��H;v�H;F�H;�H;��H;��H;��H;��H;�H;�H;G�H;��H;��H;P�H;��H;��H;�H;6�H;3�H;1 I;� I;�I;bI;�I;	I;      ~ I;� I;< I;��H;t�H;��H;��H;�H;"�H;��H;��H;��H;��H;�H;_�H;B�H;4�H;�H;�H;�H;4�H;Q�H;m�H;��H;�H;j�H;��H;k�H;��H;��H;=�H;��H;��H;��H;h�H;^�H;`�H;^�H;h�H;��H;��H;��H;=�H;��H;��H;k�H;��H;j�H;�H;��H;m�H;Q�H;2�H;�H;�H;�H;3�H;B�H;_�H;��H;��H;��H;��H;��H;"�H;�H;��H;��H;j�H;��H;< I;� I;      ��H;��H;��H;9�H;��H;�H;}�H;��H;��H;��H;��H;��H;��H;��H;��H;��H;��H;v�H;��H;��H;��H;�H;5�H;��H;��H;K�H;��H;=�H;��H;~�H;!�H;��H;��H;��H;^�H;C�H;C�H;C�H;^�H;��H;��H;��H;!�H;�H;��H;=�H;��H;I�H;��H;��H;5�H;�H;��H;��H;��H;w�H;��H;��H;��H;��H;��H;��H;��H;��H;��H;��H;}�H;#�H;��H;9�H;��H;��H;      9�H;/�H;�H;��H;$�H;r�H;��H;*�H;<�H;l�H;��H;��H;��H;h�H;W�H;Z�H;R�H;N�H;~�H;��H;��H;��H;�H;h�H;��H;;�H;��H;7�H;��H;o�H;�H;��H;��H;s�H;`�H;E�H;A�H;E�H;`�H;s�H;��H;��H;�H;p�H;��H;7�H;��H;=�H;��H;e�H;�H;��H;��H;��H;~�H;P�H;Q�H;Z�H;W�H;i�H;��H;��H;��H;o�H;?�H;)�H;��H;v�H;�H;��H;�H;'�H;      ��H;��H;��H;9�H;��H;�H;}�H;��H;��H;��H;��H;��H;��H;��H;��H;��H;��H;v�H;��H;��H;��H;�H;4�H;��H;��H;K�H;��H;=�H;��H;~�H;!�H;��H;��H;��H;^�H;C�H;C�H;C�H;^�H;��H;��H;��H;!�H;�H;��H;=�H;��H;I�H;��H;��H;5�H;�H;��H;��H;��H;w�H;��H;��H;��H;��H;��H;��H;��H;��H;��H;��H;}�H;#�H;��H;9�H;��H;��H;      } I;� I;; I;��H;r�H;��H;��H;�H;"�H;��H;��H;��H;��H;��H;_�H;B�H;4�H;�H;�H;�H;6�H;Q�H;m�H;��H;�H;j�H;��H;k�H;��H;��H;=�H;��H;��H;��H;h�H;^�H;`�H;^�H;h�H;��H;��H;��H;=�H;��H;��H;k�H;��H;j�H;�H;��H;m�H;Q�H;2�H;�H;�H;�H;3�H;B�H;^�H;�H;��H;��H;��H;��H;"�H;�H;��H;��H;j�H;��H;; I;� I;      !I;I;�I;bI;�I;� I;1 I;3�H;5�H;�H;��H;��H;P�H;��H;��H;G�H;�H;�H;��H;��H;��H;��H;�H;G�H;v�H;��H;#�H;��H;+�H;��H;o�H;/�H;��H;��H;��H;��H;n�H;��H;��H;��H;��H;2�H;o�H;��H;/�H;��H;#�H;��H;u�H;F�H;�H;��H;��H;��H;��H;�H;�H;G�H;��H;��H;P�H;��H;��H;�H;6�H;4�H;1 I;� I;�I;bI;�I;	I;      �I;jI;I;�I;�I;�I;�I;�I;XI;��H;x�H;��H;��H; �H;��H;(�H;��H;5�H;��H;��H;��H;��H;��H;��H;��H;P�H;��H;	�H;~�H;�H;��H;X�H;�H;��H;��H;��H;��H;��H;��H;��H;�H;[�H;��H;�H;�H;	�H;��H;P�H;��H;��H;��H;��H;��H;��H;��H;5�H;��H;(�H;��H; �H;��H;��H;x�H;��H;ZI;�I;�I;�I;�I;�I;I;gI;      �I;�I;WI;�I;�
I;�	I;�I;GI;�I;I;YI;} I;��H;��H;�H;s�H;��H;�H;��H;4�H;��H;��H;��H;��H;��H;��H;�H;m�H;��H;w�H;��H;��H;T�H;-�H;��H;��H;��H;��H;��H;.�H;S�H;��H;��H;x�H;��H;m�H;�H;��H;��H;��H;��H;��H;��H;3�H;��H; �H;��H;s�H;�H;��H;��H;| I;XI;I;�I;EI;�I;�	I;�
I;�I;WI;�I;      #I;I;�I;�I;�I;]I;�I;1I;BI;8	I;(I;I;�I;� I;_�H;M�H;Y�H;��H;��H;�H;j�H;��H;��H;��H;��H;��H;��H;�H;\�H;��H;X�H;��H;��H;o�H;=�H; �H;�H; �H;=�H;p�H;��H;��H;Y�H;��H;`�H;�H;��H;��H;��H;��H;��H;��H;g�H;�H;��H;��H;Y�H;M�H;_�H;� I;�I;I;&I;9	I;BI;2I;�I;^I;�I;�I;�I;I;      �I;�I;I;;I;I;hI;�I;�I;[I;�I;5I;�
I;�I;UI;�I;8 I;��H;V�H;9�H;Y�H;��H;��H;+�H;��H;��H;��H;��H;��H;�H;P�H;��H;t�H;��H;��H;��H;}�H;i�H;}�H;��H;��H;��H;w�H;��H;P�H;�H;��H;��H;��H;��H;��H;)�H;��H;��H;W�H;9�H;W�H;��H;; I;�I;SI;�I;�
I;6I;�I;\I;�I;�I;nI;I;=I;I;�I;      "I;("I;f"I;u"I;"I;G!I;�I;zI;�I;�I;�I;�I;UI;I;�I;�I;�I;�H;e�H;�H;��H;��H;��H;Y�H;��H;��H;��H;}�H;��H;�H;^�H;��H;z�H;+�H;��H;��H;��H;��H;��H;,�H;z�H;��H;`�H;�H;��H;}�H;��H;��H;��H;[�H;��H;��H;��H;�H;g�H;�H;�I;�I;�I;I;TI;�I;�I;�I;�I;}I;�I;H!I;"I;q"I;i"I;'"I;      �H;|�H;�I;�	I;I;�I;�I;� I;�!I;� I;�I;�I;�I;%I;6I;n
I;�I;�I;g I;b�H;��H;g�H;A�H;J�H;b�H;��H;��H;��H;}�H;��H;�H;j�H;�H;��H;i�H;<�H;3�H;<�H;k�H;��H;�H;k�H;�H;��H;{�H;��H;��H;��H;b�H;L�H;A�H;h�H;��H;c�H;h I;�I;�I;q
I;7I;$I;�I;�I;�I;� I;�!I;� I;~I;�I;I;�	I;�I;��H;      �NH;�TH;�dH;�}H;��H;p�H;��H;��H;�I;@I;, I;@!I;�I;aI;�I;LI;�I;�I;I;�I;:�H;=�H;��H;~�H;M�H;��H;��H;��H;��H;��H;��H;�H;��H;%�H;��H;��H;��H;��H;��H;%�H;��H;�H;��H;��H;��H;��H;��H;��H;M�H;~�H;��H;=�H;7�H;�I;I;�I;�I;JI;�I;aI;�I;@!I;- I;@I;�I;��H;��H;p�H;��H;�}H;�dH;�TH;      �IF;�YF;�F;�F;�'G;�G;��G;;CH;V�H;w�H;��H;I;I;!I;I;*I;I;4I;�
I;=I;rI;��H;��H;��H;��H;y�H;��H;��H;��H;��H;��H;��H;P�H;��H;m�H;P�H;A�H;P�H;o�H;��H;O�H;��H;��H;��H;��H;��H;��H;|�H;��H;��H;��H;��H;pI;?I;�
I;6I;
I;+I;!I;!I;I;I;��H;u�H;X�H;:CH;��G;�G;�'G;�F;�F;�YF;      EA;0lA;n�A;��B; kC;qaD;�\E;JF;�G;��G;�NH;[�H;��H; I;�I;� I;I;mI;I;�I;-I;I;R�H;��H;�H;��H;P�H;d�H;��H;��H;��H;��H;��H;z�H;�H;��H;��H;��H;�H;z�H;��H;��H;��H;��H;��H;f�H;P�H;��H;�H;��H;P�H;I;,I;�I;I;pI;I;� I;�I;�I; �H;[�H;�NH;��G;�G;JF;�\E;qaD;�jC;��B;n�A;.lA;      �J6;%�6;ݗ7;�9;_;;+.=;gj?;s�A;D�C;u2E;އF;y�G;�<H;��H;�H;�I;w I;II;VI;mI;�I;�I;nI;d�H;��H;��H;{�H;H�H;V�H;��H;��H;��H;��H;B�H;��H;��H;e�H;��H;��H;C�H;��H;��H;��H;��H;U�H;I�H;{�H;��H;��H;d�H;mI;�I;�I;nI;WI;NI;w I;�I;�H;��H;�<H;y�G;݇F;r2E;F�C;v�A;gj?;,.=;p;;�9;��7;�6;      Rp ;�!;#;&;*;p.;�3;ݘ7;��;;<j?;gkB;8�D;�xF;�G;"dH;3�H;�
I;�I;�I;�I;OI;QI;�I;oI;N�H;��H;��H;A�H; �H;/�H;��H;��H;��H;�H;p�H;6�H;!�H;6�H;p�H;�H;��H;��H;��H;,�H; �H;C�H;��H;��H;N�H;mI;�I;QI;LI;�I;�I;�I;�
I;3�H;#dH;�G;�xF;8�D;ikB;9j?;��;;ޘ7;�3;p.;*;&;#;�!;      �t�:� �:ol�:F�;� 
;��;Iz;)P$;l�,;��3;/�9;+�>;:�B;D2E;.�F;zH;�H;��H;;I;' I;WI;�I;PI;�I;I;��H;=�H;g�H;��H;��H;��H;��H;��H;��H;O�H;�H;��H;�H;Q�H;��H;��H;��H;��H;��H;��H;g�H;9�H;��H;I;�I;MI;�I;VI;* I;;I;��H;�H;{H;/�F;D2E;:�B;-�>;-�9;��3;n�,;*P$;Gz;��;� 
;F�;ql�:� �:      ��>:��G:�b:���:J��:�4�:+�:�i;[�;b;.*;dr3;��:;�!@;��C;�IF;пG;܎H;=�H;�I;. I;WI;PI;�I;*I;tI;7�H;��H;��H;��H;c�H;��H;��H;��H;-�H;��H;��H;��H;-�H;��H;��H;��H;d�H;��H;��H;��H;6�H;uI;*I;�I;OI;XI;. I;�I;<�H;ߎH;οG;�IF;��C;�!@;��:;br3;.*;b;\�;�i;+�:�4�:V��:���:�b:��G:      ����^���\tk�d� ����0/69�!:�Ȋ:�4�:�:��;;k�,;ݡ6;��=;��B;��E;��G;}H;��H;�I;& I;�I;pI;�I;?I;�I;_�H;�H;U�H;��H;)�H;��H;��H;�H;��H;��H;��H;�H;��H;��H;,�H;��H;S�H;��H;_�H;�I;?I;�I;kI;�I;' I;�I;��H;	}H;��G;��E;��B;��=;ۡ6;k�,;;��;�:�4�:�Ȋ:�!:�/69���`� �`tk�x���      &/������x���X���/�� ������n�H:�9�k:��:ko�:�B;&;d3;�<;H�A;�pE;otG;
}H;<�H;;I;�I;WI;I;�
I;I;h I;e�H;;�H;��H;��H;��H;��H;�H;��H;~�H;��H;�H;��H;��H;��H;��H;8�H;b�H;h I;	I;�
I;I;TI;�I;;I;9�H;}H;otG;�pE;G�A;�<;f3;&;�B;ko�:��:�k:P:�9�n������� ���/���X��x����      ������q
� ���9�׻,��Ʈ���;��lۺ�� ��P�9�Ȋ:I��:�;<!;��0;7;;ʓA;�pE;��G;ގH;��H;�I;II;jI;6I;�I;�I;�H;Y�H;��H;�H;7�H;�H;�H;z�H;T�H;z�H;�H;�H;5�H;�H;��H;W�H;�H;�I;�I;7I;kI;GI;�I;��H;ێH;��G;�pE;˓A;7;;��0;=!;�;I��:�Ȋ:�P�9�� ��lۺ�;�Ʈ���+��6�׻ ����q
���      ����p8����@�k���O��3/�-B��׻µ��X�@�,P��p ����>:(5�:��;pb;��/;7;;H�A;��E;οG;�H;�
I;w I;I;I;�I;�I;�I;��H;R�H;��H;��H;�H;,�H;��H;J�H;��H;,�H;�H;��H;��H;R�H;��H;�I;�I;�I;I;I;s I;�
I;�H;ͿG;��E;H�A;9;;��/;pb;��;(5�:��>:p ��,P��Z�@�µ���׻.B��3/���O�@�k���q8��      @��}�4�ݼ��˼d���,���}��G����A�һ����U��T/��:Z׳:
�;tb;��0;�<;��B;�IF;{H;6�H;�I;� I;*I;LI;n
I;�I;4 I;C�H;h�H;!�H;<�H;8�H;��H;R�H;��H;8�H;<�H;�H;i�H;C�H;5 I;�I;n
I;II;-I;� I;�I;2�H;{H;�IF;��B;�<;��0;tb;
�;Z׳:�:T/�U������B�һ����G��}��,��d����˼4�ݼ}�      I�B�PR?��5���&��3��J��׮Ҽ$F����?=�"?�
.����/�pnk����9P׳:��;;!;b3;��=;��C;+�F;#dH;�H;�I;I;�I;6I;�I;�I;X�H;�H;��H;��H;Z�H;��H;P�H;��H;X�H;��H;��H;�H;X�H;�I;�I;6I;�I;"I;�I;�H;dH;,�F;��C;��=;b3;=!;��;P׳:���9pnk���/�
.��!?�@=���$F��׮Ҽ�J���3���&��5�PR?�      +��'W��뒐�&�����j�T`I���&����Gϼ�,���T[�k�hI��V;�\nk��:,5�:�;&;ߡ6;�!@;B2E;�G;��H;�I;!I;_I;!I;I;JI;� I;��H;�H;��H;u�H;��H;\�H;��H;u�H;��H;�H;��H;� I;LI;I;!I;]I;!I;�I;��H;�G;B2E;�!@;ߡ6;&;�;(5�:�:dnk�V;�hI��k��T[��,��Gϼ�����&�T`I���j�&���뒐�'W��      �J�����D��ͽ ���)�������L�'��(��;���k����hI����/�T/���>:K��:�B;l�,;��:;8�B;�xF;�<H;��H;I;�I;�I;TI;�I;�I;��H;��H;J�H;��H;��H;��H;��H;��H;J�H;��H;��H;�I;�I;QI;�I;�I;I; �H;�<H;�xF;:�B;��:;l�,;�B;O��:��>:T/���/�hI������k�;��(��'����L����)�� ����ͽ�D����      T�:��*7���,�+���	�u�齅���#W����j�A�/��J���I���k�l�.��W��p ���Ȋ:io�:;br3;)�>;7�D;u�G;V�H;I;<!I;�I;�I;�
I;	I;r I;��H;��H;��H;��H;u�H;��H;��H;��H;��H;r I;	I;�
I;�I;�I;9!I;I;Y�H;t�G;4�D;*�>;er3;;io�:�Ȋ:x ��X��.��l��k��I���J��A�/���j�#W������u�齄�	�+���,��*7�      ^���p����4�l���M���,�Zl�U9ݽ�A���{��5��J��;���T[�!?�����,P���P�9��:��;+*;*�9;gkB;݇F;�NH;��H;, I;�I;�I;-I;I;QI;r�H;��H;��H;��H;}�H;��H;��H;��H;q�H;RI;I;-I;�I;�I;) I;��H;�NH;؇F;dkB;*�9;,*;��;��:�P�9.P������!?��T[�;���J���5��{��A��U9ݽZl���,���M�4�l����p��      7m־S�Ѿ�>ľ����՗����{��I�+�����V���{�A�/�)���,��@=�B�һZ�@��� ��k:�:b;��3;<j?;t2E;��G;x�H;@I;� I;�I;�I;1	I;I;��H;�H;��H;��H;i�H;��H;��H;�H;��H;I;1	I;�I;�I;� I;=I;x�H;��G;r2E;9j?;��3;b;�:�k:� �\�@�C�һ?=��,��)��A�/��{��V�����+��I���{�՗�������>ľS�Ѿ      E\�î�s5��z ��E۾	ֳ�^��|�Z�N?#����A����j�(��Hϼ�����µ���lۺ0:�9�4�:Y�;g�,;��;;@�C;�G;Y�H;�I;�!I;�I;NI;7I;�I;QI;.�H;�H;��H;3�H;��H;�H;.�H;NI;�I;9I;NI;�I;�!I;�I;Y�H;�G;>�C;��;;h�,;\�;�4�: :�9�lۺĵ�������Hϼ(����j��A�����N?#�|�Z�^��ֳ��E۾�z �s5�î�      H�b��>]���M�Ŏ6�î�%���>ľ$q��|�Z�+�U9ݽ#W����L����$F���G��׻�;��n��Ȋ:�i;"P$;ޘ7;s�A;JF;>CH;��H;� I;yI;�I;(I;=I;�I;*�H;��H;��H;!�H;��H;��H;*�H;�I;=I;(I;�I;vI;� I;��H;=CH;JF;p�A;ݘ7;#P$;�i;�Ȋ:�n��;�	�׻�G�$F�������L�#W��U9ݽ+�|�Z�$q���>ľ%��î�Ŏ6���M��>]�      p��򲗿���9�y�~�R���)�ov��>ľ^���I�[l����������&�خҼ�}�0B�Ǯ�������!:	+�:?z;�3;ej?;�\E;��G;��H;{I;�I;�I;�I;�I;�I;- I;��H;s�H;��H;s�H;��H;, I;�I;�I;�I;�I;�I;zI;��H;��G;�\E;bj?;�3;?z;+�:�!:����Ʈ��0B��}�خҼ��&��������Zl��I�^���>ľov���)�~�R�9�y����򲗿      �˿�<ƿrL��B1����>]���)�%��	ֳ���{���,�u��*��U`I��J���,���3/��+��� �`/69�4�:�;p.;*.=;laD;��G;p�H;�I;M!I;iI;]I;�	I;�I;� I;��H;$�H;u�H;&�H;��H;� I;�I;�	I;]I;gI;J!I;�I;n�H;��G;naD;%.=;p.;�;�4�:P/69� ��+���3/��,���J��U`I�*��u�齧�,���{�	ֳ�%����)��>]��B1��rL���<ƿ      ����>���X[忸˿�T���~�R�î��E۾՗����M���	� �����j��3�d����O�9�׻��/���R��:� 
;*;b;;�jC;�'G;�H; I;"I;I;�I;�
I;�I;�I;V�H;��H;�H;��H;U�H;�I;�I;�
I;�I;�I;"I; I;�H;�'G;�jC;_;;*;� 
;X��:����/�8�׻��O�d���3���j� �����	���M�՗���E۾î�~�R���T���˿X[�>���      O�7��v����˿B1��9�y�Ǝ6��z �����5�l�+��ͽ&�����&���˼B�k�#�����X�`� ����:O�;&;�9;��B;�F;�}H;�	I;s"I;>I;�I;�I;�I;XI;��H;6�H;��H;5�H;��H;XI;I;�I;�I;;I;q"I;�	I;�}H;�F;��B;�9;&;O�;���:d� ���X�"���B�k���˼��&�&����ͽ+�5�l������z �Ǝ6�9�y�B1���˿���v�7��      ��*��g&��#�v�X[�rL�������M�t5��>ľ����,��D�쒐��5�6�ݼ���q
��x��tk���b:Sl�:#;ϗ7;��A;�F;�dH;�I;h"I;I;xI;OI; I;�I;0 I;��H;��H;��H;0 I;�I;�I;OI;xI;I;e"I;�I;�dH;�F;��A;˗7;#;Sl�:��b:�tk��x��q
���6�ݼ�5�쒐��DὬ�,����>ľt5���M����rL��X[�v��#��g&�      ��8��4��g&�7��>����<ƿ򲗿�>]�î�S�Ѿ�p���*7����(W��PR?�}�r8�������������G:� �:�!;�6;#lA;�YF;�TH;x�H;("I;�I;�I;�I;VI; I;r I;��H;!�H;��H;s I; I;UI;�I;�I;�I;%"I;x�H;�TH;�YF;#lA;�6;�!;� �:��G:���������r8��}�PR?�(W�����*7��p��S�Ѿî��>]�򲗿�<ƿ>���7���g&��4�      ��!$������꿱�ſ�ޞ�(3s��2�@����� j���}Hͽȸ����'�G<ͼt�n�k���<Q^�d-.�h��:|W;�S%;do8;��A;cDF;�H;��H;��H;��H;S�H;J�H;R�H;��H;��H;��H;8�H;��H;��H;��H;P�H;K�H;S�H;��H;��H;��H;�H;aDF;��A;co8;�S%;|W;l��:l-.�<Q^�j���u�n�G<ͼ��'�ȸ��}Hͽ�� j���@����2�(3s��ޞ���ſ������!$�      !$�������忊�����"cm�X�-�����Sh��Zde�$-�۪ɽ�v��+�$���ɼ|mj�>���X�����ņ:wx;D�%;1�8;pB;qRF;H;4�H;[�H;�H;v�H;N�H;D�H;��H;��H;��H;3�H;��H;��H;��H;B�H;O�H;v�H;�H;X�H;4�H;H;pRF;pB;/�8;I�%;wx;�ņ:���X�=���}mj���ɼ+�$��v��۪ɽ$-�Zde�Sh������X�-�"cm��������忞����      ��������� �ԿNw�����=�\�"����n��]0X�����;����w����������]�&���F�����ɒ:��;;�';��9;"pB;�zF;�!H;��H;>�H;#�H;��H;T�H;I�H;��H;��H;��H;�H;��H;��H;��H;H�H;T�H;��H; �H;;�H;��H;�!H;�zF;"pB;��9;=�';��;�ɒ:����F�$�黯�]����������w��;�����]0X�n�����"�=�\����Nw�� �Կ��𿞏�      ����� �Կp���ޞ�bF�j�C�/E�%�;�I���D���!"��k�c���֯���J��ѻɢ)��}K�$��:�
;�M*;u�:;�C;�F;�8H;\�H;��H;{�H;��H;M�H;I�H;��H;��H;��H;
�H;��H;��H;��H;H�H;M�H;��H;z�H;��H;\�H;�8H;�F;�C;r�:;�M*;�
;&��:�}K�ɢ)��ѻ��J��֯��k�c�!"�����D��I��%�;/E�j�C�bF��ޞ�p�� �Կ��      ��ſ���Nw���ޞ�����A�W�7�%�����jɰ��|x�i{+�ֱ� ���J��  �Ѷ��\�1�+���+�p"
9��:��;�-;��<;��C;�G;�TH;T�H;�H;��H;��H;c�H;A�H;��H;��H;��H;��H;��H;��H;��H;@�H;d�H;��H;��H;�H;T�H;�TH;�G;��C;��<;�-;��; �:p"
9+�*���\�1�Ѷ���  ��J� ��ֱ�i{+��|x�jɰ�����7�%�A�W������ޞ�Nw�����      �ޞ�������bF�A�W�Y�-����BKɾ�G����O����ƽɸ��҄-���ۼㄼ64�ǐ��ζ��]:��:�;��1;�c>;q�D;�\G;HsH;��H;q�H;j�H;.�H;��H;7�H;{�H;��H;��H;��H;��H;��H;{�H;7�H;��H;.�H;g�H;m�H;��H;GsH;�\G;q�D;�c>;��1;�;��:�]:�ζ�ǐ�64�ㄼ��ۼ҄-�ɸ��ƽ�����O��G��BKɾ���Y�-�A�W�bF�������      (3s�"cm�=�\�j�C�7�%�����TҾm�� j��C(����aP����[�������Y�:��bX�8�<���k:M��: � ;�5;HR@;huE;
�G;8�H;N�H;��H;	�H;Q�H;{�H;3�H;r�H;��H;g�H;��H;g�H;��H;r�H;3�H;|�H;Q�H;	�H;��H;N�H;7�H;
�G;fuE;ER@;�5; � ;Q��:��k:8�<�_X�:����Y�������[�aP����콭C(� j�m���TҾ���7�%�j�C�=�\�"cm�      �2�X�-�"�/E�����BKɾm����s�;�5���z㻽�v��z0��;��+���*����+6��=S��M�:]�	;��(;�9;�/B;zDF;XH;׫H;��H;��H;��H;�H;��H;�H;A�H;O�H;K�H;j�H;K�H;O�H;A�H;�H;��H;�H;��H;��H;��H;ԫH;WH;vDF;�/B;�9;��(;_�	;�M�:�=S�(6�����*��+���;�z0��v��z㻽��;�5���s�m��BKɾ����/E�"�X�-�      @����������$�;jɰ��G�� j�;�5��	�Ҫɽ\����J�v���沼��]�����	x�@	��dn:Ϥ�:�v;��/;�-=;��C;J�F;&IH;��H;,�H;��H;*�H;��H;��H;��H;�H;�H;%�H;4�H;%�H;�H;�H;��H;��H;��H;)�H;��H;,�H;��H;&IH;G�F;��C;�-=;��/;�v;ͤ�:hn:<	���	x������]��沼v���J�\���Ҫɽ�	�;�5� j��G��jɰ�$�;��徺���      ��Sh��m���I���|x���O��C(���Ҫɽ����WDX�K��+<ͼㄼ�X!��s���W��tK�F��:�y;�#;
I6;9R@;�PE;��G;��H;��H;7�H;��H;��H;��H;��H;��H;��H;��H;��H;��H;��H;��H;��H;��H;��H;��H;��H;��H;7�H;��H;��H;��G;�PE;7R@;
I6;�#;�y;F��:�tK��W��s���X!�ㄼ+<ͼK��WDX�����Ҫɽ���C(���O��|x��I��m��Sh��       j�Zde�]0X��D�i{+�������y㻽\���WDX������ۼξ����;�G>ۻX��y� ?":��:��;ܷ-;��;;��B;�zF;�H;��H;��H;,�H;��H;��H;��H;~�H;��H;��H;��H;��H;��H;��H;��H;��H;��H;��H;��H;��H;��H;,�H;�H;��H;�H;�zF;��B;��;;ڷ-;��;��:,?":$�y�X�G>ۻ��;�ξ����ۼ���WDX�\���z㻽��콅��j{+��D�]0X�Zde�      ��$-������ֱ�ƽaP���v���J�K����ۼ��f�J������+��rrѺp)
9�M�:��;� $;�5;��?;��D;g\G;fH;��H;��H;��H;��H;*�H;�H;d�H;��H;n�H;g�H;t�H;M�H;t�H;i�H;n�H;��H;g�H;��H;+�H;��H;��H;��H;��H;fH;d\G;��D;��?;�5;� $;��;�M�:`)
9vrѺ�+������f�J�����ۼK���J��v��aP��ƽֱ轆����$-�      }Hͽڪɽ�;��!"�� ��ɸ����[�z0�u��+<ͼξ��f�J�����j��q*�����:Zb�:V�;��/;�L<;C;4mF;��G;�H;�H;�H;�H;P�H;b�H;��H;7�H;D�H;0�H;+�H;�H;�H;�H;+�H;/�H;C�H;9�H;��H;b�H;P�H;�H;�H;�H;�H;��G;/mF;C;�L<;��/;V�;`b�:��:��q*��j�����f�J�ξ��+<ͼu��z0���[�ɸ�� ��!"���;��ڪɽ      Ǹ���v����w�j�c��J�҄-�~��;缉沼ㄼ��;������j���5� ��<?Q:m��:fi;�M*;��8;��@;�PE;�uG;EiH;��H;��H;�H;2�H;��H;��H;��H;	�H;��H;��H;��H;��H;��H;��H;��H;��H;��H;�H;��H;��H;��H;2�H;�H;��H;��H;BiH;�uG;�PE;��@;��8;�M*;hi;k��:<?Q:��깛5��j��������;�ㄼ�沼�;�~�ф-��J�j�c���w��v��      ��'�+�$������  ���ۼ����+����]��X!�G>ۻ�+��r*����>:���:�;:�%;�5;��>;�(D;�F;�!H;?�H;`�H; �H;��H;��H;��H;�H;��H;��H;��H;��H;~�H;c�H;��H;c�H;�H;��H;��H;��H;��H;~�H;��H;��H;��H; �H;_�H;9�H;�!H;�F;�(D;��>;�5;<�%;�;���:�>:��r*��+��H>ۻ�X!���]��+�������ۼ�  �����+�$�      F<ͼ��ɼ�����֯�ж��ㄼ��Y��*�����s��X�rrѺ��8?Q:���:��
;T�#;i�3;�c=;$C;0DF;�G;�H;��H; �H;I�H;	�H;i�H;8�H;z�H;��H;v�H;M�H;h�H;!�H; �H; �H;�H;!�H;h�H;L�H;w�H;��H;z�H;4�H;i�H;�H;I�H;�H;��H;�H;�G;,DF;$C;�c=;j�3;Q�#;��
;���:@?Q:��rrѺX��s������*���Y�ㄼж���֯�������ɼ      t�n�ymj���]���J�\�1�64�6������	x��W��y�`)
9��:k��:�;P�#;\�2;�<;upB;3�E;��G;�eH;�H;F�H;��H;�H;��H;��H;Q�H;_�H;N�H;&�H;�H;��H;��H;��H;��H;��H;��H;��H;�H;'�H;N�H;^�H;N�H;��H;��H;	�H;��H;B�H;��H;�eH;��G;4�E;upB;�<;^�2;O�#;�;k��:��:p)
9$�y��W��	x����5��54�\�1���J���]�|mj�      l���=���"���ѻ,���ǐ�aX�,6�<	�� uK�,?":�M�:Zb�:di;;�%;g�3;�<;M0B;��E;�\G;�HH;U�H;��H;p�H;�H;K�H;S�H;��H;.�H;1�H;��H;��H;��H;z�H;l�H;k�H;H�H;k�H;l�H;y�H;��H;��H;��H;/�H;+�H;��H;O�H;L�H;�H;l�H;��H;U�H;�HH;�\G;��E;N0B;�<;f�3;;�%;fi;Zb�:�M�:0?":�tK�:	��-6�aX�ǐ�(����ѻ!��B���      1Q^�X��F�Ƣ)�+��ζ� �<��>S�pn:B��:��:��;V�;�M*;�5;�c=;tpB;��E;�JG;b8H;|�H;��H;%�H;A�H;��H;��H;��H;��H;�H;��H;��H;��H;p�H;�H;�H;�H;��H;�H;�H;�H;n�H;��H;��H;��H; �H;��H;��H;��H;��H;:�H; �H;��H;z�H;c8H;�JG;��E;tpB;�c=;��5;�M*;T�;��;��:B��:pn:�>S� �<��ζ�+�Ƣ)��F�X�      T-.�L����깐}K�P"
9�]:��k:�M�:ˤ�:�y;��;� $;��/;��8;��>;$C;2�E;�\G;_8H;֥H;�H;4�H;��H;K�H;��H;k�H;��H;��H;��H;��H;T�H;-�H;��H;��H;��H;��H;��H;��H;��H;��H;��H;-�H;T�H;��H;��H;��H;��H;i�H;��H;D�H;��H;4�H;�H;֥H;_8H;�\G;2�E;$C;��>;��8;��/;� $;��;�y;ˤ�:�M�:��k:�]:�"
9�}K����p��      |��:Ɔ:�ɒ:��:��:��:Q��:]�	;�v;�#;ܷ-;�5;�L<;��@;�(D;-DF;��G;�HH;|�H;�H;��H;a�H;��H;v�H;8�H;��H;��H;��H;z�H;<�H; �H;��H;��H;}�H;N�H;@�H;@�H;@�H;N�H;|�H;��H;��H;�H;:�H;w�H;��H;��H;��H;7�H;q�H;��H;`�H;��H;�H;{�H;�HH;��G;,DF;�(D;��@;�L<;�5;ٷ-;�#;�v;\�	;Q��:��:��:��:�ɒ:�ņ:      �W;�x;�;�
;��;�;� ;��(;��/;
I6;��;;�?;C;�PE;�F;�G;�eH;U�H;��H;6�H;a�H;��H;H�H;�H;}�H;��H;��H;��H;�H;��H;��H;d�H;;�H;)�H;��H;��H;��H;��H;��H;)�H;9�H;c�H;��H;��H;�H;��H;��H;��H;}�H;�H;E�H;��H;^�H;7�H;��H;U�H;�eH;�G;�F;�PE;C;�?;��;;I6;��/;��(;� ;�;ƅ;�
;�;�x;      �S%;G�%;;�';�M*;�-;��1;�5;�9;�-=;7R@;��B;��D;2mF;�uG;�!H;�H;�H;��H;%�H;��H;��H;I�H;�H;~�H;��H;��H;V�H;�H;��H;��H;D�H;�H;��H;��H;��H;��H;u�H;��H;��H;��H;��H;�H;B�H;��H;��H;�H;Q�H;��H;��H;z�H;�H;I�H;��H;��H;%�H;��H;�H;�H;�!H;�uG;2mF;��D;��B;7R@;�-=;�9;�5;��1;�-;�M*;=�';:�%;      yo8;B�8;ŏ9;u�:;��<;�c>;RR@;�/B;��C;�PE;�zF;h\G;��G;HiH;?�H;��H;C�H;q�H;?�H;J�H;r�H;�H;}�H;��H;��H;h�H;�H;��H;��H;3�H;��H;��H;��H;Q�H;K�H;?�H;�H;?�H;M�H;O�H;�H;��H;��H;/�H;��H;��H;�H;h�H;��H;��H;z�H;�H;n�H;H�H;>�H;q�H;C�H;��H;?�H;HiH;��G;g\G;�zF;�PE;��C;�/B;OR@;�c>;��<;u�:;ȏ9;4�8;      ��A;{B;pB;�C;��C;t�D;huE;xDF;J�F;��G;�H;fH;�H;��H;c�H;$�H;��H;�H;��H;��H;;�H;��H;��H;��H;H�H;��H;��H;��H;)�H;��H;��H;g�H;5�H;�H;��H;��H;��H;��H;��H;�H;3�H;g�H;��H;��H;&�H;��H;��H;��H;I�H;��H;��H;��H;8�H;��H;��H;�H;��H;!�H;c�H;��H;�H;fH;�H;��G;H�F;xDF;huE;t�D;��C;�C;pB;|B;      nDF;RF;�zF;�F;�G;�\G;�G;QH;&IH;��H;��H;��H;�H;��H; �H;I�H;	�H;K�H;��H;i�H;��H;��H;��H;g�H;��H;��H;��H;"�H;��H;��H;C�H;�H;��H;��H;��H;��H;��H;��H;��H;��H;��H;�H;A�H;��H;��H;!�H;��H;��H;��H;e�H;��H;��H;��H;i�H;��H;K�H;�H;H�H; �H;��H;�H;��H;��H;��H;&IH;QH;�G;�\G;�G;�F;�zF;sRF;      �H;	H;�!H;�8H;�TH;MsH;>�H;ثH;��H;��H;��H;��H;�H; �H;��H;
�H;��H;P�H;��H;��H;��H;��H;T�H;�H;��H;��H;�H;��H;r�H;A�H;��H;��H;��H;q�H;X�H;4�H;G�H;4�H;W�H;p�H;��H;��H;��H;?�H;p�H;��H;�H;��H;��H;�H;Q�H;��H;��H;��H;��H;Q�H;��H;	�H;��H; �H;�H;��H;��H;��H;��H;׫H;?�H;HsH;�TH;�8H;�!H;H;      ��H;7�H;��H;X�H;U�H;��H;T�H;��H;1�H;>�H;2�H;��H;�H;7�H;��H;k�H;��H;��H;��H;��H;��H;��H;
�H;��H;��H;#�H;��H;��H;2�H;��H;��H;t�H;N�H;�H;�H;�H;�H; �H;�H;�H;L�H;t�H;��H;��H;0�H;��H;��H;"�H;��H;��H;�H;��H;��H;��H;��H;��H;��H;k�H;��H;6�H;�H;��H;2�H;=�H;3�H;��H;U�H;��H;_�H;X�H;��H;C�H;      �H;_�H;8�H;��H;�H;q�H;��H;��H;��H;��H;��H;��H;Q�H;��H;��H;9�H;T�H;-�H;�H;��H;|�H;�H;��H;��H;"�H;��H;n�H;2�H;��H;��H;f�H;/�H;��H;��H;��H;��H;��H;��H;��H;��H;��H;1�H;f�H;��H;��H;2�H;p�H;��H;#�H;��H;��H;�H;y�H;��H;�H;-�H;Q�H;8�H;��H;��H;Q�H;��H;��H;��H;��H;��H;��H;p�H;
�H;��H;;�H;U�H;      �H;�H;-�H;}�H;�H;p�H;�H;��H;4�H;��H;�H;6�H;i�H;��H;��H;~�H;c�H;.�H;��H;��H;<�H;��H;��H;3�H;��H;��H;?�H;��H;��H;^�H;.�H;��H;��H;��H;��H;}�H;r�H;~�H;��H;��H;��H;��H;-�H;\�H;��H;��H;<�H;��H;��H;3�H;��H;��H;:�H;��H;��H;/�H;b�H;}�H;��H;��H;i�H;6�H;�H;��H;5�H;��H;�H;p�H;�H;}�H;(�H;�H;      V�H;��H;��H;��H;�H;/�H;\�H;��H;��H;��H;��H;�H;�H;�H;��H;��H;U�H;��H;��H;[�H;&�H;��H;B�H;��H;��H;D�H;��H;��H;e�H;1�H;��H;��H;��H;u�H;Q�H;Z�H;Z�H;Z�H;P�H;s�H;��H;��H;��H;.�H;f�H;��H;��H;C�H;��H;��H;@�H;��H;#�H;Z�H;��H;��H;U�H;��H;��H;��H;�H;�H;��H;��H;��H;��H;[�H;/�H;��H;��H;��H;��H;      U�H;_�H;[�H;V�H;j�H;��H;�H;��H;��H;��H;��H;n�H;<�H;�H;��H;��H;1�H;��H;��H;5�H;��H;h�H;�H;��H;d�H;�H;��H;v�H;/�H;��H;��H;��H;v�H;B�H;-�H;,�H;.�H;,�H;-�H;B�H;s�H;��H;��H;��H;/�H;v�H;��H;�H;f�H;��H;�H;h�H;��H;5�H;��H;��H;/�H;��H;��H;�H;?�H;n�H;��H;��H;��H;��H;�H;��H;g�H;U�H;Y�H;[�H;      W�H;Y�H;S�H;U�H;O�H;7�H;7�H;)�H;��H;��H;��H;��H;J�H;��H;��H;T�H;�H;��H;s�H;�H;��H;;�H;��H;��H;/�H;��H;��H;Q�H;��H;��H;��H;w�H;0�H;%�H;%�H; �H;��H; �H;%�H;%�H;-�H;z�H;��H;��H;��H;Q�H;��H;��H;0�H;��H;��H;;�H;��H;�H;s�H;��H;�H;T�H;��H;��H;H�H;��H;��H;��H;��H;)�H;7�H;:�H;G�H;S�H;S�H;P�H;      ��H;��H;��H;��H;��H;v�H;y�H;L�H;�H;��H;��H;w�H;5�H;��H;��H;p�H;��H;z�H; �H;��H;��H;*�H;��H;U�H;�H;��H;m�H;�H;��H;��H;s�H;C�H; �H;�H;�H;��H;��H;��H;�H;�H;�H;F�H;s�H;��H;��H;�H;m�H;��H;�H;T�H;��H;*�H;��H;��H; �H;|�H;��H;p�H;��H;��H;5�H;w�H;��H;��H;�H;L�H;y�H;y�H;��H;��H;��H;��H;      ��H;�H;��H;��H;��H;��H;��H;]�H;(�H;��H;��H;w�H;5�H;��H;��H;-�H;��H;i�H;�H;��H;U�H;��H;��H;O�H;��H;��H;U�H;�H;��H;��H;P�H;1�H;#�H;�H;��H;��H;��H;��H;��H;�H;"�H;4�H;P�H;��H;��H;�H;S�H;��H;��H;N�H;��H;��H;R�H;��H;�H;k�H;��H;-�H;��H;��H;5�H;w�H;��H;��H;(�H;\�H;��H;��H;��H;��H;��H;��H;      ��H;��H;��H;��H;��H;��H;q�H;Y�H;3�H;��H;��H;��H;!�H;��H;j�H;�H;��H;g�H;�H;��H;E�H;��H;��H;D�H;��H;��H;2�H;�H;��H;��H;[�H;0�H;��H;��H;��H;��H;��H;��H;��H;��H;��H;4�H;[�H;��H;��H;�H;1�H;��H;��H;A�H;��H;��H;D�H;��H;�H;h�H;��H;�H;l�H;��H;!�H;��H;��H;��H;3�H;W�H;q�H;��H;��H;��H;��H;��H;      ;�H;A�H;1�H;�H;�H;��H;��H;t�H;=�H;��H;��H;X�H;�H;��H;��H;(�H;��H;A�H;��H;��H;A�H;��H;q�H;�H;��H;��H;D�H;�H;��H;w�H;]�H;5�H;��H;��H;��H;��H;��H;��H;��H;��H;��H;7�H;]�H;w�H;��H;�H;C�H;��H;��H;�H;r�H;��H;A�H;��H;��H;B�H;��H;(�H;��H;��H;�H;Y�H;��H;��H;@�H;r�H;��H;��H;�H;�H;0�H;8�H;      ��H;��H;��H;��H;��H;��H;q�H;Y�H;3�H;��H;��H;��H;!�H;��H;l�H;�H;��H;g�H;�H;��H;G�H;��H;��H;C�H;��H;��H;2�H;�H;��H;��H;[�H;1�H;��H;��H;��H;��H;��H;��H;��H;��H;��H;3�H;[�H;��H;��H;�H;1�H;��H;��H;A�H;��H;��H;D�H;��H;�H;h�H;��H;�H;j�H;��H;!�H;��H;��H;��H;3�H;W�H;q�H;��H;��H;��H;��H;��H;      ��H;�H;��H;��H;��H;��H;��H;]�H;(�H;��H;��H;w�H;5�H;��H;��H;-�H;��H;i�H;�H;��H;V�H;��H;��H;O�H;��H;��H;T�H;�H;��H;��H;P�H;1�H;#�H;�H;��H;��H;��H;��H;��H;�H;"�H;5�H;P�H;��H;��H;�H;T�H;��H;��H;M�H;��H;��H;R�H;��H;�H;k�H;��H;-�H;��H;��H;5�H;w�H;��H;��H;(�H;\�H;��H;��H;��H;��H;��H;��H;      ��H;��H;��H;��H;��H;u�H;y�H;L�H;�H;��H;��H;w�H;5�H;��H;��H;p�H;��H;z�H; �H;��H;��H;*�H;��H;U�H;�H;��H;m�H;�H;��H;��H;s�H;C�H; �H;�H;�H;��H;��H;��H;�H;�H;�H;F�H;s�H;��H;��H;�H;o�H;��H;�H;T�H;��H;*�H;��H;��H; �H;|�H;��H;p�H;��H;��H;5�H;w�H;��H;��H;�H;L�H;y�H;{�H;��H;��H;��H;��H;      Z�H;V�H;U�H;V�H;L�H;7�H;9�H;(�H;��H;��H;��H;��H;H�H;��H;��H;T�H;�H;��H;s�H;�H;��H;;�H;��H;��H;0�H;��H;��H;Q�H;��H;��H;��H;w�H;.�H;#�H;%�H; �H;��H; �H;%�H;#�H;-�H;|�H;��H;��H; �H;Q�H;��H;��H;/�H;��H;��H;;�H;��H;�H;s�H;��H;�H;T�H;��H;��H;H�H;��H;��H;��H; �H;&�H;9�H;:�H;G�H;W�H;P�H;V�H;      U�H;_�H;[�H;T�H;i�H;��H;��H;��H;��H;��H;��H;n�H;=�H;�H;��H;��H;/�H;��H;��H;7�H;��H;h�H;�H;��H;f�H;�H;��H;v�H;-�H;��H;��H;��H;u�H;B�H;-�H;,�H;.�H;,�H;-�H;B�H;s�H;��H;��H;��H;1�H;v�H;��H;�H;d�H;��H;�H;h�H;��H;5�H;��H;��H;/�H;��H;��H;�H;<�H;n�H;��H;��H;��H;��H;��H;��H;i�H;U�H;[�H;[�H;      V�H;��H;��H;��H; �H;-�H;[�H;��H;��H;��H;��H;�H;�H;�H;��H;��H;T�H;��H;��H;Z�H;'�H;��H;A�H;��H;��H;D�H;��H;��H;e�H;/�H;��H;��H;��H;s�H;P�H;Z�H;Z�H;Z�H;Q�H;u�H;��H;��H;��H;/�H;f�H;��H;��H;C�H;��H;��H;@�H;��H;#�H;[�H;��H;��H;U�H;��H;��H;�H;�H;�H;��H;��H;��H;��H;\�H;1�H;��H;��H;��H;��H;       �H;�H;+�H;{�H;�H;j�H;�H;��H;5�H;��H;�H;6�H;i�H;��H;��H;~�H;c�H;.�H;��H;��H;>�H;��H;��H;3�H;��H;��H;?�H;��H;��H;^�H;-�H;��H;��H;��H;��H;~�H;r�H;}�H;��H;��H;��H;��H;.�H;\�H;��H;��H;<�H;��H;��H;3�H;��H;��H;;�H;��H;��H;/�H;b�H;�H;��H;��H;i�H;6�H;�H;��H;7�H;��H;�H;n�H;�H;{�H;+�H;�H;      �H;[�H;>�H;��H;	�H;l�H;��H;��H;��H;��H;��H;��H;Q�H;��H;��H;8�H;S�H;+�H;�H;��H;}�H;�H;��H;��H;#�H;��H;n�H;2�H;��H;��H;f�H;.�H;��H;��H;��H;��H;��H;��H;��H;��H;��H;1�H;f�H;��H;��H;2�H;p�H;��H;"�H;��H;��H;�H;z�H;��H;�H;.�H;T�H;;�H;��H;��H;Q�H;��H;��H;��H;��H;��H;��H;p�H;�H;��H;A�H;[�H;      ��H;8�H;��H;X�H;U�H;��H;U�H;��H;1�H;=�H;3�H;��H;�H;6�H;��H;k�H;��H;��H;��H;��H;��H;��H;�H;��H;��H;"�H;��H;��H;2�H;��H;��H;t�H;M�H;�H;�H; �H;�H;�H;�H;�H;M�H;v�H;��H;��H;2�H;��H;��H;#�H;��H;��H;�H;��H;��H;��H;��H;��H;��H;l�H;��H;4�H;�H;��H;0�H;>�H;4�H;��H;T�H;��H;b�H;X�H;��H;A�H;      �H;H;�!H;�8H;�TH;GsH;>�H;ثH;��H;��H;��H;��H;�H; �H;��H;
�H;��H;P�H;��H;��H;��H;��H;S�H;
�H;��H;��H;�H;��H;p�H;@�H;��H;��H;��H;p�H;W�H;4�H;G�H;2�H;X�H;p�H;��H;��H;��H;@�H;q�H;��H;�H;��H;��H;�H;S�H;��H;��H;��H;��H;Q�H;��H;	�H;��H; �H;�H;��H;��H;��H;��H;ثH;<�H;GsH;�TH;�8H;�!H;H;      sDF;{RF;�zF;�F;�G;�\G;
�G;TH;%IH;��H;��H;��H;�H;��H;��H;I�H;	�H;I�H;��H;i�H;��H;��H;��H;g�H;��H;��H;��H;!�H;��H;��H;A�H;�H;��H;��H;��H;��H;��H;��H;��H;��H;��H;�H;C�H;��H;��H;"�H;��H;��H;��H;e�H;��H;��H;��H;i�H;��H;L�H;�H;I�H; �H;��H;�H;��H;��H;��H;%IH;SH;�G;�\G;�G;�F;�zF;nRF;      ��A;|B;pB;�C;��C;t�D;huE;xDF;H�F;��G;�H;fH;�H;��H;c�H;#�H;��H;�H;��H;��H;;�H;��H;��H;��H;I�H;��H;��H;��H;&�H;��H;��H;f�H;3�H;�H;��H;��H;��H;��H;��H;�H;3�H;j�H;��H;��H;&�H;��H;��H;��H;H�H;��H;��H;��H;:�H;��H;��H;�H;��H;$�H;c�H;��H;�H;fH;�H;��G;J�F;yDF;huE;t�D;��C;�C;pB;{B;      |o8;?�8;͏9;r�:;��<;�c>;KR@;�/B;��C;�PE;�zF;g\G;��G;HiH;?�H;��H;C�H;o�H;>�H;H�H;r�H;�H;|�H;��H;��H;g�H;�H;��H;��H;2�H;��H;��H;��H;N�H;J�H;@�H;�H;?�H;M�H;Q�H;��H;��H;��H;0�H;��H;��H;�H;h�H;��H;��H;|�H;�H;o�H;J�H;?�H;s�H;B�H;��H;?�H;HiH;��G;h\G;�zF;�PE;��C;�/B;LR@;�c>;��<;p�:;Џ9;2�8;      �S%;V�%;J�';�M*;�-;��1;�5;�9;�-=;7R@;��B;��D;1mF;�uG;�!H;�H;�H;��H;%�H;��H;��H;I�H;�H;}�H;��H;��H;V�H;�H;��H;��H;B�H;�H;��H;��H;��H;��H;u�H;��H;��H;��H;��H;�H;D�H;��H;��H;�H;S�H;��H;��H;|�H;�H;I�H;��H;��H;%�H;��H;�H;�H;�!H;�uG;1mF;��D;��B;5R@;�-=;�9;�5;��1;�-;�M*;B�';D�%;      �W;�x;�;�
;��;�;� ;��(;��/;I6;��;;�?;C;�PE;�F;�G;�eH;S�H;��H;6�H;`�H;��H;G�H;�H;}�H;��H;��H;��H;�H;��H;��H;c�H;:�H;)�H;��H;��H;��H;��H;��H;)�H;:�H;d�H;��H;��H;�H;��H;��H;��H;}�H;
�H;E�H;��H;`�H;7�H;��H;V�H;�eH;�G;�F;�PE;C;�?;��;;
I6;��/;��(;� ;�;ȅ;�
;�;�x;      r��:Ɔ: ʒ:��:��:��:W��:_�	;�v;�#;ڷ-;�5;�L<;��@;�(D;,DF;��G;�HH;{�H;�H;��H;`�H;��H;u�H;7�H;��H;��H;��H;z�H;<�H;�H;��H;��H;{�H;N�H;@�H;@�H;@�H;N�H;}�H;��H;��H; �H;:�H;w�H;��H;��H;��H;8�H;r�H;��H;a�H;��H;�H;|�H;�HH;��G;-DF;�(D;��@;�L<;�5;ڷ-;�#;�v;`�	;W��:��:��:��:ʒ:�ņ:      X-.�H��x�깠}K��"
9�]:��k:�M�:ͤ�:�y;��;� $;��/;��8;��>;$C;0�E;�\G;_8H;ԥH;�H;4�H;��H;J�H;��H;i�H;��H;��H;��H;��H;T�H;,�H;��H;��H;��H;��H;��H;��H;��H;��H;��H;.�H;T�H;��H;��H;��H;��H;k�H;��H;F�H;��H;4�H;�H;ץH;a8H;�\G;3�E;$C;��>;��8;��/;� $;��;�y;Ϥ�:�M�:��k:�]: #
9�}K����x��      1Q^�X��F�Ƣ)�+��ζ� �<� >S�hn:B��:��:��;T�;�M*;�5;�c=;upB;��E;�JG;b8H;|�H;��H;%�H;>�H;��H;��H;��H;��H;�H;��H;��H;��H;o�H;�H;�H;
�H;��H;�H;�H;�H;o�H;��H;��H;��H; �H;��H;��H;��H;��H;;�H; �H;��H;z�H;e8H;�JG;��E;tpB;�c=;��5;�M*;V�;��;��:B��:tn: >S� �<��ζ�+�Ƣ)��F�X�      k���>���"���ѻ,���ǐ�_X�,6�<	���tK�,?":�M�:Zb�:di;;�%;f�3;�<;M0B;��E;�\G;�HH;U�H;��H;p�H;�H;I�H;Q�H;��H;.�H;1�H;��H;��H;��H;y�H;l�H;k�H;H�H;k�H;l�H;z�H;��H;��H;��H;/�H;+�H;��H;P�H;L�H;�H;j�H;��H;U�H;�HH;�\G;��E;N0B;�<;g�3;;�%;di;Zb�:�M�:,?": uK�8	��,6�_X�ǐ�(����ѻ"��B���      t�n�zmj���]���J�\�1�64�4������	x��W��y�`)
9��:k��:�;O�#;^�2;�<;upB;4�E;��G;�eH;�H;F�H;��H;�H;��H;��H;P�H;_�H;N�H;'�H;�H;��H;��H;��H;��H;��H;��H;��H;�H;'�H;N�H;^�H;N�H;��H;��H;	�H;��H;B�H;��H;�eH;��G;6�E;upB;�<;\�2;P�#;�;k��:��:`)
9�y��W��	x����5��54�\�1���J���]�|mj�      F<ͼ��ɼ�����֯�ж��ㄼ��Y��*�����s��X�rrѺ��<?Q:���:��
;S�#;i�3;�c=;$C;-DF;�G;�H;��H;�H;H�H;	�H;i�H;8�H;x�H;��H;v�H;M�H;h�H;!�H;�H; �H; �H;!�H;h�H;L�H;w�H;��H;z�H;4�H;i�H;�H;J�H; �H;��H;�H;�G;-DF;$C;�c=;j�3;S�#;��
;���:8?Q:��rrѺX��s������*���Y�ㄼж���֯�������ɼ      ��'�+�$������  ���ۼ����+����]��X!�H>ۻ�+��r*����>:���:�;:�%;�5;��>;�(D;�F;�!H;=�H;_�H; �H;��H;��H;��H;~�H;��H;��H;��H;��H;�H;c�H;��H;c�H;�H;��H;��H;��H;��H;~�H;��H;��H;��H;�H;`�H;;�H;�!H;�F;�(D;��>;�5;<�%;�;���:�>:��r*��+��G>ۻ�X!���]��+�������ۼ�  �����+�$�      Ǹ���v����w�j�c��J�҄-�~��;缉沼ㄼ��;������j���5����<?Q:m��:fi;�M*;��8;��@;�PE;�uG;EiH;��H;��H;�H;2�H;��H;��H;��H;	�H;��H;��H;��H;��H;��H;��H;��H;��H;��H;�H;��H;��H;��H;2�H;�H;��H;��H;BiH;�uG;�PE;��@;��8;�M*;hi;k��:<?Q: �깝5��j��������;�ㄼ�沼�;�~�ф-��J�j�c���w��v��      }Hͽڪɽ�;��!"�� ��ɸ����[�z0�u��+<ͼξ��f�J�����j��q*�����:^b�:V�;��/;�L<;C;4mF;��G;�H;�H;�H;�H;P�H;b�H;��H;7�H;C�H;/�H;+�H;�H;�H;�H;+�H;0�H;C�H;7�H;��H;b�H;M�H;�H;�H;�H;�H;��G;/mF;C;�L<;��/;V�;`b�:��:��p*��j�����f�J�ξ��+<ͼu��z0���[�ɸ�� ��!"���;��ڪɽ      ��$-������ֱ�ƽaP���v���J�K����ۼ��f�J������+��vrѺp)
9�M�:��;� $;�5;��?;��D;g\G;fH;��H;��H;��H;��H;+�H;��H;d�H;��H;p�H;i�H;u�H;M�H;u�H;g�H;n�H;�H;f�H;�H;+�H;��H;��H;��H;��H;fH;d\G;��D;��?;�5;� $;��;�M�:`)
9vrѺ�+������f�J�����ۼK���J��v��aP��ƽֱ轆����$-�       j�Zde�]0X��D�i{+�������z㻽\���WDX������ۼξ����;�G>ۻX��y�(?":��:��;ٷ-;��;;��B;�zF;�H;��H;��H;,�H;��H;��H;��H;~�H;��H;��H;��H;��H;��H;��H;��H;��H;��H;�H;��H;��H;��H;,�H;��H;��H;�H;�zF;��B;��;;ڷ-;��;��:,?":$�y�X�F>ۻ��;�ξ����ۼ���WDX�\���z㻽��콅��i{+��D�]0X�Zde�      ��Sh��m���I���|x���O��C(���Ҫɽ����WDX�K��+<ͼㄼ�X!��s���W��tK�F��:�y;�#;
I6;9R@;�PE;��G;��H;��H;7�H;��H;��H;��H;��H;��H;��H;��H;��H;��H;��H;��H;��H;��H;��H;��H;��H;��H;7�H;��H;��H;��G;�PE;7R@;
I6;�#;�y;F��:�tK��W��s���X!�ㄼ+<ͼK��WDX�����Ҫɽ���C(���O��|x��I��m��Sh��      @����������$�;jɰ��G�� j�;�5��	�Ҫɽ\����J�v���沼��]�����	x�@	��hn:Ϥ�:�v;��/;�-=;��C;G�F;&IH;��H;,�H;��H;)�H;��H;��H;��H;�H;�H;%�H;4�H;%�H;�H;�H;��H;��H;��H;)�H;��H;,�H;��H;&IH;J�F;��C;�-=;��/;�v;ͤ�:dn:<	���	x������]��沼v���J�\���Ҫɽ�	�;�5� j��G��jɰ�$�;��徺���      �2�X�-�"�/E�����BKɾm����s�;�5���z㻽�v��z0��;��+���*����+6��=S��M�:\�	;��(;�9;�/B;vDF;WH;իH;��H;��H;��H;�H;��H;�H;B�H;P�H;K�H;j�H;N�H;O�H;B�H;�H;��H;�H;��H;��H;��H;իH;VH;zDF;�/B;�9;��(;_�	;�M�:�=S�)6�����*��+���;�z0��v��z㻽��;�5���s�m��BKɾ����/E�"�X�-�      (3s�"cm�=�\�j�C�7�%�����TҾm�� j��C(����aP����[�������Y�8��aX�8�<���k:K��: � ;�5;HR@;fuE;
�G;8�H;N�H;��H;
�H;Q�H;{�H;4�H;t�H;��H;g�H;��H;g�H;��H;r�H;2�H;{�H;Q�H;�H;��H;N�H;7�H;
�G;huE;GR@;�5; � ;Q��:��k:8�<�_X�:����Y�������[�aP����콭C(� j�m���TҾ���7�%�j�C�=�\�"cm�      �ޞ�������bF�A�W�Y�-����BKɾ�G����O����ƽɸ��҄-���ۼㄼ64�ǐ��ζ��]:���:�;��1;�c>;q�D;�\G;HsH;��H;q�H;j�H;.�H;��H;9�H;{�H;��H;��H;��H;��H;��H;{�H;6�H;��H;.�H;g�H;m�H;��H;GsH;�\G;q�D;�c>;��1;�;	��:�]:�ζ�ǐ�64�ㄼ��ۼ҄-�ɸ��ƽ�����O��G��BKɾ���Y�-�A�W�bF�������      ��ſ���Nw���ޞ�����A�W�7�%�����jɰ��|x�i{+�ֱ� ���J��  �Ѷ��\�1�+���+�p"
9��:��;�-;��<;��C;�G;�TH;T�H;�H;��H;��H;c�H;A�H;��H;��H;��H;��H;��H;��H;��H;@�H;d�H;��H;��H;�H;T�H;�TH;�G;��C;��<;�-;��; �:P"
9+�*���\�1�Ѷ���  ��J� ��ֱ�i{+��|x�jɰ�����7�%�A�W������ޞ�Nw�����      ����� �Կp���ޞ�bF�j�C�/E�%�;�I���D���!"��k�c���֯���J��ѻɢ)��}K� ��:�
;�M*;u�:;�C;�F;�8H;\�H;��H;}�H;��H;M�H;I�H;��H;��H;��H;
�H;��H;��H;��H;H�H;K�H;��H;z�H;��H;\�H;�8H;�F;�C;p�:;�M*;�
;&��:�}K�ɢ)��ѻ��J��֯��k�c�!"�����D��I��%�;/E�j�C�bF��ޞ�p�� �Կ��      ��������� �ԿNw�����=�\�"����n��]0X�����;����w����������]�%���F�����ɒ:��;;�';��9;"pB;�zF;�!H;��H;>�H;#�H;��H;T�H;I�H;��H;��H;��H;�H;��H;��H;��H;H�H;T�H;��H; �H;;�H;��H;�!H;�zF;"pB;��9;=�';��;�ɒ:����F�$�黯�]����������w��;�����]0X�n�����"�=�\����Nw�� �Կ��𿞏�      !$�������忊�����"cm�X�-�����Sh��Zde�$-�۪ɽ�v��+�$���ɼ|mj�>���X�����ņ:wx;D�%;2�8;pB;qRF;H;4�H;[�H;�H;v�H;N�H;D�H;��H;��H;��H;3�H;��H;��H;��H;B�H;O�H;v�H;�H;X�H;4�H;H;pRF;pB;.�8;I�%;wx;�ņ:���X�=���}mj���ɼ+�$��v��۪ɽ$-�Zde�Sh������X�-�"cm��������忞����      gܿ6�ֿ�aǿ@^��1���\o���7����iþ�(���-=��` �A���_�4]�3p����I�Y�ѻ��)���R���::�
;�*;�:;գB;BIF;/�G;�lH;5�H;��H;k�H;��H;��H;|�H;��H;5�H;��H;5�H;��H;|�H;��H;��H;k�H;��H;2�H;�lH;0�G;BIF;գB;�:;�*;:�
;��:��R���)�X�ѻ��I�3p��4]��_�A���` ��-=��(���iþ����7�\o�1���@^���aǿ6�ֿ      6�ֿFpѿ�¿������bXi�ҕ3��
�XD��Hl��D�9��.���R��'\� �ix��5�E��ͻ�$�@  �Ǎ�:H�;��*;5�:;�B;#UF;��G;UnH;ѡH;޷H;��H;��H;��H;��H;��H;J�H;��H;J�H;��H;��H;��H;��H;��H;۷H;ΡH;UnH;��G;"UF;�B;1�:;��*;H�;ˍ�:`  ��$��ͻ5�E�ix�� �'\��R���.��D�9�Hl��XD���
�ҕ3�bXi��������¿Fpѿ      �aǿ�¿����������"Y��f'�����:o���.}��k/����(ڟ�'<Q�1#�ע��(;�4���8�� D7���:��;�,;��;;�C;CwF;#�G;�rH;\�H;¸H;A�H;&�H;"�H;��H;��H;x�H;��H;x�H;��H;��H; �H;'�H;A�H;��H;Y�H;�rH;#�G;AwF;�C;��;;�,;��;��: E7�7��3����(;�ע�1#�'<Q�(ڟ�����k/��.}�:o�������f'��"Y�����������¿      @^������m���\o���@�+�'�޾����<ce�3��ïڽ����g@������R���O*�NG������E^9(��:;�d.;�<;��C;7�F;��G;�yH;ȥH;9�H;O�H;��H;��H;�H;�H;��H;C�H;��H;�H;�H;��H;��H;O�H;7�H;ťH;�yH;��G;7�F;��C;��<;�d.;;*��:�E^9���LG���O*��R������g@�����ïڽ3��<ce�����'�޾+���@�\o�m�������      1����������\o��!J�M�#��\��YD������~PH�����b��"C��� +���ټ,����򿐻����:)��:W�;�Y1;>;�0D;��F;uH;o�H;��H;-�H;��H;��H;6�H;��H;|�H;��H;��H;��H;z�H;��H;5�H;��H;��H;*�H;��H;o�H;wH;��F;�0D;>;�Y1;W�;+��:�:���𿐻��+����ټ� +�"C���b�����~PH�����YD���\��M�#��!J�\o��������      \o�bXi��"Y���@�N�#��
��о�A���i���(����zr���_��5��ɺ�w�`��<��k�d�L�\�ВX:�P�:�`;��4;˧?;��D;�8G;�0H;ċH;��H;��H;3�H;��H;��H;(�H;��H;<�H;��H;<�H;��H;(�H;��H;��H;3�H;��H;��H;ċH;�0H;�8G;��D;ħ?;��4;�`;�P�:ȒX:T�\�i�d��<��x�`��ɺ��5��_�zr�������(��i��A���о�
�N�#���@��"Y�bXi�      ��7�ҕ3��f'�+��\���о�����.}��-=�~
���Ľ^��0:����������7�%GĻŃ$��N�����:�{;�D&;,8;*JA;"�E;�G;�LH;�H;��H;U�H;�H;4�H;��H;��H;M�H;��H;E�H;��H;M�H;��H;��H;5�H;�H;T�H;��H;�H;�LH;�G;�E;&JA;,8;�D&;�{;���:�N��$�%GĻ�7���������0:�^����Ľ~
��-=��.}������о�\��+��f'�ҕ3�      ���
�����'�޾YD���A���.}�,�D�kt���ڽ�!��\����a�ļ�
v�A��ɿ���IɺXS�9���:'(;�-;��;;��B;�IF;��G;<fH;ʝH;�H;P�H;��H;��H;��H;��H;��H;�H;��H;�H;��H;��H;��H;��H;��H;P�H;�H;ȝH;:fH;��G;�IF;��B;��;;�-;)(;���:XS�9�Iɺʿ��A���
v�a�ļ���\��!����ڽkt�,�D��.}��A��YD��'�޾�����
�      �iþXD��:o�����������i��-=�kt����R��nys�~ +���}񗼘(;�0�ѻ�s@���!�D4j:�P�:��;�D3;]�>;0FD;��F;�	H;\|H;��H;��H;Z�H;!�H;#�H;��H;L�H;b�H;��H;�H;��H;b�H;J�H;��H;%�H; �H;Y�H;��H;��H;Y|H;�	H;��F;-FD;\�>;�D3;��;�P�:D4j:��!��s@�0�ѻ�(;�}���~ +�nys��R����kt��-=��i���������:o��XD��      �(��Hl���.}�<ce�~PH���(�~
���ڽ�R���{�G�6�� �1p��f�`�Ш��,��2IҺ�L^9���:��;�~(;K�8;JA;"|E;=jG;�=H;i�H;�H;R�H;��H;V�H;��H;��H;�H;��H; �H;z�H; �H;��H;�H;��H;��H;W�H;��H;N�H;�H;g�H;�=H;:jG; |E;JA;K�8;�~(;��;���:�L^96IҺ�,��Ш�f�`�1p��� �G�6��{��R����ڽ~
���(�~PH�<ce��.}�Hl��      �-=�C�9��k/�3��������Ľ�!��nys�G�6�(#��ɺ��vz����D^��f�$�X~�l�r:(��: �;�Y1;I=;SxC;HwF;L�G;/fH;o�H;��H;��H;��H;��H;�H;�H;��H;��H;��H;��H;��H;��H;��H;
�H;�H;��H;��H;��H;��H;o�H;.fH;H�G;DwF;QxC;I=;�Y1;��;(��:x�r:h~�g�$�D^������vz��ɺ�(#�G�6�nys��!����Ľ����3���k/�C�9�      �` ��.�����ïڽ�b��zr��^��\�~ +�� ��ɺ�C��O*�Iͻ�5R�ǅ��:E��:��;�);u8;��@;�*E;�8G;o$H;r�H;i�H;"�H;V�H;��H;��H;��H;.�H;��H;"�H;�H;Q�H;�H;"�H;��H;.�H;��H;��H;��H;U�H;"�H;h�H;p�H;l$H;�8G;�*E;��@;u8;�);��;K��:�:ǅ��5R�Hͻ�O*�C��ɺ�� �~ +�\�^��zr���b��ïڽ��.��      A���R��(ڟ�����"C���_�0:������1p���vz��O*��4ֻk� �����09\�:1;m� ;�D3;e�=;̐C;lF;��G;�\H;ǗH;y�H;0�H;o�H;��H;��H;�H;+�H;;�H;��H;��H;��H;��H;��H;;�H;+�H;�H;��H;��H;n�H;0�H;v�H;ǗH;�\H;��G;	lF;̐C;c�=;�D3;m� ;1;Z�:��09 ���k��4ֻ�O*��vz�0p���輨��0:��_�#C������(ڟ��R��      �_�&\�&<Q�g@�� +��5�����`�ļ|�e�`����Hͻk��Hɺ |6�\�:Q�:<�;�d.;m�:;A�A;O|E;�NG;n'H;-�H;��H;��H;��H;\�H;{�H;��H;d�H;)�H;��H;@�H;��H;2�H;��H;@�H;��H;)�H;g�H;��H;{�H;Y�H;��H;��H;��H;+�H;k'H;�NG;O|E;A�A;m�:;�d.;?�; Q�:X�: {6��Hɺk�Hͻ���d�`�|�a�ļ�����5�� +�g@�&<Q�&\�      4]� �0#�������ټ�ɺ������
v��(;�Ш�D^���5R�&��� }6����:��:�;<�*;�+8;�!@;~�D;��F;$�G;fH;��H;��H;пH;��H;�H;��H;T�H;��H;��H;��H;��H;[�H;��H;[�H;��H;��H;��H;��H;T�H;��H;�H;��H;ϿH;��H;��H;�eH;�G;��F;|�D;�!@;�+8;=�*;�;��:���: }6�&����5R�D^��Ш��(;��
v������ɺ���ټ����0#� �      2p��hx��ע��R��+��w�`��7�A��.�ѻ�,��d�$�ǅ���09X�:��:�;�~(;�Z6;��>;��C;IF;�G;EH;x�H;�H;ܹH;A�H;\�H;G�H;,�H;�H;��H;��H;C�H;�H;��H;��H;��H;�H;B�H;��H;��H;�H;,�H;C�H;\�H;?�H;ܹH;�H;s�H;EH;�G;IF;��C;��>;�Z6;�~(;�;��:X�:��09ǅ�d�$��,��-�ѻB���7�w�`�+���R��ע�ix��      ��I�2�E��(;��O*����<��"GĻȿ���s@�0IҺP~��:V�:�P�:�;�~(;*�5;�>;]C;_�E;�cG;i$H;(|H;j�H;P�H;��H;��H;m�H;�H;S�H;��H;��H;��H;��H;t�H; �H;&�H; �H;t�H;��H;��H;��H;��H;Q�H;	�H;m�H;��H;��H;O�H;e�H;#|H;i$H;�cG;`�E;]C;�>;+�5;�~(;�; Q�:V�:�:h~�0IҺ�s@�ɿ��"GĻ�<�����O*��(;�5�E�      Z�ѻ�ͻ0���LG��򿐻u�d�Ń$��Iɺ��!��L^9x�r:E��:1;;�;=�*;�Z6;�>;Y�B;��E;9G;�	H;/nH;I�H;x�H;ؽH;��H;��H;	�H;��H;6�H;��H;��H;4�H;/�H;��H;:�H;]�H;9�H;��H;/�H;2�H;��H;��H;4�H;}�H;�H;��H;��H;ؽH;s�H;E�H;.nH;�	H;9G;��E;Y�B;�>;�Z6;<�*;<�;1;E��:x�r:�L^9��!��Iɺă$�q�d�𿐻KG��0����ͻ      {�)��$�/��������H�\��N��PS�9H4j:���:.��:��;l� ;�d.;�+8;��>;ZC;��E;�)G;��G;CdH;��H;ȫH;��H;��H;m�H;�H;�H;��H;��H;��H;z�H;��H;��H;4�H;j�H;��H;j�H;4�H;��H;��H;|�H;��H;��H;��H;�H;��H;k�H;��H;��H;īH;��H;=dH;��G;�)G;��E;ZC;��>;�+8;�d.;l� ;��;(��:���:P4j:PS�9�N��0�\����
���/���$�      P�R�0�� B7��E^9�:ĒX:���:���:�P�:��; �;�);�D3;i�:;�!@;�C;]�E;9G;��G;�`H;��H;K�H;M�H;��H;v�H;k�H;��H;��H;��H;�H;��H;?�H; �H;��H;c�H;��H;��H;��H;c�H;��H;�H;@�H;��H;�H;��H;��H;��H;h�H;u�H;��H;J�H;K�H;��H;�`H;��G;9G;\�E;�C;�!@;i�:;�D3;�);��;��;�P�:���:���:ВX:�:�E^9 B7����      ��:퍨:��:��:��:�P�:�{;&(;��;�~(;�Y1;u8;c�=;A�A;|�D;IF;�cG;�	H;CdH;��H;z�H;�H;d�H;)�H;�H;u�H;��H;��H;[�H;�H;��H;��H;��H;�H;|�H;��H;��H;��H;|�H;�H;��H;��H;��H;�H;X�H;��H;}�H;t�H;�H;#�H;d�H;�H;w�H;��H;AdH;�	H;�cG;IF;|�D;A�A;c�=;u8;�Y1;�~(;��;&(;�{;�P�:��: ��:��:ˍ�:      A�
;e�;�;	;X�;a;�D&;�-;�D3;M�8; I=;��@;͐C;R|E;��F;�G;i$H;1nH;��H;M�H;�H;��H;n�H;T�H;��H;��H;�H;��H;��H;A�H;X�H;.�H;��H;V�H;��H;��H;��H;��H;��H;V�H;��H;,�H;W�H;;�H;��H;��H;�H;��H;��H;N�H;k�H;��H;
�H;N�H;��H;/nH;i$H;�G;��F;Q|E;͐C;��@; I=;N�8;�D3;�-;�D&;a;l�;	;�;`�;      �*;��*;�,;�d.;�Y1;��4;!,8;��;;`�>;JA;UxC;�*E;lF;�NG;#�G;EH;'|H;I�H;ȫH;Q�H;g�H;p�H;��H;0�H;.�H;��H;C�H;!�H;��H;�H;��H;��H;�H;r�H;��H;��H;��H;��H;��H;r�H;�H;��H;��H;	�H;��H;!�H;A�H;��H;.�H;,�H;��H;p�H;b�H;Q�H;ȫH;I�H;$|H;EH;#�G;�NG;lF;�*E;SxC;JA;`�>;��;;!,8;��4;�Y1;�d.;�,;z�*;      2�:;B�:;��;;�<;>;ȧ?;1JA;��B;1FD;!|E;JwF;�8G;��G;p'H;fH;v�H;i�H;z�H;��H;��H;%�H;S�H;/�H;�H;P�H;��H;��H;j�H;��H;��H;O�H;��H;U�H;��H;��H;��H;��H;��H;��H;��H;P�H;��H;N�H;��H;��H;j�H;��H;��H;Q�H;�H;,�H;S�H;"�H;��H;��H;{�H;g�H;v�H;fH;p'H;��G;�8G;HwF;!|E;1FD;��B;0JA;ȧ?;>;�<;��;;5�:;      ߣB;!�B;�C;ĐC;�0D;��D;"�E;�IF;��F;;jG;K�G;q$H;�\H;2�H;��H;�H;V�H;ܽH;��H;|�H;�H;��H;3�H;U�H;��H;��H;2�H;y�H;b�H;/�H;��H;
�H;g�H;��H;��H;��H;��H;��H;��H;��H;e�H;
�H;��H;,�H;^�H;y�H;0�H;��H;��H;T�H;0�H;��H;�H;|�H;��H;޽H;S�H;�H;��H;1�H;�\H;q$H;K�G;8jG;��F;�IF;"�E;��D;�0D;ĐC;�C;"�B;      NIF;0UF;6wF;3�F;��F;�8G;��G;��G;�	H;�=H;/fH;u�H;ǗH;��H;��H;ܹH;��H;��H;j�H;j�H;r�H;��H;��H;��H;��H;/�H;^�H;B�H;��H;�H;��H;Y�H;n�H;��H;��H;��H;��H;��H;��H;��H;k�H;Y�H;��H;|�H;��H;B�H;[�H;0�H;��H;��H;��H;��H;n�H;j�H;j�H;��H;��H;ٹH;��H;��H;ǗH;u�H;/fH;�=H;�	H;��G;��G;�8G;��F;4�F;9wF;#UF;      <�G;��G;$�G;��G;{H;�0H;�LH;?fH;_|H;k�H;p�H;m�H;v�H;��H;ҿH;D�H;��H;��H;�H;��H;��H;�H;B�H;��H;,�H;a�H;5�H;��H;��H;��H;�H;g�H;��H;��H;��H;��H;��H;��H;��H;��H;��H;g�H;�H;��H;��H;��H;2�H;`�H;0�H;��H;A�H;�H;�H;��H;�H;��H;��H;A�H;ҿH;��H;v�H;m�H;p�H;i�H;`|H;=fH;�LH;�0H;�H;��G;$�G;��G;      �lH;XnH;�rH;�yH;r�H;ȋH;�H;ҝH;ťH;	�H;��H;)�H;1�H;��H;��H;^�H;n�H;�H;�H;��H;��H;��H;"�H;n�H;u�H;C�H;��H;k�H;��H;#�H;A�H;q�H;��H;��H;��H;��H;��H;��H;��H;��H;��H;q�H;A�H;�H;��H;j�H;��H;C�H;u�H;m�H;!�H;��H;��H;��H;�H;�H;m�H;^�H;��H;��H;1�H;(�H;��H;�H;ƥH;ҝH;�H;ǋH;{�H;�yH;�rH;anH;      J�H;֡H;X�H;̥H;��H;��H;��H;!�H;��H;U�H;��H;\�H;r�H;]�H;�H;H�H;�H;�H;��H;��H;\�H;��H;��H;��H;[�H;��H;��H;��H;�H;H�H;d�H;��H;��H;��H;��H;��H;��H;��H;��H;��H;��H;��H;d�H;G�H;�H;��H;��H;��H;\�H;��H;��H;��H;X�H;��H;��H;�H;�H;H�H;�H;]�H;r�H;Z�H;��H;R�H;��H; �H;��H;��H;�H;̥H;[�H;̡H;      ��H;�H;̸H;<�H;<�H;��H;^�H;W�H;d�H;��H;��H;��H;��H;��H;��H;0�H;W�H;3�H;��H;�H;�H;>�H;�H;��H;%�H;|�H;��H;!�H;G�H;\�H;{�H;y�H;��H;��H;��H;��H;��H;��H;��H;��H;��H;{�H;{�H;Z�H;E�H;!�H;��H;|�H;%�H;��H;�H;<�H;�H;	�H;��H;3�H;T�H;/�H;��H;��H;��H;��H;��H;��H;e�H;Z�H;\�H;��H;:�H;<�H;ǸH;�H;      q�H;��H;N�H;X�H;��H;3�H;�H; �H;+�H;^�H;��H;��H;��H;��H;Z�H;�H;��H;��H;��H;��H;��H;X�H;��H;T�H;��H;��H;�H;B�H;d�H;}�H;��H;��H;v�H;y�H;��H;��H;h�H;��H;��H;y�H;t�H;��H;��H;|�H;e�H;B�H;�H;��H;��H;Q�H;��H;W�H;��H;��H;��H;��H;��H;�H;X�H;��H;��H;��H;��H;^�H;-�H; �H;�H;6�H;��H;[�H;O�H;��H;      ��H;��H;.�H;��H;��H;��H;8�H;��H;*�H;��H;�H;��H;�H;m�H;��H;��H;��H;��H;��H;J�H;��H;2�H;��H;��H;�H;Y�H;e�H;r�H;��H;|�H;��H;��H;x�H;r�H;��H;j�H;`�H;j�H;��H;r�H;u�H;��H;��H;|�H;��H;r�H;e�H;W�H;
�H;��H;��H;0�H;��H;I�H;��H;��H;��H;��H;��H;n�H;�H;��H;�H;��H;,�H;��H;8�H;��H;��H;��H;/�H;��H;      ��H;��H;,�H;��H;C�H;��H;��H;��H;��H;��H;�H;:�H;1�H;0�H;�H;��H;��H;1�H;��H;%�H;��H;��H;�H;Y�H;a�H;n�H;��H;��H;��H;��H;v�H;{�H;|�H;{�H;Y�H;Y�H;��H;Y�H;Y�H;{�H;y�H;|�H;v�H;��H;��H;��H;��H;m�H;c�H;W�H;�H;��H;��H;%�H;��H;4�H;��H;��H;�H;0�H;/�H;8�H;�H;��H;��H;��H;��H;��H;;�H;��H;,�H;��H;      ��H;��H;��H;�H;��H;$�H;��H;��H;Q�H;�H;��H;��H;@�H; �H;��H;M�H;��H;2�H;��H;��H;#�H;W�H;q�H;��H;��H;��H;��H;��H;��H;��H;x�H;t�H;v�H;d�H;U�H;Z�H;^�H;Z�H;U�H;d�H;u�H;v�H;x�H;��H;��H;��H;��H;��H;��H;��H;o�H;V�H;"�H;��H;��H;3�H;��H;M�H;��H; �H;@�H;��H;��H;	�H;T�H;��H;��H;(�H;��H;	�H;��H;��H;      ��H;��H;��H;)�H;��H;��H;X�H;��H;k�H;��H;��H;0�H;��H;J�H;��H;)�H;~�H;��H;6�H;k�H;��H;��H;��H;��H;��H;��H;��H;��H;��H;��H;��H;��H;W�H;U�H;`�H;U�H;9�H;U�H;`�H;V�H;U�H;��H;��H;��H;��H;��H;��H;��H;��H;��H;��H;��H;��H;k�H;6�H;��H;|�H;)�H;��H;J�H;��H;0�H;��H;��H;k�H;��H;X�H;��H;��H;*�H;��H;��H;      2�H;X�H;��H;��H;��H;7�H;��H;,�H;��H;#�H;��H;�H;��H;��H;c�H;��H;	�H;4�H;m�H;��H;��H;��H;��H;��H;��H;��H;��H;��H;��H;��H;��H;n�H;W�H;^�H;V�H;R�H;A�H;R�H;V�H;\�H;V�H;q�H;��H;��H;��H;��H;��H;��H;��H;��H;��H;��H;��H;��H;m�H;6�H;�H;��H;b�H;��H;��H;�H;��H;&�H;��H;*�H;��H;<�H;��H;��H;��H;P�H;      ��H;��H;�H;G�H;��H;��H;L�H;��H;�H;}�H;��H;^�H;��H;<�H;��H;��H;/�H;V�H;��H;��H;��H;��H;��H;��H;��H;��H;��H;��H;��H;��H;k�H;g�H;��H;a�H;9�H;B�H;=�H;B�H;9�H;a�H;��H;h�H;k�H;��H;��H;��H;��H;��H;��H;��H;��H;��H;��H;��H;��H;W�H;-�H;��H;��H;<�H;��H;^�H;��H;��H;�H;��H;L�H;��H;��H;G�H;�H;��H;      2�H;X�H;��H;��H;��H;7�H;��H;,�H;��H;#�H;��H;�H;��H;��H;b�H;��H;	�H;4�H;m�H;��H;��H;��H;��H;��H;��H;��H;��H;��H;��H;��H;��H;n�H;W�H;^�H;V�H;R�H;A�H;R�H;V�H;\�H;V�H;q�H;��H;��H;��H;��H;��H;��H;��H;��H;��H;��H;��H;��H;m�H;6�H;�H;��H;c�H;��H;��H;�H;��H;%�H;��H;*�H;��H;<�H;��H;��H;��H;N�H;      ��H;��H;��H;*�H;��H;��H;W�H;��H;k�H;��H;��H;0�H;��H;J�H;��H;)�H;~�H;��H;6�H;k�H;��H;��H;��H;��H;��H;��H;��H;��H;��H;��H;��H;��H;W�H;V�H;`�H;U�H;9�H;U�H;`�H;U�H;U�H;��H;��H;��H;��H;��H;��H;��H;��H;��H;��H;��H;��H;k�H;6�H;��H;|�H;)�H;��H;J�H;��H;0�H;��H;��H;k�H;��H;X�H;��H;��H;*�H;��H;��H;      ��H;��H;��H;	�H;��H;$�H;��H;��H;Q�H;	�H;��H;��H;@�H; �H;��H;M�H;��H;2�H;��H;��H;%�H;V�H;o�H;��H;��H;��H;��H;��H;��H;��H;x�H;t�H;v�H;d�H;U�H;Z�H;^�H;Z�H;U�H;d�H;u�H;v�H;x�H;��H;��H;��H;��H;��H;��H;��H;q�H;W�H;#�H;��H;��H;3�H;��H;M�H;��H; �H;@�H;��H;��H;�H;S�H;��H;��H;(�H;��H;�H;��H;��H;      ��H;��H;-�H;��H;B�H;��H;��H;��H;��H;��H;�H;8�H;/�H;0�H;�H;��H;��H;1�H;��H;$�H;��H;��H;�H;W�H;c�H;n�H;��H;��H;��H;��H;v�H;{�H;{�H;y�H;Y�H;Y�H;��H;W�H;Y�H;y�H;y�H;}�H;v�H;��H;��H;��H;��H;m�H;a�H;W�H;�H;��H;��H;'�H;��H;2�H;��H;��H;�H;0�H;/�H;:�H;�H;��H;��H;��H;��H;��H;;�H;��H;)�H;��H;      ��H;��H;/�H;��H;��H;��H;<�H;��H;*�H;��H;�H;��H;�H;m�H;��H;��H;��H;��H;��H;I�H;��H;0�H;��H;��H;
�H;Y�H;e�H;r�H;��H;{�H;��H;��H;u�H;r�H;��H;j�H;`�H;j�H;��H;r�H;u�H;��H;��H;}�H;��H;r�H;e�H;W�H;�H;��H;��H;2�H;��H;J�H;��H;��H;��H;��H;��H;m�H;�H;��H;�H;��H;,�H;��H;;�H;��H;��H;��H;/�H;��H;      q�H;��H;N�H;[�H;��H;3�H;�H; �H;-�H;]�H;��H;��H;��H;��H;X�H;�H;��H;��H;��H;��H;��H;W�H;��H;T�H;��H;��H;�H;B�H;c�H;}�H;��H;��H;u�H;y�H;��H;��H;h�H;��H;��H;y�H;t�H;��H;��H;|�H;e�H;B�H;�H;��H;��H;R�H;��H;X�H;��H;��H;��H;��H;��H;�H;Z�H;��H;��H;��H;��H;`�H;-�H;�H;�H;6�H;��H;X�H;N�H;��H;      ��H;�H;ʸH;:�H;:�H;��H;_�H;Z�H;d�H;��H;��H;��H;��H;��H;��H;/�H;U�H;2�H;��H;�H;�H;<�H;�H;��H;%�H;|�H;��H;!�H;E�H;\�H;{�H;y�H;��H;��H;��H;��H;��H;��H;��H;��H;��H;{�H;{�H;Z�H;G�H;!�H;��H;|�H;%�H;��H;�H;>�H;�H;�H;��H;4�H;U�H;2�H;��H;��H;��H;��H;��H;��H;g�H;[�H;_�H;��H;8�H;<�H;ʸH;�H;      C�H;ҡH;^�H;˥H;�H;��H;��H;!�H;��H;R�H;��H;\�H;r�H;]�H;�H;H�H;�H;}�H;��H;��H;^�H;��H;��H;��H;\�H;��H;��H;��H;�H;H�H;d�H;��H;��H;��H;��H;��H;��H;��H;��H;��H;��H;��H;d�H;G�H;�H;��H;��H;��H;[�H;��H;��H;��H;[�H;��H;��H;��H;�H;J�H;�H;]�H;r�H;\�H;��H;T�H;��H;!�H;��H;��H;�H;ƥH;b�H;ϡH;      �lH;WnH;�rH;�yH;r�H;ǋH;�H;ҝH;ťH;�H;��H;(�H;1�H;��H;��H;^�H;n�H;�H;�H;��H;��H;��H;!�H;m�H;u�H;B�H;��H;j�H;��H;"�H;A�H;q�H;��H;��H;��H;��H;��H;��H;��H;��H;��H;r�H;A�H;!�H;��H;k�H;��H;C�H;u�H;n�H;!�H;��H;��H;��H;�H;�H;m�H;`�H;��H;��H;1�H;(�H;��H;	�H;ƥH;ԝH;�H;ƋH;~�H;�yH;�rH;bnH;      6�G;��G;$�G;��G;zH;�0H;�LH;?fH;_|H;j�H;p�H;m�H;v�H;��H;ҿH;C�H;��H;��H;�H;��H;��H;�H;B�H;��H;0�H;`�H;4�H;��H;��H;��H;�H;g�H;��H;��H;��H;��H;��H;��H;��H;��H;��H;h�H;�H;��H;��H;��H;4�H;a�H;,�H;��H;A�H;�H;��H;��H;�H;��H;��H;C�H;ҿH;��H;v�H;m�H;s�H;j�H;`|H;?fH;�LH;�0H;|H;��G;#�G;��G;      SIF;-UF;AwF;6�F;��F;�8G;�G;��G;�	H;�=H;/fH;r�H;ǗH;��H;��H;۹H;��H;��H;j�H;j�H;t�H;��H;��H;��H;��H;/�H;^�H;B�H;��H;~�H;��H;W�H;m�H;��H;��H;��H;��H;��H;��H;��H;k�H;Z�H;��H;|�H;��H;B�H;]�H;0�H;��H;��H;��H;��H;o�H;j�H;j�H;��H;��H;ܹH;��H;��H;ƗH;u�H;/fH;�=H;�	H;��G;��G;�8G;��F;4�F;AwF;UF;      ߣB;!�B;�C;ĐC;�0D;��D;"�E;�IF;��F;:jG;L�G;q$H;�\H;1�H;��H;�H;T�H;ٽH;��H;|�H;�H;��H;2�H;U�H;��H;��H;2�H;y�H;a�H;.�H;��H;	�H;e�H;��H;��H;��H;��H;��H;��H;��H;e�H;�H;��H;.�H;_�H;y�H;0�H;��H;��H;U�H;2�H;��H;�H;}�H;��H;߽H;S�H;�H;��H;1�H;�\H;q$H;K�G;:jG;��F;�IF;"�E;��D;�0D;ĐC;�C;!�B;      4�:;A�:;��;;�<;>;̧?;-JA;��B;2FD;$|E;JwF;�8G;��G;p'H;fH;v�H;i�H;x�H;��H;��H;%�H;S�H;.�H;�H;Q�H;��H;��H;j�H;��H;��H;N�H;��H;R�H;��H;��H;��H;��H;��H;��H;��H;S�H;��H;O�H;��H;��H;j�H;��H;��H;P�H;�H;.�H;S�H;#�H;��H;��H;{�H;g�H;v�H;fH;n'H;��G;�8G;HwF; |E;2FD;��B;,JA;ͧ?;>;��<;��;;2�:;      �*;��*;�,;�d.;�Y1;��4;%,8;��;;`�>;JA;SxC;�*E;
lF;�NG;#�G;EH;%|H;F�H;ȫH;P�H;g�H;p�H;��H;/�H;.�H;��H;C�H;!�H;��H;�H;��H;��H;�H;r�H;��H;��H;��H;��H;��H;r�H;�H;��H;��H;	�H;��H;!�H;A�H;��H;.�H;.�H;��H;p�H;c�H;S�H;ȫH;K�H;'|H;EH;$�G;�NG;lF;�*E;SxC; JA;`�>;��;;',8;��4;�Y1;�d.;�,;��*;      A�
;e�;�;	;Z�;a;�D&;�-;�D3;N�8; I=;��@;͐C;Q|E;��F;�G;h$H;.nH;��H;M�H;�H;��H;m�H;S�H;��H;��H;�H;��H;��H;?�H;W�H;,�H;��H;V�H;��H;��H;��H;��H;��H;V�H;��H;.�H;X�H;<�H;��H;��H;�H;��H;��H;Q�H;k�H;��H;�H;N�H;��H;2nH;h$H;�G;��F;R|E;͐C;��@; I=;M�8;�D3;�-;�D&;a;o�;	;�;`�;      ��:፨:�: ��:��:�P�:�{;)(;��;�~(;�Y1;u8;b�=;A�A;|�D;IF;�cG;�	H;AdH;��H;y�H;�H;f�H;(�H;�H;t�H;��H;��H;Z�H;�H;��H;��H;��H;�H;|�H;��H;��H;��H;|�H;�H;��H;��H;��H;�H;X�H;��H;}�H;u�H;�H;%�H;c�H;�H;w�H;��H;CdH;�	H;�cG;IF;|�D;A�A;e�=;u8;�Y1;�~(;��;)(;�{;�P�:%��:��:�:Ǎ�:      p�R�0�� >7��E^9��:��X:���:���:�P�:��;��;�);�D3;i�:;�!@;�C;\�E;
9G;��G;�`H;��H;K�H;M�H;��H;u�H;h�H;��H;��H;��H;�H;��H;?�H; �H;��H;c�H;��H;��H;��H;c�H;��H;�H;@�H;��H;�H;��H;��H;��H;k�H;v�H;��H;J�H;K�H;��H;�`H;��G;9G;]�E;�C;�!@;i�:;�D3;�);��;��;�P�:���:���:ВX:�:�E^9 >7����      {�)��$�.��
������H�\��N��PS�9H4j:���:*��:��;l� ;�d.;�+8;��>;ZC;��E;�)G;��G;@dH;��H;ȫH;��H;��H;j�H; �H;�H;��H;��H;��H;z�H;��H;��H;4�H;j�H;��H;j�H;4�H;��H;��H;|�H;��H;��H;��H;�H;��H;m�H;��H;��H;īH;��H;@dH;��G;�)G;��E;YC;��>;�+8;�d.;l� ;��;.��:���:P4j:XS�9�N��0�\�������/���$�      Z�ѻ�ͻ1���LG��򿐻v�d�ă$��Iɺ��!��L^9x�r:E��:1;;�;<�*;�Z6;�>;X�B;��E;9G;�	H;.nH;I�H;x�H;ؽH;��H;��H;�H;��H;6�H;��H;��H;4�H;/�H;��H;:�H;]�H;:�H;��H;/�H;2�H;��H;��H;4�H;}�H;	�H;��H;��H;ؽH;t�H;F�H;/nH;�	H;9G;��E;Y�B;�>;�Z6;=�*;;�;1;E��:x�r:�L^9��!��Iɺă$�q�d��LG��0����ͻ      ��I�2�E��(;��O*����<��"GĻȿ���s@�.IҺP~��:V�: Q�:�;�~(;+�5;�>;\C;_�E;�cG;i$H;(|H;i�H;O�H;��H;��H;m�H;�H;S�H;��H;��H;��H;��H;t�H;�H;&�H; �H;t�H;��H;��H;��H;��H;Q�H;	�H;m�H;��H;��H;P�H;f�H;#|H;i$H;�cG;a�E;]C;�>;+�5;�~(;�;�P�:V�:�:X~�4IҺ�s@�ȿ��"GĻ�<�����O*��(;�5�E�      3p��hx��ע��R��+��x�`��7�A��.�ѻ�,��d�$�ǅ���09V�:��:�;�~(;�Z6;��>;��C;IF;�G;EH;w�H;�H;۹H;A�H;\�H;G�H;,�H;�H;��H;��H;B�H;�H;��H;��H;��H;�H;C�H;��H;��H;�H;,�H;C�H;\�H;?�H;ܹH;�H;t�H;EH;�G;IF;��C;��>;�Z6;�~(;�;��:X�:��09ǅ�d�$��,��.�ѻA���7�v�`�+���R��ע�ix��      4]� �0#�������ټ�ɺ������
v��(;�Ш�D^���5R�&��� }6����:��:�;9�*;�+8;�!@;|�D;��F;$�G;fH;��H;��H;пH;��H;�H;��H;T�H;��H;��H;��H;��H;[�H;��H;[�H;��H;��H;��H;��H;T�H;��H;�H;��H;ϿH;��H;��H;�eH;�G;��F;|�D;�!@;�+8;>�*;�;��:���: }6�&����5R�D^��Ш��(;��
v������ɺ���ټ����0#� �      �_�&\�&<Q�g@�� +��5�����a�ļ|�d�`����Iͻk��Hɺ {6�X�:Q�:=�;�d.;m�:;?�A;O|E;�NG;n'H;+�H;��H;��H;��H;Z�H;{�H;��H;d�H;+�H;��H;@�H;��H;2�H;��H;@�H;��H;(�H;e�H;��H;{�H;Z�H;��H;��H;��H;-�H;k'H;�NG;O|E;B�A;m�:;�d.;?�; Q�:\�: |6��Hɺk�Hͻ���d�`�|�`�ļ�����5�� +�g@�&<Q�&\�      A���R��(ڟ�����"C���_�0:������0p���vz��O*��4ֻk� �����09\�:1;m� ;�D3;b�=;̐C;lF;��G;�\H;ǗH;y�H;0�H;o�H;��H;��H;�H;+�H;;�H;��H;��H;��H;��H;��H;;�H;*�H;�H;��H;��H;m�H;0�H;v�H;ɗH;�\H;��G;	lF;̐C;e�=;�D3;m� ;1;Z�:��09 ���k��4ֻ�O*��vz�1p���輨��0:��_�"C������(ڟ��R��      �` ��.�����ïڽ�b��zr��^��\�~ +�� ��ɺ�C��O*�Iͻ�5R�ǅ��:I��:��;�);u8;��@;�*E;�8G;l$H;q�H;k�H;"�H;V�H;��H;��H;��H;0�H;��H;"�H;�H;Q�H;�H;"�H;��H;-�H;��H;��H;��H;U�H;"�H;h�H;q�H;o$H;�8G;�*E;��@;u8;�);��;K��:��:ǅ��5R�Iͻ�O*�C��ɺ�� �~ +�\�^��zr���b��ïڽ��.��      �-=�C�9��k/�3��������Ľ�!��nys�G�6�(#��ɺ��vz����D^��g�$�X~�p�r:(��: �;�Y1;I=;SxC;HwF;H�G;/fH;p�H;��H;��H;��H;��H;�H;�H;��H;��H;��H;��H;��H;��H;��H;
�H;�H;��H;��H;��H;��H;m�H;/fH;L�G;DwF;QxC;I=;�Y1;��;(��:x�r:h~�g�$�D^������vz��ɺ�(#�G�6�nys��!����Ľ����3���k/�D�9�      �(��Hl���.}�<ce�~PH���(�~
���ڽ�R���{�G�6�� �1p��f�`�Ш��,��2IҺ�L^9���:��;�~(;K�8;JA;"|E;:jG;�=H;i�H;�H;Q�H;��H;W�H;��H;��H;�H;��H; �H;z�H; �H;��H;�H;��H;��H;V�H;��H;N�H;�H;g�H;�=H;=jG; |E;JA;K�8;�~(;��;���:�L^96IҺ�,��Ш�f�`�1p��� �G�6��{��R����ڽ~
���(�~PH�<ce��.}�Hl��      �iþXD��:o�����������i��-=�kt����R��nys�~ +���}񗼘(;�0�ѻ�s@���!�D4j:�P�:��;�D3;]�>;0FD;��F;�	H;\|H;��H;��H;Y�H; �H;#�H;��H;J�H;b�H;��H;�H;��H;b�H;L�H;��H;#�H;!�H;Y�H;��H;��H;Y|H;�	H;��F;.FD;\�>;�D3;��;�P�:D4j:��!��s@�0�ѻ�(;�}���~ +�nys��R����kt��-=��i���������:o��XD��      ���
�����'�޾YD���A���.}�,�D�kt���ڽ�!��\����a�ļ�
v�A��ɿ���IɺXS�9���:&(;�-;��;;��B;�IF;��G;<fH;ȝH;�H;P�H;��H;��H;��H;��H;��H;�H;��H;!�H;��H;��H;��H;��H;��H;P�H;�H;ʝH;:fH;��G;�IF;��B;��;;�-;)(;���:XS�9�Iɺʿ��A���
v�a�ļ���\��!����ڽkt�,�D��.}��A��YD��'�޾�����
�      ��7�ҕ3��f'�+��\���о�����.}��-=�~
���Ľ^��0:����������7�%GĻă$��N�����:�{;�D&;,8;*JA;�E;�G;�LH;�H;��H;U�H;�H;4�H;��H;��H;M�H;��H;E�H;��H;M�H;��H;��H;4�H;�H;T�H;��H;�H;�LH;�G;"�E;(JA;,8;�D&;�{;���:�N��$�&GĻ�7���������0:�^����Ľ~
��-=��.}������о�\��+��f'�ҕ3�      \o�bXi��"Y���@�M�#��
��о�A���i���(����zr���_��5��ɺ�x�`��<��j�d�T�\�ȒX:�P�:�`;��4;ȧ?;��D;�8G;�0H;ċH;��H;��H;3�H;��H;��H;(�H;��H;<�H;��H;=�H;��H;(�H;��H;��H;3�H;��H;��H;ċH;�0H;�8G;��D;Ƨ?;��4;�`;�P�:ȒX:L�\�i�d��<��x�`��ɺ��5��_�zr�������(��i��A���о�
�M�#���@��"Y�bXi�      1����������\o��!J�M�#��\��YD������~PH�����b��"C��� +���ټ,����򿐻����:#��:W�;�Y1;>;�0D;��F;uH;o�H;�H;-�H;��H;��H;6�H;��H;|�H;��H;��H;��H;z�H;��H;5�H;��H;��H;*�H;��H;o�H;wH;��F;�0D;>;�Y1;W�;+��:�:���񿐻��,����ټ� +�"C���b�����~PH�����YD���\��M�#��!J�\o��������      @^������m���\o���@�+�'�޾����<ce�3��ïڽ����g@������R���O*�NG������E^9$��:;�d.;�<;��C;7�F;��G;�yH;ƥH;:�H;O�H;��H;��H;�H;�H;��H;C�H;��H;�H;�H;��H;��H;O�H;7�H;ťH;�yH;��G;7�F;��C;�<;�d.;;*��:�E^9���MG���O*��R������g@�����ïڽ3��<ce�����'�޾+���@�\o�m�������      �aǿ�¿����������"Y��f'�����:o���.}��k/����(ڟ�'<Q�1#�ע��(;�4���8�� E7���:��;�,;��;;�C;CwF;#�G;�rH;\�H;¸H;A�H;&�H;"�H;��H;��H;x�H;��H;x�H;��H;��H; �H;'�H;A�H;��H;Y�H;�rH;#�G;AwF;�C;��;;�,;��;��: E7�8��3����(;�ע�1#�'<Q�(ڟ�����k/��.}�:o�������f'��"Y�����������¿      6�ֿFpѿ�¿������bXi�ҕ3��
�XD��Hl��D�9��.���R��'\� �ix��5�E��ͻ�$�P  �Ǎ�:H�;��*;5�:;�B;#UF;��G;UnH;ѡH;޷H;��H;��H;��H;��H;��H;J�H;��H;J�H;��H;��H;��H;��H;��H;۷H;ΡH;UnH;��G;"UF;�B;2�:;��*;H�;ˍ�:`  ��$��ͻ5�E�ix�� �'\��R���.��D�9�Hl��XD���
�ҕ3�bXi��������¿Fpѿ      �?��~h��?v��� ��:�X��O/�1y�D�;㰖��+X����ѽ����en;�d�������B(�䚩�d���e9�:�;�Y.;R�<;�WC;%[F;�G;*0H;sjH;V�H;u�H;��H;Q�H;��H;��H;��H;��H;��H;��H;��H;O�H;��H;u�H;T�H;pjH;*0H;�G;$[F;�WC;O�<;�Y.;�;�:Рe9d��䚩��B(�����d��en;������ѽ���+X�㰖�D�;1y��O/�:�X�� ��?v��~h��      h��1���c�����y�YvS�sM+��v�9ɾ�����T�#]�\ν����~\8�����x��	%�Y������(�9Y-�:p�;��.;�<;�nC;�dF;�G;�1H; kH;ǌH;ӤH;�H;��H;��H;��H;��H;��H;��H;��H;��H;��H;�H;ӤH;ÌH;kH;�1H;�G;�dF;�nC;�<;��.;p�;]-�:�9���X���
%��x�����~\8�����\ν#]��T�����9ɾ�v�sM+�YvS���y�c���1���      ?v��c���X ��c�h�9E�Z��m���㼾����nH�ֈ�~�ý�Ȅ��s/��o��#�����.J��2к8
�9Dg�:�l;S0;!]=;��C;�F;|�G;F6H;]mH;H�H;ѥH;��H;(�H;n�H;��H;1�H;�H;1�H;��H;n�H;&�H;��H;ѥH;C�H;ZmH;F6H;|�G;�F;��C;]=;V0;�l;Dg�: 
�92к.J������#���o��s/��Ȅ�~�ýֈ��nH����㼾m���Z��9E�c�h�X ��c���      � ����y�c�h��N��O/����E�߾B���*|��6�s}�䳽pSt�A�!�wrμLF{��_� Y��֓���:��:�Z;�2;�O>;�D;j�F;��G;B=H;�pH;��H;x�H;�H;�H;�H;��H;��H;��H;��H;��H;�H;�H;�H;v�H;��H;�pH;B=H;��G;g�F;�D;�O>;�2;�Z; ��:�:ؓ�� Y���_�LF{�wrμA�!�pSt�䳽s}��6��*|�B��E�߾����O/��N�c�h���y�      :�X�YvS�9E��O/��S�KW����������PS\��� ���>����Y���׃����]�����2�b���Y���Y:��:r`;b�4;�?;a�D;
�F;�G;/FH;}uH;�H;��H;��H;?�H;��H;O�H;D�H;'�H;D�H;N�H;��H;=�H;��H;��H;ޓH;zuH;/FH;!�G;�F;`�D;�?;f�4;r`;��:��Y:��Y�2�b�������]�׃�����Y�>����彔� �PS\���������KW���S��O/�9E�YvS�      �O/�sM+�Z�����KW��9ɾD���Mw�� :�l��|�ýM��bn;�f���zv���E<��˻��-�(���y�:�^;�%;��7;��@;<5E;�"G; �G;cPH;3{H;�H;��H;��H;��H;$�H;>�H;�H;��H;�H;>�H;"�H;��H;��H;��H;ޗH;/{H;cPH;�G;�"G;:5E;}�@;��7;�%;�^;�y�:(����-��˻�E<�zv��f���bn;�M��|�ýl��� :��Mw�D��9ɾKW�����Z��sM+�      1y��v�m���E�߾����D��A����nH���Hὡu����d�4O�qrμO"�����
	�����pr89�;�:c�;�+;}|:;�7B;�E;5bG;�H;[H;��H;L�H;ȯH;%�H;r�H;t�H;7�H;�H;��H;�H;7�H;r�H;r�H;'�H;ȯH;J�H;��H;[H;�H;4bG;�E;�7B;||:;�+;d�;�;�:pr89���
	�����O"��qrμ4O���d��u��H����nH�A���D������E�߾m����v�      D�;9ɾ㼾B�������Mw��nH�����Z�䳽Ε��w\8�w#������^N�V���b�Ix�X5:��:6�;��0;E]=;T�C;�[F;�G;�)H;fH;��H;F�H;m�H;��H;F�H;��H;\�H;��H;��H;��H;\�H;��H;D�H;��H;k�H;F�H;��H;fH;�)H;�G;�[F;P�C;D]=;��0;7�;��:P5:Ix��b�V��^N�����w#��v\8�Ε��䳽�Z񽳯��nH��Mw�����B��㼾9ɾ      㰖��������*|�PS\�� :����Z�p$�������K�z���Oļ����������A&����V/�:�^;��#;�G6;a�?;�D;t�F;��G;#@H;�pH;�H;��H;>�H;}�H;W�H;��H;��H;�H;��H;�H;��H;��H;W�H;�H;>�H;��H;�H;�pH; @H;��G;p�F;�D;`�?;�G6;��#;�^;V/�:���B&������������Oļz���K�����p$���Z���� :�PS\��*|�������      �+X��T��nH��6��� �l��H�䳽�����mR����ټ�����E<��?ݻ@d\����� !:�d�:��;6�,;��:;�7B;��E;�LG;aH;SH;�{H;��H;�H;@�H;k�H;~�H;<�H;��H; �H;��H; �H;��H;;�H;|�H;p�H;@�H;�H;��H;�{H;~SH;`H;�LG;��E;7B;��:;6�,;��;�d�:!:����Ad\��?ݻ�E<�����ټ����mR�����䳽H�l���� ��6��nH��T�      ��#]�ֈ�s}���|�ý�u��Ε���K�����o�ov���&R�%��\^����� x>���:nB;Z";~�4;��>;gD;��F;�G;�)H;�dH;��H;>�H;��H;W�H;[�H;��H;��H;N�H;;�H;��H;:�H;N�H;��H;��H;^�H;V�H;��H;;�H;��H;�dH;�)H;�G;��F;eD;��>;z�4;W";nB;
��: |>����\^��%���&R�ov���o�����K�Ε���u��|�ý��s}�ֈ�#]�      �ѽ\ν}�ý䳽>���M����d�v\8�z��ټov����Y��_����B���[���Y:m��:^m;�r-;!�:;��A;XoE;�"G;y�G;�GH;�sH;�H;��H;�H;W�H;F�H;��H;��H;��H;T�H;�H;T�H;��H;��H;��H;H�H;V�H;�H;��H;�H;�sH;�GH;v�G;�"G;ToE;��A;!�:;�r-;\m;s��:��Y:�[�C��
����_���Y�ov��ټz��v\8���d� M��>���䳽}�ý\ν      ���������Ȅ�pSt��Y�bn;�4O�w#���Oļ�����&R��_������N3�؅Y� 4:"�:ޯ;�?&;�G6;�X?;�D;QxF;ޚG;]!H;�^H;��H;�H;��H;k�H;2�H;)�H;��H;=�H;�H;~�H;<�H;~�H;�H;<�H;��H;*�H;2�H;k�H;��H;�H;��H;�^H;X!H;ٚG;MxF;�D;�X?;�G6;�?&;߯;�:�3:܅Y��N3������_��&R������Oļw#��4O�an;��Y�pSt��Ȅ�����      en;�}\8��s/�@�!���e���prμ��������E<�$��
����N3�PHx���9�:�^;a ;D2;��<;�B;˲E;W5G;+�G;ZFH;�qH;ʎH;s�H;�H;v�H;��H;��H;)�H;��H;G�H;��H;6�H;��H;G�H;��H;)�H;��H;��H;w�H;ߴH;r�H;ȎH;�qH;XFH;(�G;S5G;˲E;�B;��<;B2;b ;�^;�:��9LHx��N3�
���$���E<��������prμe�����@�!��s/�~\8�      c������o�wrμ׃��yv��O"��^N�����?ݻ\^��E����Y���9��:��:��;b�.;�|:;?A;��D;M�F;׶G;*H;CaH;@�H;��H;�H;d�H;F�H;d�H;��H;$�H;E�H;��H;��H;�H;��H;��H;E�H;$�H;��H;c�H;D�H;`�H;�H;��H;@�H;@aH;*H;ѶG;K�F;��D;?A;�|:;b�.;��;��:��:��9��Y�E��\^���?ݻ���^N�O"��yv��׃��wrμ�o����      �����x���#��JF{���]��E<����W�뻮���>d\���뺬[� 4:�:���:�[;z�,;��8;:!@;�0D;�[F;C{G;H;lPH;?vH;�H;i�H;&�H;W�H;��H;��H;�H;�H;��H;��H;��H;��H;��H;��H;��H;�H;�H;��H;��H;Q�H;&�H;f�H;�H;<vH;ePH;H;C{G;�[F;�0D;9!@;��8;z�,;�[;���:�: 4:�[����=d\�����X�뻩���E<���]�JF{��#���x��      �B(�%�����_������˻	���b�A&����� p>���Y: �:�^;��;x�,;%`8;v�?;�C;�F;GG;n�G;@H;OkH;)�H;/�H;�H;~�H;��H;��H;��H;D�H;��H;	�H;��H;��H;��H;��H;��H;
�H;��H;F�H;��H;��H;��H;}�H;�H;/�H;'�H;KkH;@H;n�G;GG;�F;�C;x�?;&`8;x�,;��;�^; �:��Y: |>�����?&��b�	���˻�����_����	%�      嚩�X���+J���X��4�b��-����Ix���� !:��:k��:ޯ;_ ;`�.;��8;v�?;�C;��E;[#G;�G;2H;bH;p�H;��H;��H;ԷH;
�H;��H;C�H;a�H;c�H;�H;B�H;��H;d�H;��H;d�H;��H;A�H;�H;c�H;a�H;A�H;��H;�H;ҷH;��H;��H;l�H;bH;2H;
�G;\#G;��E;�C;s�?;��8;`�.;b ;ܯ;k��:��:!:���(Ix�����-�.�b��X��+J��]���      P����� кғ����Y����r89P5:Z/�:�d�:nB;^m;�?&;D2;�|:;6!@;�C;��E;�G;��G;~(H;![H;�zH;f�H;�H;˳H;��H;��H;��H;��H;��H;$�H;y�H;X�H;w�H;(�H;��H;(�H;w�H;X�H;x�H;&�H;��H;��H;��H;��H;��H;˳H;�H;b�H;�zH;![H;z(H; �G;�G;��E;߳C;6!@;�|:;D2;�?&;`m;nB;�d�:`/�:D5:�r89�����Y�ғ�� к���       �e9��9H
�9�:��Y:�y�:�;�:��:�^;��;W";�r-;�G6;��<;?A;�0D;�F;X#G;��G;%H;�WH;�vH;��H;l�H;r�H;��H;:�H;��H;��H;e�H; �H;��H;��H;U�H;;�H;��H;%�H;��H;9�H;U�H;��H;��H; �H;b�H;��H;��H;6�H;��H;o�H;f�H;��H;�vH;~WH;%H;��G;Y#G;�F;�0D;?A;��<;�G6;�r-;W";��;�^;��:�;�:�y�:��Y:�:@
�9h�9      �:}-�:Ng�:��:��:�^;g�;6�;��#;8�,;|�4;�:;�X?;�B;��D;�[F;GG;�G;�(H;�WH;�uH;��H;@�H;'�H;O�H;&�H;��H;�H;�H;��H;��H;�H;��H;�H;��H;��H;��H;��H;��H;�H;��H;�H;��H;��H;�H;�H;��H;%�H;M�H;!�H;=�H;��H;�uH;�WH;~(H;�G;GG;�[F;��D;�B;�X?;�:;z�4;6�,;��#;4�;g�;�^;��:��:Ng�:]-�:      ;��; m;�Z;s`;�%;�+;��0;�G6;��:;��>;��A;�D;˲E;N�F;B{G;n�G;2H;#[H;�vH;��H;z�H;�H;��H;��H;��H;��H;��H;��H;�H;m�H;h�H;��H;��H;��H;��H;�H;��H;��H;��H;��H;f�H;k�H;�H;��H;��H;��H;��H;��H;�H;�H;x�H;��H;�vH;![H;2H;l�G;A{G;N�F;̲E;�D;��A;��>;��:;�G6;��0;�+;�%;�`;�Z; m;��;      �Y.;��.;T0;�2;^�4;��7;�|:;D]=;d�?;�7B;iD;XoE;PxF;W5G;ֶG;H;@H;bH;�zH;��H;@�H;�H;w�H;��H;��H;��H;��H;$�H;M�H;��H;��H;��H;��H;v�H;�H;P�H;x�H;N�H;�H;v�H;��H;��H;��H;��H;J�H;$�H;��H;��H;��H;��H;u�H;�H;:�H;��H;�zH;bH;@H;H;ֶG;W5G;PxF;YoE;gD;�7B;d�?;D]=;�|:;��7;h�4;�2;V0;��.;      d�<;&�<;(]=;�O>;��?;~�@;�7B;R�C;�D;��E;��F;�"G;ٚG;+�G;*H;iPH;MkH;s�H;f�H;j�H;"�H;��H;��H;c�H;a�H;h�H;y�H;��H;R�H;l�H;+�H;@�H;<�H;�H;s�H;��H;��H;��H;t�H;�H;8�H;@�H;)�H;h�H;N�H;��H;w�H;h�H;c�H;a�H;��H;��H;�H;i�H;d�H;s�H;LkH;iPH;*H;+�G;ٚG;�"G;��F;��E;�D;R�C;�7B;��@;��?;�O>;)]=;�<;      �WC;	oC;�C;�D;c�D;?5E;�E;�[F;t�F;�LG;�G;|�G;[!H;_FH;FaH;AvH;.�H;��H;�H;w�H;R�H;��H;��H;h�H;&�H;8�H;r�H;��H;�H;��H;�H;��H;��H;h�H;��H;�H;�H;�H;��H;f�H;��H;��H;
�H;��H;�H;��H;o�H;8�H;'�H;g�H;��H;��H;O�H;y�H;�H;��H;,�H;@vH;FaH;]FH;Z!H;|�G;�G;�LG;v�F;�[F;�E;?5E;d�D;�D;�C;
oC;      2[F;�dF;�F;g�F;�F;�"G;7bG;�G;��G;bH;�)H;�GH;�^H;�qH;=�H;�H;/�H;��H;ɳH;��H;#�H;��H;��H;g�H;1�H;Z�H;��H;��H;��H;��H;��H;��H;W�H;��H;�H;F�H;F�H;F�H;�H;��H;T�H;��H;��H;��H;��H;��H;��H;\�H;4�H;e�H;��H;��H;�H;��H;ȳH;��H;,�H;�H;=�H;�qH;�^H;�GH;�)H;aH;��G;�G;7bG;�"G;�F;i�F;�F;�dF;      �G;��G;|�G;��G;#�G;#�G;�H;*H;$@H;�SH;�dH;�sH;��H;ʎH;��H;j�H;�H;ӷH;��H;=�H;��H;��H;��H;|�H;k�H;��H;��H;q�H;��H;��H;��H;-�H;��H;�H;6�H;i�H;��H;i�H;5�H;�H;��H;-�H;��H;��H;��H;q�H;��H;��H;n�H;z�H;��H;��H;��H;=�H;��H;ӷH;�H;h�H;��H;ʎH;��H;�sH;�dH;SH;'@H; *H;�H;"�G;)�G;��G;}�G;��G;      "0H;�1H;O6H;@=H;0FH;fPH;[H;fH;�pH;�{H;��H;�H;�H;w�H;�H;(�H;~�H;�H;��H;��H;�H;��H;&�H;��H;��H;��H;p�H;��H;��H;��H;2�H;��H;��H;C�H;u�H;��H;z�H;��H;u�H;A�H;��H;��H;2�H;��H;��H;��H;p�H;��H;��H;��H;$�H;��H;�H;��H;��H;�H;}�H;(�H;�H;v�H;�H;�H;��H;�{H;�pH;fH;[H;fPH;:FH;>=H;O6H;�1H;      �jH;#kH;ZmH;�pH;}uH;2{H;��H;��H;�H;��H;>�H;��H;��H;�H;e�H;X�H;��H;��H;��H;��H;
�H;��H;J�H;U�H;�H;��H;��H;��H;��H; �H;��H;��H;(�H;f�H;��H;��H;��H;��H;��H;f�H;%�H;��H;��H;�H;��H;��H;��H;��H;�H;T�H;I�H;��H;�H;��H;��H;��H;��H;X�H;d�H;�H;��H;��H;=�H;��H;�H;��H;��H;5{H;�uH;�pH;[mH;kH;      a�H;͌H;Q�H;��H;�H;�H;T�H;N�H;��H;�H;��H;!�H;r�H;�H;J�H;��H;��H;?�H;��H;i�H;��H;�H;��H;l�H;��H;��H;��H;��H;�H;}�H;��H;/�H;d�H;��H;��H;��H;��H;��H;��H;��H;b�H;0�H;��H;{�H;�H;��H;��H;��H;��H;k�H;��H;�H;��H;h�H;��H;@�H;��H;��H;J�H;~�H;r�H;!�H;��H;�H;��H;P�H;T�H;�H;�H;��H;N�H;ʌH;      y�H;�H;ޥH;��H;ͩH;��H;ӯH;v�H;H�H;H�H;`�H;c�H;9�H;��H;i�H;��H;��H;a�H;��H;�H;��H;n�H;��H;/�H;�H;��H;��H;4�H;��H;��H;)�H;]�H;��H;��H;��H;��H;��H;��H;��H;��H;��H;]�H;)�H;��H;��H;4�H;��H;��H;�H;.�H;��H;m�H;��H;�H;��H;a�H;��H;��H;i�H;��H;9�H;a�H;^�H;H�H;H�H;v�H;ӯH;��H;ʩH;��H;ߥH;�H;      ǵH;�H;��H;�H;��H;��H;+�H;��H;��H;p�H;c�H;O�H;-�H;��H;��H;�H;M�H;e�H;+�H;��H;�H;l�H;��H;D�H;��H;��H;*�H;��H;��H;0�H;Y�H;w�H;��H;��H;��H;��H;��H;��H;��H;��H;��H;w�H;Y�H;2�H;��H;��H;*�H;��H;��H;B�H;��H;j�H;�H;��H;*�H;e�H;M�H;�H;��H;��H;-�H;P�H;c�H;p�H;��H;��H;)�H;��H;��H;�H;öH;�H;      X�H;��H;2�H;�H;L�H;��H;w�H;Q�H;a�H;��H;��H;��H;�H;0�H;*�H;�H;��H;�H;}�H;��H;��H;��H;��H;B�H;��H;W�H;��H;��H;+�H;k�H;��H;��H;��H;��H;��H;��H;��H;��H;��H;��H;��H;��H;��H;k�H;,�H;��H;��H;U�H;��H;?�H;��H;��H;��H;��H;|�H;�H;��H;�H;(�H;0�H; �H;��H;��H;��H;a�H;O�H;w�H;��H;C�H;�H;2�H;��H;      ��H;�H;k�H;�H; �H;!�H;|�H;�H;��H;?�H;��H;��H;@�H;��H;L�H;��H;�H;C�H;^�H;\�H;"�H;��H;s�H;�H;_�H;��H;�H;@�H;f�H;��H;��H;��H;��H;��H;��H;��H;��H;��H;��H;��H;��H;��H;��H;��H;g�H;@�H;�H;��H;a�H;�H;r�H;��H;!�H;\�H;\�H;E�H;�H;��H;J�H;��H;@�H;��H;��H;?�H;��H;�H;|�H;%�H;��H;�H;k�H;�H;      ��H;��H;�H;��H;m�H;:�H;B�H;j�H;��H;��H;U�H;��H;�H;N�H;��H;��H;��H;��H;z�H;B�H; �H;��H;�H;w�H;��H;�H;3�H;u�H;��H;��H;��H;��H;��H;��H;��H;��H;��H;��H;��H;��H;��H;��H;��H;��H;��H;u�H;0�H;�H;��H;t�H;�H;��H;��H;B�H;z�H;��H;��H;��H;��H;N�H;�H;��H;T�H;��H;��H;i�H;B�H;>�H;b�H;��H;�H;��H;      ��H;�H;<�H;��H;W�H;�H;�H;�H;�H;!�H;D�H;`�H;��H;��H;��H;��H;��H;b�H;,�H;��H;��H;��H;M�H;��H;�H;C�H;g�H;��H;��H;��H;��H;��H;��H;��H;��H;��H;��H;��H;��H;��H;��H;��H;��H;��H;��H;��H;f�H;A�H;�H;��H;M�H;��H;��H;��H;,�H;c�H;��H;��H;��H;��H;��H;`�H;B�H;$�H;�H;�H;�H;�H;L�H;��H;<�H;��H;      ��H;��H;!�H;��H;:�H;��H;��H;��H;��H;��H;�H;$�H;A�H;@�H;�H;��H;��H;��H;��H;*�H;��H;�H;t�H;��H;��H;C�H;��H;~�H;��H;��H;��H;��H;��H;��H;��H;��H;��H;��H;��H;��H;��H;��H;��H;��H;��H;~�H;��H;D�H;��H;��H;t�H;�H;��H;,�H;��H;��H;��H;��H;�H;@�H;A�H;$�H;�H;��H;��H;��H;��H;��H;.�H;��H; �H;��H;      ��H;�H;<�H;��H;X�H;�H;�H;�H;�H;!�H;D�H;`�H;��H;��H;��H;��H;��H;b�H;,�H;��H;��H;��H;M�H;��H;�H;C�H;g�H;��H;��H;��H;��H;��H;��H;��H;��H;��H;��H;��H;��H;��H;��H;��H;��H;��H;��H;��H;f�H;C�H;�H;��H;M�H;��H;��H;��H;,�H;c�H;��H;��H;��H;��H;��H;`�H;D�H;"�H;�H;�H;�H;�H;L�H;��H;:�H;��H;      ��H;��H;�H;��H;m�H;:�H;B�H;l�H;��H;��H;T�H;��H;�H;N�H;��H;��H;��H;��H;z�H;B�H; �H;��H;�H;v�H;��H;�H;2�H;u�H;��H;��H;��H;��H;��H;��H;��H;��H;��H;��H;��H;��H;��H;��H;��H;��H;��H;u�H;0�H;�H;��H;t�H;�H;��H;��H;B�H;z�H;��H;��H;��H;��H;N�H;�H;��H;T�H;��H;��H;i�H;B�H;>�H;c�H;��H;�H;��H;      ��H;�H;k�H;�H; �H;!�H;|�H;�H;��H;?�H;��H;��H;@�H;��H;J�H;��H;�H;C�H;\�H;\�H;%�H;��H;r�H;�H;a�H;��H;�H;@�H;d�H;��H;��H;��H;��H;��H;��H;��H;��H;��H;��H;��H;��H;��H;��H;��H;i�H;@�H;�H;��H;_�H;�H;s�H;��H;!�H;\�H;^�H;E�H;�H;��H;J�H;��H;@�H;��H;��H;?�H;��H;�H;|�H;%�H;��H;�H;j�H;�H;      Y�H;��H;2�H;�H;I�H;��H;w�H;O�H;a�H;��H;��H;��H; �H;0�H;(�H;�H;��H;�H;|�H;��H;��H;��H;��H;?�H;��H;W�H;��H;��H;+�H;j�H;��H;��H;��H;��H;��H;��H;��H;��H;��H;��H;��H;��H;��H;m�H;,�H;��H;��H;U�H;��H;?�H;��H;��H;��H;��H;}�H;�H;��H;�H;*�H;0�H; �H;��H;��H;��H;a�H;M�H;w�H;��H;C�H;�H;/�H;��H;      ǵH;�H;ĶH;�H;��H;��H;.�H;��H;��H;n�H;b�H;O�H;-�H;��H;��H;�H;M�H;d�H;*�H;��H;�H;j�H;��H;B�H;��H;��H;*�H;��H;��H;0�H;Y�H;u�H;��H;��H;��H;��H;��H;��H;��H;��H;��H;x�H;Y�H;2�H;��H;��H;*�H;��H;��H;D�H;��H;l�H;�H;��H;+�H;g�H;M�H;�H;��H;��H;-�H;P�H;b�H;p�H;��H;��H;/�H;��H;��H;�H;öH;�H;      y�H;�H;ߥH;��H;ͩH;��H;ӯH;v�H;H�H;G�H;`�H;a�H;9�H;��H;i�H;��H;��H;`�H;��H;�H;��H;m�H;��H;/�H;�H;��H;��H;4�H;��H;��H;)�H;\�H;��H;��H;��H;��H;��H;��H;��H;��H;��H;_�H;)�H;��H;��H;4�H;��H;��H;�H;/�H;��H;n�H;��H;�H;��H;a�H;��H;��H;i�H;��H;9�H;c�H;^�H;I�H;H�H;v�H;ӯH;��H;ʩH;��H;ߥH;�H;      Z�H;͌H;Q�H;��H;�H;�H;W�H;P�H;��H;�H;��H;!�H;r�H;�H;J�H;��H;��H;?�H;��H;i�H;��H;�H;��H;k�H;��H;��H;��H;��H;�H;}�H;��H;/�H;c�H;��H;��H;��H;��H;��H;��H;��H;c�H;0�H;��H;{�H;�H;��H;��H;��H;��H;l�H;��H;�H;��H;i�H;��H;@�H;��H;��H;J�H;~�H;r�H;!�H;��H;�H;��H;Q�H;V�H;�H;�H;��H;O�H;̌H;      �jH;kH;amH;�pH;�uH;/{H;��H;��H;�H;��H;>�H;��H;��H;�H;d�H;X�H;��H;��H;��H;��H;�H;��H;J�H;T�H;�H;��H;��H;��H;��H; �H;��H;��H;'�H;f�H;��H;��H;��H;��H;��H;f�H;'�H;��H;��H;�H;��H;��H;��H;��H;�H;U�H;I�H;��H;�H;��H;��H;��H;��H;Z�H;d�H;�H;��H;��H;>�H;��H;�H;��H;��H;1{H;�uH;�pH;bmH;kH;      "0H;�1H;M6H;>=H;0FH;fPH;[H;fH;�pH;�{H;��H;�H;�H;w�H;�H;(�H;~�H;�H;��H;��H;�H;��H;&�H;��H;��H;��H;p�H;��H;��H;��H;2�H;��H;��H;@�H;t�H;��H;z�H;��H;u�H;C�H;��H;��H;2�H;��H;��H;��H;p�H;��H;��H;��H;$�H;��H;�H;��H;��H;�H;}�H;*�H;�H;u�H;�H;�H;��H;�{H;�pH;fH;[H;cPH;=FH;@=H;P6H;�1H;      �G;��G;}�G;��G;"�G;�G;�H; *H;$@H;�SH;�dH;�sH;��H;ʎH;��H;i�H;�H;зH;��H;=�H;��H;��H;��H;|�H;n�H;��H;��H;q�H;��H;��H;��H;-�H;��H;�H;5�H;i�H;��H;g�H;6�H;�H;��H;.�H;��H;��H;��H;q�H;��H;��H;k�H;z�H;��H;��H;��H;=�H;��H;ԷH;�H;i�H;��H;ʎH;��H;�sH;�dH;�SH;&@H;*H;�H;�G;#�G;��G;|�G;�G;      7[F;�dF;�F;l�F;�F;�"G;7bG;�G;��G;bH;�)H;�GH;�^H;�qH;<�H;�H;.�H;��H;ȳH;��H;#�H;��H;��H;g�H;4�H;Z�H;��H;��H;��H;��H;��H;��H;U�H;��H;�H;F�H;F�H;F�H;�H;��H;T�H;��H;��H;��H;��H;��H;��H;\�H;1�H;e�H;��H;��H;�H;��H;ɳH;��H;.�H;�H;=�H;�qH;�^H;�GH;�)H;aH;��G;
�G;8bG;�"G;�F;i�F;�F;�dF;      �WC;	oC;�C;�D;d�D;>5E;�E;�[F;t�F;�LG; �G;|�G;Z!H;]FH;FaH;AvH;-�H;��H;�H;w�H;R�H;��H;��H;h�H;'�H;7�H;r�H;��H;�H;��H;
�H;��H;��H;f�H;��H;�H;�H;�H;��H;f�H;��H;��H;�H;��H;�H;��H;o�H;8�H;&�H;h�H;��H;��H;Q�H;z�H;�H;��H;,�H;AvH;FaH;]FH;[!H;|�G;�G;�LG;t�F;�[F;�E;>5E;c�D;�D;�C;	oC;      g�<;$�<;/]=;�O>;�?;��@;�7B;U�C;�D;��E;��F;�"G;ۚG;+�G;*H;iPH;MkH;p�H;d�H;i�H;"�H;��H;��H;b�H;c�H;g�H;y�H;��H;Q�H;k�H;)�H;>�H;:�H;�H;q�H;��H;��H;��H;t�H;�H;;�H;A�H;+�H;i�H;O�H;��H;w�H;h�H;a�H;c�H;��H;��H; �H;j�H;f�H;u�H;LkH;iPH;*H;+�G;ٚG;�"G;��F;��E;�D;U�C;�7B;��@; �?;�O>;0]=;�<;      �Y.;��.;f0;�2;^�4;��7;�|:;D]=;d�?;�7B;gD;YoE;NxF;W5G;ֶG;H;@H;bH;�zH;��H;@�H;�H;v�H;��H;��H;��H;��H;$�H;L�H;��H;��H;��H;��H;v�H;�H;P�H;x�H;N�H;�H;v�H;��H;��H;��H;��H;J�H;$�H;��H;��H;��H;��H;v�H;�H;;�H;��H;�zH;bH;@H;H;׶G;W5G;NxF;YoE;gD;7B;d�?;D]=;�|:;��7;d�4;�2;[0;��.;      ;��;�l;�Z;v`;�%;�+;��0;�G6;��:;��>;��A;�D;̲E;M�F;B{G;l�G;2H;![H;�vH;��H;x�H;�H;��H;��H;�H;��H;��H;��H;�H;k�H;f�H;��H;��H;��H;��H;�H;��H;��H;��H;��H;h�H;m�H;�H;��H;��H;��H;��H;��H;��H;�H;z�H;��H;�vH;#[H;2H;l�G;B{G;P�F;˲E;�D;��A;��>;��:;�G6;��0;�+;�%;�`;�Z; m;��;      �:o-�:Vg�:��:��:�^;j�;7�;��#;8�,;|�4;�:;�X?;�B;��D;�[F;GG;�G;~(H;�WH;�uH;��H;>�H;%�H;M�H;#�H;��H;�H;�H;��H;��H;�H;��H;�H;��H;��H;��H;��H;��H;�H;��H;�H;��H;��H;�H;�H;��H;&�H;O�H;"�H;>�H;��H;�uH;�WH;�(H;�G;GG;�[F;��D;�B;�X?;�:;z�4;6�,;��#;7�;i�;�^;��:��:Vg�:Y-�:      �e9��9h
�9�:��Y:�y�:�;�:��:�^;��;W";�r-;�G6;��<;?A;�0D;�F;X#G;��G;%H;�WH;�vH;��H;j�H;o�H;��H;9�H;��H;��H;e�H; �H;��H;��H;U�H;9�H;��H;%�H;��H;;�H;U�H;��H;��H; �H;b�H;��H;��H;7�H;��H;r�H;h�H;��H;�vH;�WH;%H;��G;Y#G;�F;�0D;?A;��<;�G6;�r-;V";��;�^;��:�;�:�y�:��Y:�:X
�9`�9      P����� кғ����Y� ���r89L5:Z/�:�d�:nB;^m;�?&;D2;�|:;6!@;߳C;��E;�G;��G;}(H;![H;�zH;f�H;�H;ɳH;��H;��H;��H;��H;��H;$�H;y�H;X�H;w�H;(�H;��H;(�H;w�H;X�H;x�H;&�H;��H;��H;��H;��H;��H;̳H;�H;b�H;�zH;![H;{(H; �G;�G;��E;߳C;6!@;�|:;D2;�?&;^m;nB;�d�:`/�:L5:�r89�����Y�ғ�� к~��      嚩�Y���+J���X��4�b��-���� Ix����!:
��:k��:ܯ;_ ;`�.;��8;u�?;�C;��E;[#G;�G;2H;bH;o�H;��H;��H;ԷH;�H;��H;C�H;a�H;a�H;�H;A�H;��H;d�H;��H;d�H;��H;B�H;�H;d�H;a�H;A�H;��H;
�H;ҷH;��H;��H;n�H;bH;2H;
�G;\#G;��E;�C;u�?;��8;`�.;_ ;ޯ;k��:��: !:��� Ix�����-�.�b��X��+J��]���      �B(�%�����_������˻	���b�A&����� t>���Y: �:�^;��;x�,;&`8;u�?;�C;�F;GG;n�G;@H;OkH;'�H;.�H;�H;}�H;��H;��H;��H;F�H;��H;
�H;��H;��H;��H;��H;��H;
�H;��H;F�H;��H;��H;��H;~�H;�H;/�H;)�H;KkH;@H;n�G;GG;�F;�C;y�?;%`8;x�,;��;�^; �:��Y: p>�����?&��b�	���˻�����_����
%�      �����x���#��JF{���]��E<����W�뻮���=d\���뺰[� 4: �:���:�[;z�,;��8;9!@;�0D;�[F;C{G;H;iPH;<vH;�H;i�H;&�H;U�H;��H;��H;�H;�H;��H;��H;��H;��H;��H;��H;��H;�H;�H;��H;��H;Q�H;&�H;f�H;�H;?vH;hPH;H;C{G;�[F;�0D;:!@;��8;z�,;�[;���:�: 4:�[����?d\�����W�뻩���E<���]�JF{��#���x��      c������o�wrμ׃��yv��O"��^N�����?ݻ\^��E����Y���9��:��:��;_�.;�|:;?A;��D;K�F;׶G;*H;@aH;?�H;��H;�H;d�H;F�H;c�H;��H;&�H;E�H;��H;��H;�H;��H;��H;F�H;$�H;��H;d�H;D�H;a�H;�H;��H;@�H;CaH;*H;ѶG;M�F;��D;?A;�|:;c�.;��;��:��:��9��Y�E��\^���?ݻ���^N�O"��yv��׃��wrμ�o����      en;�}\8��s/�@�!�~��e���prμ��������E<�$��
����N3�THx���9�:�^;a ;B2;��<;�B;˲E;W5G;+�G;XFH;�qH;ʎH;r�H;�H;w�H;��H;��H;*�H;��H;G�H;��H;6�H;��H;G�H;��H;(�H;��H;��H;v�H;ߴH;s�H;ȎH;�qH;ZFH;(�G;S5G;˲E;�B;��<;D2;c ;�^;�:��9PHx��N3�
���$���E<��������prμe���~��@�!��s/�}\8�      ���������Ȅ�pSt��Y�bn;�4O�w#���Oļ�����&R��_������N3�؅Y��3: �:ޯ;�?&;�G6;�X?;�D;QxF;ޚG;X!H;�^H;��H;�H;��H;k�H;2�H;)�H;��H;<�H;�H;~�H;<�H;~�H;�H;=�H;��H;)�H;2�H;k�H;��H;�H;��H;�^H;]!H;ؚG;MxF;�D;�X?;�G6;�?&;�; �: 4:؅Y��N3������_��&R������Oļw#��4O�an;��Y�pSt��Ȅ�����      �ѽ\ν}�ý䳽>���M����d�v\8�z��ټov����Y��_����B���[���Y:k��:\m;�r-;�:;��A;VoE;�"G;v�G;�GH;�sH;�H;��H;�H;V�H;E�H;��H;��H;��H;V�H;�H;V�H;��H;��H;��H;H�H;W�H;�H;��H;�H;�sH;�GH;y�G;�"G;ToE;��A;!�:;�r-;^m;s��:��Y:�[�A������_���Y�ov��ټz��v\8���d� M��>���䳽}�ý\ν      ��#]�ֈ�s}���|�ý�u��Ε���K�����o�ov���&R�&��\^����� |>���:nB;Z";x�4;��>;gD;��F;�G;�)H;�dH;��H;>�H;��H;V�H;[�H;��H;��H;N�H;:�H;��H;;�H;N�H;��H;��H;^�H;W�H;��H;;�H;��H;�dH;�)H;�G;��F;eD;��>;|�4;X";nB;
��: |>����\^��%���&R�ov���o�����K�Ε���u��|�ý��s}�ֈ�#]�      �+X��T��nH��6��� �l��H�䳽�����mR����ټ�����E<��?ݻAd\������ :�d�:��;6�,;��:;�7B;��E;�LG;aH;SH;�{H;��H;�H;@�H;n�H;~�H;;�H;��H; �H;��H; �H;��H;<�H;|�H;k�H;@�H;�H;��H;�{H;SH;aH;�LG;��E;�7B;��:;6�,;��;�d�:!:����@d\��?ݻ�E<�����ټ����mR�����䳽H�l���� ��6��nH��T�      㰖��������*|�PS\�� :����Z�p$�������K�z���Oļ����������A&����V/�:�^;��#;�G6;a�?;�D;p�F;��G;"@H;�pH;�H;��H;>�H;}�H;X�H;��H;��H;�H;��H;�H;��H;��H;V�H;}�H;>�H;��H;�H;�pH; @H;��G;t�F;�D;`�?;�G6;��#;�^;V/�:���C&������������Oļz���K�����p$���Z���� :�PS\��*|�������      D�;9ɾ㼾B�������Mw��nH�����Z�䳽Ε��v\8�w#������^N�W���b�Ix�P5:��:4�;��0;D]=;R�C;�[F;�G;�)H;fH;��H;F�H;k�H;��H;F�H;��H;^�H;��H;��H;��H;\�H;��H;D�H;��H;m�H;F�H;��H;fH;�)H;
�G;�[F;P�C;E]=;��0;7�;��:X5:Ix��b�V��^N�����w#��v\8�Ε��䳽�Z񽳯��nH��Mw�����B��㼾9ɾ      1y��v�m���E�߾����D��A����nH���Hὡu����d�4O�qrμO"�����		�����pr89�;�:b�;�+;}|:;�7B;�E;4bG;�H;[H;��H;L�H;ȯH;$�H;s�H;t�H;7�H;�H;��H;�H;7�H;t�H;p�H;%�H;ȯH;J�H;��H;[H;�H;4bG;�E;�7B;||:;�+;d�;�;�:pr89���
	�����O"��qrμ4O���d��u��H����nH�A���D������E�߾m����v�      �O/�sM+�Z�����KW��9ɾD���Mw�� :�l��|�ýM��bn;�f���yv���E<��˻��-�(���y�:�^;�%;��7;��@;:5E;�"G; �G;cPH;2{H;�H;��H;��H;��H;"�H;>�H;�H;��H;�H;>�H;$�H;��H;��H;��H;ޗH;/{H;cPH;�G;�"G;<5E;~�@;��7;�%;�^;�y�:(����-��˻�E<�yv��f���bn;�M��|�ýl��� :��Mw�D��9ɾKW�����Z��sM+�      :�X�YvS�9E��O/��S�KW����������PS\��� ���>����Y���׃����]�����3�b���Y���Y:��:r`;b�4;�?;`�D;
�F;�G;/FH;}uH;�H;��H;��H;?�H;��H;O�H;D�H;'�H;D�H;N�H;��H;=�H;��H;��H;ޓH;|uH;/FH;!�G;�F;a�D;�?;f�4;r`;��:��Y:��Y�1�b�������]�׃�����Y�>����彔� �PS\���������KW���S��O/�9E�YvS�      � ����y�c�h��N��O/����E�߾B���*|��6�s}�䳽pSt�A�!�wrμLF{��_� Y��ؓ���:��:�Z;�2;�O>;�D;i�F;��G;B=H;�pH;��H;v�H;�H;�H;�H;��H;��H;��H;��H;��H;�H;�H;�H;x�H;��H;�pH;B=H;��G;i�F;�D;�O>;�2;�Z; ��:�:֓�� Y���_�LF{�wrμA�!�pSt�䳽s}��6��*|�B��E�߾����O/��N�c�h���y�      ?v��c���X ��c�h�9E�Z��m���㼾����nH�ֈ�~�ý�Ȅ��s/��o��#�����.J��2к 
�9@g�:�l;S0;!]=;��C;�F;|�G;F6H;]mH;G�H;ѥH;��H;(�H;n�H;��H;0�H;�H;1�H;��H;n�H;&�H;��H;ѥH;D�H;ZmH;F6H;|�G;�F;��C;]=;V0;�l;Dg�:0
�92к.J������#���o��s/��Ȅ�~�ýֈ��nH����㼾m���Z��9E�c�h�X ��c���      h��1���d�����y�YvS�sM+��v�9ɾ�����T�#]�\ν����~\8�����x��	%�Y������(�9Y-�:p�;��.;�<;�nC;�dF;�G;�1H;kH;ǌH;ӤH;�H;��H;��H;��H;��H;��H;��H;��H;��H;��H;�H;ӤH;ŌH;kH;�1H;�G;�dF;�nC;�<;��.;p�;]-�:�9���X���
%��x�����~\8�����\ν#]��T�����9ɾ�v�sM+�YvS���y�c���1���      IEb�c]��N���7����v� ���˾��-�j��!,�u���P��Km�1��@,˼˪x�b���1��$�����:Q�:�;B�1;2,>;��C;�wF;��G;� H;�>H;�hH;Z�H;|�H;C�H;#�H;��H;4�H;��H;5�H;��H;#�H;B�H;}�H;Z�H;�hH;�>H;� H;��G;�wF;��C;/,>;F�1;�;U�:��:$����1��c��˪x�@,˼1��Km�P��u����!,�-�j�����˾v� ������7��N�c]�      c]�g�W��TI�v3� E�������Ǿy����f�;)�*��x;���Fi��k���Ǽ�[t�U�	�8Ȅ�4X���:���:��;WJ2;OZ>;H	D;F;D�G;H;�?H;�iH;��H;�H;|�H;A�H;��H;`�H;��H;`�H;��H;A�H;z�H;�H;��H;�iH;�?H;H;D�G;~F;H	D;KZ>;]J2;��;���:�:4X��8Ȅ�U�	��[t���Ǽ�k��Fi�x;��*��;)��f�y�����Ǿ���� E�v3��TI�g�W�      �N��TI���;�1�'�l��쾃���{󐾷Z��K ��s�E����&^���"����g�����u�!��3<:���: ;dg3;��>;xBD;��F;�G;�H;OBH;{kH;\�H;�H;4�H;�H;v�H;��H;N�H;��H;u�H;߼H;2�H;�H;\�H;xkH;KBH;�H;�G;��F;xBD;��>;gg3; ;��:3<:!���u������g��"����&^�E����s潨K ��Z�{󐾃�����l�1�'���;��TI�      ��7�v3�1�'����v� ��{Ծ"���J���}�F�����ӽ���e�L�Ov��뮼\T�����PV���=��)i:^��:�z ;�$5;��?;�D;ϺF;��G;�H;�FH;�nH;��H;��H;w�H;�H;=�H;\�H;��H;\�H;=�H;�H;u�H;��H;��H;�nH;�FH;�H;��G;ϺF;�D;��?;�$5;�z ;b��:�)i:��=��PV����\T��뮼Ov�e�L�����ӽ���}�F�J���"����{Ծv� ����1�'�v3�      ��� E�l�v� �Y�ݾm���X͓��f��>/�����'���섽U�6��t�w��h�:�2Tʻ�.�p۷�ht�:�;��$;�Y7;Y�@;�	E;�F;;�G;�H;ALH;�rH;��H;ѤH;)�H;#�H;7�H;Q�H;��H;O�H;6�H;#�H;'�H;ӤH;��H;�rH;>LH;�H;<�G;�F;�	E;U�@;�Y7;��$;�;ft�:p۷��.�2Tʻh�:�w���t�U�6��섽�'������>/��f�X͓�m���Y�ݾv� �l� E�      v� ��������{Ծm���y���^�x��SC��^���޽D����e�-��L�Ѽ,G������R�� ���`ݤ8뇲:�Y;P�);��9;��A;��E;�G; �G;k!H;DSH;�wH;y�H;��H;F�H;��H;}�H;��H;��H;��H;}�H;��H;F�H;��H;y�H;�wH;@SH;k!H;�G;�G;��E;��A;��9;P�);�Y;釲:@ݤ8 ����R�����,G��K�Ѽ-���e�D�����޽�^��SC�^�x�y���m����{Ծ�쾤���      ��˾��Ǿ����#���X͓�^�x���J��K �r���"������?����뮼6�[�.���&3|��W��x�:j�:�';n/;fg<;�C;oF;�NG;��G;2-H;r[H;�}H;˗H;ΪH;��H;��H;�H;��H;�H;��H;�H;��H;��H;ϪH;˗H;�}H;o[H;2-H;��G;�NG;lF;�C;dg<;n/;�';d�:x�:�W��&3|�.���6�[��뮼���?����"��r����K ���J�^�x�X͓�#���������Ǿ      ��y���{�J����f��SC��K �tn���Ž����Z��k�&}ռ3X��ky-�9���|.����P�:�+�:��;4;9�>; D;�wF;5�G;��G;�9H;[dH;w�H;��H;f�H;t�H;��H;��H;Y�H;v�H;Y�H;��H;��H;r�H;g�H;��H;w�H;XdH;�9H;��G;5�G;�wF;�D;9�>;4;��;�+�:�P�:���}.�9���ky-�3X��'}ռ�k��Z�����Žtn���K ��SC��f�J���{�y���      -�j��f��Z�}�F��>/��^�r����ŽJ ���Fi��Q+��t�vT��y�W�����1��:Ⱥ�W�9�P�:�Y;��(;
�8;�A;�E;
�F;m�G;�H;�FH;�mH;��H;ơH;D�H;q�H;��H;��H;��H;��H;��H;��H;��H;q�H;F�H;ġH;��H;�mH;�FH;�H;m�G;�F;�E;�A;
�8;��(;�Y;�P�: X�98Ⱥ�1�����z�W�vT���t�Q+��Fi�J ���Žr����^��>/�}�F��Z��f�      �!,�;)��K ���������޽"������Fi��0����鷼��x�����.��b�(� ���*i:���:@�;��0;O�<;�C;��E;=G;��G;�$H;gTH;�wH;�H;�H;R�H;��H;C�H;��H;��H;��H;��H;��H;C�H;��H;T�H;�H;�H;�wH;gTH;�$H;��G;=G;��E;�C;O�<;��0;>�;���:�*i:��b�(��.�������x�鷼����0��Fi����"����޽�������K �;)�      u���*��s��ӽ�'��D�������Z��Q+�����"��#G��ʻ0��׻ޕb�NW���X�9С�:,`;�*';�Y7;$@;+�D;��F;�G;��G;;8H;bH;�H;]�H;��H;x�H;��H;��H;��H;U�H;A�H;U�H;��H;��H;��H;{�H;��H;]�H;�H;bH;:8H;��G;�G;��F;(�D;$@;�Y7;�*';,`;֡�:�X�9NW��ߕb��׻ʻ0�#G���"������Q+��Z����D����'���ӽ�s�*��      P��x;��E�������섽�e��?��k��t�鷼#G���e7�Ƙ�
Ȅ��0�@�t�&u�:,�:z;�1;X�<;f�B;,�E;G;��G;eH;wJH;aoH;�H;��H;�H;��H;��H;%�H;��H;�H;��H;�H;��H;$�H;��H;��H;�H;��H;�H;coH;uJH;dH;��G;G;(�E;f�B;X�<;�1;z;,�:"u�:��t��0�
Ȅ�Ř껎e7�#G��鷼�t��k��?��e��섽���E���x;��      Km��Fi��&^�d�L�U�6�-����&}ռvT����x�ɻ0�Ƙ����$���ط��n`:��:�;+�*;>�8;�@;<�D;m�F;�}G;��G;�1H;�[H;u|H;ƕH;ߨH;��H;��H;��H;��H;��H;��H;{�H;��H;��H;��H;��H;��H;��H;ߨH;ÕH;u|H;�[H;�1H;��G;�}G;i�F;<�D;�@;<�8;+�*;�;��:�n`:�ط�#�����Ƙ�ɻ0���x�uT��'}ռ��-��V�6�d�L��&^��Fi�      0���k��Nv��t�J�Ѽ�뮼3X��x�W�����׻	Ȅ�"��P���4<:a��:�Y;�t%;�$5;�Z>;aC;��E;9*G;l�G;H;HH;ulH;��H;�H;ɯH;׼H;��H;��H;�H;~�H;v�H;6�H;v�H;~�H;�H;��H;��H;ؼH;ȯH;	�H;��H;rlH;HH;H;h�G;5*G;��E;aC;�Z>;�$5;�t%;�Y;[��:�4<:H��#��	Ȅ��׻���x�W�3X���뮼J�Ѽ�t�Nv���k�      @,˼��Ǽ�"���뮼w��+G��5�[�ky-�����.��ޕb��0��ط��4<:�L�:�\;��!;�J2;�g<;U0B;2CE;0�F;U�G;��G;�4H;�\H;|H;��H;��H;`�H;��H;H�H;��H;W�H;X�H;�H;��H;�H;Z�H;X�H;��H;K�H;��H;]�H;��H;��H;|H;�\H;�4H;��G;N�G;0�F;1CE;U0B;�g<;�J2;��!;�\;�L�:�4<:�ط��0�ޕb��.�����ly-�5�[�+G��w���뮼�"����Ǽ      ʪx��[t���g�[T�h�:����*���9����1��_�(�LW����t��n`:_��:�\;{ ;��0;a;;	=A;�D;�wF;�cG;[�G;�!H;�MH;�oH;|�H;��H;̯H;��H;n�H;��H;c�H;v�H;�H;��H;-�H;��H;�H;u�H;a�H;��H;m�H;��H;ƯH;��H;x�H;�oH;�MH;�!H;V�G;�cG;�wF;�D;=A;b;;��0;{ ;�\;_��:�n`: �t�NW��_�(��1��:���+������h�:�[T���g��[t�      b��R�	�������2Tʻ�R��3|�{.�6Ⱥ����X�9&u�:��:�Y;��!;��0;�:;��@;CD;�2F;8G;��G;�H;q@H;-dH;̀H;}�H;M�H;P�H;U�H;��H;��H;��H;v�H;��H;�H;��H;�H;��H;v�H;��H;��H;��H;R�H;L�H;L�H;x�H;̀H;-dH;k@H;�H;��G;|8G;�2F;CD;��@;�:;��0;��!;�Y;��:&u�:�X�9���4Ⱥ}.�3|��R��2Tʻ������T�	�      �1��7Ȅ��u��PV��.�����W������W�9�*i:֡�:,�:�;�t%;�J2;^;;��@;sD;F;/G;��G;�H;�5H;�ZH;<xH;H�H;2�H;�H;�H;a�H;w�H;#�H;8�H;2�H;F�H;b�H;��H;b�H;F�H;0�H;7�H;%�H;u�H;`�H;�H;�H;/�H;H�H;;xH;�ZH;�5H;�H;�G;.G;F;tD;��@;^;;�J2;�t%;�;,�:֡�: +i:X�9���W������.��PV��u�;Ȅ�      ���4X��� ����=��۷��ݤ8��:�P�:�P�:���:,`;{;*�*;�$5;�g<;=A;CD;F;�G;��G;n�G;�-H;"SH;aqH;�H;ǝH;��H;�H;C�H;��H;��H;��H;]�H;��H;��H;��H;��H;��H;��H;��H;[�H;��H;��H;��H;>�H;�H;��H;ɝH;�H;\qH;SH;�-H;i�G;��G;�G;F;CD;=A;�g<;�$5;*�*;};,`;���:�P�:�P�:��:`ޤ8X۷���=�� ��4X��      ��:d�: 3<:�)i:ft�:釲:d�:�+�:�Y;B�;�*';�1;:�8;�Z>;R0B;�D;�2F;,G;��G;#�G;�)H;�NH;|lH;S�H;p�H;��H;��H;8�H;��H;�H;B�H;2�H;;�H;c�H;��H;��H;��H;��H;��H;c�H;:�H;4�H;B�H;�H;��H;5�H;��H;��H;m�H;N�H;ylH;�NH;�)H;#�G;��G;+G;�2F;�D;R0B;�Z>;:�8;�1;�*';@�;�Y;�+�:d�::zt�:�)i: 3<:@�:      k�:
��:��:T��:�;�Y;�';��;��(;��0;�Y7;T�<;�@;aC;1CE;�wF;8G;��G;n�G;�)H;�LH;jH;=�H;f�H;��H;۳H;žH;m�H;0�H;��H;�H;^�H;��H;��H;��H;��H;��H;��H;��H;��H;��H;`�H;�H;��H;,�H;k�H;þH;ڳH;��H;`�H;<�H;jH;�LH;�)H;n�G;��G;|8G;�wF;/CE;aC;�@;T�<;�Y7;��0;��(;��;�';�Y;�;V��:��:���:      �;��;;�z ;��$;[�);x/;(4;�8;P�<;$@;i�B;?�D;��E;2�F;�cG;��G;�H;�-H;�NH;jH;Q�H;��H;��H;�H;ʼH;��H;��H;U�H;��H;��H;9�H;V�H;��H;��H;u�H;��H;u�H;��H;��H;S�H;9�H;��H;��H;Q�H;��H;��H;ʼH;�H;��H;��H;P�H;jH;�NH;�-H;�H;��G;�cG;3�F;��E;?�D;i�B;$@;R�<;�8;%4;x/;[�);��$;�z ;;��;      M�1;]J2;gg3;�$5;�Y7;��9;jg<;:�>;A;�C;-�D;.�E;l�F;;*G;S�G;Y�G;�H;�5H;"SH;}lH;=�H;��H;5�H;�H;��H;u�H;m�H;?�H;��H;��H;��H;��H;��H;��H;��H;7�H;��H;6�H;��H;��H;��H;��H;��H;��H;��H;?�H;h�H;u�H;��H;߰H;1�H;��H;9�H;~lH;!SH;�5H;�H;X�G;R�G;;*G;l�F;.�E;-�D;�C;�A;9�>;lg<;��9;�Y7;�$5;jg3;MJ2;      G,>;ZZ>;��>;��?;Z�@;��A;�C;�D;�E;��E;��F;G;�}G;j�G;��G;�!H;n@H;�ZH;_qH;S�H;b�H;��H;�H;(�H;��H;��H;W�H;!�H; �H;�H;u�H;F�H;��H;��H;q�H;��H;�H;��H;r�H;��H;��H;F�H;t�H;�H;��H;!�H;T�H;��H;��H;#�H;߰H;��H;]�H;S�H;_qH;�ZH;k@H;�!H;��G;j�G;�}G;G;��F;��E;�E;�D;�C;��A;a�@;��?;��>;OZ>;      ��C;P	D;hBD;�D;�	E;��E;mF;�wF;
�F;=G;�G;��G;��G;H;�4H;�MH;3dH;>xH;�H;w�H;��H;�H;��H;��H;V�H;�H;��H;��H;��H;��H;��H;��H;��H;j�H;�H;l�H;v�H;l�H;�H;g�H;��H;��H;��H;��H;��H;��H;��H;�H;V�H;��H;��H;�H;��H;w�H;�H;AxH;0dH;�MH;�4H;H;��G;��G;�G;=G;
�F;�wF;mF;ÄE;�	E;�D;hBD;R	D;      �wF;�F;��F;ϺF;!�F;�G;�NG;2�G;n�G; �G;��G;fH;�1H;HH;�\H;�oH;ʀH;F�H;ƝH;��H;ٳH;ɼH;r�H;��H;�H;}�H;I�H;D�H;��H;��H;B�H;~�H;`�H;#�H;��H;��H;��H;��H;��H;#�H;]�H;~�H;@�H;��H;��H;D�H;F�H;~�H;�H;��H;p�H;ǼH;ӳH;��H;ĝH;F�H;ʀH;�oH;�\H;HH;�1H;fH;��G;��G;o�G;2�G;�NG;�G;(�F;кF;��F;�F;      �G;I�G;�G;��G;?�G;'�G;��G;��G;�H;�$H;>8H;{JH;�[H;slH;|H;|�H;�H;0�H;��H;��H;ǾH;��H;k�H;Z�H;��H;L�H;-�H;��H;u�H;#�H;b�H;=�H;�H;��H;��H;2�H;@�H;2�H;��H;��H;
�H;:�H;`�H; �H;r�H;��H;*�H;J�H;��H;X�H;j�H;��H;þH;��H;��H;0�H;|�H;{�H;|H;slH;�[H;{JH;>8H;�$H;�H;��G;��G;$�G;F�G;��G;�G;J�G;      � H; H;�H;�H;�H;n!H;9-H;�9H;�FH;nTH;	bH;hoH;v|H;��H;��H;��H;M�H;�H;�H;;�H;m�H;��H;@�H;$�H;}�H;G�H;��H;��H;�H;3�H;3�H;�H;��H;�H;F�H;��H;��H;��H;F�H;�H;��H;�H;2�H;/�H;�H;��H;��H;E�H;~�H;$�H;?�H;��H;j�H;9�H;�H;�H;J�H;��H;��H;��H;u|H;hoH;bH;lTH;�FH;�9H;9-H;k!H;�H;�H;�H;(H;      ?H;�?H;NBH;�FH;ALH;DSH;x[H;`dH;�mH;�wH;�H;�H;ƕH;�H;��H;ͯH;S�H;�H;B�H;��H;0�H;T�H;��H;�H;��H;��H;r�H;�H;O�H;!�H;��H;��H;�H;e�H;��H;��H;��H;��H;��H;e�H;��H;��H;��H;�H;N�H;�H;q�H;��H;��H;�H;��H;T�H;.�H;��H;B�H;�H;R�H;ͯH;��H;�H;ƕH;�H;�H;�wH;�mH;^dH;x[H;ESH;HLH;�FH;NBH;�?H;       iH;�iH;�kH;�nH;�rH;�wH;�}H;~�H;��H;��H;f�H;áH;�H;үH;d�H;��H;X�H;]�H;��H;�H;��H;��H;��H;�H;��H;��H; �H;2�H;�H;��H;��H;�H;S�H;��H;��H;��H;��H;��H;��H;��H;N�H;�H;��H;��H;�H;/�H;�H;��H;��H;�H;��H;��H;��H;�H;��H;^�H;V�H;��H;d�H;ЯH;�H;��H;f�H;��H;��H;��H;�}H;�wH;�rH;�nH;�kH;�iH;      ^�H;�H;i�H;��H;ȏH;y�H;ԗH;��H;ΡH;#�H;��H;'�H;��H;�H;��H;u�H;��H;w�H;��H;I�H;#�H;��H;��H;x�H;��H;D�H;_�H;4�H;��H;��H;	�H;a�H;��H;��H;�H;�H;�H;�H;�H;��H;��H;b�H;	�H;��H;��H;4�H;]�H;@�H;��H;x�H;��H;��H; �H;G�H;��H;u�H;��H;t�H;��H;߼H;��H;%�H;��H;#�H;ΡH;��H;ԗH;|�H;ŏH;��H;j�H;�H;      ��H;��H;�H;��H;פH;��H;ҪH;p�H;J�H;U�H;��H;��H;��H;��H;O�H;��H;�H;%�H;��H;;�H;d�H;@�H;��H;J�H;��H;~�H;;�H;�H;��H;�H;\�H;��H;��H;�H;�H;6�H;R�H;6�H;�H;�H;��H;��H;^�H;�H;��H;�H;:�H;z�H;��H;I�H;��H;=�H;c�H;;�H;��H;&�H; �H;��H;N�H;��H;��H;��H;��H;U�H;K�H;m�H;ҪH;��H;֤H;��H;�H;�H;      J�H;��H;=�H;~�H;3�H;G�H;ƸH;�H;z�H;��H;��H;��H;��H;��H;��H;g�H;��H;4�H;`�H;B�H;��H;V�H;��H;��H;��H;a�H;�H;��H;�H;X�H;��H;��H;�H;+�H;O�H;D�H;7�H;D�H;O�H;+�H;��H;��H;��H;X�H;�H;��H;�H;^�H;��H;��H;��H;U�H;��H;B�H;_�H;5�H;��H;g�H;��H;��H;��H;��H;��H;��H;z�H;}�H;ƸH;K�H;,�H;�H;?�H;��H;      5�H;Q�H;ݼH;�H;0�H;��H;��H;��H;��H;G�H;��H;+�H;��H;�H;\�H;�H;}�H;2�H;��H;k�H;��H;��H;��H;��H;a�H;#�H;��H;�H;c�H;��H;��H;�H;$�H;7�H;b�H;p�H;N�H;p�H;b�H;7�H;"�H;�H;��H;��H;f�H;�H;��H; �H;a�H;��H;��H;��H;��H;k�H;��H;3�H;{�H;�H;\�H;�H;��H;+�H;��H;G�H;��H;��H;��H;��H;&�H;�H;ݼH;I�H;      ��H;�H;��H;G�H;U�H;{�H;�H;��H;��H;��H;��H;��H;��H;��H;`�H;�H;��H;D�H;��H;��H;��H;��H;��H;u�H;�H;��H;��H;F�H;��H;��H;��H;�H;M�H;d�H;G�H;d�H;��H;d�H;G�H;d�H;J�H;�H;��H;��H;��H;F�H;��H;��H;�H;r�H;��H;��H;��H;��H;��H;F�H;��H;�H;^�H;��H;��H;��H;��H;��H;��H;��H;�H;��H;J�H;I�H;��H; �H;      1�H;k�H;��H;b�H;c�H;�H;��H;f�H;
�H;��H;]�H;�H;��H;��H;�H;��H;�H;]�H;��H;��H;��H;w�H;6�H;��H;g�H;��H;1�H;��H;��H;��H;�H;:�H;C�H;r�H;d�H;\�H;k�H;\�H;d�H;p�H;A�H;=�H;�H;��H;��H;��H;/�H;��H;h�H;��H;6�H;w�H;��H;��H;��H;_�H;�H;��H;�H;}�H;��H;�H;\�H;��H;
�H;c�H;��H;��H;V�H;b�H;��H;a�H;      ��H;��H;`�H;��H;��H;��H;�H;�H;�H;��H;H�H;��H;�H;?�H;��H;4�H;��H;��H;��H;��H;��H;��H;��H;�H;o�H;��H;?�H;��H;��H;��H;�H;Y�H;7�H;R�H;��H;m�H;Y�H;m�H;��H;R�H;5�H;[�H;�H;��H;��H;��H;=�H;��H;o�H;�H;��H;��H;��H;��H;��H;��H;��H;4�H;��H;?�H;�H;��H;H�H;��H;�H;}�H;�H;��H;��H;��H;`�H;��H;      1�H;k�H;��H;c�H;d�H;�H;��H;f�H;
�H;��H;]�H;�H;��H;��H;�H;��H;�H;]�H;��H;��H;��H;w�H;6�H;��H;h�H;��H;1�H;��H;��H;��H;�H;:�H;C�H;r�H;d�H;\�H;k�H;\�H;d�H;p�H;A�H;=�H;�H;��H;��H;��H;/�H;��H;g�H;��H;6�H;w�H;��H;��H;��H;_�H;�H;��H;�H;}�H;��H;�H;]�H;��H;
�H;c�H;��H;��H;X�H;b�H;��H;a�H;      ��H;�H;��H;I�H;U�H;{�H;�H;��H;��H;��H;��H;��H;��H;��H;^�H;�H;��H;D�H;��H;��H;��H;��H;��H;t�H;�H;��H;��H;F�H;��H;��H;��H;�H;M�H;d�H;G�H;d�H;��H;d�H;G�H;d�H;J�H;�H;��H;��H;��H;F�H;��H;��H;�H;r�H;��H;��H;��H;��H;��H;F�H;��H;�H;^�H;��H;��H;��H;��H;��H;��H;��H;�H;��H;J�H;G�H;��H; �H;      7�H;Q�H;޼H;�H;0�H;��H;��H;��H;��H;G�H;��H;+�H;��H;�H;\�H;�H;}�H;2�H;��H;j�H;��H;��H;��H;��H;a�H;"�H;��H;�H;c�H;��H;��H;�H;$�H;7�H;b�H;p�H;N�H;n�H;b�H;7�H;"�H;�H;��H;��H;f�H;�H;��H;#�H;a�H;��H;��H;��H;��H;k�H;��H;3�H;{�H;�H;\�H;�H;��H;+�H;��H;G�H;��H;��H;��H;��H;%�H;�H;ݼH;I�H;      M�H;��H;?�H;��H;1�H;H�H;ƸH;}�H;z�H;��H;��H;��H;��H;��H;��H;g�H;��H;4�H;_�H;A�H;��H;U�H;��H;��H;��H;`�H;�H;��H;�H;X�H;��H;��H;�H;)�H;O�H;D�H;7�H;D�H;O�H;)�H;��H;��H;��H;Z�H;�H;��H;
�H;`�H;��H;��H;��H;V�H;��H;C�H;`�H;4�H;��H;g�H;��H;��H;��H;��H;��H;��H;z�H;{�H;ƸH;M�H;)�H;�H;<�H;��H;      ��H;��H;�H;��H;ؤH;��H;֪H;p�H;K�H;U�H;�H;��H;��H;��H;N�H;��H;�H;%�H;��H;<�H;g�H;=�H;��H;I�H;��H;{�H;:�H;�H;��H;�H;^�H;��H;��H;�H;�H;6�H;R�H;6�H;�H;�H;��H;��H;\�H;�H;��H;�H;:�H;|�H;��H;J�H;��H;@�H;c�H;;�H;��H;&�H; �H;��H;N�H;��H;��H;��H;�H;V�H;M�H;n�H;֪H;��H;֤H;��H;�H;�H;      ^�H;�H;i�H;��H;ȏH;x�H;ԗH;��H;ΡH;"�H;��H;%�H;��H;�H;��H;u�H;��H;t�H;��H;G�H;%�H;��H;��H;z�H;��H;B�H;]�H;4�H;��H;��H;	�H;a�H;��H;��H;�H;�H;�H;�H;�H;��H;��H;b�H;	�H;��H;��H;4�H;_�H;C�H;��H;x�H;��H;��H; �H;I�H;��H;w�H;��H;u�H;��H;�H;��H;'�H;��H;%�H;ΡH;��H;ԗH;|�H;ŏH;��H;i�H;�H;      �hH;�iH;�kH;�nH;�rH;�wH;�}H;��H;��H;��H;f�H;áH;�H;үH;d�H;��H;X�H;]�H;��H;�H;��H;��H;��H;
�H;��H;��H;�H;/�H;�H;��H;��H;�H;P�H;��H;��H;��H;��H;��H;��H;��H;P�H;�H;��H;��H;�H;2�H;�H;��H;��H;�H;��H;��H;��H;�H;��H;^�H;V�H;��H;d�H;ЯH;�H;áH;f�H;��H;��H;��H;�}H;�wH;�rH;�nH;�kH;�iH;      ?H;�?H;UBH;�FH;HLH;ASH;|[H;adH;�mH;�wH;�H;�H;ƕH;�H;��H;ͯH;S�H;�H;B�H;��H;3�H;T�H;��H;�H;��H;��H;q�H;�H;N�H;�H;��H;��H; �H;e�H;��H;��H;��H;��H;��H;e�H; �H;��H;��H;�H;O�H;�H;t�H;��H;��H;�H;��H;T�H;.�H;��H;B�H;�H;R�H;ϯH;��H;�H;ƕH;�H;�H;�wH;�mH;`dH;|[H;DSH;CLH;�FH;VBH;�?H;      � H;H;�H;�H;�H;k!H;9-H;�9H;�FH;lTH;	bH;hoH;u|H;��H;��H;��H;L�H;�H;�H;9�H;o�H;��H;@�H;$�H;~�H;E�H;��H;��H;�H;2�H;2�H;�H;��H;�H;D�H;��H;��H;��H;F�H;�H;��H;�H;3�H;0�H;�H;��H;��H;H�H;}�H;$�H;?�H;��H;j�H;;�H;�H;�H;L�H;��H;��H;��H;v|H;hoH;bH;nTH;�FH;�9H;9-H;k!H;�H;�H;�H;+H;      ��G;J�G;�G;��G;?�G;#�G;��G;��G;�H;�$H;>8H;{JH;�[H;slH;|H;|�H;}�H;/�H;��H;��H;ȾH;��H;k�H;X�H;��H;J�H;-�H;��H;t�H;!�H;`�H;:�H;�H;��H;��H;2�H;@�H;1�H;��H;��H;�H;>�H;b�H;!�H;t�H;��H;,�H;L�H;��H;X�H;j�H;��H;ľH;��H;��H;2�H;}�H;{�H;|H;slH;�[H;{JH;?8H;�$H;�H;��G;��G;!�G;@�G;��G;�G;B�G;      �wF;�F;��F;ӺF;$�F;�G;�NG;5�G;m�G;��G;��G;eH;�1H;HH;�\H;�oH;ʀH;E�H;ĝH;��H;ٳH;ǼH;r�H;��H;�H;}�H;I�H;D�H;��H;��H;@�H;|�H;^�H;#�H;��H;��H;��H;��H;��H;#�H;]�H;�H;B�H;��H;��H;D�H;H�H;~�H;�H;��H;r�H;ɼH;ԳH;��H;ƝH;F�H;ɀH;�oH;�\H;HH;�1H;fH;��G;��G;n�G;4�G;�NG;�G;(�F;кF;��F;|F;      ��C;P	D;gBD;�D;�	E;��E;mF;�wF;	�F;=G;�G;��G;��G;H;�4H;�MH;1dH;>xH;�H;v�H;��H;�H;��H;��H;V�H;�H;��H;��H;��H;��H;��H;��H;��H;g�H;�H;n�H;v�H;l�H;�H;h�H;��H;��H;��H;��H;��H;��H;��H;�H;V�H;��H;��H;�H;��H;x�H;�H;AxH;0dH;�MH;�4H;H;��G;��G;�G;=G;
�F;�wF;mF;��E;�	E;�D;hBD;P	D;      J,>;YZ>;�>;��?;V�@; �A;�C;D;�E;��E;��F;G;�}G;j�G;��G;�!H;m@H;�ZH;_qH;S�H;b�H;��H;�H;&�H;��H;��H;W�H;!�H; �H;�H;t�H;E�H;��H;��H;o�H;��H;�H;��H;r�H;��H;��H;H�H;u�H;
�H;��H;!�H;V�H;��H;��H;(�H;�H;��H;_�H;S�H;_qH;�ZH;m@H;�!H;��G;j�G;�}G;G;��F;��E;�E; D;�C;�A;f�@;��?;�>;NZ>;      F�1;jJ2;yg3;�$5;�Y7;��9;pg<;:�>;�A;�C;-�D;/�E;j�F;;*G;S�G;Y�G;�H;�5H;!SH;}lH;?�H;��H;4�H;�H;��H;s�H;m�H;?�H;��H;��H;��H;��H;��H;��H;��H;6�H;��H;7�H;��H;��H;��H;��H;��H;��H;��H;?�H;j�H;v�H;��H;�H;3�H;��H;9�H;~lH;"SH;�5H;�H;Y�G;U�G;;*G;j�F;.�E;-�D;�C;A;9�>;pg<;��9;�Y7;�$5;ng3;ZJ2;      �;��;;�z ;��$;Z�);x/;(4;�8;R�<;$@;i�B;?�D;��E;2�F;�cG;��G;�H;�-H;�NH;jH;P�H;��H;��H;�H;ɼH;��H;��H;T�H;��H;��H;9�H;U�H;��H;��H;u�H;��H;u�H;��H;��H;U�H;;�H;��H;��H;Q�H;��H;��H;̼H;�H;��H;��H;Q�H;jH;�NH;�-H;�H;��G;�cG;3�F;��E;?�D;j�B;$@;P�<;�8;'4;x/;[�);��$;�z ;;��;      ]�:���:��:V��:�;�Y;�';��;��(;��0;�Y7;T�<;�@;aC;1CE;�wF;}8G;��G;n�G;�)H;�LH;jH;=�H;c�H;��H;ٳH;ľH;k�H;/�H;��H;�H;^�H;��H;��H;��H;��H;��H;��H;��H;��H;��H;a�H;�H;��H;,�H;m�H;ľH;۳H;��H;b�H;<�H;jH;�LH;�)H;n�G;��G;}8G;�wF;1CE;aC;�@;T�<;�Y7;��0;��(;��;�';�Y;�;V��:��:���:      ��:h�:43<:�)i:pt�:凲:j�:�+�:�Y;B�;�*';�1;:�8;�Z>;R0B;�D;�2F;)G;��G;"�G;�)H;�NH;|lH;S�H;m�H;��H;��H;5�H;��H;�H;B�H;2�H;;�H;c�H;��H;��H;��H;��H;��H;c�H;:�H;4�H;B�H;�H;��H;8�H;��H;��H;p�H;P�H;ylH;�NH;�)H;$�G;��G;.G;�2F;�D;R0B;�Z>;:�8;�1;�*';@�;�Y;�+�:j�::~t�:�)i: 3<:<�:      ���4X��� ����=��۷��ݤ8��:�P�:�P�:���:,`;{;*�*;�$5;�g<;=A;CD;F;�G;��G;l�G;�-H;!SH;_qH;�H;ǝH;��H;�H;A�H;��H;��H;��H;\�H;��H;��H;��H;��H;��H;��H;��H;\�H;��H;��H;��H;A�H;�H;��H;ɝH;�H;\qH;SH;�-H;l�G;��G;�G;F;CD;=A;�g<;�$5;*�*;};,`;���:�P�:�P�:��:`ޤ8X۷���=�� ��4X��      �1��7Ȅ��u��PV��.�����W������W�9 +i:֡�:,�:�;�t%;�J2;^;;��@;sD;F;.G;��G;�H;�5H;�ZH;;xH;F�H;2�H;�H;�H;a�H;u�H;#�H;8�H;0�H;F�H;b�H;��H;b�H;F�H;2�H;7�H;%�H;w�H;`�H;�H;�H;/�H;I�H;<xH;�ZH;�5H;�H;�G;0G;F;tD;��@;^;;�J2;�t%;�;,�:֡�:�*i:X�9���W������.��PV��u�;Ȅ�      b��R�	�������2Tʻ�R��3|�{.�8Ⱥ����X�9&u�:��:�Y;��!;��0;�:;��@;CD;�2F;8G;��G;�H;p@H;-dH;ʀH;|�H;L�H;O�H;T�H;��H;��H;��H;v�H;��H;�H;��H;�H;��H;w�H;��H;��H;��H;T�H;N�H;M�H;y�H;̀H;-dH;m@H;�H;��G;}8G;�2F;CD;��@;�:;��0;��!;�Y;��:&u�:�X�9���2Ⱥ{.�3|��R��1Tʻ������T�	�      ʪx��[t���g�[T�g�:����+���:����1��_�(�NW�� �t��n`:[��:�\;{ ;��0;a;;=A;�D;�wF;�cG;Y�G;�!H;�MH;�oH;{�H;��H;˯H;��H;m�H;��H;c�H;u�H;�H;��H;-�H;��H;�H;v�H;a�H;��H;n�H;��H;ȯH;��H;z�H;�oH;�MH;�!H;V�G;�cG;�wF;�D;	=A;b;;��0;{ ;�\;_��:�n`: �t�LW��a�(��1��9���*������h�:�[T���g��[t�      @,˼��Ǽ�"���뮼w��,G��5�[�ky-�����.����b��0��ط��4<:�L�:�\;��!;�J2;�g<;S0B;1CE;0�F;S�G;��G;�4H;�\H;|H;��H;��H;_�H;��H;G�H;��H;X�H;Z�H;�H;��H;�H;X�H;X�H;��H;K�H;��H;_�H;��H;��H;|H;�\H;�4H;��G;O�G;0�F;1CE;V0B;�g<;�J2;��!;�\;�L�:�4<:�ط��0�ޕb��.�����ky-�5�[�+G��w���뮼�"����Ǽ      0���k��Nv��t�K�Ѽ�뮼3X��x�W�����׻
Ȅ�#��P���4<:[��:�Y;�t%;�$5;�Z>;aC;��E;9*G;j�G;H;HH;slH;��H;
�H;ɯH;ؼH;��H;��H;�H;~�H;v�H;6�H;v�H;~�H;�H;��H;��H;׼H;ɯH;
�H;��H;slH;HH;H;h�G;5*G;��E;aC;�Z>;�$5;�t%;�Y;a��:�4<:P��"��	Ȅ��׻���x�W�3X���뮼J�Ѽ�t�Nv���k�      Km��Fi��&^�d�L�U�6�-����'}ռuT����x�ɻ0�Ƙ����$���ط��n`:��:�;+�*;<�8;�@;<�D;m�F;�}G;��G;�1H;�[H;u|H;ĕH;ߨH;��H;��H;��H;��H;��H;��H;{�H;��H;��H;��H;��H;��H;��H;ߨH;ÕH;u|H;�[H;�1H;��G;�}G;i�F;<�D;�@;>�8;+�*;�;��:�n`:�ط�$�����Ƙ�ɻ0���x�uT��&}ռ��-��U�6�d�L��&^��Fi�      P��x;��E�������섽�e��?��k��t�鷼#G���e7�Ƙ�
Ȅ��0㺀�t�$u�:,�:z;�1;T�<;f�B;+�E;G;��G;dH;wJH;coH;�H;��H;�H;��H;��H;%�H;��H;�H;��H;�H;��H;%�H;��H;��H;�H;��H;�H;aoH;wJH;dH;��G;G;)�E;f�B;X�<;�1;z;,�:$u�:��t��0�
Ȅ�Ƙ껍e7�#G��鷼�t��k��?��e��섽���E���x;��      u���*��s��ӽ�'��D�������Z��Q+�����"��#G��ʻ0��׻ߕb�NW���X�9ҡ�:,`;�*';�Y7;$@;+�D;��F;�G;��G;;8H;bH;�H;]�H;��H;w�H;��H;��H;��H;U�H;A�H;U�H;��H;��H;��H;z�H;��H;]�H;�H;bH;;8H;��G;�G;��F;(�D;$@;�Y7;�*';,`;֡�:�X�9RW��ޕb��׻ʻ0�#G���"������Q+��Z����D����'���ӽ�s�*��      �!,�;)��K ���������޽"������Fi��0����鷼��x�����.��b�(� ���*i:���:@�;��0;O�<;�C;��E;=G;��G;�$H;gTH;�wH;�H;�H;Q�H;��H;C�H;��H;��H;��H;��H;��H;C�H;��H;R�H;�H;�H;�wH;gTH;�$H;��G;=G;��E;�C;O�<;��0;>�;���:�*i:��b�(��.�������x�鷼����0��Fi����"����޽�������K �;)�      -�j��f��Z�}�F��>/��^�r����ŽJ ���Fi��Q+��t�vT��z�W�����1��6Ⱥ�W�9�P�:�Y;��(;
�8;�A;�E;�F;k�G;�H;�FH;�mH;��H;ġH;C�H;r�H;��H;��H;��H;��H;��H;��H;��H;p�H;D�H;ơH;��H;�mH;�FH;�H;k�G;
�F;�E;�A;
�8;��(;�Y;�P�: X�9<Ⱥ�1�����y�W�vT���t�Q+��Fi�J ���Žr����^��>/�}�F��Z��f�      ��y���{�J����f��SC��K �tn���Ž����Z��k�'}ռ3X��ky-�9���{.����P�:�+�:�;4;9�>;�D;�wF;5�G;��G;�9H;[dH;w�H;��H;f�H;t�H;��H;��H;Y�H;v�H;[�H;��H;��H;r�H;f�H;��H;w�H;XdH;�9H;��G;4�G;�wF;�D;:�>;4;��;�+�:�P�:���~.�9���ky-�3X��&}ռ�k��Z�����Žtn���K ��SC��f�J���{�y���      ��˾��Ǿ����#���X͓�^�x���J��K �r���"������?����뮼6�[�.���%3|��W��x�:f�:�';n/;fg<;�C;lF;�NG;��G;2-H;r[H;�}H;˗H;ΪH;¸H;��H;�H;��H;�H;��H;�H;��H;��H;ΪH;˗H;�}H;q[H;2-H;��G;�NG;oF;�C;dg<;n/;�';d�:x�:�W��&3|�.���6�[��뮼���?����"��r����K ���J�^�x�X͓�#���������Ǿ      v� ��������{Ծm���y���^�x��SC��^���޽D����e�-��K�Ѽ,G������R�����@ݤ8釲:�Y;P�);��9;��A;��E;�G; �G;k!H;DSH;�wH;y�H;��H;G�H;��H;}�H;��H;��H;��H;}�H;��H;D�H;��H;y�H;�wH;@SH;k!H;�G;�G;��E;��A;��9;P�);�Y;釲:`ݤ8 ����R�����,G��K�Ѽ-���e�D�����޽�^��SC�^�x�y���m����{Ծ�쾤���      ��� E�l�v� �Y�ݾm���X͓��f��>/�����'���섽U�6��t�w��h�:�2Tʻ�.�p۷�ft�:�;��$;�Y7;Y�@;�	E;�F;;�G;�H;ALH;�rH;��H;ѤH;)�H;#�H;7�H;O�H;��H;Q�H;6�H;#�H;'�H;ӤH;��H;�rH;?LH;�H;<�G;�F;�	E;V�@;�Y7;��$;�;ft�:p۷��.�3Tʻh�:�w���t�U�6��섽�'������>/��f�X͓�m���Y�ݾv� �l� E�      ��7�v3�1�'����v� ��{Ծ"���J���}�F�����ӽ���e�L�Ov��뮼\T�����PV���=��)i:\��:�z ;�$5;��?;�D;ϺF;��G;�H;�FH;�nH;��H;��H;w�H;�H;=�H;\�H;��H;\�H;=�H;�H;u�H;��H;��H;�nH;�FH;�H;��G;ϺF;�D;��?;�$5;�z ;b��:�)i:��=��PV����\T��뮼Ov�e�L�����ӽ���}�F�J���"����{Ծv� ����1�'�v3�      �N��TI���;�1�'�l��쾃���{󐾷Z��K ��s�E����&^���"����g�����u�!��3<:���: ;dg3;��>;xBD;��F;�G;�H;NBH;{kH;\�H;�H;4�H;߼H;v�H;��H;N�H;��H;v�H;�H;2�H;�H;\�H;xkH;LBH;�H;�G;��F;xBD;��>;hg3; ;��:3<:!���u������g��"����&^�E����s潨K ��Z�{󐾃�����l�1�'���;��TI�      c]�g�W��TI�v3� E�������Ǿy����f�;)�*��x;���Fi��k���Ǽ�[t�U�	�8Ȅ�4X���:���:��;WJ2;OZ>;H	D;~F;D�G;H;�?H;�iH;��H;�H;|�H;A�H;��H;`�H;��H;`�H;��H;A�H;z�H;�H;��H;�iH;�?H;H;C�G;~F;H	D;KZ>;]J2;��;���:�:4X��8Ȅ�U�	��[t���Ǽ�k��Fi�x;��*��;)��f�y�����Ǿ���� E�v3��TI�g�W�      4�$��� ����%��C��+�þ�*��6Dx���=�����Pν���+'K��c�(��}�V����/E^���S��w[:���:e;T�4;@`?;�mD;��F;TvG;;�G;{H;OH;�sH;�H;��H;��H;"�H;|�H;P�H;|�H;"�H;��H;��H;�H;�sH;}OH;xH;;�G;TvG;��F;�mD;<`?;W�4;e;���:�w[:��S�-E^����}�V�(���c�+'K�����Pν�����=�6Dx��*��+�þC��%������� �      �� ����T��P��3������0��9�s�ۀ:�j9�"�ʽ6Z���G��8�.���5S����0X���D��Bd:�B�: ;�4;È?;�~D;K�F;yG;��G;� H;FPH;EtH;>�H;��H;��H;`�H;��H;b�H;��H;b�H;��H;��H;A�H;EtH;CPH;� H;��G;yG;J�F;�~D;��?;!�4; ;�B�:�Bd:��D�0X���껻5S�.���8��G�6Z��"�ʽj9�ۀ:�9�s��0�����3��Q��T�����      ���T��;�
������Yؾ"���ᥒ���f���0�^[�T8��Ԑ����>�����TȤ��6H�r�ܻ$rF����L�}:҆�:c";U�5;��?;x�D;֮F;�G;��G;k#H;~RH;�uH;��H;�H;��H;��H;�H;��H;�H;��H;��H;�H;��H;�uH;{RH;h#H;��G;�G;ӮF;x�D;��?;X�5;c";҆�:D�}:���"rF�s�ܻ�6H�TȤ�������>�Ԑ��T8��^[���0���f�ᥒ�"����Yؾ����;�
�T��      %��Q������AI�+�þ S��>���xS��Q"��s������}��0� 켑�����6�V�ƻR}*�p�����:ox;[%;�l7;ڳ@;��D;��F;��G;��G;.(H;VH;�xH;��H;q�H;βH;�H;��H;��H;��H;�H;ϲH;p�H;��H;�xH;VH;*(H;��G;��G;��F;��D;ճ@;�l7;[%;ox;��:x���P}*�W�ƻ��6����� ��0���}�����s��Q"�xS�>��� S��+�þAIᾧ���Q��      C��3�很Yؾ+�þĪ�~쏾�k�ۀ:�����ؽ�����c�cy���Ҽ���O� �v�D�� (7e�:��
;��(;�_9;��A;�\E;��F;͝G;��G;�.H;�ZH;|H;!�H;u�H;��H;@�H;�H;��H;�H;?�H;��H;t�H;#�H;|H;�ZH;�.H;��G;ϝG;��F;�\E;��A;�_9;��(;��
;_�: (7B��v�N� ������Ҽcy��c�������ؽ��ۀ:��k�~쏾Ī�+�þ�Yؾ3��      *�þ���"����R��~쏾:�s��H�����������Ӑ����D��c�����L�f�],�����P���9��:�;+j-;t�;;|�B;�E;�G;��G;��G;�6H;�`H;��H;��H;��H;~�H;վH;}�H;�H;}�H;վH;�H;��H;��H;��H;�`H;�6H;��G;��G;�G;�E;x�B;t�;;+j-;�;��:�9�P�����],�L�f������c���D�Ӑ�������������H�:�s�~쏾�R��"������      �*���0��॒�>����k��H��#%�][��Pνt��h�f�9/%���伎�����=��?ػ�FL���D�R�R:�:1�;?2;��=;ǚC;�0F;zGG;��G;LH;@H;�gH;��H;a�H;ڬH;øH;��H;�H;��H;�H;��H;øH;ڬH;b�H;��H;�gH;@H;JH;��G;zGG;�0F;ÚC;��=;>2;1�;�:N�R:��D��FL��?ػ��=��������9/%�h�f�t���Pν^[��#%��H��k�>���ᥒ��0��      6Dx�9�s���f�xS�ڀ:����][��7ս�榽��}���;��8�^�����r����IG�����ά�#��:�;�}$;҄6;#�?;�D;�F;�pG;��G;H;UJH;`oH;m�H;��H;*�H;h�H;��H;��H;W�H;��H;��H;h�H;)�H;��H;m�H;`oH;RJH;H;��G;�pG;�F; �D;#�?;҄6;�}$;�;!��:�ά���IG�������r�^����8���;���}��榽�7ս][����ۀ:�xS���f�9�s�      ��=�ۀ:���0��Q"��������Pν�榽D���G�7����Ҽ ��VE:�N�ܻ�D^�и��<i:D��:�;?|,;��:;t�A;ViE;��F;I�G;��G;�(H;eUH;�wH;��H;W�H;��H;$�H;�H;��H;D�H;��H;�H;"�H;��H;X�H;��H;�wH;bUH;�(H;��G;I�G;��F;RiE;q�A;��:;@|,;�;D��:<i:θ���D^�N�ܻVE:� ����Ҽ7���G�D���榽�Pν�������Q"���0�ۀ:�      ���j9�^[��s��ؽ���t����}��G������8c��c�V�P,��*�����P����:��:g ;o�3;�0>;�C;�F;9G;]�G;�H;8H;�`H;-�H;�H;+�H;v�H;�H;{�H;�H;E�H;�H;{�H;�H;t�H;.�H;�H;-�H;�`H;8H;�H;]�G;9G;�F;�C;�0>;m�3;f ;��:��:p������*��P,�c�V�8c��������G���}�t�������ؽ�s�^[�j9�      �Pν"�ʽT8���������Ӑ��h�f���;�7�����KȤ�A�f�3��^ߵ�mo5��D�.�-:?��:�>;�+;�_9;�A;��D;>�F;�vG;�G;CH;�GH;�lH;�H;ĞH;%�H;Z�H;&�H;��H;4�H;X�H;4�H;��H;%�H;Y�H;(�H;ĞH;�H;�lH;�GH;BH;�G;�vG;9�F;��D;�A;�_9;�+;�>;C��:&�-:�D�no5�]ߵ�3��A�f�KȤ����7����;�h�f�Ӑ���������T8��"�ʽ      
���6Z��Ӑ����}��c���D�9/%��8���Ҽ8c��@�f����'�ƻ�/X�|���P��9	�:;�;�";��3;N>;_YC;��E;�G;�G;��G;�,H;0WH;BxH;��H;b�H;�H;@�H;�H;d�H;r�H;b�H;r�H;e�H;�H;@�H;�H;b�H;��H;AxH;0WH;�,H;��G;�G;�G;��E;_YC;N>;��3;�";>�;�:P��9|����/X�'�ƻ���@�f�7c����Ҽ�8�9/%���D��c���}�Ӑ��6Z��      +'K��G���>��0�cy��c����^��� ��c�V�2��'�ƻ�od���º t(7�4�:���:��;�P.;�:;'zA;L�D;�F;rnG;h�G;H;�@H;RfH;��H;[�H;�H;�H;�H;�H;��H;��H;n�H;��H;��H;�H;�H;�H;�H;[�H;��H;QfH;�@H;H;d�G;lnG;�F;L�D;'zA;�:;�P.;��;���:�4�: t(7��º�od�(�ƻ2��c�V� ��^�����伛c�dy��0���>��G�      �c��8���������Ҽ����������r�UE:�O,�[ߵ��/X���º@Ȭ�\�}:�:�;O�);8m7;/�?;��C;&F;�)G;8�G;u�G;2*H;�SH;�tH;��H;��H;"�H;޽H;��H;�H;C�H;��H;��H;��H;C�H;�H;��H;�H;"�H;��H;��H;�tH;�SH;2*H;t�G;4�G;})G;&F;��C;-�?;8m7;Q�);�;�:`�}: Ȭ���º�/X�[ߵ�N,�TE:���r�����������Ҽ�������8�      (��.��SȤ��������K�f���=����N�ܻ�*��mo5�|��� t(7\�}:�n�:0�;�>&;��4;��=;��B;�E;4�F;��G;�G;]H;�AH;�eH;m�H;	�H;��H;�H;��H;T�H;��H;��H;��H;��H;��H;��H;��H;R�H;��H;�H;��H;�H;m�H;�eH;�AH;ZH;�G;��G;4�F;�E;��B;��=;��4;�>&;0�;�n�:X�}: t(7|���mo5��*��N�ܻ�����=�J�f��������SȤ�.��      {�V��5S��6H���6�N� �^,��?ػJG���D^�����D�P��9�4�:�:2�;�%;��3;,�<;pB;�E; �F;�XG;-�G;r H;�0H;�WH;�vH;!�H;��H;�H;ĽH;��H;��H;��H;��H;��H;n�H;��H;��H;��H;��H;��H;��H;�H;��H;!�H;�vH;WH;�0H;l H;)�G;�XG;�F;�E;pB;,�<;��3;�%;2�;�:�4�:P��9�D�����D^�KG���?ػ],�N� ���6��6H��5S�      ��ﻹ��q�ܻV�ƻv�����FL���̸�� ��6�-:	�:���:�;�>&;��3;h9<;'�A;��D;iZF;E5G;$�G;�G;�!H;bJH;akH;ԅH;�H;��H;͸H;�H;��H;��H;�H;��H;��H;'�H;��H;��H;�H;��H;��H;�H;ʸH;��H;�H;ЅH;akH;_JH;�!H;�G;$�G;B5G;iZF;��D;(�A;h9<;��3;�>&;�;���:	�:.�-: ��ȸ�����FL����u�V�ƻq�ܻ���      0E^�0X�rF�M}*�D��Q����D��ά�@i:��:G��:<�;��;N�);��4;)�<;%�A;:�D;�9F;�G;��G;n�G;iH;H?H;�aH;D}H;��H;��H;˳H;�H;��H;��H;��H;O�H;��H;V�H;��H;V�H;��H;N�H;��H;��H;��H;�H;ȳH;��H;��H;F}H;�aH;B?H;eH;n�G;��G;�G;�9F;;�D;$�A;(�<;��4;O�);��;>�;G��:��:Li: Ϭ���D�Q��>��L}*�rF�$0X�      ��S���D�̖�h��� (7 �9j�R:!��:J��: ��:�>;�";�P.;9m7;��=;nB;��D;�9F;CG;F�G;��G;�H;�6H;�YH;vH;Q�H; �H;2�H;4�H;��H;V�H;��H;M�H;j�H;��H;��H;*�H;��H;��H;j�H;K�H;��H;T�H;��H;0�H;/�H;�H;S�H;vH;�YH;�6H;�H;}�G;G�G;AG;�9F;��D;mB;��=;8m7;�P.;�";�>; ��:P��:��:n�R:X�9 (7`���̖���D�      �w[:�Bd:X�}:��:c�:��:�:�;�;h ;�+;��3;�:;(�?;��B;�E;dZF;�G;C�G;��G;mH;�1H;TH;�pH;�H;}�H;�H;��H;��H;��H;1�H;��H;��H;U�H;(�H;H�H;��H;H�H;(�H;S�H;��H;��H;1�H;��H;��H;��H;�H;|�H;�H;�pH;�SH;�1H;iH;��G;C�G;�G;dZF;�E;��B;(�?;�:;��3;�+;g ;�;�;�:��:w�:��:X�}:�Bd:      ���:�B�:���:hx;��
;�;5�;�}$;?|,;p�3;�_9;M>;%zA;��C;�E;�F;C5G;��G;��G;oH;�/H;!QH;4mH;}�H;ϗH;ƧH;��H;/�H;��H;K�H;��H;��H;��H;�H;��H;x�H;��H;x�H;��H;�H;��H;��H;��H;H�H;��H;-�H;��H;ŧH;͗H;y�H;1mH; QH;�/H;oH;��G;��G;@5G;�F;�E;��C;%zA;M>;�_9;o�3;B|,;�}$;5�;�;��
;kx;܆�:�B�:      e;$ ;u";V%;��(;5j-;L2;ۄ6;ġ:;�0>;�A;_YC;L�D;'F;5�F;�XG;"�G;p�G;�H;�1H; QH;�kH;��H;��H;j�H;b�H;�H;��H;��H;C�H;��H;�H;��H;��H;��H;��H;��H;��H;��H;��H;��H;�H;��H;?�H;��H;��H;�H;b�H;i�H;��H;��H;�kH;QH;�1H;�H;p�G;"�G;�XG;7�F;&F;N�D;_YC;�A;�0>;ǡ:;ڄ6;I2;6j-;�(;V%;t"; ;      `�4;!�4;X�5;�l7;�_9;v�;;��=;&�?;t�A;�C;��D;��E;�F;�)G;��G;+�G;
�G;kH;�6H;TH;4mH;��H;�H;<�H;�H;��H;[�H;g�H;�H;��H;L�H; �H;i�H;��H;��H;��H;��H;��H;��H;��H;f�H; �H;L�H;��H;�H;g�H;W�H;��H;�H;:�H;ޔH;��H;/mH;TH;�6H;kH;
�G;)�G;��G;�)G;�F;��E;��D;�C;u�A;$�?;��=;x�;;�_9;�l7;[�5;�4;      U`?;ψ?;��?;س@;��A;y�B;КC;�D;ViE;�F;;�F;�G;mnG;7�G;�G;o H;�!H;I?H;�YH;�pH;y�H;��H;<�H;w�H;úH;^�H;z�H;;�H;��H;��H;��H;��H;��H;�H;��H;m�H;��H;j�H;��H;�H;��H;��H;��H;��H;��H;;�H;w�H;]�H;úH;u�H;8�H;��H;v�H;�pH;�YH;H?H;�!H;o H;�G;7�G;lnG;�G;;�F;�F;ViE;�D;ΚC;{�B;��A;ڳ@;��?;ň?;      �mD;�~D;h�D;��D;�\E;	�E;�0F;�F;��F;	9G;�vG;�G;g�G;x�G;]H;�0H;fJH;�aH;vH;�H;ӗH;o�H;��H;˺H;!�H;��H;��H;F�H;�H;/�H;��H;u�H;��H;�H;��H;�H;`�H;�H;��H;�H;��H;u�H;��H;-�H;�H;F�H;��H;��H;!�H;ǺH;�H;m�H;ЗH;�H;vH;�aH;cJH;�0H;]H;w�G;f�G;�G;�vG;9G;��F;�F;�0F;	�E;�\E;��D;g�D;�~D;      ��F;Z�F;ˮF;��F;��F;�G;}GG;�pG;I�G;_�G;�G;��G;H;2*H;�AH;WH;`kH;B}H;N�H;{�H;ħH;`�H;��H;]�H;��H;k�H;��H;��H;��H;J�H;G�H;��H;��H;��H;n�H;��H;�H;��H;o�H;��H;��H;��H;E�H;G�H;��H;��H;��H;m�H;��H;Z�H;��H;_�H;��H;|�H;N�H;C}H;^kH;}WH;�AH;0*H;H;��G;�G;]�G;J�G;�pG;}GG;�G;��F;��F;ˮF;O�F;      dvG;yG;�G;��G;ѝG;��G;��G;��G;��G;�H;BH;�,H;�@H;�SH;�eH;�vH;ԅH;��H;�H;�H;��H;�H;[�H;|�H;��H;��H;��H;��H;�H;�H;��H;��H;��H;{�H;�H;[�H;[�H;[�H;
�H;y�H;��H;��H;��H;�H;�H;��H;��H;��H;��H;|�H;X�H;�H;��H;�H; �H;��H;ԅH;�vH;�eH;�SH;�@H;�,H;BH;�H;��G;��G;��G;��G;םG;��G;�G;yG;      2�G;��G;��G;��G;��G;��G;QH;H;�(H; 8H;�GH;7WH;TfH;�tH;n�H;!�H;�H;��H;/�H;��H;/�H;��H;h�H;>�H;B�H;��H;��H;��H;��H;��H;��H;��H;��H;�H;��H;��H;��H;��H;��H;�H;��H;��H;��H;��H;��H;��H;��H;��H;C�H;?�H;g�H;��H;*�H;��H;-�H;��H;�H;"�H;n�H;�tH;RfH;7WH;�GH; 8H;�(H;H;QH;��G;��G;��G;��G;��G;      �H;� H;k#H;3(H;�.H;�6H;@H;XJH;hUH;�`H;�lH;FxH;��H;��H;�H;��H;��H;ɳH;4�H;��H;��H;��H;�H;��H;�H;��H;�H;��H;k�H;��H;��H;��H;&�H;��H;��H;	�H;(�H;	�H;��H;��H;#�H;��H;��H;��H;h�H;��H;�H;��H;�H;��H;�H;��H;��H;��H;3�H;ȳH;��H;��H;	�H;��H;��H;ExH;�lH;�`H;jUH;XJH;@H;�6H;�.H;3(H;k#H;� H;      �OH;OPH;�RH;VH;�ZH;�`H;�gH;hoH;�wH;5�H;�H;ƑH;b�H;��H;��H;�H;иH;�H;��H;��H;K�H;@�H;��H;��H;%�H;G�H;�H;��H;��H;��H;��H;#�H;��H;�H;5�H;X�H;m�H;X�H;5�H;�H;��H;#�H;��H;��H;��H;��H;
�H;C�H;&�H;��H;��H;@�H;J�H;��H;��H;�H;θH;�H;��H;��H;b�H;đH;�H;5�H;�wH;joH;�gH;�`H;�ZH;VH;�RH;LPH;      �sH;XtH;�uH;�xH;)|H;��H;��H;v�H;��H;#�H;˞H;o�H;�H;)�H;�H;˽H;"�H;��H;W�H;8�H;��H;��H;L�H;��H;��H;H�H;��H;��H;��H;��H;�H;��H; �H;I�H;��H;��H;��H;��H;��H;I�H;��H;��H;�H;��H;��H;��H;��H;E�H;��H;��H;G�H;��H;��H;8�H;W�H;��H;!�H;ʽH;�H;(�H;�H;m�H;˞H;%�H;��H;u�H;��H;��H;&|H;�xH;�uH;XtH;      ��H;K�H;��H;��H;(�H;��H;g�H;��H;\�H;.�H;-�H;#�H;	�H;�H;��H;�H;��H;��H;��H;�H;��H;�H;"�H;��H;q�H;��H;��H;��H;��H;%�H;��H;�H;D�H;��H;��H;��H;��H;��H;��H;��H;B�H;�H;��H;&�H;��H;��H;��H;��H;r�H;��H;�H;�H;��H;�H;��H;��H;��H;�H;��H;�H;	�H;%�H;-�H;.�H;^�H;��H;g�H;��H;&�H;��H;��H;G�H;      ��H;�H;��H;z�H;�H;�H;ݬH;5�H;ȳH;x�H;]�H;I�H;�H;��H;V�H;��H;��H;��H;N�H;��H;��H;��H;j�H;��H;��H;��H;��H;��H;*�H;��H;�H;I�H;��H;��H;��H;��H;�H;��H;��H;��H;��H;J�H;�H;��H;,�H;��H;��H;��H;��H;��H;g�H;��H;��H;��H;N�H;��H;��H;��H;U�H;��H;�H;H�H;]�H;y�H;ȳH;3�H;ެH;�H;v�H;z�H;��H;��H;      ��H;�H;��H;ղH;��H;~�H;̸H;t�H;+�H;�H;-�H;%�H;!�H;�H;��H;��H;�H;N�H;m�H;]�H;�H;��H;��H;�H;�H;��H;v�H;�H;��H;�H;F�H;��H;��H;��H;��H;��H;�H;��H;��H;��H;��H;��H;D�H;�H;��H;�H;v�H;��H;�H;�H;��H;��H;�H;]�H;m�H;O�H;�H;��H;��H;�H;!�H;%�H;,�H;�H;,�H;r�H;̸H;��H;��H;ֲH;��H;��H;      $�H;x�H;�H;�H;\�H;ӾH;��H;��H;�H;�H;��H;p�H;��H;J�H;��H;��H;��H;��H;��H;1�H;��H;��H;��H;��H;��H;m�H;�H;��H;��H;9�H;��H;��H;��H;��H;�H;�H;�H;�H;�H;��H;��H;��H;��H;8�H;��H;��H;�H;m�H;��H;��H;��H;��H;��H;1�H;��H;��H;��H;��H;��H;J�H;��H;p�H;��H;��H;�H;��H;��H;ؾH;Q�H;�H;�H;p�H;      {�H;��H;'�H;��H;!�H;{�H;*�H;��H;��H;�H;<�H;}�H;��H;��H;��H;��H;��H;P�H;��H;T�H;��H;��H;��H;p�H;�H;��H;Z�H;��H;�H;[�H;��H;��H;��H;�H;�H;+�H;"�H;+�H;�H;��H;��H;��H;��H;[�H;�H;��H;X�H;��H;�H;n�H;��H;��H;��H;R�H;��H;R�H;��H;��H;��H;��H;��H;}�H;<�H;	�H;��H;��H;*�H;��H;�H;��H;)�H;��H;      U�H;l�H;��H;��H;��H;�H;��H;`�H;N�H;F�H;`�H;n�H;r�H;��H;��H;u�H;.�H;��H;-�H;��H;��H;��H;��H;��H;Z�H;�H;Z�H;��H;*�H;v�H;��H;��H;�H;	�H;�H;$�H;.�H;$�H;�H;	�H;�H;��H;��H;v�H;-�H;��H;X�H;�H;Z�H;��H;��H;��H;��H;��H;-�H;��H;,�H;u�H;��H;��H;r�H;n�H;`�H;I�H;O�H;]�H;��H;�H;��H;��H;��H;b�H;      {�H;��H;'�H;��H;!�H;|�H;*�H;��H;��H;�H;<�H;}�H;��H;��H;��H;��H;��H;P�H;��H;R�H;��H;��H;��H;p�H;�H;��H;Z�H;��H;�H;Z�H;��H;��H;��H;�H;�H;+�H;"�H;+�H;�H;��H;��H;��H;��H;\�H;�H;��H;X�H;��H;�H;p�H;��H;��H;��H;T�H;��H;R�H;��H;��H;��H;��H;��H;}�H;=�H;	�H;��H;��H;+�H;��H;�H;��H;&�H;��H;      "�H;x�H;�H;�H;\�H;ӾH;��H;��H;�H;�H;��H;p�H;��H;J�H;��H;��H;��H;��H;��H;1�H;��H;��H;��H;��H;��H;m�H;�H;��H;��H;8�H;��H;��H;��H;��H;�H;�H;�H;�H;�H;��H;��H;��H;��H;;�H;��H;��H;�H;n�H;��H;��H;��H;��H;��H;1�H;��H;��H;��H;��H;��H;J�H;��H;p�H;��H;��H;�H;��H;��H;ؾH;Q�H;�H;�H;n�H;      °H;�H;��H;ֲH;��H;~�H;̸H;t�H;+�H;�H;-�H;%�H;!�H;�H;��H;��H;�H;N�H;m�H;\�H;!�H;��H;��H;�H;�H;��H;v�H;�H;��H;�H;D�H;��H;��H;��H;��H;��H;�H;��H;��H;��H;��H;��H;F�H;�H;��H;�H;v�H;��H;�H;�H;��H;��H;�H;]�H;m�H;P�H;�H;��H;��H;�H;!�H;%�H;-�H;�H;,�H;r�H;̸H;��H;��H;ղH;��H;��H;      ��H;�H;��H;{�H;}�H;�H;ެH;4�H;ȳH;x�H;]�H;H�H;�H;��H;U�H;��H;��H;��H;N�H;��H;��H;��H;i�H;��H;��H;��H;��H;��H;*�H;��H;�H;I�H;��H;��H;��H;��H;�H;��H;��H;��H;��H;L�H;�H;��H;,�H;��H;��H;��H;��H;��H;i�H;��H;��H;��H;N�H;��H;��H;��H;V�H;��H;�H;I�H;]�H;y�H;ȳH;1�H;ݬH;�H;u�H;{�H;��H;�H;      ��H;K�H;��H;��H;(�H;��H;i�H;��H;\�H;/�H;-�H;#�H;	�H;�H;��H;�H;��H;��H;��H;�H;��H;�H;"�H;��H;r�H;��H;��H;��H;��H;%�H;��H;�H;C�H;��H;��H;��H;��H;��H;��H;��H;B�H;�H;��H;&�H;��H;��H;��H;��H;q�H;��H; �H;�H;��H;�H;��H;��H;��H;�H;��H;�H;	�H;%�H;-�H;/�H;^�H;��H;i�H;��H;$�H;��H;��H;G�H;      �sH;XtH;�uH;�xH;)|H;��H;��H;v�H;��H;#�H;˞H;m�H;�H;)�H;�H;˽H;!�H;��H;W�H;8�H;��H;��H;L�H;��H;��H;G�H;��H;��H;��H;��H;�H;��H;��H;I�H;��H;��H;��H;��H;��H;I�H;��H;��H;�H;��H;��H;��H;��H;G�H;��H;��H;I�H;��H;��H;8�H;W�H;��H;!�H;˽H;�H;)�H;�H;o�H;ʞH;%�H;��H;v�H;��H;��H;&|H;�xH;�uH;WtH;      �OH;MPH;�RH;VH;�ZH;�`H;�gH;koH;�wH;4�H;�H;đH;b�H;��H;��H;�H;иH;�H;��H;��H;N�H;@�H;��H;��H;&�H;D�H;�H;��H;��H;��H;��H;#�H;��H;�H;5�H;X�H;m�H;X�H;5�H;�H;��H;%�H;��H;��H;��H;��H;�H;F�H;%�H;��H;��H;@�H;J�H;��H;��H;�H;θH;��H;��H;��H;b�H;ƑH;�H;4�H;�wH;koH;�gH;�`H;�ZH;VH;�RH;MPH;      �H;� H;r#H;1(H;�.H;�6H;@H;YJH;hUH;�`H;�lH;FxH;��H;��H;	�H;��H;��H;ƳH;3�H;��H;��H;��H;�H;��H;�H;��H;�H;��H;h�H;��H;��H;��H;%�H;��H;��H;	�H;(�H;	�H;��H;��H;%�H;��H;��H;��H;i�H;��H;�H;��H;�H;��H;�H;��H;��H;��H;4�H;˳H;��H;��H;�H;��H;��H;FxH;�lH;�`H;iUH;XJH;@H;�6H;�.H;.(H;r#H;� H;      2�G;��G;��G;��G;��G;��G;QH;H;�(H; 8H;�GH;7WH;RfH;�tH;n�H;"�H;�H;��H;-�H;��H;0�H;��H;h�H;>�H;C�H;��H;��H;��H;��H;��H;��H;��H;��H;�H;��H;��H;��H;��H;��H;�H;��H;��H;��H;��H;��H;��H;��H;��H;B�H;?�H;g�H;��H;-�H;��H;/�H;��H;�H;"�H;n�H;�tH;TfH;7WH;�GH; 8H;�(H;H;QH;��G;��G;��G;��G;��G;      ^vG;yG;�G;��G;НG;��G;��G;��G;��G;�H;BH;�,H;�@H;�SH;�eH;�vH;ԅH;��H; �H;�H;��H;�H;Z�H;|�H;��H;��H;��H;��H;�H;�H;��H;��H;��H;y�H;
�H;[�H;[�H;Z�H;�H;y�H;��H;��H;��H;�H;�H;��H;��H;��H;��H;|�H;Z�H;�H;��H;�H;�H;��H;҅H;�vH;�eH;�SH;�@H;�,H;CH;�H;��G;��G;��G;��G;ӝG;��G;�G;yG;      ��F;V�F;ծF;��F;��F;�G;{GG;�pG;I�G;_�G;�G;��G;H;0*H;�AH;WH;`kH;B}H;N�H;{�H;ħH;_�H;��H;Z�H;��H;k�H;��H;��H;��H;I�H;E�H;��H;��H;��H;m�H;��H;�H;��H;o�H;��H;��H;��H;G�H;G�H;��H;��H;��H;m�H;��H;\�H;��H;`�H;��H;{�H;N�H;C}H;^kH;WH;�AH;2*H;H;��G;�G;]�G;I�G;�pG;}GG;�G;��F;��F;ծF;L�F;      �mD;�~D;g�D;��D;�\E;	�E;�0F;�F;��F;	9G;�vG;�G;f�G;w�G;]H;�0H;cJH;�aH;vH;�H;ӗH;m�H;��H;ȺH;!�H;��H;��H;F�H;�H;/�H;��H;t�H;��H;�H;��H;�H;`�H;�H;��H;�H;��H;x�H;��H;-�H;�H;F�H;��H;��H;!�H;ʺH;��H;o�H;җH;�H;vH;�aH;cJH;�0H;]H;w�G;g�G;�G;�vG;9G;��F;�F;�0F;�E;�\E;��D;g�D;�~D;      Z`?;͈?;�?;׳@;��A;~�B;̚C;�D;WiE; F;=�F;�G;mnG;7�G;�G;o H;�!H;E?H;�YH;�pH;z�H;��H;;�H;v�H;úH;\�H;x�H;;�H;��H;��H;��H;��H;��H;�H;��H;k�H;��H;k�H;��H;�H;��H;��H;��H;��H;��H;;�H;x�H;^�H;úH;w�H;:�H;��H;v�H;�pH;�YH;K?H;�!H;o H;�G;7�G;mnG;�G;:�F;�F;WiE;�D;̚C;�B;ƘA;׳@;�?;?;      Y�4;,�4;j�5;�l7;�_9;z�;;��=;&�?;u�A;�C;��D;��E;�F;�)G;��G;*�G;
�G;gH;�6H;TH;5mH;��H;�H;;�H;�H;��H;Z�H;g�H;�H;��H;L�H; �H;i�H;��H;��H;��H;��H;��H;��H;��H;g�H; �H;L�H;��H;�H;g�H;Z�H;��H;�H;;�H;ޔH;��H;/mH;TH;�6H;lH;
�G;+�G;��G;�)G;�F;��E;��D;�C;u�A;$�?;��=;|�;;�_9;�l7;_�5;�4;      e;" ;u";V%;��(;5j-;I2;ۄ6;ġ:;�0>;�A;_YC;N�D;'F;5�F;�XG;!�G;n�G;�H;�1H; QH;�kH;��H;��H;i�H;`�H;�H;��H;��H;C�H;��H;�H;��H;��H;��H;��H;��H;��H;��H;��H;��H;�H;��H;?�H;��H;��H;	�H;c�H;j�H;��H;��H;�kH; QH;�1H;�H;q�G;!�G;�XG;7�F;&F;L�D;`YC;�A;�0>;ǡ:;ۄ6;L2;5j-;�(;V%;t"; ;      ���:�B�:��:kx;��
;�;8�;�}$;?|,;o�3;�_9;M>;%zA;��C;�E;�F;B5G;��G;��G;mH;�/H; QH;2mH;|�H;͗H;ħH;��H;-�H;��H;K�H;��H;��H;��H;�H;��H;x�H;��H;x�H;��H;�H;��H;��H;��H;H�H;��H;/�H;��H;ƧH;ϗH;y�H;2mH;!QH;�/H;pH;��G;��G;B5G;�F;�E;��C;%zA;M>;�_9;m�3;@|,;�}$;9�;�;��
;ix;��:�B�:      �w[:�Bd:l�}:��:k�:��:�:�;�;h ;�+;��3;�:;(�?;��B;�E;dZF;�G;C�G;��G;mH;�1H;TH;�pH;�H;{�H;�H;��H;��H;��H;1�H;��H;��H;S�H;(�H;J�H;��H;J�H;(�H;U�H;��H;��H;1�H;��H;��H;��H;�H;}�H;�H;�pH; TH;�1H;lH;��G;C�G;�G;dZF;�E;��B;(�?;�:;��3;�+;h ;�;�;�:��:y�:��:\�}:�Bd:      ��S���D�̖�`��� (7 �9n�R:!��:J��: ��:�>;�";�P.;8m7;��=;mB;��D;�9F;AG;F�G;��G;�H;�6H;�YH;vH;P�H;�H;/�H;3�H;��H;T�H;��H;M�H;j�H;��H;��H;*�H;��H;��H;j�H;K�H;��H;V�H;��H;2�H;2�H;�H;S�H;vH;�YH;�6H;�H;}�G;G�G;CG;�9F;��D;nB; �=;8m7;�P.;�";�>; ��:N��:!��:j�R:`�9 (7h���̖���D�      .E^�0X�rF�M}*�F��Q����D��ά�@i:��:E��:>�;��;N�);��4;(�<;%�A;:�D;�9F;�G;��G;n�G;hH;G?H;�aH;C}H;��H;��H;ɳH;�H;��H;��H;��H;N�H;��H;V�H;��H;V�H;��H;O�H;��H;��H;��H;�H;ȳH;��H;��H;F}H;�aH;D?H;gH;n�G;��G;�G;�9F;;�D;$�A;)�<;��4;N�);��;<�;G��:��:Li: Ϭ���D�Q��?��N}*�rF�$0X�      ��ﻺ��r�ܻW�ƻv�����FL���̸�� ��2�-:	�:���:�;�>&;��3;h9<;%�A;��D;iZF;B5G;$�G;�G;�!H;_JH;`kH;ԅH;�H;��H;͸H;�H;��H;��H;�H;��H;��H;'�H;��H;��H;�H;��H;��H;�H;̸H;��H;�H;ЅH;ckH;bJH;�!H;�G;$�G;C5G;jZF;��D;(�A;h9<;��3;�>&;�;���:	�:2�-:@��ȸ�����FL����u�V�ƻq�ܻ���      |�V��5S��6H���6�N� �^,��?ػJG���D^�����D�P��9�4�:�:2�;�%;��3;*�<;pB;�E;�F;�XG;+�G;p H;�0H;}WH;�vH;!�H;��H;�H;��H;��H;��H;��H;��H;��H;n�H;��H;��H;��H;��H;��H;ĽH;�H;��H;!�H;�vH;�WH;�0H;m H;)�G;�XG;�F;�E;pB;-�<;��3;�%;3�;�:�4�:P��9�D�����D^�JG���?ػ\,�N� ���6��6H��5S�      (��.��SȤ��������K�f���=����O�ܻ�*��no5�|��� t(7X�}:�n�:0�;�>&;��4;��=;��B;�E;4�F;��G;�G;ZH;�AH;�eH;m�H;�H;��H;�H;��H;U�H;��H;��H;��H;��H;��H;��H;��H;T�H;��H;�H;��H;�H;m�H;�eH;�AH;]H;�G;��G;4�F;�E;��B;��=;��4;�>&;0�;�n�:X�}: t(7|���mo5��*��N�ܻ�����=�J�f��������SȤ�.��      �c��8���������Ҽ����������r�UE:�N,�[ߵ��/X���º`Ȭ�`�}:�:�;O�);8m7;+�?;��C;&F;�)G;7�G;t�G;0*H;�SH;�tH;��H;��H;"�H;޽H;��H;�H;C�H;��H;��H;��H;C�H;�H;��H;߽H;"�H;��H;��H;�tH;�SH;2*H;u�G;5�G;})G;&F;��C;-�?;8m7;R�);�;�:\�}:`Ȭ���º�/X�[ߵ�N,�TE:���r�����������Ҽ�������8�      +'K��G���>��0�cy��c����^��� ��c�V�3��(�ƻ�od���º t(7�4�:���:��;�P.;�:;%zA;L�D;�F;rnG;d�G;H;�@H;QfH;��H;[�H;�H;�H;�H;�H;��H;��H;n�H;��H;��H;�H;�H;�H;�H;[�H;��H;QfH;�@H; H;h�G;knG;�F;L�D;'zA;�:;�P.;��;���:�4�: u(7��º�od�'�ƻ2��c�V� ��^�����会c�cy��0���>��G�      ���6Z��Ӑ����}��c���D�9/%��8���Ҽ7c��@�f����(�ƻ�/X�z���P��9�:<�;�";��3;K>;_YC;��E;�G;�G;��G;�,H;0WH;BxH;��H;b�H;�H;A�H;�H;e�H;t�H;b�H;t�H;d�H;�H;>�H;�H;b�H;��H;AxH;0WH;�,H;��G;�G;�G;��E;_YC;O>;��3;�";>�;�:@��9z����/X�'�ƻ���@�f�7c����Ҽ�8�9/%���D��c���}�Ӑ��6Z��      �Pν"�ʽT8���������Ӑ��h�f���;�7�����KȤ�A�f�3��^ߵ�no5��D�*�-:A��:�>;�+;�_9;�A;��D;>�F;�vG;�G;CH;�GH;�lH;�H;ĞH;%�H;Z�H;%�H;��H;4�H;X�H;4�H;��H;&�H;Y�H;&�H;ĞH;�H;�lH;�GH;BH;�G;�vG;9�F;��D;�A;�_9;�+;�>;E��:&�-:�D�mo5�^ߵ�3��A�f�KȤ����7����;�h�f�Ӑ���������T8��"�ʽ      ���j9�^[��s��ؽ���t����}��G������8c��c�V�P,��*�����`����:��:g ;l�3;�0>;�C;�F;9G;]�G;�H;8H;�`H;-�H;�H;+�H;v�H;�H;{�H;�H;E�H;�H;{�H;�H;u�H;,�H;�H;-�H;�`H;8H;�H;]�G;9G;�F;�C;�0>;o�3;f ;��:��:p������*��P,�c�V�8c��������G���}�t�������ؽ�s�^[�j9�      ��=�ۀ:���0��Q"��������Pν�榽D���G�7����Ҽ ��VE:�N�ܻ�D^�̸��8i:D��:�;>|,;��:;s�A;ViE;��F;I�G;��G;�(H;eUH;�wH;��H;W�H;³H;"�H;�H;��H;D�H;��H;�H;$�H;��H;W�H;��H;�wH;bUH;�(H;��G;I�G;��F;RiE;s�A;��:;@|,;�;D��:@i:Ҹ���D^�N�ܻVE:� ����Ҽ7���G�D���榽�Pν�������Q"���0�ۀ:�      6Dx�9�s���f�xS�ڀ:����^[��7ս�榽��}���;��8�^�����r����IG�����ά�!��:�;�}$;҄6;#�?;�D;�F;�pG;��G;H;UJH;`oH;m�H;��H;*�H;j�H;��H;��H;W�H;��H;��H;j�H;)�H;��H;m�H;`oH;RJH;H;��G;�pG;�F; �D;#�?;҄6;�}$;�;#��:�ά���IG�������r�^����8���;���}��榽�7ս^[����ڀ:�xS���f�9�s�      �*���0��॒�>����k��H��#%�^[��Pνt��h�f�9/%���伎�����=��?ػ�FL���D�N�R:�:.�;>2;��=;ǚC;�0F;zGG;��G;JH;@H;�gH;��H;a�H;۬H;ŸH;��H;�H;��H;�H;��H;øH;جH;a�H;��H;�gH;@H;LH;��G;zGG;�0F;ŚC;��=;?2;2�;�:R�R:��D��FL��?ػ��=��������9/%�h�f�t���Pν^[��#%��H��k�>���॒��0��      *�þ���"����R��~쏾:�s��H�����������Ӑ����D��c�����L�f�],�����P���9��:�;+j-;r�;;|�B;�E;�G;��G;��G;�6H;�`H;��H;��H;�H;�H;վH;}�H;�H;��H;վH;~�H;��H;��H;��H;�`H;�6H;��G;��G;�G;�E;x�B;t�;;+j-;�;��:�9�P�����],�L�f������c���D�Ӑ�������������H�:�s�~쏾�R��"������      C��3�很Yؾ+�þĪ�~쏾�k�ۀ:�����ؽ�����c�cy���Ҽ���N� �v�D�� (7_�:��
;��(;�_9;��A;�\E;��F;͝G;��G;�.H;�ZH;|H;!�H;u�H;��H;@�H;�H;��H;�H;?�H;��H;t�H;#�H;|H;�ZH;�.H;��G;ϝG;��F;�\E;��A;�_9;��(;��
;a�: (7B��w�O� ������Ҽcy��c�������ؽ��ۀ:��k�~쏾Ī�+�þ�Yؾ3��      %��Q������AI�+�þ S��>���xS��Q"��s������}��0� 켑�����6�V�ƻQ}*�x�����:lx;[%;�l7;ڳ@;��D;��F;��G;��G;-(H;	VH;�xH;��H;q�H;ϲH;�H;��H;��H;��H;�H;βH;p�H;��H;�xH;VH;,(H;��G;��G;��F;��D;ճ@;�l7;[%;px;��:p���P}*�W�ƻ��6����� ��0���}�����s��Q"�xS�>��� S��+�þAIᾧ���Q��      ���T��;�
������Yؾ"���॒���f���0�^[�T8��Ԑ����>�����TȤ��6H�r�ܻ$rF����H�}:Ά�:c";U�5;��?;x�D;ӮF;�G;��G;k#H;~RH;�uH;��H;�H;��H;��H;�H;��H;�H;��H;��H;�H;��H;�uH;{RH;h#H;��G;�G;ծF;x�D;��?;X�5;c";҆�:H�}:���"rF�s�ܻ�6H�TȤ�������>�Ԑ��T8��^[���0���f�॒�"����Yؾ����;�
�T��      �� ����T��Q��3������0��9�s�ۀ:�j9�"�ʽ6Z���G��8�.���5S����0X���D��Bd:�B�: ;�4;È?;�~D;K�F;yG;��G;� H;FPH;EtH;>�H;��H;��H;`�H;��H;b�H;��H;b�H;��H;��H;A�H;EtH;CPH;� H;��G;yG;J�F;�~D;��?;"�4; ;�B�:�Bd:��D�0X���껻5S�.���8��G�6Z��"�ʽj9�ۀ:�9�s��0�����3��Q��T�����      IF�Zh����ZVھ:�������~���S��#��o��>S��t₽9�6�|���sy��dFB��Eֻ�A?��	�Y�:z��:c�";�46;V@;}�D;ɩF;�nG;�G;5H;0@H;gH;y�H;[�H;��H;�H;��H;�H;��H;�H;��H;Y�H;|�H;gH;.@H;2H;�G;�nG;ɩF;}�D;R@;�46;c�";|��:}Y�:�	��A?��EֻdFB�sy��|���9�6�t₽>S���o���#��S��~������:��ZVھ��Zh��      Zh���b���쾪*־�v��+���*��+�O�Y� �s��r���؀�N�3����Iݜ�J�>�e�ѻ �9�X���4o�:)% ;oM#;g�6;GA@;�D;ïF;qG;m�G;KH;�@H;�gH;�H;��H;�H;F�H;"�H;�H;"�H;F�H;�H;��H;�H;�gH;�@H;HH;m�G;qG;ïF;�D;AA@;l�6;oM#;*% ;0o�:X�����9�f�ѻJ�>�Iݜ����N�3��؀��r��s�Y� �+�O�*��+����v���*־���b��      ���쾷�޾35ʾP;���:��-�v��E�c'����w����u���+��W��A����4���Ļ>9)��j���W�:N�;%;
l7; �@;�D;�F;�wG;w�G;mH;\CH;UiH;G�H;��H;ѪH;�H;��H;��H;��H;�H;ѪH;��H;G�H;UiH;WCH;jH;w�G;�wG;�F;�D;�@;l7;%;M�;�W�:�j��=9)���Ļ��4��A���W缊�+���u�w�����c'��E�-�v��:��P;��35ʾ��޾��      ZVھ�*־25ʾu��������M���9b��5�����ս����Xc���֖ռ�I��b�$�}T���Z��^��$�:��;j�';A�8;RA;�9E;��F;ςG;�G;{H;%GH;<lH;|�H;f�H;�H;��H;��H;�H;��H;��H;�H;e�H;|�H;<lH;#GH;xH;�G;ςG;��F;�9E;RA;D�8;j�';��;"�:�^���Z�}T��b�$��I��֖ռ���Xc������ս���5��9b��M������u���25ʾ�*־      :���v��P;������UP��J�r�~�H�Y� ���:@��֓����K�g�־���s������ܺ04u9'&�:�;2�+;��:;�"B;��E;	�F;�G;�G;fH;TLH;'pH;r�H;��H;ЭH;h�H;�H;��H;�H;g�H;ѭH;��H;t�H;&pH;PLH;eH;�G;�G;�F;��E;�"B;��:;2�+;�;#&�:04u9�ܺ������s�־�g���K�֓��:@����Y� �~�H�J�r�VP������P;���v��      ����+����:���M��J�r�+�O�#,�[�
��gٽuĥ���u�1�u���4Ϥ���P�[��.o��p��:}��:�P;C�/;\�<;C;<�E;�!G;H�G;'�G;�%H;�RH;�tH;*�H;q�H;�H;5�H;��H;3�H;��H;5�H;�H;q�H;-�H;�tH;�RH;�%H;'�G;G�G;�!G;;�E;C;\�<;C�/;�P;y��::�p���.o�[򻹎P�3Ϥ�u���1���u�vĥ��gٽ\�
�#,�+�O�J�r��M���:��+���      �~��*��-�v� :b�~�H�#,�PZ����<S��|^����N������μ�I��&+�(����.�(����j~:j��:(m;��3;=�>;G�C;dPF;�FG;g�G;�G;�/H;"ZH;�zH;y�H;��H;��H;R�H;W�H;�H;V�H;R�H;��H;��H;{�H;�zH;!ZH;�/H;�G;f�G;�FG;aPF;A�C;=�>;��3;)m;d��:�j~:����.�)���&+��I����μ�����N�|^��<S�����PZ�#,�~�H� :b�-�v�*��      �S�+�O��E��5�Y� �[�
���罪9��,l���Xc���(��������[�����ݎ�hܺP:9��:@�	;Fd';q 8;_�@;��D;�F;HjG;��G;vH;�:H;cbH;�H;:�H;^�H;s�H;��H;f�H;�H;f�H;��H;s�H;\�H;;�H;�H;bbH;�:H;vH;��G;HjG;	�F;��D;_�@;o 8;Gd';?�	;��:`:9lܺ�ݎ������[��������(��Xc�,l���9�����[�
�Y� ��5��E�+�O�      �#�Y� �c'������gٽ<S��,l��W�j�J�3��i��վ�����(���Ļ|A?���B���@:�[�:Q;
�.;��;;�tB;/�E;��F;X�G;�G;H;�FH;IkH;��H;S�H;<�H;��H;?�H;��H;'�H;��H;>�H;��H;<�H;T�H;��H;HkH;�FH;
H;�G;X�G;��F;,�E;�tB;��;;�.;Q;�[�:��@:��B�|A?���Ļ(������վ��i�J�3�V�j�,l��<S���gٽ����c'�Y� �       p��s��罰�ս:@��vĥ�|^���Xc�J�3���	�ӌ˼�]��`FB�[򻾜���Ӻ ��8��:��;�M#;}=5;)?;q�C;�@F;0:G;�G;C�G;]'H;�RH;�tH;��H;��H;X�H;޻H;��H;��H;s�H;��H;��H;޻H;W�H;��H;��H;�tH;�RH;]'H;A�G;�G;-:G;�@F;p�C;)?;}=5;�M#;��;��: ��8�Ӻ����[�`FB��]��Ԍ˼��	�J�3��Xc�|^��vĥ�;@����ս���s�      >S���r��w�����֓����u���N���(��i�ӌ˼�A����P�rs��T|������\:(�:x�;�n-;��:;�A;�,E;��F;VoG;�G;�H;�7H;o_H;3~H;�H;3�H;��H;A�H;��H;l�H;��H;j�H;��H;@�H;��H;5�H;�H;0~H;m_H;�7H;�H;�G;SoG;��F;�,E;�A;�:;�n-;x�;,�:�\:����T|��rs���P��A��ӌ˼�i���(���N���u�֓�����w���r��      t₽�؀���u��Xc���K�1�������վ��]����P����QT����9�L�o�X3�9y&�:\�	;f%;d�5;��>;»C;�F;�!G;ʚG;��G;mH;�HH;�kH;͇H;}�H;íH;߹H;��H;~�H;��H;�H;��H;��H;��H;޹H;ƭH;}�H;͇H;�kH;�HH;kH;��G;ƚG;�!G;�F;»C;��>;_�5;f%;_�	;u&�:X3�9L�o���9�QT�������P��]���վ�����1���K��Xc���u��؀�      9�6�N�3���+���g�u�����μ�������_FB�qs�QT��@�D��{���9u9�q�:���:~Y;�t0;�;;�B;:E;�F;$hG;�G;6�G;�0H;�XH;^xH;P�H;��H;3�H;)�H;�H;E�H;\�H;k�H;\�H;D�H;�H;)�H;4�H;��H;P�H;[xH;�XH;�0H;7�G;�G; hG;�F;:E;�B;�;;�t0;�Y;���:�q�:�9u9�{��@�D�QT��qs�_FB����������μt���h�����+�N�3�      {������W�Ֆռ־�3Ϥ��I����[�(�[����9��{���:9FX�:[X�:FQ;E,;��8;�A@;%BD;�@F;�,G;��G;��G;�H;�DH;PhH;e�H;��H;��H;��H;T�H;S�H;�H;��H;��H;��H;�H;P�H;T�H;��H;��H;��H;b�H;MhH;�DH;�H;��G;��G;�,G;�@F;%BD;�A@;��8;H,;CQ;YX�:HX�:�:9�{����9��[�(���[��I��2Ϥ�־�Ֆռ�W����      ry��Iݜ��A���I����s���P�&+������Ļ����R|�L�o��9u9FX�:�+�:\;�);݄6;��>;�PC;��E;�F;�xG;W�G;�H;�1H;HXH;3wH;�H;G�H;5�H;��H;J�H;u�H;��H;�H;��H;�H;��H;s�H;J�H;��H;5�H;E�H;��H;2wH;EXH;�1H;�H;Q�G;�xG;�F;��E;�PC;��>;��6;�);[;�+�:FX�:�9u9L�o�R|�������Ļ���&+���P���s��I���A��Jݜ�      cFB�I�>���4�b�$��� [�%����ݎ�zA?��Ӻ����`3�9�q�:WX�:\;��';�=5;��=;�B;?GE;l�F;�UG;L�G;�G;�H;�HH;DjH;*�H;��H;x�H;e�H;z�H;�H;t�H;A�H;Q�H;��H;Q�H;A�H;r�H;�H;z�H;e�H;x�H;��H;*�H;@jH;�HH;�H;�G;F�G;�UG;g�F;=GE;�B;��=;�=5;��';^;YX�:�q�:X3�9�����ӺyA?��ݎ�&���[���b�$���4�K�>�      �Eֻ^�ѻ��Ļ}T�����.o��.�cܺ��B�`��8�\:{&�:���:EQ;�);�=5;�:=;:#B;��D; vF;7G;�G;��G;�H;�:H;D^H;�zH;,�H;��H;��H;=�H;��H;��H;O�H;��H;^�H;��H;]�H;��H;O�H;��H;��H;<�H;��H;��H;+�H;�zH;D^H;�:H;�H;��G;�G;7G; vF;��D;<#B;�:=;�=5;�);EQ;���:{&�:�\:���8��B�fܺ�.��.o���}T����Ļd�ѻ      �A?���9�89)��Z��ܺ�p�����`:9��@:��:0�:_�	;Y;E,;݄6;��=;8#B;��D;�XF;�!G;��G;H�G;�H;%/H;�SH;�qH;�H;�H;��H;�H;��H;�H;��H;�H;��H;N�H;��H;M�H;��H;�H;��H;�H;��H;�H;��H;�H;�H;�qH;�SH;/H;�H;H�G;��G;�!G;XF;��D;7#B;��=;݄6;E,;Y;_�	;0�:��:��@:0:9����p���ܺ�Z�99)��9�      ��	�X����j��@^��4u9":�j~:��:�[�:�;{�;i%;�t0;��8;��>;�B;��D;XF;ZG;��G;��G;��G;$&H;7KH;�iH;�H;��H;l�H;��H;<�H;��H;��H;��H;e�H;��H;�H;��H;�H;��H;d�H;��H;��H;��H;8�H;��H;k�H;��H;�H;�iH;3KH;&H;��G;��G;��G;ZG;�XF;��D;�B;��>;��8;�t0;h%;{�;�;�[�:��:�j~:>:�4u9 ^���j��X���      �Y�:Zo�:�W�:*�:'&�:{��:h��:?�	;Q;�M#;�n-;a�5;�;;�A@;�PC;9GE;�uF;�!G;��G;��G;C�G;| H;?EH;�cH;o}H;��H;�H;ձH;��H;��H;��H;]�H;��H;��H;��H;��H;!�H;��H;��H;��H;��H;_�H;��H;��H;�H;ұH;�H;��H;o}H;�cH;9EH;y H;@�G;��G;��G;�!G;�uF;8GE;�PC;�A@;�;;a�5;�n-;�M#;Q;?�	;f��:��:=&�:(�:�W�:Ho�:      ���:8% ;X�;��;�;�P;/m;Fd';
�.;�=5;��:;��>;�B;$BD;��E;j�F;7G;��G;��G;D�G;�H;BH;;`H;yH;��H;V�H;��H;�H;��H;�H;��H;b�H;��H;t�H;&�H;�H;��H;�H;&�H;t�H;��H;c�H;��H;�H;|�H;�H;��H;V�H;��H;}yH;8`H;BH;�H;D�G;��G;��G;7G;i�F;��E;$BD;�B;��>;�:;~=5;�.;Fd';/m;�P;�;��;T�;)% ;      p�";�M#;%;e�';6�+;N�/;��3;y 8;��;;/?;�A;ûC;:E;�@F;�F;�UG;�G;J�G;��G;} H;BH;�^H;ywH;O�H;��H;�H;ķH;b�H;4�H;\�H;T�H;�H;��H;�H;��H;y�H;��H;y�H;��H;�H;��H;�H;T�H;W�H;.�H;a�H;��H;�H;��H;J�H;vwH;�^H;BH;~ H;��G;K�G;�G;�UG;�F;�@F;:E;ûC;�A;/?;��;;y 8;��3;N�/;L�+;e�';%;�M#;      �46;n�6;l7;=�8;��:;^�<;B�>;b�@;�tB;p�C;�,E;�F;�F;�,G;�xG;J�G;��G;�H;$&H;@EH;;`H;{wH;c�H;h�H;{�H;�H;ϿH;��H;	�H;2�H;`�H;t�H;��H;��H;��H;��H;��H;��H;��H;��H;��H;r�H;`�H;/�H;�H;��H;˿H;�H;|�H;e�H;a�H;ywH;5`H;@EH;"&H;�H;��G;I�G;�xG;�,G;�F;�F;�,E;p�C;�tB;a�@;B�>;`�<;��:;=�8;l7;`�6;      k@;TA@;*�@;RA;�"B;	C;N�C;��D;/�E;�@F;��F;�!G;hG;��G;T�G;�G;�H;#/H;6KH;�cH;{yH;M�H;g�H;��H;;�H;��H;��H;�H;F�H;��H;��H;��H;q�H;��H;��H;��H;��H;��H; �H;��H;n�H;��H;��H;��H;C�H;�H;��H;��H;;�H;��H;e�H;L�H;xyH;�cH;4KH;%/H;�H;�G;T�G;��G;hG;�!G;��F;�@F;0�E;��D;M�C;
C;�"B;RA;*�@;JA@;      ��D;�D;�D;�9E;��E;A�E;aPF;�F;��F;-:G;SoG;̚G;�G;��G;�H;�H;�:H;�SH;�iH;v}H;��H;��H;��H;C�H;n�H;�H;b�H;��H;��H;c�H;�H;?�H;��H;!�H;��H;V�H;��H;U�H;��H;�H;��H;?�H;�H;b�H;��H;��H;a�H;�H;m�H;?�H;�H;��H;��H;x}H;�iH;�SH;�:H;�H;�H;��G;�G;͚G;UoG;,:G;��F;	�F;cPF;A�E;��E;�9E; �D;�D;      ۩F;үF;�F;��F;�F;�!G;�FG;GjG;X�G;�G;�G;��G;5�G;�H;�1H;�HH;C^H;�qH;�H;��H;S�H;�H;�H;��H;�H;C�H;S�H;��H;��H;��H;��H;��H;&�H;�H;��H;�H;A�H;�H;��H;�H;!�H;��H;��H;��H;��H;��H;S�H;B�H;�H;��H;�H;�H;O�H;��H;�H;�qH;A^H;�HH;�1H;�H;6�G; �G;�G;�G;Y�G;GjG;�FG;�!G;�F;��F;�F;ɯF;      �nG;"qG;�wG;ՂG;�G;N�G;n�G;��G;�G;A�G;�H;qH;�0H;�DH;FXH;DjH;�zH;�H;��H;�H;��H;ķH;ͿH;��H;]�H;W�H;t�H;��H;��H;��H;��H;�H;�H;��H;k�H;��H;��H;��H;j�H;��H;�H;�H;��H;��H;��H;��H;s�H;U�H;]�H;��H;˿H;·H;��H;�H;��H;�H;�zH;CjH;FXH;�DH;�0H;qH;�H;A�G;�G;��G;n�G;L�G;�G;ӂG;�wG;!qG;      
�G;s�G;��G;�G;�G;*�G;�G;H;H;d'H;�7H;�HH;�XH;QhH;3wH;*�H;+�H;�H;h�H;رH;�H;b�H;��H;�H;��H;��H;��H;q�H;��H;|�H;��H;��H;��H;��H;�H;;�H;L�H;:�H;�H;��H;��H;��H;��H;x�H;��H;o�H;��H;��H;��H;�H;��H;a�H;�H;رH;i�H;�H;)�H;*�H;4wH;PhH;�XH;�HH;�7H;d'H;H;H;�G;*�G;�G;�G;��G;|�G;      NH;JH;oH;H;hH;�%H;�/H;�:H;�FH;�RH;o_H;lH;]xH;d�H;�H;��H;��H;��H;��H;��H;��H;2�H;�H;J�H;��H;��H;��H;��H;Y�H;��H;�H;��H;��H;�H;|�H;��H;��H;��H;|�H;�H;��H;��H;��H;��H;W�H;��H;��H;��H;��H;J�H;�H;1�H;}�H;��H;��H;��H;��H;��H;�H;d�H;^xH; lH;n_H;�RH;�FH;�:H;�/H;�%H;mH;H;mH;@H;      <@H;AH;eCH;,GH;gLH;�RH;)ZH;jbH;RkH;�tH;:~H;ڇH;W�H;��H;K�H;|�H;��H;�H;8�H;��H;�H;Y�H;-�H;��H;Z�H;��H;��H;y�H;��H;��H;��H;��H;1�H;��H;��H;	�H;�H;�H;��H;��H;-�H;��H;��H;��H;��H;x�H;��H;��H;[�H;��H;,�H;Y�H;�H;��H;:�H;�H;��H;|�H;K�H;��H;U�H;هH;<~H;�tH;UkH;kbH;)ZH;�RH;bLH;,GH;`CH; AH;      gH;�gH;ciH;IlH;5pH;�tH;�zH;�H;��H;�H;$�H;��H;��H;��H;9�H;n�H;C�H;��H;��H;��H;��H;T�H;`�H;��H;�H;��H;��H;��H;��H;��H;��H;<�H;��H;��H;�H;C�H;_�H;C�H;�H;��H;��H;>�H;��H;��H;�H;��H;��H;��H;�H;��H;]�H;T�H;��H;��H;��H;��H;A�H;l�H;9�H;��H;��H;��H;%�H;�H;��H;�H;�zH; uH;3pH;JlH;ciH;�gH;      ��H;��H;T�H;��H;y�H;0�H;�H;C�H;X�H;��H;:�H;ͭH;9�H;��H;��H;��H;�H;�H;��H;g�H;j�H;"�H;u�H;��H;:�H;��H;�H;��H;��H;��H;:�H;��H;��H;5�H;_�H;~�H;z�H;~�H;^�H;5�H;��H;��H;:�H;��H;��H;��H;�H;��H;<�H;��H;r�H;"�H;h�H;g�H;��H;�H;�H;��H;��H;��H;9�H;ͭH;;�H;��H;Z�H;A�H;��H;3�H;x�H;��H;U�H;�H;      b�H;ǚH;ɛH;m�H;��H;t�H;��H;i�H;C�H;Z�H;��H;�H;.�H;Y�H;O�H;	�H;��H;��H;��H;��H;��H;��H;��H;x�H;��H;(�H;�H;��H;��H;8�H;��H;��H;8�H;q�H;��H;��H;��H;��H;��H;p�H;5�H;��H;��H;:�H;��H;��H;�H;&�H;��H;w�H;��H;��H;��H;��H;��H;��H;��H;	�H;M�H;Y�H;,�H;�H;��H;[�H;C�H;h�H;��H;w�H;��H;m�H;ɛH;��H;      ͩH;�H;̪H;�H;ܭH;�H;��H;��H;��H;�H;H�H;��H;�H;W�H;y�H;|�H;V�H;�H;h�H;��H;|�H;�H;��H;��H;�H;�H;��H;��H;�H;��H;��H;5�H;j�H;��H;��H;��H;��H;��H;��H;��H;h�H;8�H;��H;��H;�H;��H;��H;�H;�H;��H;��H;�H;y�H;��H;h�H;�H;U�H;|�H;y�H;W�H;�H;��H;G�H;�H;��H;~�H;��H;�H;ҭH;�H;ΪH;�H;      �H;]�H;��H;��H;��H;5�H;\�H;��H;H�H;��H;��H;��H;L�H;�H;��H;I�H;��H;��H;��H;��H;1�H;��H;��H;�H;��H;��H;g�H;�H;|�H;��H;�H;b�H;��H;��H;��H;��H;��H;��H;��H;��H;��H;c�H;�H;��H;~�H;�H;e�H;��H;��H;�H;��H;��H;.�H;��H;��H;��H;��H;I�H;��H;�H;K�H;��H;��H;��H;H�H;��H;\�H;9�H;y�H;��H;��H;T�H;      ��H;,�H;ʺH;ĻH;�H;��H;b�H;r�H;��H; �H;t�H;��H;b�H;��H;�H;X�H;e�H;I�H;�H;��H; �H;|�H;��H;��H;Q�H;�H;��H;:�H;��H;�H;B�H;�H;��H;��H;��H;��H;��H;��H;��H;��H;��H;��H;B�H;�H;��H;:�H;��H;�H;R�H;��H;��H;|�H;�H;��H;�H;J�H;d�H;X�H;�H;��H;b�H;��H;s�H;�H;��H;p�H;a�H;��H;	�H;ĻH;̺H;$�H;      �H;�H;��H;��H;þH;5�H;�H;
�H;2�H;u�H;��H;�H;n�H;��H;��H;�H;��H;��H;��H;*�H;��H;��H;��H;��H;��H;=�H;��H;P�H;��H;�H;b�H;�H;��H;��H;��H;��H;��H;��H;��H;��H;��H;��H;b�H;�H;��H;P�H;��H;>�H;��H;��H;��H;��H;��H;*�H;��H;��H;��H;�H;��H;��H;n�H;�H;��H;w�H;2�H;�H;�H;:�H;��H;��H;��H;�H;      ��H;.�H;ʺH;ĻH;�H;��H;b�H;r�H;��H; �H;t�H;��H;b�H;��H;�H;X�H;e�H;I�H;�H;��H;!�H;|�H;��H;��H;R�H;�H;��H;:�H;��H;�H;B�H;�H;��H;��H;��H;��H;��H;��H;��H;��H;��H;��H;B�H;�H;��H;:�H;��H;�H;Q�H;��H;��H;|�H;�H;��H;�H;J�H;d�H;X�H;�H;��H;b�H;��H;t�H;�H;��H;p�H;b�H;��H;�H;ĻH;ȺH;!�H;      �H;]�H;��H;��H;��H;5�H;\�H;��H;H�H;��H;��H;��H;L�H;�H;��H;I�H;��H;��H;��H;��H;2�H;��H;��H;�H;��H;��H;g�H;�H;}�H;��H;�H;a�H;��H;��H;��H;��H;��H;��H;��H;��H;��H;f�H;�H;��H;~�H;�H;e�H;��H;��H;�H;��H;��H;.�H;��H;��H;��H;��H;I�H;��H;�H;L�H;��H;��H;��H;H�H;��H;\�H;9�H;y�H;��H;��H;T�H;      ΩH;�H;ΪH;�H;ޭH;�H;��H;��H;��H;�H;H�H;��H;�H;W�H;y�H;|�H;V�H; �H;h�H;��H;�H;�H;��H;��H;�H;�H;��H;��H;�H;��H;��H;5�H;i�H;��H;��H;��H;��H;��H;��H;��H;i�H;8�H;��H;��H;�H;��H;��H;�H;�H;��H;��H;�H;{�H;��H;h�H;�H;U�H;|�H;y�H;W�H;�H;��H;H�H;�H;��H;�H;��H;�H;ѭH;�H;ΪH;�H;      d�H;ǚH;ɛH;o�H;��H;t�H;��H;h�H;C�H;Z�H;��H;�H;,�H;Y�H;M�H;	�H;��H;��H;��H;��H;��H;��H;��H;w�H;��H;'�H;�H;��H;��H;8�H;��H;��H;6�H;o�H;��H;��H;��H;��H;��H;p�H;5�H;��H;��H;:�H;��H;��H;�H;'�H;��H;w�H;��H;��H;��H;��H;��H;��H;��H;	�H;N�H;Y�H;,�H;�H;��H;[�H;C�H;e�H;��H;x�H;��H;o�H;țH;ÚH;      ��H;��H;U�H;��H;y�H;0�H;��H;C�H;X�H;��H;:�H;ͭH;9�H;��H;��H;��H;�H;�H;��H;i�H;m�H;"�H;u�H;��H;<�H;��H;�H;��H;��H;��H;:�H;��H;��H;5�H;^�H;~�H;z�H;~�H;_�H;5�H;��H;��H;:�H;��H;��H;��H;�H;��H;:�H;��H;t�H;"�H;i�H;g�H;��H;�H;�H;��H;��H;��H;9�H;ͭH;:�H;��H;Z�H;A�H;��H;2�H;v�H;��H;V�H;�H;      gH;�gH;ciH;JlH;5pH;�tH;�zH;�H;��H;�H;%�H;��H;��H;��H;9�H;n�H;A�H;��H;��H;��H;��H;T�H;`�H;��H;�H;��H;��H;��H;��H;��H;��H;<�H;��H;��H;�H;C�H;_�H;C�H;�H;��H;��H;>�H;��H;��H;�H;��H;��H;��H;�H;��H;]�H;T�H;��H;��H;��H;��H;A�H;n�H;9�H;��H;��H;��H;"�H;�H;��H;�H;�zH; uH;3pH;IlH;ciH;�gH;      7@H;AH;dCH;,GH;bLH;�RH;,ZH;mbH;SkH;�tH;:~H;ڇH;T�H;��H;K�H;|�H;��H;�H;8�H;��H;	�H;Y�H;-�H;��H;[�H;��H;��H;x�H;��H;��H;��H;��H;0�H;��H;��H;	�H;�H;	�H;��H;��H;0�H;��H;��H;��H;��H;y�H;��H;��H;Z�H;��H;,�H;Y�H;�H;��H;8�H;�H;��H;}�H;K�H;��H;W�H;ڇH;:~H;�tH;VkH;mbH;,ZH;�RH;aLH;-GH;cCH;AH;      GH;FH;tH;~H;lH;�%H;�/H;�:H;�FH;�RH;o_H;lH;]xH;d�H;�H;��H;��H;��H;��H;��H;��H;1�H;�H;H�H;��H;��H;��H;��H;W�H;��H;��H;��H;��H;�H;z�H;��H;��H;��H;|�H;�H;��H;��H;�H;��H;Y�H;��H;��H;��H;��H;J�H;�H;2�H;��H;��H;��H;��H;��H;��H;�H;d�H;]xH;lH;o_H;�RH;�FH;�:H;�/H;�%H;iH;{H;tH;GH;      
�G;s�G;��G;�G;�G;*�G;�G;�H;H;d'H; 8H;�HH;�XH;QhH;4wH;*�H;+�H;�H;i�H;ױH;�H;a�H;��H;�H;��H;��H;��H;o�H;��H;{�H;��H;��H;��H;��H;
�H;;�H;L�H;;�H;�H;��H;��H;��H;��H;y�H;��H;q�H;��H;��H;��H;�H;��H;b�H;�H;رH;h�H;�H;)�H;+�H;3wH;OhH;�XH;�HH;�7H;d'H;H;H;�G;'�G;�G;�G;��G;~�G;      �nG;$qG;�wG;΂G;�G;I�G;m�G;��G;�G;B�G;�H;qH;�0H;�DH;FXH;DjH;�zH;�H;��H;�H;��H;·H;̿H;��H;]�H;W�H;v�H;��H;��H;��H;��H;�H;�H;��H;j�H;��H;��H;��H;k�H;��H;�H;�H;��H;��H;��H;��H;s�H;W�H;]�H;��H;̿H;ķH;��H;�H;��H;�H;�zH;CjH;FXH;�DH;�0H;qH;�H;B�G;�G;��G;m�G;H�G;�G;΂G;�wG;qG;      ߩF;ίF;�F;��F;�F;�!G;�FG;JjG;W�G;�G;�G;��G;6�G;�H;�1H;�HH;C^H;�qH;�H;��H;T�H;�H;�H;��H;�H;B�H;T�H;��H;��H;��H;��H;��H;#�H;�H;��H;�H;A�H;�H;��H;�H;#�H;��H;��H;��H;��H;��H;S�H;C�H;�H;��H;�H;�H;O�H;��H;�H;�qH;A^H;�HH;�1H;�H;5�G;��G;�G;�G;X�G;GjG;�FG;�!G;�F;��F;�F;įF;      ��D;�D; �D;�9E;��E;A�E;cPF;�F;��F;-:G;UoG;͚G;�G;��G;�H;�H;�:H;�SH;�iH;w}H;��H;��H;��H;B�H;m�H;�H;b�H;��H;��H;c�H;�H;=�H;��H;�H;��H;U�H;��H;V�H;��H; �H;��H;A�H;�H;b�H;��H;��H;b�H;�H;n�H;B�H;��H;��H;��H;w}H;�iH;�SH;�:H;�H;�H;��G;�G;̚G;SoG;,:G;��F;�F;aPF;A�E;��E;�9E; �D;�D;      q@;QA@;0�@;RA;�"B;C;K�C;��D;0�E;�@F;��F;�!G; hG;��G;T�G;�G;�H;"/H;4KH;�cH;}yH;L�H;g�H;��H;;�H;��H;��H;�H;F�H;��H;��H;��H;p�H;��H;��H;��H;��H;��H; �H;��H;p�H;��H;��H;��H;C�H;�H;��H;��H;;�H;��H;e�H;M�H;zyH;�cH;6KH;%/H;�H;�G;T�G;��G;hG;�!G;��F;�@F;0�E;��D;K�C;C;�"B;RA;-�@;GA@;      �46;y�6;!l7;=�8;��:;c�<;F�>;b�@;�tB;p�C;�,E;�F;
�F;�,G;�xG;J�G;��G;�H;"&H;?EH;;`H;ywH;c�H;h�H;|�H;�H;ͿH;��H;�H;2�H;`�H;r�H;��H;��H;��H;��H;��H;��H;��H;��H;��H;t�H;`�H;/�H;�H;��H;̿H; �H;{�H;g�H;c�H;{wH;8`H;BEH;$&H;�H;��G;J�G;�xG;�,G;
�F;�F;�,E;m�C;�tB;a�@;H�>;c�<;��:;<�8;l7;k�6;      p�";�M#;%;e�';6�+;N�/;��3;{ 8;��;;/?;�A;ûC;:E;�@F;�F;�UG;�G;H�G;��G;| H;BH;�^H;ywH;O�H;��H;�H;·H;a�H;2�H;\�H;T�H;�H;��H;�H;��H;y�H;��H;y�H;��H;�H;��H;�H;T�H;W�H;/�H;b�H;��H;�H;��H;L�H;vwH;�^H;BH;} H;��G;K�G;�G;�UG;�F;�@F;:E;ĻC;�A;/?;�;;y 8;��3;N�/;L�+;e�';%;�M#;      ���:3% ;\�;��;�;�P;3m;Hd';
�.;�=5;�:;��>;�B;$BD;��E;i�F;7G;��G;��G;C�G;�H;BH;:`H;yH;��H;V�H;��H;�H;�H;�H;��H;b�H;��H;r�H;&�H;�H;��H;�H;&�H;t�H;��H;e�H;��H;�H;}�H;�H;��H;V�H;��H;}yH;:`H;BH;�H;D�G;��G;��G;7G;i�F;��E;$BD;�B;��>;�:;}=5;�.;Gd';2m;�P;�;��;Z�;(% ;      �Y�:Zo�:�W�:$�:/&�:y��:j��:@�	;Q;�M#;�n-;a�5;�;;�A@;�PC;8GE;�uF;�!G;��G;��G;C�G;y H;=EH;�cH;o}H;��H;�H;ұH;��H;��H;��H;]�H;��H;��H;��H;��H;!�H;��H;��H;��H;��H;_�H;��H;��H;��H;ձH;�H;��H;o}H;�cH;<EH;| H;@�G;��G;��G;�!G;�uF;9GE;�PC;�A@;�;;_�5;�n-;�M#;Q;@�	;l��:��:=&�:&�:�W�:Ho�:      ��	�X����j�� ^��4u9":�j~:��:�[�:�;{�;h%;�t0;��8;��>;�B;��D;XF;ZG;��G;��G;��G;"&H;6KH;�iH;�H;��H;k�H;��H;;�H;��H;��H;��H;d�H;��H;�H;��H;�H;��H;e�H;��H;��H;��H;:�H;��H;l�H;��H;�H;�iH;4KH; &H;��G;��G;��G;ZG;�XF;��D;�B;��>;��8;�t0;i%;{�;�;�[�:��:�j~:B:�4u9@^���j��P���      �A?���9�89)��Z��ܺ�p�����P:9��@:��:.�:_�	;Y;B,;݄6;��=;8#B;��D;XF;�!G;��G;H�G;�H;#/H;�SH;�qH;�H;�H;��H;�H;��H;�H;��H;�H;��H;M�H;��H;M�H;��H;�H;��H;�H;��H;�H;��H;�H;�H;�qH;�SH;!/H;�H;H�G;��G;�!G;�XF;��D;7#B;��=;݄6;D,;Y;_�	;0�:��:��@:0:9����p���ܺ�Z�99)��9�      �Eֻ_�ѻ��Ļ}T�����.o��.�cܺ��B����8�\:{&�:���:EQ;�);�=5;�:=;:#B;��D;�uF;7G;�G;��G;�H;�:H;C^H;�zH;+�H;��H;��H;<�H;��H;��H;O�H;��H;^�H;��H;^�H;��H;Q�H;��H;��H;=�H;��H;��H;,�H;�zH;F^H;�:H;�H;��G;�G;7G; vF;��D;<#B;�:=;�=5;�);EQ;���:{&�:�\:@��8��B�fܺ�.��.o���}T����Ļd�ѻ      cFB�I�>���4�b�$��� [�&����ݎ�zA?��Ӻ����`3�9�q�:WX�:^;��';�=5;��=;�B;=GE;i�F;�UG;I�G;�G;�H;�HH;CjH;*�H;��H;x�H;e�H;x�H;�H;r�H;A�H;Q�H;��H;Q�H;A�H;t�H;�H;{�H;e�H;x�H;��H;*�H;AjH;�HH;�H;�G;I�G;�UG;i�F;?GE;�B;��=;�=5;��';^;WX�:�q�:`3�9�����ӺzA?��ݎ�%���[���b�$���4�K�>�      ry��Iݜ��A���I����s���P�&+������Ļ����T|�L�o��9u9FX�:�+�:[;�);݄6;��>;�PC;��E;�F;�xG;V�G;�H;�1H;FXH;2wH;�H;G�H;5�H;��H;K�H;u�H;��H;�H;��H;�H;��H;v�H;J�H;��H;5�H;E�H;��H;3wH;FXH;�1H;�H;S�G;�xG;�F;��E;�PC;��>;��6;�);\;�+�:FX�:�9u9L�o�R|�������Ļ���&+���P���s��I���A��Jݜ�      {������W�Ֆռ־�3Ϥ��I����[�(�[����9��{���:9JX�:YX�:EQ;F,;��8;�A@;$BD;�@F;�,G;��G;��G;�H;�DH;MhH;d�H;��H;��H;��H;U�H;Q�H;�H;��H;��H;��H;�H;Q�H;R�H;��H;��H;��H;d�H;PhH;�DH;�H;��G;��G;�,G;�@F;&BD;�A@;��8;H,;EQ;[X�:FX�:�:9�{����9��[�(���[��I��2Ϥ�־�Ֆռ�W����      9�6�N�3���+���g�u�����μ�������_FB�qs�QT��@�D��{���9u9�q�:���:Y;�t0;�;;�B;:E;�F;$hG;�G;6�G;�0H;�XH;]xH;P�H;��H;3�H;)�H;�H;D�H;\�H;k�H;\�H;E�H;�H;(�H;4�H;��H;P�H;[xH;�XH;�0H;9�G;�G;hG;
�F;:E;�B;�;;�t0;�Y;���:�q�:�9u9�{��@�D�QT��qs�_FB����������μt���g�����+�N�3�      t₽�؀���u��Xc���K�1�������վ��]����P����QT����9�L�o�X3�9w&�:^�	;f%;a�5;��>;»C;�F;�!G;ƚG;��G;mH;�HH;�kH;͇H;}�H;íH;�H;��H;��H;��H;�H;��H;~�H;��H;޹H;ĭH;}�H;͇H;�kH;�HH;mH;��G;ʚG;�!G;�F;»C;��>;b�5;f%;_�	;u&�:H3�9L�o���9�QT�������P��]���վ�����1���K��Xc���u��؀�      >S���r��w�����֓����u���N���(��i�ӌ˼�A����P�rs��T|������\:*�:x�;�n-;�:;�A;�,E;��F;SoG;�G;�H;�7H;o_H;2~H;�H;1�H;��H;@�H;��H;l�H;��H;l�H;��H;A�H;��H;5�H;�H;2~H;m_H;�7H;�H;�G;VoG;��F;�,E;�A;�:;�n-;x�;,�:�\:����T|��rs���P��A��ӌ˼�i���(���N���u�֓�����w���r��       p��s��罰�ս:@��vĥ�|^���Xc�J�3���	�Ԍ˼�]��`FB�[򻾜���Ӻ ��8��:��;�M#;{=5;)?;q�C;�@F;-:G;�G;B�G;]'H;�RH;�tH;��H;��H;X�H;޻H;��H;��H;s�H;��H;��H;޻H;W�H;��H;��H;�tH;�RH;]'H;B�G;�G;0:G;�@F;p�C;)?;}=5;�M#;��;��:���8�Ӻ����[�`FB��]��Ԍ˼��	�J�3��Xc�|^��vĥ�:@����ս���s�      �#�Y� �c'������gٽ<S��,l��V�j�J�3��i��վ�����(���Ļ|A?���B���@:�[�:Q;	�.;��;;�tB;/�E;��F;X�G;�G;
H;�FH;HkH;��H;S�H;=�H;��H;>�H;��H;'�H;��H;>�H;��H;;�H;S�H;��H;HkH;�FH;H;�G;X�G;��F;,�E;�tB;��;;�.;Q;�[�:��@:��B�|A?���Ļ(������վ��i�J�3�V�j�,l��<S���gٽ����c'�Y� �      �S�+�O��E��5�Y� �[�
���罪9��,l���Xc���(��������[�����ݎ�hܺ@:9��:@�	;Dd';o 8;_�@;��D;	�F;HjG;��G;vH;�:H;cbH;�H;:�H;_�H;t�H;��H;f�H;�H;g�H;��H;t�H;\�H;:�H;�H;cbH;�:H;vH;��G;GjG;�F;��D;_�@;q 8;Gd';?�	;��:`:9lܺ�ݎ������[��������(��Xc�,l���9�����[�
�Y� ��5��E�+�O�      �~��*��-�v� :b�~�H�#,�PZ����<S��|^����N������μ�I��&+�)����.� ����j~:f��:'m;��3;=�>;G�C;aPF;�FG;g�G;�G;�/H;"ZH;�zH;y�H;��H;��H;R�H;V�H;�H;W�H;R�H;��H;��H;y�H;�zH;!ZH;�/H;�G;f�G;�FG;dPF;C�C;=�>;��3;)m;d��:�j~:����.�)���&+��I����μ�����N�|^��<S�����PZ�#,�~�H� :b�-�v�*��      ����+����:���M��J�r�+�O�#,�\�
��gٽuĥ���u�1�u���4Ϥ���P� [��.o��p��:y��:�P;C�/;[�<;C;;�E;�!G;H�G;'�G;�%H;�RH;�tH;*�H;r�H;�H;5�H;��H;3�H;��H;5�H;�H;p�H;-�H;�tH;�RH;�%H;'�G;G�G;�!G;<�E;C;\�<;C�/;�P;y��::�p���.o� [򻹎P�4Ϥ�u���1���u�uĥ��gٽ\�
�#,�+�O�J�r��M���:��+���      :���v��P;������UP��J�r�~�H�X� ���:@��֓����K�g�־���s������ܺ04u9%&�:�;2�+;��:;�"B;��E;	�F;�G;�G;hH;TLH;&pH;r�H;��H;ѭH;h�H;�H;��H;�H;g�H;ЭH;��H;t�H;'pH;QLH;eH;�G;�G;�F;��E;�"B;��:;2�+;�;%&�:04u9�ܺ������s�־�g���K�֓��:@����X� �~�H�J�r�UP������P;���v��      ZVھ�*־25ʾu��������M���9b��5�����ս����Xc���֖ռ�I��b�$�}T���Z��^��$�:��;j�';@�8;RA;�9E;��F;ςG;�G;{H;&GH;<lH;|�H;f�H;�H;��H;��H;�H;��H;��H;�H;e�H;z�H;<lH;#GH;xH;�G;ςG;��F;�9E;RA;F�8;j�';��;"�:�^���Z�~T��b�$��I��֖ռ���Xc������ս���5��9b��M������u���25ʾ�*־      ���쾷�޾35ʾP;���:��,�v��E�c'����w����u���+��W��A����4���Ļ>9)��j���W�:L�;%;
l7; �@;�D;�F;�wG;w�G;mH;ZCH;UiH;G�H;��H;ѪH;�H;��H;��H;��H;�H;ѪH;��H;G�H;UiH;WCH;jH;w�G;�wG;�F;�D;�@;l7;%;N�;�W�:�j��<9)���Ļ��4��A���W缊�+���u�w�����c'��E�,�v��:��P;��35ʾ��޾��      Zh���b���쾪*־�v��+���*��+�O�Y� �s��r���؀�N�3����Iݜ�J�>�e�ѻ �9�X���4o�:)% ;oM#;g�6;HA@;�D;ïF;qG;m�G;KH;�@H;�gH;�H;��H;�H;F�H;"�H;�H;"�H;H�H;�H;��H;�H;�gH;�@H;HH;m�G;qG;ïF;�D;CA@;l�6;oM#;*% ;0o�:X�����9�f�ѻJ�>�Iݜ����N�3��؀��r��s�Y� �+�O�*��+����v���*־���b��      ���
^�X_ݾ��ɾm*���{x�*G�T,�����b��f@{���/����噼�J;�`�ͻ�4��W���:!;��#;?�6;[@;L�D;̱F;�lG;��G;qH;�:H;�bH;�H;W�H;^�H;�H; �H;�H; �H;�H;^�H;V�H;�H;�bH;�:H;nH;��G;�lG;̱F;L�D;[@;B�6;��#;#;��:�W� �4�b�ͻ�J;�噼����/�f@{��b�����T,�*G�{x��m*����ɾX_ݾ
^�      
^�7���:پ�žj�����	9t�t�C������ꪫ�``w�N-����4`����7�HSɻ�K/�xyƹ§�:�/;�f$;�7;�~@;g�D;��F;�nG;�G;ZH;�;H;�cH;��H;��H;��H;=�H;W�H;O�H;W�H;?�H;��H;��H;��H;�cH;�;H;WH;�G;�nG;��F;g�D;�~@;�7;�f$;�/;���:xyƹ�K/�ISɻ��7�4`�����N-�``w�ꪫ������t�C�	9t���j����ž�:پ8��      X_ݾ�:پ�V;+���Ƥ�Oa����g��$:��Z�uݽ�ƣ��l�m.%��߼q���9.�ܴ��pV�p2p�A�: x;J(&;V�7;6�@;E;�F;suG;E�G;�H;�=H;xeH;��H;��H;~�H;�H;�H;�H;�H;߲H;}�H;��H;��H;xeH;�=H;�H;E�G;suG;�F;E;1�@;Y�7;H(&; x;A�:p2p�oV�ݴ���9.�q���߼m.%��l��ƣ�uݽ�Z��$:���g�Oa���Ƥ�+���V;�:پ      ��ɾ�ž+��tת��#�����T��J+�>��2̽�s���yZ����Xμoy��%��mϨ�l,� ��6'��:�
;^�(;xN9;��A;�NE;f�F;�G;��G;�H;�AH;`hH;�H;j�H;�H;�H;ҹH;��H;ҹH;�H;�H;i�H;�H;^hH;�AH;�H;��G;�G;f�F;�NE;��A;|N9;[�(;�
;#��: ��6l,�mϨ�&��oy��Xμ����yZ��s���2̽>��J+���T�#����tת�+���ž      l*��j����Ƥ���/��C�c��G=����zｖж��ɇ�Y�C���."���;k��&��-����˺�X�9���:9;�h,;�	;;�PB;��E;� G;�G;��G;�H;,GH;|lH;4�H;ǜH;ūH;m�H;2�H;�H;2�H;l�H;īH;ƜH;5�H;|lH;)GH;�H;��G;�G;� G;��E;�PB;�	;;�h,;9;���:�X�9��˺�-���&��;k�."����Y�C��ɇ��ж��z����G=�C�c��/����Ƥ�j���      ���Oa��$���C�c�t�C�~#�!��XvϽ�����l�kg*����
���I�����\c�9퀺�t,:��:�;�_0;��<;�1C;�E;�#G;f�G;3�G;B H;�MH;eqH;ۋH;��H;�H;^�H;̼H;��H;̼H;`�H;�H;��H;ދH;eqH;�MH;< H;3�G;e�G;�#G;�E;�1C;��<;�_0;�;��:�t,:8퀺�\c�����I��
�����kg*��l�����XvϽ!��~#�t�C�C�c�$���Oa����      {x�	9t���g���T��G=�~#�6�tݽ�b������JG�����Ǽpy��W�$�w���4�$�pvƹ@��:�&�:�� ;T4;��>;[D;�[F;�FG;��G;*�G;3*H;UH;&wH;.�H;�H;��H;��H;��H;[�H;��H;��H;��H;�H;0�H;&wH;~UH;0*H;*�G;��G;�FG;�[F;TD;��>;T4;�� ;�&�:@��:`vƹ4�$�x���W�$�py���Ǽ���JG������b��tݽ6�~#��G=���T���g�	9t�      *G�t�C��$:��J+��� ��tݽb���2I���yZ���"����ܫ��rT��� �,M��̃˺pm94ٶ:x�;
`(;�8;��@;��D;�F;shG;��G;�H;c5H;^H;�}H;�H;�H;��H;��H;��H;i�H;��H;��H;��H;�H; �H;�}H;^H;_5H;�H;��G;shG; �F;��D;��@;�8;`(;v�;4ٶ:�m9Ѓ˺+M���� �rT�ܫ�������"��yZ�2I��b���tݽ �����J+��$:�t�C�      S,����Z�>��z�XvϽ�b��2I��n]a�M-�n� �+"����{�Q�!�������4��P(��nQ:�L�:�;܊/;�'<;�B;�E;	�F;��G;��G;_H;oAH;;gH;|�H;g�H;��H;ȶH;��H;)�H;��H;)�H;��H;ȶH;��H;i�H;|�H;:gH;lAH;\H;��G;��G;�F;�E;��B;�'<;ފ/;�;�L�:�nQ:�P(���4�����Q�!���{�+"��n� �M-�n]a�2I���b��XvϽ�z�>��Z���      ������uݽ�2̽�ж����������yZ�N-�۷�8aļaO���J;���軚�|���º�M@9���:B�;�f$;��5;�N?;^D;�LF;#;G;ͤG;�G;�!H;NH;�pH;��H;�H;Z�H; �H;t�H;��H;��H;��H;t�H; �H;Y�H;�H;��H;�pH;NH;�!H;�G;ΤG; ;G;�LF;\D;�N?;��5;�f$;B�;���:�M@9��º��|�����J;�`O��8aļ۷�N-��yZ����������ж��2̽uݽ���      �b��ꪫ��ƣ��s���ɇ��l�JG���"�n� �8aļj���I��C��ۙ�[��uƹD�k:���:�;W>.;)
;;��A;�AE;z�F;9mG;��G;��G;�2H;[H;�zH;
�H;��H;ĳH;��H;a�H;.�H;D�H;.�H;a�H;��H;³H;��H;
�H;�zH;[H;�2H;��G;��G;5mG;v�F;�AE;��A;&
;;V>.;�;���:@�k:�uƹ[��ۙ��C��I�j��8aļn� ���"�JG��l��ɇ��s���ƣ�ꪫ�      f@{�``w��l��yZ�Y�C�kg*�������+"��`O���I�I|�IϨ��K/��$T�
Q:W��:��;�(&; $6;�%?;��C;�#F;$G;J�G;��G;�H;WCH;hH;��H;��H;��H;�H;#�H;S�H;��H;��H;��H;U�H;!�H;�H;��H;��H;��H;hH;WCH;�H;��G;F�G;$G;�#F;��C;�%?;�#6;�(&;��;S��:
Q:�$T��K/�IϨ�H|��I�`O��+"����鼴��kg*�Y�C��yZ��l�``w�      ��/�N-�l.%����������Ǽܫ����{��J;��C�IϨ�bO:�� [�9���:w;��;K.1;(<;�5B;�NE;6�F;VfG;�G;a�G;"+H;TH;uH;N�H;�H;P�H;~�H;��H;�H;.�H;T�H;.�H;�H;��H;}�H;Q�H;�H;N�H; uH;TH;+H;b�G;
�G;RfG;1�F;�NE;�5B;(<;K.1;��;u;���: [�9�bO:�IϨ��C��J;���{�ܫ���Ǽ��������l.%�N-�      ������߼Wμ-"���
��oy��qT�P�!�����ۙ��K/�� m9�A�:���::�;H�,;�N9;`@;�^D;�LF;�.G;�G;��G;�H;�?H;IdH;I�H;��H;;�H;˶H;��H;�H;��H;��H;��H;��H;��H;
�H;��H;ζH;;�H;��H;F�H;IdH;�?H;�H;��G;�G;|.G;�LF;�^D;_@;�N9;J�,;8�;���:�A�:0m9��K/��ۙ����P�!�qT�py���
��-"��Wμ�߼���       噼4`��q��oy���;k��I�W�$��� �������|�Z��$T� [�9�A�:`��:'�;%�);37;��>;�tC;5�E;�F;vG;D�G;��G;1,H;�SH;�sH;��H;��H;A�H;��H;��H;j�H;��H;'�H;�H;%�H;��H;j�H;��H;��H;A�H;��H;��H;�sH;�SH;3,H;��G;@�G;
vG;�F;4�E;�tC;��>;47;$�);%�;`��:�A�: [�9�$T�Z���|������� �W�$��I��;k�oy��q��5`��      �J;���7��9.�%���&����t���,M����4���º�uƹQ:���:���:'�;��(;��5;��=;��B;�[E;d�F;UG;ѩG;��G;�H;�CH;DfH;��H;��H;$�H;��H;��H;��H;��H;,�H;n�H;U�H;l�H;,�H;��H;��H;��H;��H;$�H;��H;��H;@fH;�CH;�H;��G;̩G;UG;`�F;�[E;��B;��=;��5;��(;'�;���:���:Q:�uƹ��º��4�,M��t�����軳&�%���9.���7�      ^�ͻBSɻ۴��nϨ��-���\c�+�$�Ƀ˺�P(�N@9L�k:Y��:w;8�;(�);��5;^�=;7QB;�E;�F;J8G;f�G;v�G;�	H;�5H;�YH;uwH;	�H;�H;�H;żH;��H;��H;U�H;��H;��H;W�H;��H;��H;W�H;��H;��H;żH;�H;�H;	�H;qwH;�YH;�5H;�	H;o�G;f�G;I8G;�F;�E;:QB;]�=;��5;&�);8�;v;Y��:H�k: N@9�P(�̃˺+�$��\c��-��nϨ�ܴ��HSɻ      �4��K/�kV�f,���˺M퀺`vƹpm9�nQ:���:���:��;��;F�,;37;��=;4QB;��D;�cF;D$G;�G;�G;�G;�)H;�NH;nH;�H;��H;Z�H;F�H;F�H;�H;��H;�H;��H;��H;G�H;��H;��H;�H;��H;�H;D�H;C�H;W�H;��H;
�H;nH;�NH;�)H; �G;�G;�G;F$G;�cF;��D;4QB;��=;37;H�,;��;��;���:���:�nQ:`m9`vƹD퀺��˺f,�lV��K/�      XW�hyƹ�1p�  �6�X�9�t,:N��:6ٶ:�L�:D�;�;�(&;L.1;�N9;��>;��B;�E;�cF;G;W�G;�G;��G;� H;FH;�eH;�H;�H;�H;�H;��H;D�H;�H;��H;��H;!�H;x�H;��H;x�H;!�H;��H;��H;�H;A�H;��H;�H;�H;�H;�H;�eH;FH;� H;��G;�G;W�G;G;�cF;�E;��B;��>;�N9;L.1;�(&;�;C�;�L�:4ٶ:P��:�t,:�X�9  �6�1p�hyƹ      "��:觎:A�:-��:���:��:�&�:v�;�;�f$;V>.;�#6;(<;Y@;�tC;�[E;�F;@$G;S�G;�G;G�G;�H;
@H;�_H;%zH;��H;S�H;�H;h�H;��H;��H;��H;��H;��H;�H;0�H;��H;0�H;
�H;��H;��H;��H;��H;��H;a�H;�H;P�H;��H;%zH;�_H;@H;�H;D�G;�G;R�G;B$G;�F;�[E;�tC;Y@;(<;�#6;W>.;�f$;�;x�;�&�:��:���:-��:A�:ا�:      /;�/;
x;�
; 9;�;�� ;`(;܊/;��5;&
;;�%?;�5B;�^D;4�E;c�F;I8G;�G;�G;I�G;�H;�<H;�[H;vH;��H;��H;n�H;s�H;��H;��H;��H;��H;A�H;��H;��H;��H;�H;��H;��H;��H;?�H;��H;��H;��H;��H;p�H;l�H;��H;��H;vH;�[H;�<H;�H;I�G;�G;�G;G8G;c�F;3�E;�^D;�5B;�%?;%
;;��5;ߊ/;
`(;�� ;��;9;�
;x;�/;      ��#;�f$;^(&;Y�(;�h,;�_0;b4;$�8;�'<;�N?;��A;��C;�NE;�LF;�F;UG;h�G;�G;��G;�H;�<H;�ZH;tH;-�H;ӚH;��H;�H;��H;��H;M�H;t�H;g�H;��H;��H;!�H;�H;I�H;�H;!�H;��H;��H;e�H;t�H;G�H;��H;��H;�H;��H;՚H;(�H;tH;�ZH;�<H;�H;��G;�G;e�G;UG;�F;�LF;�NE;��C;��A;�N?;�'<;$�8;b4;�_0;i,;Y�(;[(&;�f$;      L�6;�7;]�7;uN9;�	;;��<;��>;��@;�B;^D;�AE;�#F;4�F;.G;vG;ѩG;q�G;�G;� H;@H;�[H;tH;i�H;��H;%�H;^�H;6�H;[�H;1�H;Y�H;��H;��H;y�H;b�H;o�H;&�H;g�H;&�H;n�H;b�H;w�H;��H;��H;U�H;-�H;X�H;2�H;^�H;%�H;��H;h�H;tH;�[H;@H;� H;�G;p�G;ΩG;vG;.G;5�F;�#F;�AE;^D;�B;��@;��>;��<;�	;;uN9;]�7;�7;      "[@;�~@;C�@;��A; QB;�1C;bD;��D;�E;�LF;y�F;$G;QfG;�G;C�G;��G;�	H;�)H;FH;�_H;vH;*�H;��H;��H;n�H;P�H;_�H;��H;��H;��H;B�H;��H;�H;��H;��H;/�H;x�H;/�H;��H;��H;	�H;��H;@�H;��H;��H;��H;^�H;P�H;n�H;��H;��H;*�H;vH;�_H;FH;�)H;�	H;��G;A�G;�G;QfG;$G;y�F;�LF;�E;��D;`D;�1C;	QB;��A;B�@;�~@;      a�D;o�D;E;�NE;��E;�E;�[F;�F;�F;";G;6mG;L�G;�G;��G;��G;�H;�5H;�NH;�eH;,zH;��H;ؚH;*�H;v�H;ؼH;��H;`�H;��H;.�H;��H;��H;��H;��H;��H;��H;(�H;D�H;%�H;��H;��H;��H;��H;��H;��H;*�H;��H;\�H;��H;ؼH;t�H;'�H;ؚH;��H;,zH;�eH;�NH;�5H;�H;��G;��G;�G;M�G;6mG; ;G;�F;�F;�[F;�E;��E;�NE;E;o�D;      �F;��F;�F;i�F;� G;�#G;�FG;shG;��G;ΤG;��G;��G;`�G;�H;0,H;�CH;�YH;nH;�H;��H;��H;��H;[�H;P�H;��H;)�H;l�H;��H;J�H;U�H;��H;=�H;��H;��H;��H;��H;��H;��H;��H;��H;��H;=�H;��H;S�H;I�H;��H;k�H;(�H;��H;M�H;Z�H;��H;��H;��H;�H;nH;�YH;�CH;.,H;�H;a�G;��G;��G;ͤG;��G;qhG;�FG;�#G;� G;i�F;�F;��F;      �lG;�nG;tuG;�G;�G;l�G;��G;��G;��G;�G;��G;�H;"+H;�?H;�SH;DfH;uwH;
�H;�H;U�H;o�H;�H;6�H;c�H;Y�H;o�H;��H;�H;��H;a�H;U�H;��H;��H;��H;7�H;��H;��H;��H;6�H;��H;��H;��H;S�H;_�H;��H;�H;��H;n�H;Y�H;a�H;3�H;�H;l�H;U�H;�H;�H;uwH;DfH;�SH;�?H;"+H;�H;��G;�G;��G;��G;��G;j�G;��G;�G;tuG;�nG;      ��G;�G;P�G;��G;��G;6�G;2�G;�H;bH;�!H;�2H;]CH;TH;MdH;�sH;��H;�H;��H;�H;�H;r�H;��H;[�H;��H;��H;��H;�H;��H;F�H;�H;��H;��H;��H;r�H;��H;��H;P�H;��H;��H;r�H;��H;��H;��H;	�H;D�H;��H;�H;��H;��H;��H;X�H;��H;o�H;�H;�H;��H;�H;��H;�sH;JdH;TH;]CH;�2H;�!H;cH;�H;2�G;6�G;�G;��G;O�G;'�G;      �H;[H;�H;�H;�H;E H;9*H;f5H;pAH;NH;[H;hH;uH;G�H;��H;��H;�H;Y�H;�H;h�H;��H;��H;/�H;��H;'�H;L�H;��H;F�H;�H;��H;��H;��H;m�H;��H;L�H;��H;��H;��H;L�H;��H;j�H;��H;��H;��H;�H;F�H;��H;J�H;(�H;��H;-�H;��H;��H;h�H;�H;Y�H;�H;��H;��H;G�H;uH;hH;[H;NH;sAH;e5H;9*H;E H;�H;�H;�H;QH;      �:H;�;H;>H;�AH;>GH;�MH;�UH;"^H;GgH;�pH;�zH;��H;T�H;��H;��H;(�H;�H;B�H;��H;��H;��H;J�H;V�H;��H;��H;R�H;_�H;
�H;��H;��H;��H;c�H;��H;l�H;��H;��H;��H;��H;��H;l�H;��H;c�H;��H;��H;��H;
�H;^�H;P�H;��H;��H;U�H;J�H;��H;��H;��H;B�H;�H;'�H;��H;��H;T�H;��H;�zH;�pH;IgH;%^H;�UH;�MH;:GH;�AH;>H;�;H;      �bH;�cH;�eH;lhH;�lH;iqH;0wH;�}H;��H;H;�H;��H;��H;B�H;E�H;ǶH;̼H;D�H;D�H;��H;��H;t�H;��H;D�H;��H;��H;S�H;��H;��H;��H;x�H;��H;`�H;��H;��H;'�H;I�H;'�H;��H;��H;]�H;��H;v�H;��H;��H;��H;R�H;��H;��H;D�H;��H;t�H;��H;��H;D�H;D�H;ʼH;ŶH;E�H;@�H;��H;��H;�H;ċH;��H;�}H;0wH;jqH;�lH;nhH;�eH;�cH;      +�H;��H;�H;'�H;<�H;�H;4�H;'�H;m�H;�H;ǥH;��H;U�H;ӶH;�H; �H;��H;�H;�H;��H;��H;j�H;��H; �H;��H;=�H;��H;��H;��H;d�H;��H;v�H;��H;$�H;J�H;w�H;f�H;v�H;J�H;$�H;��H;v�H;��H;e�H;��H;��H;��H;:�H;��H; �H;��H;j�H;��H;��H;�H;�H;��H;��H;�H;ӶH;U�H;��H;ǥH;�H;n�H;$�H;4�H;�H;;�H;&�H;�H;��H;      ^�H;��H;��H;r�H;ќH;��H;�H;��H; �H;\�H;ƳH; �H;��H;��H;��H;��H;��H;��H;��H;��H;H�H;��H;z�H;�H;��H;��H;��H;��H;q�H; �H;a�H;��H;2�H;L�H;��H;��H;i�H;��H;��H;L�H;/�H;��H;a�H;�H;r�H;��H;��H;��H;��H;�H;w�H;��H;F�H;��H;��H;��H;��H;��H;��H;��H;~�H;�H;ƳH;]�H;�H;�H;�H;��H;ʜH;r�H;��H;��H;      n�H;��H;z�H;�H;ЫH;�H;��H;��H;϶H;$�H;��H;(�H;��H;�H;n�H;��H;\�H;�H;��H;��H;��H;��H;c�H;��H;��H;��H;��H;q�H;��H;l�H;��H;$�H;D�H;��H;��H;��H;��H;��H;��H;��H;C�H;&�H;��H;n�H;��H;q�H;��H;��H;��H;��H;b�H;��H;��H;��H;��H;�H;[�H;��H;n�H;�H;��H;(�H;��H;$�H;϶H;��H;��H;�H;ƫH;�H;|�H;��H;      �H;T�H;�H;
�H;��H;`�H;��H;�H;��H;z�H;k�H;^�H; �H;��H;��H;5�H;��H;��H;$�H;�H;��H;%�H;o�H;��H;��H;��H;3�H;��H;L�H;��H;��H;M�H;��H;��H;��H;��H;��H;��H;��H;��H;��H;P�H;��H;��H;M�H;��H;2�H;��H;��H;��H;n�H;$�H;��H;�H;$�H;��H;��H;5�H;��H;��H; �H;^�H;i�H;{�H;��H;�H;��H;d�H;}�H;�H;�H;K�H;      �H;`�H;�H;׹H;D�H;ʼH;��H;��H;7�H;��H;8�H;��H;6�H;��H;+�H;u�H;��H;��H;~�H;:�H;��H;�H;)�H;6�H;!�H;��H;��H;��H;��H;��H;&�H;x�H;��H;��H;��H;��H;��H;��H;��H;��H;��H;{�H;&�H;��H;��H;��H;��H;��H;"�H;5�H;)�H;�H;��H;:�H;~�H;��H;��H;u�H;)�H;��H;6�H;��H;8�H;��H;7�H;��H;��H;μH;7�H;عH;��H;W�H;      �H;Y�H;��H;��H;�H;��H;d�H;q�H;��H;��H;N�H;��H;Y�H;��H;�H;_�H;]�H;?�H;��H;��H;�H;N�H;g�H;~�H;@�H;��H;��H;T�H;��H;��H;J�H;l�H;h�H;��H;��H;��H;��H;��H;��H;��H;e�H;m�H;J�H;��H;��H;T�H;��H;��H;@�H;{�H;g�H;N�H;�H;��H;��H;@�H;\�H;_�H;�H;��H;Y�H;��H;N�H;��H;��H;n�H;d�H;��H;�H;��H;��H;Q�H;      �H;a�H;�H;عH;D�H;ʼH;��H;��H;7�H;��H;8�H;��H;6�H;��H;)�H;u�H;��H;��H;~�H;:�H;��H;�H;)�H;6�H;"�H;��H;��H;��H;��H;��H;&�H;x�H;��H;��H;��H;��H;��H;��H;��H;��H;��H;{�H;&�H;��H;��H;��H;��H;��H;!�H;5�H;)�H;�H;��H;:�H;~�H;��H;��H;u�H;)�H;��H;6�H;��H;:�H;��H;9�H;��H;��H;μH;7�H;عH;�H;V�H;      �H;T�H;�H;
�H;��H;`�H;��H;�H;��H;z�H;h�H;^�H; �H;��H;��H;5�H;��H;��H;$�H;�H;��H;$�H;n�H;��H;��H;��H;3�H;��H;L�H;��H;��H;M�H;��H;��H;��H;��H;��H;��H;��H;��H;��H;Q�H;��H;��H;M�H;��H;2�H;��H;��H;��H;o�H;%�H;��H;�H;$�H;��H;��H;5�H;��H;��H; �H;^�H;i�H;{�H;��H;�H;��H;c�H;~�H;
�H;�H;K�H;      o�H;��H;|�H;�H;ЫH;�H;��H;��H;϶H;$�H;��H;(�H;��H;�H;n�H;��H;\�H;�H;��H;��H;��H;��H;b�H;��H;��H;��H;��H;q�H;��H;l�H;��H;#�H;D�H;��H;��H;��H;��H;��H;��H;��H;C�H;'�H;��H;n�H;��H;q�H;��H;��H;��H;��H;c�H;��H;��H;��H;��H;�H;[�H;��H;n�H;�H;��H;(�H;��H;$�H;ѶH;��H;��H;�H;ūH;�H;}�H;��H;      a�H;��H;��H;t�H;МH;��H;�H;�H;�H;\�H;ƳH;�H;~�H;��H;��H;��H;��H;��H;��H;��H;I�H;��H;z�H;�H;��H;��H;��H;��H;q�H; �H;a�H;��H;1�H;J�H;��H;��H;i�H;��H;��H;J�H;/�H;��H;a�H;�H;r�H;��H;��H;��H;��H;�H;y�H;��H;F�H;��H;��H;��H;��H;��H;��H;��H;~�H; �H;ƳH;]�H; �H;�H;�H;��H;ǜH;t�H;��H;��H;      +�H;��H;�H;$�H;<�H;�H;7�H;'�H;m�H;�H;ǥH;��H;U�H;ӶH;�H;��H;��H;�H;�H;��H;��H;j�H;��H; �H;��H;;�H;��H;��H;��H;d�H;��H;v�H;��H;$�H;J�H;w�H;f�H;v�H;J�H;$�H;��H;w�H;��H;e�H;��H;��H;��H;;�H;��H; �H;��H;j�H;��H;��H;�H;�H;��H; �H;�H;ӶH;T�H;��H;ǥH;�H;n�H;$�H;7�H;�H;:�H;$�H;�H;��H;      �bH;�cH;�eH;nhH;�lH;iqH;0wH;�}H;��H;H;�H;��H;��H;B�H;E�H;ǶH;ʼH;C�H;D�H;��H;��H;t�H;��H;F�H;��H;��H;R�H;��H;��H;��H;v�H;��H;^�H;��H;��H;'�H;I�H;'�H;��H;��H;]�H;��H;x�H;��H;��H;��H;S�H;��H;��H;D�H;��H;t�H;��H;��H;D�H;D�H;ʼH;ǶH;E�H;B�H;��H;��H;�H;ċH;��H;�}H;0wH;lqH;�lH;lhH;�eH;�cH;      �:H;�;H;>H;�AH;9GH;�MH;�UH;%^H;HgH;�pH;�zH;��H;T�H;��H;��H;'�H;�H;A�H;��H;��H;��H;J�H;V�H;��H;��H;R�H;_�H;
�H;��H;��H;��H;a�H;��H;k�H;��H;��H;��H;��H;��H;l�H;��H;d�H;��H;��H;��H;
�H;^�H;P�H;��H;��H;U�H;J�H;��H;��H;��H;C�H;�H;*�H;��H;��H;T�H;��H;�zH;�pH;IgH;%^H;�UH;�MH;7GH;�AH;>H;�;H;      �H;XH;�H;�H;�H;? H;<*H;h5H;qAH;NH;[H;hH;uH;G�H;��H;��H;�H;W�H;�H;j�H;��H;��H;.�H;��H;(�H;L�H;��H;F�H;�H;��H;��H;��H;k�H;��H;J�H;��H;��H;��H;L�H;��H;k�H;��H;��H;��H;�H;F�H;��H;J�H;'�H;��H;.�H;��H;��H;h�H;�H;Z�H;�H;��H;��H;G�H;uH;hH;[H;NH;sAH;f5H;<*H;C H;�H;�H;�H;XH;      ��G;�G;P�G;��G;��G;6�G;2�G;�H;bH;�!H;�2H;]CH;TH;MdH;�sH;��H;	�H;�H;�H;�H;u�H;��H;Y�H;��H;��H;��H;�H;��H;F�H;�H;��H;��H;��H;q�H;��H;��H;P�H;��H;��H;r�H;��H;��H;��H;
�H;D�H;��H;�H;��H;��H;��H;Y�H;��H;o�H;�H;�H;��H;�H;��H;�sH;JdH;TH;]CH;�2H;�!H;cH;�H;2�G;3�G;�G;��G;P�G;(�G;      �lG;�nG;wuG;�G;�G;g�G;��G;��G;��G;�G;��G;�H;"+H;�?H;�SH;FfH;vwH;
�H;�H;W�H;r�H;�H;5�H;b�H;Y�H;o�H;��H;�H;��H;a�H;S�H;��H;��H;��H;6�H;��H;��H;��H;7�H;��H;��H;��H;U�H;_�H;��H;�H;��H;o�H;Y�H;b�H;5�H;�H;l�H;U�H;�H;�H;twH;DfH;�SH;�?H;"+H;�H;��G;�G;��G;��G;��G;f�G;�G;�G;tuG;�nG;      �F;��F;�F;j�F;� G;�#G;�FG;thG;��G;ΤG;��G;��G;a�G;�H;.,H;�CH;�YH;	nH;�H;��H;��H;��H;[�H;N�H;��H;)�H;k�H;��H;J�H;U�H;��H;;�H;��H;��H;��H;��H;��H;��H;��H;��H;��H;>�H;��H;R�H;I�H;��H;k�H;)�H;��H;P�H;[�H;��H;��H;��H;�H;nH;�YH;�CH;0,H;�H;`�G;��G;��G;ͤG;��G;qhG;�FG;�#G;� G;j�F;�F;��F;      a�D;q�D;E;�NE;��E;�E;�[F;�F;�F;";G;8mG;M�G;�G;��G;��G;�H;�5H;�NH;�eH;,zH;��H;ؚH;*�H;v�H;ؼH;��H;]�H;��H;-�H;��H;��H;��H;��H;��H;��H;%�H;D�H;(�H;��H;��H;��H;��H;��H;��H;+�H;��H;]�H;��H;ؼH;u�H;'�H;ؚH;��H;.zH;�eH;�NH;�5H;�H;��G;��G;�G;L�G;6mG; ;G;�F;�F;�[F;�E;��E;�NE;E;o�D;      ([@;�~@;F�@;��A;�PB;�1C;_D;��D;�E;�LF;z�F;$G;RfG;�G;A�G;��G;�	H;�)H;FH;�_H;vH;*�H;��H;��H;n�H;P�H;_�H;��H;��H;��H;@�H;��H;�H;��H;��H;/�H;x�H;/�H;��H;��H;�H;��H;B�H;��H;��H;��H;_�H;P�H;n�H;��H;��H;*�H;vH;�_H;FH;�)H;�	H;��G;C�G;�G;QfG;$G;w�F;�LF;�E;��D;_D;�1C;QB;��A;D�@;�~@;      F�6;�7;m�7;uN9;�	;;��<;��>;��@;�B;^D;�AE;�#F;4�F;.G;vG;ϩG;q�G;�G;� H;@H;�[H;tH;i�H;��H;%�H;]�H;5�H;X�H;.�H;X�H;��H;��H;y�H;b�H;n�H;&�H;g�H;&�H;o�H;b�H;w�H;��H;��H;V�H;.�H;[�H;5�H;^�H;%�H;��H;h�H;tH;�[H;@H;� H;�G;q�G;ѩG;vG;~.G;2�F;�#F;�AE;[D;�B;��@;��>;��<;�	;;tN9;a�7;�7;      ��#;�f$;^(&;Y�(;�h,;�_0;b4;%�8;�'<;�N?;��A;��C;�NE;�LF;�F;UG;e�G;�G;��G;�H;�<H;�ZH;tH;-�H;՚H;��H;�H;��H;��H;K�H;t�H;g�H;��H;��H;!�H;�H;I�H;�H;!�H;��H;��H;g�H;t�H;H�H;��H;��H;�H;��H;ӚH;*�H;tH;�ZH;�<H;�H;��G;�G;f�G;UG;�F;�LF;�NE;��C;��A;�N?;�'<;$�8;b4;�_0;i,;Y�(;\(&;�f$;      ';�/;x;�
; 9;�;�� ;`(;܊/;��5;(
;;�%?;�5B;�^D;3�E;c�F;I8G;�G;�G;H�G;�H;�<H;�[H;vH;��H;��H;n�H;p�H;��H;��H;��H;��H;A�H;��H;��H;��H;�H;��H;��H;��H;A�H;��H;��H;��H;��H;s�H;l�H;��H;��H;vH;�[H;�<H;�H;I�G;�G;�G;G8G;c�F;4�E;�^D;�5B;�%?;&
;;��5;ފ/;`(;�� ;��;9;�
;x;�/;       ��:꧎:A�:)��:���:��:�&�:x�;�;�f$;W>.;�#6;(<;Y@;�tC;�[E;�F;@$G;R�G;�G;H�G;�H;@H;�_H;%zH;��H;S�H;�H;g�H;��H;��H;��H;��H;��H;
�H;1�H;��H;1�H;�H;��H;��H;��H;��H;��H;c�H;�H;Q�H;��H;%zH;�_H;@H;�H;E�G;�G;S�G;B$G;�F;�[E;�tC;Y@;(<;�#6;T>.;�f$;�;x�;�&�:��:���:)��:A�:֧�:      XW�pyƹ�1p�  �6�X�9�t,:P��:4ٶ:�L�:C�;�;�(&;L.1;�N9;��>;��B;�E;�cF;G;V�G;�G;��G;� H;FH;�eH;�H;�H;�H;�H;��H;A�H;	�H;��H;��H; �H;x�H;��H;x�H;!�H;��H;��H;�H;D�H;��H;�H;�H;�H;�H;�eH;FH;� H;��G;�G;Y�G;G;�cF;�E;��B;��>;�N9;L.1;�(&;�;D�;�L�:4ٶ:N��:�t,:�X�9  �6�1p�hyƹ       �4��K/�jV�f,���˺Q퀺`vƹpm9�nQ:���:���:��;��;E�,;37;��=;4QB;��D;�cF;D$G;�G;�G;�G;�)H;�NH;nH;�H;��H;Z�H;E�H;D�H;�H;��H;�H;��H;��H;G�H;��H;��H;�H;��H;�H;F�H;E�H;Y�H;��H;
�H;nH;�NH;�)H; �G;�G;��G;F$G;�cF;��D;3QB;��=;37;F�,;��;��;���:���:�nQ:Pm9`vƹF퀺��˺f,�lV��K/�      _�ͻBSɻ۴��nϨ��-���\c�+�$�Ƀ˺�P(� N@9L�k:Y��:v;8�;&�);��5;^�=;6QB;�E;�F;J8G;f�G;s�G;�	H;�5H;�YH;uwH;	�H;�H;�H;żH;��H;��H;W�H;��H;��H;W�H;��H;��H;W�H;��H;��H;żH;�H;�H;	�H;rwH;�YH;�5H;�	H;p�G;f�G;I8G;�F;�E;9QB;^�=;��5;(�);8�;w;Y��:L�k: N@9�P(�̃˺,�$��\c��-��nϨ�ܴ��HSɻ      �J;���7��9.�%���&����t���,M����4���º�uƹQ:���:���:'�;��(;��5;��=;��B;�[E;a�F;UG;ΩG;��G;�H;�CH;CfH;��H;��H;$�H;��H;��H;��H;��H;,�H;l�H;U�H;n�H;,�H;��H;��H;��H;��H;$�H;��H;��H;AfH;�CH;�H;��G;ΩG;UG;c�F;�[E;��B;��=;��5;��(;'�;���:���:Q:�uƹ��º��4�,M��t�����軳&�%���9.���7�       噼4`��q��oy���;k��I�W�$��� �������|�Z��$T� [�9�A�:`��:%�;%�);17;��>;�tC;4�E;�F;vG;D�G;��G;1,H;�SH;�sH;��H;��H;A�H;��H;��H;j�H;��H;%�H;�H;'�H;��H;k�H;��H;��H;A�H;��H;��H;�sH;�SH;3,H;��G;@�G;vG;�F;5�E;�tC;��>;57;$�);'�;`��:�A�: [�9�$T�Z���|������� �W�$��I��;k�oy��q��5`��      ������߼Wμ-"���
��py��qT�P�!�����ۙ��K/�� m9�A�:���:8�;I�,;�N9;]@;�^D;�LF;.G;�G;��G;�H;�?H;IdH;G�H;��H;;�H;˶H;��H;�H;��H;��H;��H;��H;��H;
�H;��H;̶H;;�H;��H;G�H;IdH;�?H;�H;��G;�G;|.G;�LF;�^D;_@;�N9;J�,;8�;���:�A�: m9��K/��ۙ����P�!�qT�oy���
��-"��Xμ�߼���      ��/�N-�l.%����������Ǽܫ����{��J;��C�IϨ�bO:�� [�9���:v;��;K.1;(<;�5B;�NE;5�F;VfG;
�G;`�G;"+H;TH;uH;N�H;�H;P�H;~�H;��H;�H;.�H;T�H;.�H;�H;��H;}�H;P�H;�H;N�H; uH;TH;+H;e�G;�G;QfG;2�F;�NE;�5B;(<;K.1;��;u;���: [�9�bO:�IϨ��C��J;���{�ܫ���Ǽ��������l.%�N-�      f@{�``w��l��yZ�Y�C�kg*�������+"��`O���I�H|�IϨ��K/��$T�
Q:W��:��;�(&;�#6;�%?;��C;�#F;$G;F�G;��G;�H;WCH;hH;��H;��H;��H;�H;#�H;U�H;��H;��H;��H;S�H;#�H;�H;��H;��H;��H;hH;WCH;�H;��G;J�G;$G;�#F;��C;�%?;�#6;�(&;��;Q��:Q:�$T��K/�IϨ�H|��I�`O��+"����鼴��kg*�Y�C��yZ��l�``w�      �b��ꪫ��ƣ��s���ɇ��l�JG���"�n� �8aļj���I��C��ۙ�[��uƹD�k:���:�;W>.;%
;;��A;�AE;z�F;5mG;��G;��G;�2H;[H;�zH;
�H;��H;ĳH;��H;a�H;.�H;D�H;.�H;a�H;��H;³H;��H;
�H;�zH;[H;�2H;��G;��G;9mG;v�F;�AE;��A;(
;;V>.;�;���:<�k:�uƹ[��ۙ��C��I�j��8aļn� ���"�JG��l��ɇ��s���ƣ�ꪫ�      ������uݽ�2̽�ж����������yZ�N-�۷�8aļaO���J;���軚�|���º�M@9���:B�;�f$;��5;�N?;^D;�LF; ;G;ͤG;�G;�!H;NH;�pH;��H;�H;Z�H; �H;t�H;��H;��H;��H;t�H; �H;Y�H;�H;��H;�pH;NH;�!H;�G;ΤG;#;G;�LF;\D;�N?;��5;�f$;B�;���:�M@9��º��|�����J;�aO��8aļ۷�N-��yZ����������ж��2̽uݽ���      S,����Z�>��z�XvϽ�b��2I��n]a�M-�n� �+"����{�Q�!�������4��P(��nQ:�L�:�;ۊ/;�'<;�B;�E;�F;��G;��G;\H;oAH;:gH;|�H;g�H;��H;ȶH;��H;)�H;��H;)�H;��H;ȶH;��H;g�H;|�H;:gH;lAH;_H;��G;��G;	�F;�E;��B;�'<;ފ/;�;�L�:�nQ:�P(���4�����Q�!���{�+"��n� �M-�n]a�2I���b��XvϽ�z�>��Z���      *G�t�C��$:��J+��� ��tݽb���2I���yZ���"����ܫ��rT��� �,M��̃˺pm94ٶ:x�;`(;�8;��@;��D; �F;shG;��G;�H;c5H;^H;�}H;�H;�H;��H;��H;��H;i�H;��H;��H;��H;�H;�H;�}H;^H;a5H;�H;��G;qhG;�F;��D;��@;�8;`(;v�;4ٶ:�m9Ѓ˺,M���� �rT�ܫ�������"��yZ�2I��b���tݽ �����J+��$:�t�C�      {x�	9t���g���T��G=�~#�6�tݽ�b������JG�����Ǽpy��W�$�x���2�$�hvƹ@��:�&�:�� ;T4;��>;YD;�[F;�FG;��G;*�G;3*H;UH;&wH;.�H;�H;��H;��H;��H;[�H;��H;��H;��H;�H;.�H;&wH;~UH;2*H;*�G;��G;�FG;�[F;WD;��>;T4;�� ;�&�:@��:`vƹ5�$�x���W�$�py���Ǽ���JG������b��tݽ6�~#��G=���T���g�	9t�      ���Oa��$���C�c�t�C�~#�!��XvϽ�����l�kg*����
���I�����\c�9퀺�t,:��:�;�_0;��<;�1C;�E;�#G;f�G;3�G;A H;�MH;eqH;ۋH;��H;�H;`�H;̼H;��H;μH;^�H;�H;��H;ދH;eqH;�MH;> H;3�G;e�G;�#G;�E;�1C;��<;�_0;�;��:�t,:6퀺�\c�����I��
�����kg*��l�����XvϽ!��~#�t�C�C�c�$���Oa����      l*��j����Ƥ���/��C�c��G=����zｖж��ɇ�Y�C���."���;k��&��-����˺�X�9���: 9;�h,;�	;;�PB;��E;� G;�G;��G;�H;,GH;|lH;4�H;ǜH;īH;m�H;2�H;�H;2�H;l�H;ūH;ƜH;5�H;|lH;)GH;�H;��G;�G;� G;��E;�PB;�	;;�h,;9;���:�X�9��˺�-���&��;k�."����Y�C��ɇ��ж��z����G=�C�c��/����Ƥ�j���      ��ɾ�ž+��tת��#�����T��J+�>��2̽�s���yZ����Xμoy��&��mϨ�l,� ��6%��:�
;[�(;xN9;��A;�NE;f�F;�G;��G;�H;�AH;^hH;�H;j�H;�H;�H;ҹH;��H;ҹH;�H;�H;i�H;�H;`hH;�AH;�H;��G;�G;f�F;�NE;��A;|N9;^�(;�
;%��: ��6l,�nϨ�%��oy��Xμ����yZ��s���2̽>��J+���T�#����tת�+���ž      X_ݾ�:پ�V;+���Ƥ�Oa����g��$:��Z�uݽ�ƣ��l�m.%��߼q���9.�ܴ��pV�p2p�A�:�w;H(&;U�7;6�@;E;�F;suG;E�G;�H;�=H;xeH;��H;��H;}�H;�H;�H;�H;�H;�H;~�H;��H;��H;xeH;�=H;�H;E�G;suG;�F;E;2�@;Y�7;J(&; x;A�:p2p�nV�ݴ���9.�q���߼m.%��l��ƣ�uݽ�Z��$:���g�Oa���Ƥ�+���V;�:پ      
^�7���:پ�žj�����	9t�t�C������ꪫ�``w�N-����4`����7�HSɻ�K/�xyƹ§�:�/;�f$;�7;�~@;g�D;��F;�nG;�G;ZH;�;H;�cH;��H;��H;��H;=�H;W�H;O�H;W�H;?�H;��H;��H;��H;�cH;�;H;WH;�G;�nG;��F;g�D;�~@;�7;�f$;�/;���:xyƹ�K/�ISɻ��7�4`�����N-�``w�ꪫ������t�C�	9t���j����ž�:پ7��      IF�Zh����YVھ:�������~���S��#��o��=S��t₽9�6�{���ry��dFB��Eֻ�A?��	�Y�:z��:c�";�46;V@;y�D;ɩF;�nG;�G;2H;.@H;gH;y�H;Y�H;��H;�H;��H;�H;��H;�H;��H;X�H;z�H;gH;-@H;/H;�G;�nG;ʩF;y�D;S@;�46;c�";~��:}Y�:�	��A?��EֻdFB�ry��{���9�6�t₽=S���o���#��S��~������:��YVھ��Zh��      Zh���b���쾪*־�v��,���*��+�O�Y� �s��r���؀�N�3���Hݜ�J�>�c�ѻ �9�X���4o�:(% ;oM#;h�6;GA@;�D;ïF;qG;n�G;GH;�@H;�gH;�H;��H;�H;F�H;"�H;�H;"�H;H�H;�H;��H;�H;�gH;�@H;DH;n�G;qG;ïF;�D;CA@;n�6;oM#;(% ;0o�:X�����9�e�ѻJ�>�Iݜ���N�3��؀��r��s�Y� �+�O�*��,����v���*־���b��      ���쾷�޾25ʾP;���:��-�v��E�c'����v����u���+��W��A����4���Ļ>9)��j���W�:N�;%;l7;"�@;�D;�F;�wG;x�G;jH;ZCH;UiH;F�H;��H;ΪH;�H;��H;��H;��H;�H;ΪH;��H;F�H;UiH;WCH;hH;x�G;�wG;�F;�D;�@;l7;%;N�;�W�:�j��=9)���Ļ��4��A���W缊�+���u�v�����c'��E�-�v��:��P;��25ʾ��޾��      YVھ�*־25ʾu��������M���9b��5�����ս����Xc���֖ռ�I��a�$�|T���Z�`^��"�:��;i�';C�8;RA;�9E;��F;̂G;�G;xH;%GH;<lH;z�H;c�H;�H;��H;��H;�H;��H;��H;�H;b�H;|�H;>lH;"GH;uH;�G;̂G;��F;�9E;RA;F�8;i�';��;�:�^���Z�}T��b�$��I��֖ռ���Xc������ս���5��9b��M������u���25ʾ�*־      :���v��P;������UP��J�r��H�X� ���:@��֓����K�g�־���s�~�����ܺ 4u9%&�:�;2�+;��:;�"B;��E;	�F;�G;�G;cH;VLH;&pH;o�H;��H;ѭH;j�H;�H;��H;�H;g�H;ЭH;��H;r�H;&pH;SLH;bH;�G;�G;�F;��E;�"B;��:;2�+;�;#&�:04u9�ܺ��~����s�־�g���K�֓��:@����X� ��H�J�r�VP������P;���v��      ����,����:���M��J�r�*�O�#,�[�
��gٽuĥ���u�~1�t���3Ϥ���P�[��.o��p��:}��:�P;D�/;\�<;
C;<�E;�!G;G�G;'�G;�%H;�RH;�tH;*�H;q�H;�H;5�H;��H;3�H;��H;5�H;�H;p�H;,�H;�tH;�RH;�%H;'�G;E�G;�!G;;�E;C;[�<;C�/;�P;y��::�p���.o�[򻹎P�3Ϥ�t���~1���u�uĥ��gٽ[�
�#,�*�O�J�r��M���:��,���      �~��*��-�v��9b��H�#,�PZ����<S��|^����N������μ�I��&+�'����.� ����j~:j��:)m;��3;>�>;F�C;dPF;�FG;g�G;�G;�/H;"ZH;�zH;y�H;��H;��H;R�H;W�H;�H;W�H;R�H;��H;��H;{�H;�zH;!ZH;�/H;�G;f�G;�FG;aPF;@�C;=�>;��3;+m;b��:�j~:����.�(���&+��I����μ�����N�|^��<S�����PZ�#,��H��9b�-�v�*��      �S�+�O��E��5�X� �[�
���罪9��,l���Xc���(��������[�����ݎ�fܺ`:9��:@�	;Gd';o 8;_�@;��D;�F;JjG;��G;uH;�:H;bbH;�H;7�H;^�H;v�H;��H;f�H;�H;f�H;��H;t�H;\�H;:�H;�H;bbH;�:H;uH;��G;HjG;	�F;��D;_�@;o 8;Gd';?�	;��:�:9gܺ�ݎ������[��������(��Xc�,l���9�����[�
�X� ��5��E�+�O�      �#�Y� �c'������gٽ<S��,l��V�j�J�3��i��վ�����(���Ļ{A?���B���@:�[�:Q;�.;��;;�tB;-�E;��F;X�G;�G;
H;�FH;IkH;��H;S�H;<�H;��H;>�H;��H;'�H;��H;>�H;��H;<�H;T�H;��H;GkH;�FH;
H;�G;X�G;��F;*�E;�tB;��;;�.;Q;�[�:��@:��B�{A?���Ļ(������վ��i�J�3�V�j�,l��<S���gٽ����c'�Y� �       p��s��罰�ս:@��uĥ�|^���Xc�J�3���	�ӌ˼�]��_FB�[򻽜���Ӻ@��8��:��;�M#;}=5;)?;q�C;�@F;/:G;�G;B�G;^'H;�RH;�tH;��H;��H;W�H;޻H;��H;��H;s�H;��H;��H;޻H;U�H;��H;��H;�tH;�RH;]'H;?�G;�G;,:G;�@F;p�C;)?;}=5;�M#;��;��: ��8�Ӻ����[�_FB��]��ӌ˼��	�J�3��Xc�|^��uĥ�:@����ս���s�      >S���r��v�����֓����u���N���(��i�Ҍ˼�A����P�qs��R|������\:*�:x�;�n-;��:;
�A;�,E;��F;VoG;�G;�H;�7H;o_H;0~H;�H;3�H;��H;A�H;��H;j�H;��H;j�H;��H;@�H;��H;5�H;�H;0~H;m_H;�7H;�H; �G;SoG;��F;�,E;
�A;�:;�n-;x�;.�:�\:����R|��qs���P��A��Ҍ˼�i���(���N���u�֓�����v���r��      t₽�؀���u��Xc���K�1�������վ��]����P����PT����9�L�o�d3�9y&�:^�	;h%;b�5;��>;��C;�F;�!G;ʚG;��G;mH;�HH;�kH;̇H;~�H;��H;޹H;��H;~�H;��H;�H;��H;��H;��H;޹H;ĭH;~�H;̇H;�kH;�HH;kH;��G;ǚG;�!G;�F;��C;��>;a�5;h%;a�	;w&�:l3�9H�o���9�PT�������P��]���վ�����~1���K��Xc���u��؀�      9�6�M�3���+���g�t�����μ�������^FB�ps�PT��B�D��{��:u9�q�:���:~Y;�t0;�;;�B;:E;�F;$hG;�G;5�G;�0H;�XH;[xH;P�H;��H;3�H;)�H;�H;E�H;]�H;k�H;]�H;D�H;�H;)�H;4�H;��H;N�H;ZxH;�XH;�0H;7�G;�G; hG;�F;:E;�B;�;;�t0;�Y;���:�q�::u9�{��@�D�PT��ps�^FB����������μt���h�����+�N�3�      z�����W�Ֆռ־�2Ϥ��I����[�(�[����9��{���:9FX�:[X�:FQ;E,;��8;�A@;%BD;�@F;�,G;��G;��G;�H;�DH;OhH;d�H;��H;��H;��H;T�H;Q�H;�H;��H;��H;��H;�H;N�H;T�H;��H;��H;��H;a�H;MhH;�DH;�H;��G;��G;�,G;�@F;%BD;�A@;��8;H,;FQ;[X�:HX�: ;9�{����9��[�(���[��I��2Ϥ�־�Ֆռ�W���      ry��Hݜ��A���I����s���P�&+������Ļ����R|�H�o�:u9DX�:�+�:\;�);݄6;��>;�PC;��E;�F;�xG;V�G;�H;�1H;FXH;3wH;�H;H�H;5�H;��H;K�H;u�H;��H;�H;��H;�H;��H;u�H;J�H;��H;5�H;E�H;��H;2wH;EXH;�1H;�H;S�G;�xG;�F;��E;�PC;��>;��6;�);\;�+�:DX�::u9L�o�R|�������Ļ���&+���P���s��I���A��Iݜ�      cFB�I�>���4�a�$�~��[�$����ݎ�zA?��Ӻ����l3�9�q�:WX�:^;��';�=5;��=;�B;@GE;l�F;�UG;L�G;	�G;�H;�HH;CjH;*�H;��H;y�H;e�H;x�H;�H;t�H;A�H;Q�H;��H;Q�H;A�H;q�H;�H;z�H;e�H;x�H;��H;*�H;@jH;�HH;�H;�G;H�G;�UG;i�F;=GE;�B;��=;�=5;��';^;[X�:�q�:l3�9�����ӺxA?��ݎ�$���[�~��a�$���4�K�>�      �Eֻ\�ѻ��Ļ|T�����.o��.�`ܺ��B����8�\:{&�:���:EQ;�);�=5;�:=;:#B;��D;vF;7G;�G;��G;�H;�:H;D^H;�zH;,�H;��H;��H;<�H;��H;��H;O�H;��H;^�H;��H;^�H;��H;Q�H;��H;��H;<�H;��H;��H;,�H;�zH;D^H;�:H;�H;��G;�G;7G;vF;��D;<#B;�:=;�=5;�);EQ;���:{&�:�\:���8��B�aܺ�.��.o���|T����Ļb�ѻ      �A?���9�99)��Z��ܺ�p�����p:9��@:��:0�:_�	;Y;D,;݄6;��=;8#B;��D;�XF;�!G;��G;H�G;�H;#/H;�SH;�qH;�H;�H;��H;�H;��H;�H;��H;�H;��H;N�H;��H;M�H;��H;�H;��H;�H;��H;�H;��H;�H;�H;�qH;�SH;/H;�H;G�G;��G;�!G;�XF;��D;7#B;��=;݄6;E,;Y;_�	;0�:��:��@:`:9����p���ܺ�Z�:9)��9�      �	�H���xj�� ^��04u9*:�j~:��:�[�:�;|�;j%;�t0;��8;��>;�B;��D;�XF;YG;��G;��G;��G;"&H;7KH;�iH;�H;��H;k�H;��H;;�H;��H;��H;��H;e�H;��H;�H;��H;�H;��H;e�H;��H;��H;��H;8�H;��H;k�H;��H;�H;�iH;3KH;&H;��G;��G;��G;YG;�XF;��D;�B;��>;��8;�t0;i%;|�;�;�[�:��:�j~:F:�4u9 ^���j��H���      �Y�:Zo�:�W�:&�:)&�:{��:h��:?�	;Q;�M#;�n-;a�5;�;;�A@;�PC;9GE;�uF;�!G;��G;��G;C�G;w H;<EH;�cH;o}H;��H;�H;ԱH;��H;��H;��H;_�H;��H;��H;�H;��H;!�H;��H;�H;��H;��H;`�H;��H;��H;�H;ұH;�H;��H;m}H;�cH;9EH;w H;@�G;��G;��G;�!G;�uF;9GE;�PC;�A@;�;;a�5;�n-;�M#;Q;@�	;f��:���:?&�:(�:�W�:Ho�:      ���:9% ;Y�;��;�;�P;/m;Hd';�.;�=5;�:;��>;�B;$BD;��E;i�F;7G;��G;��G;D�G;�H;BH;<`H;�yH;��H;V�H;��H;�H;��H;�H;��H;e�H;��H;r�H;&�H;�H;�H;�H;&�H;r�H;��H;f�H;��H; �H;|�H;�H;��H;V�H;��H;{yH;8`H;BH;�H;F�G;��G;��G;7G;i�F;��E;$BD;�B;��>;�:;~=5;�.;Gd';0m;�P;�;��;W�;)% ;      q�";�M#;%;f�';6�+;N�/;��3;{ 8;��;;-?;�A;ûC;:E;�@F;�F;�UG;�G;J�G;��G;| H;BH;�^H;ywH;O�H;��H;�H;·H;b�H;4�H;\�H;T�H;�H;��H;�H;��H;y�H;��H;y�H;��H;�H;��H;�H;T�H;V�H;.�H;a�H;��H;�H;��H;I�H;uwH;�^H;BH;| H;��G;K�G;�G;�UG;�F;�@F;:E;ûC;�A;/?;�;;{ 8;��3;P�/;N�+;f�';%;�M#;      �46;q�6;l7;=�8;��:;`�<;B�>;b�@;�tB;q�C;�,E;�F;
�F;�,G;�xG;J�G;��G;�H;!&H;@EH;;`H;{wH;c�H;h�H;{�H;�H;ͿH;��H;�H;2�H;`�H;t�H;��H;��H;��H;��H;��H;��H;��H;��H;��H;t�H;`�H;-�H;�H;��H;˿H;�H;|�H;g�H;`�H;xwH;5`H;@EH;!&H;�H;��G;H�G;�xG;�,G;�F;�F;�,E;p�C;�tB;b�@;B�>;b�<;��:;=�8;l7;d�6;      n@;YA@;.�@;RA;�"B;C;N�C;��D;/�E;�@F;��F;�!G;!hG;��G;T�G;�G;�H;#/H;4KH;�cH;{yH;M�H;g�H;��H;9�H;��H;��H;�H;F�H;��H;��H;��H;q�H;��H;��H;��H;��H;��H; �H;��H;n�H;��H;��H;��H;A�H;�H;��H;��H;;�H;��H;e�H;J�H;wyH;�cH;4KH;%/H;�H;�G;T�G;��G; hG;�!G;��F;�@F;0�E;��D;M�C;	C;�"B;RA;-�@;NA@;      ��D;�D; �D;�9E;��E;B�E;cPF;�F;��F;/:G;UoG;̚G;�G;��G;�H;�H;�:H;�SH;�iH;w}H;��H;��H;��H;B�H;m�H;�H;a�H;��H;��H;c�H;�H;=�H;��H;!�H;��H;U�H;��H;U�H;��H;�H;��H;=�H;�H;b�H;��H;��H;`�H;�H;n�H;?�H;��H;��H;��H;v}H;�iH;�SH;�:H;�H;�H;��G;�G;͚G;UoG;-:G;��F;�F;dPF;A�E;��E;�9E;��D;�D;      ۩F;ԯF;�F;��F;�F;�!G;�FG;JjG;W�G;�G;�G;��G;5�G;�H;�1H;�HH;C^H;�qH;�H;��H;S�H;�H;�H;��H;�H;C�H;S�H;��H;��H;��H;��H;��H;'�H;�H;��H;�H;B�H;�H;��H;�H;#�H;��H;��H;��H;��H;��H;Q�H;B�H;�H;��H;�H;�H;O�H;��H;�H;�qH;@^H;�HH;�1H;�H;5�G;��G;�G;�G;X�G;HjG;�FG;�!G;�F;��F;�F;˯F;      �nG;"qG;�wG;ӂG;�G;N�G;n�G;��G;�G;B�G;�H;qH;�0H;�DH;FXH;DjH;�zH;�H;��H;�H;��H;·H;̿H;��H;]�H;U�H;t�H;��H;��H;��H;��H;�H;�H;��H;k�H;��H;��H;��H;j�H;��H;�H;�H;��H;��H;��H;��H;s�H;S�H;]�H;��H;˿H;·H;��H;�H;��H;�H;�zH;CjH;FXH;�DH;�0H;qH;�H;B�G;�G;��G;o�G;K�G;�G;ӂG;�wG;!qG;      
�G;t�G;��G;�G;�G;*�G;�G;H;H;a'H;�7H;�HH;�XH;QhH;3wH;*�H;+�H;�H;h�H;ױH;�H;a�H;��H;�H;��H;��H;��H;q�H;��H;{�H;��H;��H;��H;��H;�H;:�H;M�H;:�H;�H;��H;��H;��H;��H;v�H;��H;q�H;��H;��H;��H;�H;��H;_�H;�H;ױH;h�H;�H;)�H;*�H;4wH;PhH;�XH;�HH;�7H;a'H;H;H;�G;,�G;�G;�G;��G;��G;      NH;JH;oH;~H;fH;�%H;�/H;�:H;�FH;�RH;o_H;lH;]xH;d�H;�H;��H;��H;��H;��H;��H;��H;2�H;�H;J�H;��H;��H;��H;��H;Y�H;��H;��H;��H;��H;�H;|�H;��H;��H;��H;|�H;�H;��H;��H;��H;��H;W�H;��H;��H;��H;��H;J�H;�H;1�H;�H;��H;��H;��H;��H;��H;�H;d�H;^xH; lH;o_H;�RH;�FH;�:H;�/H;�%H;mH;~H;mH;?H;      ?@H;AH;gCH;/GH;hLH;�RH;)ZH;kbH;SkH;�tH;<~H;ڇH;U�H;��H;K�H;|�H;��H;�H;8�H;��H;�H;Y�H;-�H;��H;Z�H;��H;��H;y�H;��H;��H;��H;��H;0�H;��H;��H;	�H;�H;	�H;��H;��H;-�H;��H;��H;��H;��H;x�H;��H;��H;[�H;��H;,�H;W�H;�H;��H;7�H;�H;��H;|�H;I�H;��H;U�H;ڇH;=~H;�tH;VkH;mbH;)ZH;�RH;eLH;-GH;cCH;AH;      gH;�gH;fiH;IlH;5pH;�tH;�zH;�H;��H;�H;$�H;��H;��H;��H;9�H;n�H;C�H;��H;��H;��H;��H;T�H;a�H;��H;�H;��H;��H;��H;��H;��H;��H;<�H;��H;��H;�H;C�H;_�H;C�H;�H;��H;��H;>�H;��H;��H;�H;��H;�H;��H;�H;��H;]�H;S�H;��H;��H;��H;��H;A�H;l�H;9�H;��H;��H;��H;%�H;�H;��H;�H;�zH; uH;3pH;JlH;fiH;�gH;      ��H;��H;U�H;��H;y�H;0�H;�H;C�H;X�H;��H;:�H;ͭH;9�H;��H;��H;��H;�H;�H;��H;g�H;l�H;"�H;u�H;��H;9�H;��H;�H;��H;��H;��H;:�H;��H;��H;5�H;^�H;~�H;z�H;}�H;^�H;5�H;��H;��H;;�H;��H;��H;��H;�H;��H;<�H;��H;t�H;"�H;j�H;g�H;��H;�H;�H;��H;��H;��H;9�H;˭H;:�H;��H;Z�H;A�H;�H;3�H;x�H;��H;U�H;�H;      b�H;ǚH;țH;m�H;��H;t�H;��H;i�H;C�H;Z�H;��H;�H;.�H;[�H;O�H;	�H;��H;��H;��H;��H;��H;��H;��H;w�H;��H;'�H;�H;��H;��H;8�H;��H;��H;8�H;p�H;��H;��H;��H;��H;��H;p�H;5�H;��H;��H;8�H;��H;��H;�H;$�H;��H;w�H;��H;��H;��H;��H;��H;��H;��H;	�H;M�H;Y�H;,�H;�H;��H;[�H;C�H;h�H;��H;w�H;��H;m�H;țH;��H;      ˩H;�H;ΪH;�H;ܭH;�H;��H;��H;��H;�H;I�H;��H;�H;W�H;y�H;|�H;V�H;�H;h�H;��H;{�H;�H;��H;��H;�H;�H;��H;��H;�H;��H;��H;4�H;i�H;��H;��H;��H;��H;��H;��H;��H;h�H;6�H;��H;��H;�H;��H;��H;�H;�H;��H;��H;�H;y�H;��H;h�H;�H;U�H;|�H;y�H;W�H;�H;��H;G�H;�H;��H;�H;��H;�H;ҭH;�H;ϪH;�H;      �H;^�H;��H;��H;��H;6�H;\�H;��H;H�H;��H;��H;��H;L�H;�H;��H;K�H;��H;��H;��H;��H;/�H;��H;��H;�H;��H;��H;g�H;�H;|�H;��H;�H;a�H;��H;��H;��H;��H;��H;��H;��H;��H;��H;b�H;�H;��H;~�H;�H;e�H;��H;��H;�H;��H;��H;-�H;��H;��H;��H;��H;I�H;��H;�H;L�H;��H;��H;��H;I�H;��H;\�H;;�H;{�H;��H;��H;V�H;      ��H;.�H;̺H;ŻH;�H;��H;b�H;r�H;��H; �H;v�H;��H;c�H;��H;!�H;X�H;e�H;I�H;�H;��H;�H;{�H;��H;��H;Q�H;�H;��H;:�H;��H;�H;B�H;�H;��H;��H;��H;��H;��H;��H;��H;��H;��H;��H;B�H;�H;��H;:�H;��H;�H;R�H;��H;��H;{�H;�H;��H;�H;J�H;d�H;X�H;!�H;��H;d�H;��H;t�H;�H;��H;q�H;b�H;��H;�H;ŻH;ϺH;%�H;      �H;�H;��H;��H;ľH;5�H;�H;�H;2�H;v�H;��H;�H;o�H;��H;��H;�H;��H;��H;��H;(�H;��H;��H;��H;��H;��H;=�H;��H;Q�H;��H;�H;a�H;�H;��H;��H;��H;��H;��H;��H;��H;��H;��H;��H;a�H;�H;��H;Q�H;��H;>�H;��H;��H;��H;��H;��H;(�H;��H;��H;��H;�H;��H;��H;o�H;�H;��H;y�H;3�H;�H;�H;:�H;��H;��H;��H;�H;      ��H;.�H;̺H;ŻH;�H;��H;b�H;r�H;��H; �H;v�H;��H;d�H;��H;!�H;X�H;e�H;I�H;�H;��H; �H;{�H;��H;��H;R�H;�H;��H;:�H;��H;�H;B�H;�H;��H;��H;��H;��H;��H;��H;��H;��H;��H;��H;B�H;�H;��H;:�H;��H;�H;Q�H;��H;��H;{�H;�H;��H;�H;J�H;d�H;X�H;!�H;��H;c�H;��H;v�H;�H;��H;p�H;b�H;��H;�H;ŻH;˺H;"�H;      �H;^�H;��H;��H;��H;6�H;\�H;��H;H�H;��H;��H;��H;L�H;�H;��H;I�H;��H;��H;��H;��H;1�H;��H;��H;�H;��H;��H;g�H;�H;}�H;��H;�H;_�H;��H;��H;��H;��H;��H;��H;��H;��H;��H;e�H;�H;��H;~�H;�H;e�H;��H;��H;�H;��H;��H;-�H;��H;��H;��H;��H;K�H;��H;�H;L�H;��H;��H;��H;H�H;��H;]�H;;�H;{�H;��H;��H;V�H;      ͩH;�H;ΪH;�H;ܭH;�H;��H;��H;��H;�H;H�H;��H;�H;W�H;y�H;|�H;V�H;�H;h�H;��H;}�H;�H;��H;��H;�H;�H;��H;��H;�H;��H;��H;4�H;i�H;��H;��H;��H;��H;��H;��H;��H;h�H;6�H;��H;��H;�H;��H;��H;�H;�H;��H;��H;�H;y�H;��H;h�H;�H;U�H;|�H;y�H;W�H;�H;��H;I�H;�H;��H;�H;��H;�H;ѭH;�H;ϪH;�H;      d�H;ǚH;ɛH;o�H;��H;t�H;��H;h�H;C�H;Z�H;��H;�H;,�H;[�H;N�H;	�H;��H;��H;��H;��H;��H;��H;��H;w�H;��H;&�H;�H;��H;��H;7�H;��H;��H;6�H;o�H;��H;��H;��H;��H;��H;o�H;5�H;��H;��H;8�H;��H;��H;�H;&�H;��H;u�H;��H;��H;��H;��H;��H;��H;��H;	�H;O�H;Y�H;,�H;�H;��H;[�H;C�H;e�H;��H;x�H;��H;o�H;ƛH;ĚH;      ��H;��H;U�H;��H;y�H;0�H;��H;B�H;X�H;��H;:�H;ͭH;9�H;��H;��H;��H;�H;�H;��H;i�H;o�H;"�H;u�H;��H;<�H;��H;�H;��H;��H;��H;;�H;��H;��H;5�H;^�H;~�H;z�H;}�H;^�H;5�H;��H;��H;:�H;��H;��H;��H;�H;��H;9�H;��H;t�H;"�H;j�H;g�H;��H;�H;�H;��H;��H;��H;7�H;˭H;:�H;��H;Z�H;?�H;��H;2�H;u�H;��H;V�H;�H;      gH;�gH;eiH;JlH;5pH;�tH;�zH;�H;��H;�H;%�H;��H;��H;��H;9�H;n�H;A�H;��H;��H;��H;��H;S�H;a�H;��H;�H;��H;�H;��H;��H;��H;��H;<�H;��H;��H;�H;C�H;_�H;C�H;�H;��H;��H;>�H;��H;��H;�H;��H;��H;��H;�H;��H;^�H;T�H;��H;��H;��H;��H;A�H;n�H;9�H;��H;��H;��H;"�H;�H;��H;�H;�zH; uH;3pH;IlH;fiH;�gH;      :@H;AH;eCH;/GH;dLH;�RH;,ZH;mbH;UkH;�tH;<~H;ڇH;T�H;��H;I�H;{�H;��H;�H;7�H;��H;�H;W�H;-�H;��H;[�H;��H;��H;x�H;��H;��H;��H;��H;.�H;��H;��H;	�H;�H;	�H;��H;��H;.�H;��H;��H;��H;��H;y�H;��H;��H;Z�H;��H;,�H;Y�H;�H;��H;8�H;�H;��H;}�H;K�H;��H;U�H;ڇH;<~H;�tH;VkH;mbH;,ZH;�RH;bLH;/GH;eCH;AH;      FH;FH;tH;|H;lH;�%H;�/H;�:H;�FH;�RH;q_H;lH;]xH;d�H;�H;��H;��H;��H;��H;��H;��H;1�H;�H;J�H;��H;��H;��H;��H;W�H;��H;��H;��H;��H;�H;z�H;��H;��H;��H;|�H;�H;��H;��H;��H;��H;Y�H;��H;��H;��H;��H;J�H;�H;2�H;��H;��H;��H;��H;��H;��H;�H;d�H;]xH;lH;q_H;�RH;�FH;�:H;�/H;�%H;hH;zH;qH;DH;      
�G;u�G;��G;�G;�G;,�G;�G;�H;H;a'H; 8H;�HH;�XH;QhH;4wH;*�H;+�H;�H;h�H;ױH;�H;_�H;��H;�H;��H;��H;��H;q�H;��H;y�H;��H;��H;��H;��H;
�H;:�H;M�H;:�H;�H;��H;��H;��H;��H;x�H;��H;q�H;��H;��H;��H;�H;��H;a�H;�H;ױH;h�H;�H;)�H;+�H;3wH;OhH;�XH;�HH;�7H;a'H;H;H;�G;'�G;�G;�G;��G;�G;      �nG;"qG;�wG;΂G;�G;I�G;n�G;��G;�G;C�G;�H;qH;�0H;�DH;FXH;DjH;�zH;�H;��H;�H;��H;·H;̿H;��H;]�H;T�H;t�H;��H;��H;��H;��H;�H;�H;��H;j�H;��H;��H;��H;k�H;��H;�H;�H;��H;��H;��H;��H;s�H;U�H;]�H;��H;˿H;·H;��H;�H;��H;�H;�zH;CjH;FXH;�DH;�0H;qH;�H;B�G;�G;��G;m�G;I�G;�G;΂G;�wG;qG;      �F;ͯF;�F;��F;�F;�!G;�FG;JjG;W�G;�G;�G;��G;5�G;�H;�1H;�HH;A^H;�qH;�H;��H;T�H;�H;�H;��H;�H;B�H;Q�H;��H;��H;��H;��H;��H;$�H;�H;��H;�H;B�H;�H;��H;�H;$�H;��H;��H;��H;��H;��H;S�H;C�H;�H;��H;�H;�H;O�H;��H;�H;�qH;A^H;�HH;�1H;�H;5�G;��G;�G;�G;W�G;HjG;�FG;�!G;�F;��F;�F;ƯF;      ��D;�D; �D;�9E;��E;B�E;dPF;�F;��F;/:G;VoG;͚G;�G;��G;�H;�H;�:H;�SH;�iH;v}H;��H;��H;��H;B�H;n�H;�H;a�H;��H;��H;c�H;�H;<�H;��H;�H;��H;U�H;��H;U�H;��H; �H;��H;@�H;�H;b�H;��H;��H;a�H;�H;m�H;@�H;��H;��H;��H;w}H;�iH;�SH;�:H;�H;�H;��G;�G;̚G;UoG;-:G;��F;�F;cPF;B�E;��E;�9E;��D;�D;      s@;UA@;1�@;RA;�"B;C;K�C;��D;0�E;�@F;��F;�!G;!hG;��G;T�G;�G;�H;"/H;4KH;�cH;{yH;J�H;g�H;��H;;�H;��H;��H;�H;D�H;��H;��H;~�H;p�H;��H;��H;��H;��H;��H; �H;��H;p�H;��H;��H;��H;C�H;�H;��H;��H;9�H;��H;e�H;M�H;zyH;�cH;4KH;%/H;�H;�G;T�G;��G; hG;�!G;��F;�@F;0�E;��D;K�C;C;�"B;RA;0�@;KA@;      �46;z�6;!l7;=�8;��:;c�<;F�>;b�@;�tB;q�C;�,E;�F;
�F;�,G;�xG;I�G;��G;�H;!&H;?EH;;`H;xwH;a�H;h�H;|�H;�H;ͿH;��H;�H;0�H;`�H;t�H;��H;��H;��H;��H;��H;��H;��H;��H;��H;t�H;`�H;/�H;�H;��H;˿H;�H;{�H;g�H;a�H;{wH;8`H;BEH;!&H;�H;��G;J�G;�xG;�,G;�F;�F;�,E;n�C;�tB;b�@;F�>;e�<;��:;=�8;l7;k�6;      q�";�M#;%;f�';6�+;N�/;��3;| 8;��;;/?;�A;ûC;:E;�@F;�F;�UG;�G;H�G;��G;z H;BH;�^H;xwH;M�H;��H;�H;·H;a�H;2�H;Z�H;T�H;�H;��H;�H;��H;y�H;��H;y�H;��H;�H;��H;�H;T�H;W�H;/�H;b�H;��H;�H;��H;M�H;vwH;�^H;BH;| H;��G;K�G;�G;�UG;�F;�@F;:E;ĻC;�A;-?;�;;x 8;��3;N�/;J�+;f�';%;�M#;      ���:3% ;\�;��;�;�P;5m;Kd';�.;�=5;�:;��>;�B;$BD;��E;i�F;7G;��G;��G;D�G;�H;BH;:`H;yH;��H;V�H;��H;�H;�H;�H;��H;e�H;��H;q�H;&�H;�H;�H;�H;&�H;r�H;��H;f�H;��H;�H;�H;�H;��H;V�H;��H;}yH;;`H;BH;�H;F�G;��G;��G;7G;i�F;��E;$BD;�B;��>;�:;}=5;�.;Jd';3m;�P;�;��;[�;*% ;      �Y�:Zo�:�W�:$�:/&�:{��:j��:@�	;Q;�M#;�n-;a�5;�;;�A@;�PC;9GE;�uF;�!G;��G;��G;D�G;w H;<EH;�cH;m}H;��H;�H;ұH;��H;��H;��H;_�H;��H;��H;�H;��H;!�H;��H;�H;��H;��H;`�H;��H;��H;�H;ԱH;�H;��H;o}H;�cH;9EH;w H;@�G;��G;��G;�!G;�uF;9GE;�PC;�A@;�;;_�5;�n-;�M#;Q;@�	;j��:���:;&�:"�:�W�:Fo�:      �	�H���xj�� ^��04u9*:�j~:��:�[�:�;|�;i%;�t0;��8;��>;�B;��D;�XF;YG;��G;��G;��G;"&H;7KH;�iH;�H;��H;k�H;��H;;�H;��H;��H;��H;e�H;��H;�H;��H;�H;��H;e�H;��H;��H;��H;8�H;��H;k�H;��H;�H;�iH;3KH;&H;��G;��G;��G;YG;�XF;��D;�B;��>;��8;�t0;j%;|�;�;�[�:��:�j~:F:�4u9 ^���j��H���      �A?���9�89)��Z��ܺ�p�����`:9��@:��:0�:_�	;Y;D,;݄6;��=;8#B;��D;�XF;�!G;��G;G�G;�H;#/H;�SH;�qH;�H;�H;��H;�H;��H;�H;��H;�H;��H;M�H;��H;N�H;��H;�H;��H;�H;��H;�H;��H;�H;�H;�qH;�SH;/H;�H;H�G;��G;�!G;�XF;��D;7#B;��=;݄6;D,;Y;_�	;0�:��:��@:0:9����p���ܺ�Z�:9)��9�      �Eֻ]�ѻ��Ļ}T�����.o��.�`ܺ��B����8�\:}&�:���:FQ;�);�=5;�:=;:#B;��D;vF;7G;�G;��G;�H;�:H;C^H;�zH;,�H;��H;��H;<�H;��H;��H;Q�H;��H;^�H;��H;^�H;��H;Q�H;��H;��H;<�H;��H;��H;,�H;�zH;F^H;�:H;�H;��G;�G;7G;vF;��D;<#B;�:=;�=5;�);EQ;���:{&�:�\:���8��B�cܺ�.��.o���}T����Ļb�ѻ      cFB�H�>���4�a�$�~��[�$����ݎ�zA?��Ӻ����l3�9�q�:WX�:^;��';�=5;��=;�B;=GE;j�F;�UG;J�G;�G;�H;�HH;CjH;*�H;��H;x�H;e�H;x�H;�H;q�H;A�H;Q�H;��H;Q�H;A�H;t�H;�H;z�H;e�H;x�H;��H;*�H;@jH;�HH;�H;�G;H�G;�UG;j�F;=GE;�B;��=;�=5;��';^;WX�:�q�:l3�9�����ӺxA?��ݎ�$���[�~��a�$���4�K�>�      ry��Hݜ��A���I����s���P�&+������Ļ����R|�H�o�:u9DX�:�+�:\;�);݄6;��>;�PC;��E;�F;�xG;V�G;�H;�1H;FXH;2wH;�H;H�H;5�H;��H;M�H;u�H;��H;�H;��H;�H;��H;v�H;K�H;��H;5�H;E�H;��H;3wH;EXH;�1H;�H;S�G;�xG;�F;��E;�PC;��>;��6;�);\;�+�:DX�::u9H�o�R|�������Ļ���&+���P���s��I���A��Jݜ�      z�����W�Ֆռ־�2Ϥ��I����[�(�[����9��{���:9HX�:[X�:GQ;F,;��8;�A@;$BD;�@F;�,G;��G;��G;�H;�DH;MhH;b�H;��H;��H;��H;U�H;P�H;�H;��H;��H;��H;�H;P�H;R�H;��H;��H;��H;d�H;OhH;�DH;�H;��G;��G;�,G;�@F;%BD;�A@;��8;H,;EQ;[X�:FX�:�:9�{����9��[�(���[��I��2Ϥ�־�Ֆռ�W���      9�6�M�3���+���g�t�����μ�������^FB�ps�PT��@�D��{��:u9�q�:���:Y;�t0;�;;�B;:E;�F;$hG;�G;5�G;�0H;�XH;[xH;N�H;��H;3�H;)�H;�H;D�H;]�H;k�H;_�H;E�H;�H;(�H;3�H;��H;P�H;ZxH;�XH;�0H;9�G;�G;hG;�F;:E;�B;�;;�t0;�Y;���:�q�::u9�{��B�D�PT��ps�^FB����������μt���g�����+�N�3�      t₽�؀���u��Xc���K�~1�������վ��]����P����PT����9�H�o�l3�9y&�:_�	;h%;a�5;��>;��C;�F;�!G;ǚG;��G;mH;�HH;�kH;̇H;~�H;��H;�H;��H;��H;��H;�H;��H;~�H;��H;ܹH;ĭH;~�H;̇H;�kH;�HH;kH;��G;ʚG;�!G;�F;��C;��>;a�5;h%;a�	;u&�:\3�9L�o���9�PT�������P��]���վ�����~1���K��Xc���u��؀�      >S���r��v�����֓����u���N���(��i�Ҍ˼�A����P�qs��R|������\:,�:x�;�n-;�:;
�A;�,E;��F;SoG;�G;�H;�7H;o_H;0~H;�H;3�H;��H;@�H;��H;j�H;��H;j�H;��H;A�H;��H;4�H;�H;0~H;m_H;�7H;�H; �G;VoG;��F;�,E;
�A;�:;�n-;x�;.�:�\:����T|��qs���P��A��Ҍ˼�i���(���N���u�֓�����v���r��       p��s��罰�ս:@��uĥ�|^���Xc�J�3���	�ӌ˼�]��_FB�[򻼜���Ӻ@��8��:��;�M#;{=5;)?;p�C;�@F;,:G;�G;A�G;]'H;�RH;�tH;��H;��H;X�H;޻H;��H;��H;s�H;��H;��H;޻H;W�H;��H;��H;�tH;�RH;^'H;?�G;�G;/:G;�@F;p�C;)?;}=5;�M#;��;��: ��8�Ӻ����[�_FB��]��ӌ˼��	�J�3��Xc�|^��uĥ�:@����ս���s�      �#�Y� �c'������gٽ<S��,l��V�j�J�3��i��վ�����(���Ļ|A?���B���@:�[�:Q;
�.;��;;�tB;-�E;��F;X�G;�G;
H;�FH;HkH;��H;S�H;=�H;��H;>�H;��H;'�H;��H;>�H;��H;;�H;S�H;��H;HkH;�FH;
H;�G;X�G;��F;*�E;�tB;��;;�.;Q;�[�:��@:��B�{A?���Ļ(������վ��i�I�3�V�j�,l��<S���gٽ����c'�Y� �      �S�+�O��E��5�X� �[�
���罪9��,l���Xc���(��������[�����ݎ�dܺ`:9��:@�	;Dd';o 8;_�@;��D;	�F;HjG;��G;uH;�:H;bbH;�H;8�H;_�H;v�H;��H;f�H;�H;g�H;��H;w�H;\�H;8�H;�H;bbH;�:H;uH;��G;HjG;�F;��D;_�@;o 8;Hd';?�	;��:p:9jܺ�ݎ������[��������(��Xc�,l���9�����[�
�X� ��5��E�+�O�      �~��*��-�v��9b��H�#,�PZ����<S��|^����N������μ�I��&+�(����.�����j~:d��:(m;��3;=�>;F�C;aPF;�FG;g�G;�G;�/H;"ZH;�zH;y�H;��H;��H;R�H;W�H;�H;W�H;R�H;��H;��H;y�H;�zH;!ZH;�/H;�G;f�G;�FG;dPF;A�C;=�>;��3;+m;b��:�j~:����.�(���&+��I����μ�����N�|^��<S�����PZ�#,��H��9b�-�v�*��      ����,����:���M��J�r�*�O�#,�[�
��gٽuĥ���u�~1�t���3Ϥ���P�[��.o��p��:y��:�P;C�/;Y�<;
C;;�E;�!G;G�G;'�G;�%H;�RH;�tH;*�H;q�H;�H;5�H;��H;3�H;��H;5�H;�H;p�H;,�H;�tH;�RH;�%H;'�G;E�G;�!G;<�E;C;\�<;D�/;�P;y��::�p���.o�[򻸎P�3Ϥ�t���~1���u�uĥ��gٽ[�
�#,�*�O�J�r��M���:��,���      :���v��P;������UP��J�r��H�X� ���:@��֓����K�g�־���s�~�����ܺ04u9#&�:�;2�+;��:;�"B;��E;	�F;�G;�G;eH;VLH;&pH;o�H;��H;ЭH;h�H;�H;��H;�H;g�H;ѭH;��H;r�H;&pH;SLH;bH;�G;�G;�F;��E;�"B;��:;2�+;�;#&�: 4u9�ܺ��~����s�־�g���K�֓��:@����X� ��H�J�r�UP������P;���v��      YVھ�*־25ʾu��������M���9b��5�����ս����Xc���֖ռ�I��b�$�|T���Z��^�� �:��;i�';C�8;RA;�9E;��F;̂G;�G;xH;&GH;>lH;|�H;c�H;�H;��H;��H;�H;��H;��H;�H;b�H;z�H;<lH;#GH;uH;�G;̂G;��F;�9E;RA;F�8;i�';��;�:`^���Z�}T��a�$��I��֖ռ���Xc������ս���5��9b��M������u���25ʾ�*־      ���쾶�޾25ʾP;���:��,�v��E�c'����v����u���+��W��A����4���Ļ>9)��j���W�:M�;%;l7;"�@;�D;�F;�wG;x�G;jH;ZCH;UiH;F�H;��H;ΪH;�H;��H;��H;��H;�H;ΪH;��H;F�H;UiH;WCH;hH;x�G;�wG;�F;�D;�@;l7;%;N�;�W�:�j��=9)���Ļ��4��A���W缊�+���u�v�����c'��E�,�v��:��P;��25ʾ��޾��      Zh���b���쾪*־�v��,���*��+�O�Y� �s��r���؀�N�3���Iݜ�J�>�d�ѻ �9�X���2o�:(% ;oM#;h�6;GA@;�D;ïF;qG;n�G;GH;�@H;�gH;�H;��H;�H;F�H;"�H;�H;"�H;H�H;�H;��H;�H;�gH;�@H;DH;n�G;qG;ïF;�D;DA@;n�6;oM#;(% ;0o�:X�����9�d�ѻJ�>�Iݜ���N�3��؀��r��s�Y� �+�O�*��,����v���*־���b��      4�$��� ����%��D��+�þ�*��6Dx���=�����Pν
���*'K��c�(��|�V����-E^���S��w[:���:e;T�4;>`?;�mD;��F;RvG;;�G;xH;}OH;�sH;�H;��H;��H;!�H;|�H;Q�H;|�H; �H;��H;��H;�H;�sH;|OH;uH;;�G;PvG;��F;�mD;<`?;W�4;e;���:�w[:��S�,E^����}�V�(���c�*'K�
����Pν�����=�6Dx��*��+�þD��%������� �      �� ����T��P��2��
����0��8�s�ڀ:�j9�!�ʽ5Z���G��8�.���5S����0X���D��Bd:�B�: ;�4;?;�~D;J�F;yG;��G;� H;FPH;CtH;=�H;��H;��H;_�H;��H;b�H;��H;`�H;��H;��H;>�H;CtH;CPH;� H;��G;yG;K�F;�~D;��?;!�4; ;�B�:�Bd:��D�0X���껺5S�.���8��G�6Z��"�ʽj9�ڀ:�8�s��0��
���3��P��T�����      ���T��;�
������Yؾ"���ᥒ���f���0�][�S8��Ӑ����>�����SȤ��6H�p�ܻ"rF����N�}:І�:c";U�5;��?;u�D;ծF;�G;��G;j#H;~RH;�uH;~�H;�H;��H;��H;�H;��H;�H;��H;��H;�H;~�H;�uH;{RH;g#H;��G;�G;ծF;u�D;��?;X�5;c";І�:F�}:���"rF�r�ܻ�6H�SȤ�������>�Ӑ��S8��][���0���f�ᥒ�"����Yؾ����;�
�T��      %��P������AI�+�þ�R��=���yS��Q"��s������}��0��켐�����6�U�ƻP}*�x�����:ox;Z%;�l7;س@;��D;��F;��G;��G;,(H;VH;�xH;��H;p�H;ϲH;�H;��H;��H;��H;�H;ϲH;o�H;��H;�xH;VH;)(H;��G;��G;��F;��D;Գ@;�l7;Z%;px;��:x���P}*�V�ƻ��6��������0���}�����s��Q"�yS�=����R��+�þAIᾧ���Q��      D��3�很Yؾ+�þĪ�~쏾�k�ڀ:�����ؽ�����c�cy���Ҽ���N� �v�B�� (7f�:��
;��(;�_9;��A;�\E;��F;ʝG;��G;�.H;�ZH;|H;�H;t�H;��H;?�H;�H;��H;�H;=�H;��H;q�H;!�H;|H;�ZH;�.H;��G;̝G;��F;�\E;��A;�_9;��(;��
;b�: (7@��v�N� ������Ҽcy��c�������ؽ��ڀ:��k�~쏾Ī�+�þ�Yؾ3��      *�þ
���"����R��~쏾:�s��H�����������Ӑ����D��c�����J�f�],�����P���9��:�;+j-;r�;;{�B;�E;�G;��G;��G;�6H;�`H;��H;��H;��H;�H;ӾH;}�H;�H;}�H;ӾH;�H;��H;��H;��H;�`H;�6H;��G;��G;�G;�E;w�B;r�;;*j-;�;��:�9�P�����],�J�f������c���D�Ӑ�������������H�9�s�~쏾�R��"���
���      �*���0��ᥒ�>����k��H��#%�][��Pνt��g�f�8/%���伍�����=��?ػ�FL���D�R�R:�:/�;?2;��=;ƚC;�0F;yGG;��G;JH;@H;�gH;��H;^�H;ڬH;ŸH;��H;�H;��H;�H;��H;øH;جH;`�H;��H;�gH;@H;IH;��G;zGG;�0F;C;��=;>2;1�;�:R�R:��D��FL��?ػ��=��������8/%�h�f�t���Pν][��#%��H��k�>���ᥒ��0��      6Dx�8�s���f�xS�ڀ:����][��7ս�榽��}���;��8�]�����r����HG�����ά� ��:�;�}$;҄6;#�?;�D;�F;�pG;��G;H;UJH;aoH;k�H;��H;*�H;h�H;��H;��H;W�H;��H;��H;h�H;)�H;��H;k�H;aoH;TJH;H;��G;�pG;�F;��D;#�?;҄6;�}$;�;"��:�ά���HG�������r�]����8���;���}��榽�7ս][����ڀ:�xS���f�8�s�      ��=�ڀ:���0��Q"��������Pν�榽C���G�7����Ҽ ��TE:�M�ܻ�D^�̸��<i:F��:�;>|,;��:;t�A;UiE;��F;J�G;��G;�(H;fUH;�wH;��H;W�H;��H;$�H;�H;��H;C�H;��H;�H;$�H;��H;X�H;��H;�wH;cUH;�(H;��G;L�G;��F;RiE;s�A;��:;?|,;�;H��:@i:̸���D^�M�ܻTE:� ����Ҽ7���G�C���榽�Pν�������Q"���0�ڀ:�      ���j9�][��s��ؽ���t����}��G������7c��b�V�O,��*�����@����:��:g ;m�3;�0>;�C;�F;9G;]�G;�H;8H;�`H;,�H;�H;+�H;u�H;�H;{�H;�H;C�H;�H;{�H;�H;t�H;,�H;�H;,�H;�`H;8H;�H;_�G;9G;�F;�C;�0>;m�3;f ;��:��:P������*��O,�b�V�7c��������G���}�t�������ؽ�s�][�j9�      �Pν!�ʽS8���������Ӑ��g�f���;�7�����JȤ�@�f�2��\ߵ�jo5� �D�2�-:C��:�>;�+;�_9;�A;��D;;�F;�vG;�G;BH;�GH;�lH;�H;ĞH;&�H;Y�H;&�H;��H;4�H;X�H;4�H;��H;&�H;W�H;)�H;ĞH;�H;�lH;�GH;?H;�G;�vG;7�F;��D;�A;�_9;�+;�>;I��:*�-: �D�jo5�[ߵ�2��?�f�JȤ����7����;�g�f�Ґ���������S8��"�ʽ      
���6Z��Ӑ����}��c���D�9/%��8���Ҽ6c��?�f����&�ƻ�/X�t���`��9�:>�;�";��3;N>;\YC;��E;�G;�G;��G;�,H;0WH;AxH;��H;b�H;�H;@�H;�H;e�H;t�H;d�H;t�H;e�H;�H;@�H;�H;b�H;��H;?xH;0WH;�,H;��G;�G;�G;��E;\YC;N>;��3;�";@�;
�:`��9t����/X�&�ƻ���?�f�7c����Ҽ�8�9/%���D��c���}�Ӑ��6Z��      *'K��G���>��0�cy��c����]��� ��b�V�2��&�ƻ�od���º v(7�4�:���:��;�P.;�:;'zA;J�D;�F;pnG;g�G;H;�@H;QfH;��H;[�H;�H;�H;�H; �H;��H;��H;m�H;��H;��H;�H;�H;�H;�H;[�H;��H;QfH;�@H;H;c�G;knG;�F;J�D;'zA;�:;�P.;��;���:�4�: v(7��º�od�&�ƻ2��b�V� ��]�����会c�cy��0���>��G�      �c��8���������Ҽ����������r�SE:�N,�Zߵ��/X���º Ȭ�^�}:	�:�;O�);8m7;.�?;��C;&F;�)G;5�G;t�G;2*H;�SH;�tH;��H;��H;"�H;޽H;��H;�H;C�H;��H;��H;��H;C�H;�H;��H;�H;"�H;��H;��H;�tH;�SH;3*H;s�G;4�G;{)G;&F;��C;.�?;8m7;R�);�;	�:b�}:�Ǭ���º�/X�Zߵ�N,�RE:���r�����������Ҽ�������8�      '��.��RȤ��������J�f���=����N�ܻ�*��ho5�t��� v(7Z�}:�n�:2�;�>&;��4;��=;��B;�E;5�F;��G;�G;]H;�AH;�eH;m�H;	�H;��H;�H;��H;R�H;��H;��H;��H;��H;��H;��H;��H;Q�H;��H;�H;��H;�H;k�H;�eH;�AH;ZH;�G;��G;4�F;�E;��B;��=;��4;�>&;2�;�n�:Z�}: v(7t���ho5��*��L�ܻ�����=�I�f��������RȤ�.��      {�V��5S��6H���6�M� �],��?ػHG���D^���� �D�`��9�4�:�:3�;�%;��3;,�<;nB;�E;!�F;�XG;+�G;r H;�0H;WH;�vH;!�H;��H;�H;ýH;��H;��H;��H;��H;��H;n�H;��H;��H;��H;��H;��H;ýH;�H;��H;�H;�vH;�WH;�0H;l H;)�G;�XG;�F;�E;nB;,�<;��3;�%;3�;	�:�4�:h��9 �D�����D^�HG���?ػ\,�N� ���6��6H��5S�      ��ﻺ��p�ܻU�ƻu�����FL���ȸ�� ��6�-:�:���:�;�>&;��3;h9<;'�A;��D;jZF;C5G;$�G;�G;�!H;`JH;`kH;ԅH;�H;��H;͸H;�H;��H;��H;�H;��H;��H;'�H;��H;��H;�H;��H;��H;�H;̸H;��H;�H;΅H;akH;`JH;�!H;�G;"�G;B5G;jZF;��D;)�A;h9<;��3;�>&;�;���:�:2�-: ��ĸ�����FL����t�U�ƻp�ܻ���      ,E^�0X�rF�K}*�B��Q����D��ά�Di:��:I��:>�;��;N�);��4;)�<;%�A;;�D;�9F;�G;��G;n�G;iH;H?H;�aH;C}H;��H;��H;˳H;�H;��H;��H;��H;O�H;��H;V�H;��H;V�H;��H;O�H;��H;��H;��H;�H;ȳH;��H;��H;D}H;�aH;D?H;gH;m�G;��G;�G;�9F;;�D;$�A;)�<;��4;Q�);��;?�;I��:��:Li:�ά���D��P��<��K}*�rF�!0X�      ��S���D�Ė�P��� (78�9n�R:"��:J��:$��:�>;�";�P.;9m7;��=;mB;��D;�9F;@G;F�G;��G;�H;�6H;�YH;vH;P�H; �H;0�H;3�H;��H;V�H;��H;M�H;j�H;��H;��H;(�H;��H;��H;j�H;J�H;��H;T�H;��H;0�H;/�H;�H;Q�H;vH;�YH;�6H;�H;|�G;F�G;@G;�9F;��D;mB;�=;8m7;�P.;�";�>;$��:P��: ��:r�R:x�9 (7P���Ė���D�      �w[:�Bd:^�}:��:h�:��:�:�;�;h ;�+;��3;�:;(�?;��B;�E;dZF;�G;A�G;��G;lH;�1H;TH;�pH;�H;|�H;�H;��H;��H;��H;3�H;��H;��H;U�H;*�H;H�H;��H;J�H;*�H;U�H;��H;��H;1�H;��H;��H;��H;�H;{�H;�H;�pH; TH;�1H;iH;��G;@�G;�G;dZF;�E;��B;(�?;�:;��3;�+;h ;�;�;�:��:~�:��:Z�}:�Bd:      ���:�B�:��:kx;��
;�;5�;�}$;>|,;r�3;�_9;M>;'zA;��C;�E;�F;B5G;��G;��G;mH;�/H; QH;2mH;}�H;ϗH;ŧH;��H;/�H;��H;K�H;��H;��H;��H;�H;��H;y�H;��H;x�H;��H;�H;��H;��H;��H;G�H;��H;-�H;��H;ŧH;͗H;w�H;1mH; QH;�/H;oH;��G;��G;@5G;�F;�E;��C;'zA;M>;�_9;o�3;@|,;�}$;7�;�;��
;nx;��:�B�:      e;% ;x";V%;��(;5j-;L2;݄6;ơ:;�0>;�A;_YC;L�D;&F;7�F;�XG;"�G;n�G;�H;�1H; QH;�kH;��H;��H;i�H;`�H;�H;��H;��H;C�H;��H;�H;��H;��H;��H;��H;��H;��H;��H;��H;��H;�H;��H;=�H;��H;��H;�H;b�H;i�H;��H;��H;�kH;QH;�1H;�H;n�G;�G;�XG;8�F;&F;L�D;_YC;�A;�0>;ǡ:;ۄ6;L2;8j-;�(;W%;u"; ;      ^�4;%�4;\�5;�l7;�_9;x�;;��=;'�?;u�A;�C;��D;��E;�F;�)G;��G;*�G;�G;hH;�6H;TH;1mH;��H;�H;<�H;�H;��H;Z�H;g�H;�H;��H;L�H; �H;i�H;��H;��H;��H;��H;��H;��H;��H;f�H;�H;L�H;��H;�H;e�H;W�H;��H;�H;8�H;ޔH;��H;-mH;TH;�6H;iH;
�G;)�G;��G;~)G;�F;��E;��D;�C;x�A;&�?;��=;x�;;�_9;�l7;^�5;�4;      X`?;׈?; �?;ܳ@;��A;y�B;КC;�D;ViE;�F;;�F;�G;mnG;7�G;�G;m H;�!H;G?H;�YH;�pH;y�H;��H;;�H;w�H;��H;]�H;z�H;<�H;��H;��H;��H;��H;��H;�H;��H;k�H;��H;j�H;��H;�H;��H;��H;��H;��H;��H;:�H;w�H;\�H;úH;u�H;8�H;��H;u�H;�pH;�YH;H?H;�!H;m H;�G;7�G;mnG;�G;;�F;�F;WiE;�D;͚C;{�B;ĘA;۳@;��?;ʈ?;      �mD;�~D;h�D;��D;�\E;�E;�0F;�F;��F;	9G;�vG;�G;g�G;x�G;_H;�0H;fJH;�aH;vH;�H;җH;m�H;��H;ʺH;�H;��H;��H;H�H;�H;-�H;��H;t�H;��H;�H;��H;�H;`�H;�H;��H;	�H;��H;u�H;��H;,�H;�H;E�H;��H;��H;!�H;ǺH;�H;l�H;ϗH;�H;vH;�aH;cJH;�0H;_H;w�G;f�G;�G;�vG;	9G;��F;�F;�0F;
�E;�\E;��D;g�D;�~D;      ��F;]�F;ϮF;��F;��F;�G;{GG;�pG;J�G;]�G;�G;��G;H;2*H;�AH;WH;`kH;B}H;M�H;|�H;§H;]�H;��H;\�H;��H;k�H;��H;��H;��H;G�H;E�H;��H;��H;��H;n�H;��H;�H;��H;n�H;��H;��H;��H;E�H;G�H;��H;��H;��H;j�H;��H;Z�H;��H;]�H;��H;{�H;M�H;B}H;]kH;|WH;�AH;2*H;H;��G;�G;\�G;L�G;�pG;{GG;�G;��F;��F;̮F;S�F;      hvG;yG;�G;��G;֝G;��G;��G;��G;��G;�H;CH;�,H;�@H;�SH;�eH;�vH;ԅH;��H;�H;�H;��H;�H;X�H;~�H;��H;��H;��H;��H;�H;�H;��H;��H;��H;{�H;�H;[�H;[�H;Z�H;�H;y�H;��H;��H;��H;�H;�H;��H;��H;��H;��H;z�H;W�H;	�H;��H;�H;�H;��H;҅H;�vH;�eH;�SH;�@H;�,H;EH;�H;��G;��G;��G;��G;۝G;��G;�G;yG;      4�G;��G;��G;��G;��G;��G;QH;H;�(H;8H;�GH;6WH;TfH;�tH;n�H;!�H;�H;��H;-�H;��H;-�H;��H;h�H;?�H;B�H;��H;��H;��H;��H;��H;��H;��H;��H;�H;��H;��H;��H;��H;��H;�H;��H;��H;��H;��H;��H;��H;��H;��H;C�H;>�H;e�H;��H;*�H;��H;-�H;��H;�H;!�H;n�H;�tH;RfH;7WH;�GH;8H;�(H;H;QH;��G;��G;��G;��G;��G;      �H;� H;n#H;3(H;�.H;�6H;@H;[JH;hUH;�`H;�lH;FxH;��H;��H;�H;��H;��H;ƳH;3�H;��H;��H;��H;�H;��H;�H;��H;�H;��H;k�H;��H;��H;��H;&�H;��H;��H;�H;(�H;�H;��H;��H;"�H;��H;��H;��H;h�H;��H;�H;��H;�H;��H;�H;��H;��H;��H;3�H;ɳH;��H;��H;�H;��H;��H;CxH;�lH;�`H;jUH;YJH;@H;�6H;�.H;3(H;m#H;� H;      �OH;QPH;�RH;VH;�ZH;�`H;�gH;koH;�wH;7�H;�H;đH;b�H;��H;��H;�H;θH;�H;��H;��H;K�H;@�H;��H;��H;%�H;D�H;�H;��H;��H;��H;��H;"�H;��H;�H;4�H;X�H;m�H;X�H;4�H;�H;��H;#�H;��H;��H;��H;��H;
�H;C�H;&�H;��H;��H;@�H;J�H;��H;��H;�H;͸H;�H;��H;��H;b�H;ÑH;�H;7�H;�wH;moH;�gH;�`H;�ZH;VH;�RH;OPH;      �sH;XtH;�uH;�xH;)|H;��H;��H;y�H;��H;#�H;ʞH;m�H;�H;)�H;�H;˽H;"�H;��H;V�H;8�H;��H;��H;L�H;��H;��H;H�H;��H;��H;��H;��H;�H;��H; �H;J�H;��H;��H;��H;��H;��H;J�H;��H;��H;�H;��H;��H;��H;��H;E�H;��H;��H;I�H;��H;��H;8�H;V�H;��H;!�H;ʽH;�H;(�H;�H;l�H;˞H;&�H;��H;x�H;��H;��H;%|H;�xH;�uH;XtH;       �H;O�H;��H;��H;(�H;��H;e�H;��H;^�H;/�H;/�H;%�H;	�H;�H;��H;�H;��H;��H;��H;�H;��H;�H;"�H;��H;o�H;��H;��H;��H;��H;%�H;��H;�H;F�H;��H;��H;��H;��H;��H;��H;��H;C�H;	�H;��H;&�H;��H;��H;��H;��H;r�H;��H; �H;�H;��H;�H;��H;��H;��H;�H;��H;�H;	�H;#�H;/�H;/�H;_�H;��H;e�H;��H;'�H;��H;��H;K�H;      ��H;�H;��H;z�H;�H;�H;ެH;5�H;ɳH;y�H;]�H;I�H;�H;��H;U�H;��H;��H;��H;O�H;��H;��H;��H;i�H;��H;��H;��H;��H;��H;*�H;��H;�H;J�H;��H;��H;��H;��H;�H;��H;��H;��H;��H;J�H;�H;��H;,�H;��H;��H;��H;��H;��H;g�H;��H;��H;��H;O�H;��H;��H;��H;U�H;��H;�H;H�H;^�H;{�H;ɳH;4�H;ެH;�H;x�H;{�H;��H;��H;      °H;�H;��H;ڲH;��H;�H;̸H;v�H;,�H; �H;.�H;&�H;"�H;�H;��H;��H;�H;N�H;m�H;]�H;�H;��H;��H;�H;�H;��H;v�H;�H;��H;�H;F�H;��H;��H;��H;��H;��H;�H;��H;��H;��H;��H;��H;F�H;�H;��H;�H;v�H;��H;�H;�H;��H;��H;�H;\�H;m�H;O�H;�H;��H;��H;�H;"�H;&�H;-�H; �H;,�H;u�H;̸H;��H;��H;ڲH;��H; �H;      "�H;x�H;�H;�H;[�H;վH;��H;��H;�H;��H;��H;r�H;��H;L�H;��H;��H;��H;��H;��H;2�H;��H;��H;��H;��H;��H;k�H;�H;��H;��H;6�H;��H;��H;��H;��H;�H;�H;�H;�H;�H;��H;��H;��H;��H;8�H;��H;��H;�H;k�H;��H;��H;��H;��H;��H;1�H;��H;��H;��H;��H;��H;J�H;��H;r�H;��H;��H;�H;��H;��H;پH;Q�H;�H;�H;p�H;      {�H;��H;)�H;��H;"�H;}�H;*�H;��H;��H;�H;?�H;�H;��H;��H;��H;��H;��H;R�H;��H;R�H;��H;��H;��H;q�H;�H;��H;X�H;��H;	�H;Z�H;��H;��H;��H;��H;�H;)�H; �H;)�H;�H;��H;��H;��H;��H;Z�H;�H;��H;W�H;��H;�H;n�H;��H;��H;��H;R�H;��H;S�H;��H;��H;��H;��H;��H;�H;=�H;
�H;��H;��H;*�H;��H;�H;��H;*�H;��H;      W�H;m�H;��H;��H;��H;�H;��H;a�H;N�H;H�H;b�H;n�H;r�H;��H;��H;w�H;/�H;��H;+�H;��H;��H;��H;��H;��H;Z�H;�H;X�H;��H;*�H;s�H;��H;��H;�H;	�H;�H;"�H;.�H;"�H;�H;	�H;��H;��H;��H;t�H;-�H;��H;W�H;�H;Z�H;��H;��H;��H;��H;��H;+�H;��H;.�H;w�H;��H;��H;r�H;n�H;b�H;J�H;O�H;^�H;��H;�H;��H;��H;��H;c�H;      {�H;��H;)�H;��H;"�H;}�H;*�H;��H;��H;�H;?�H;�H;��H;��H;��H;��H;��H;R�H;��H;R�H;��H;��H;��H;p�H;�H;��H;X�H;��H;	�H;Z�H;��H;��H;��H;��H;�H;)�H; �H;)�H;�H;��H;��H;��H;��H;Z�H;�H;��H;W�H;��H;�H;p�H;��H;��H;��H;R�H;��H;S�H;��H;��H;��H;��H;��H;�H;?�H;	�H;��H;��H;*�H;��H;�H;��H;'�H;��H;      !�H;x�H;�H;�H;[�H;վH;��H;��H;�H;��H;��H;r�H;��H;L�H;��H;��H;��H;��H;��H;2�H;��H;��H;��H;��H;��H;k�H;�H;��H;��H;6�H;��H;��H;��H;��H;�H;�H;�H;�H;�H;��H;��H;��H;��H;8�H;��H;��H;�H;k�H;��H;��H;��H;��H;��H;1�H;��H;��H;��H;��H;��H;L�H;��H;r�H;��H;��H;�H;��H;��H;پH;Q�H;�H;�H;n�H;      ðH;�H;��H;ڲH;��H;��H;̸H;u�H;+�H; �H;.�H;&�H;"�H;�H;��H;��H;�H;N�H;m�H;]�H;!�H;��H;��H;�H;�H;��H;v�H;�H;��H;�H;F�H;��H;��H;��H;��H;��H;�H;��H;��H;��H;��H;��H;F�H;�H;��H;�H;v�H;��H;�H;�H;��H;��H;�H;\�H;m�H;O�H;�H;��H;��H;�H;"�H;&�H;.�H; �H;,�H;t�H;̸H;��H;��H;ڲH;��H; �H;      ��H;�H;��H;{�H;}�H;�H;ެH;4�H;ɳH;y�H;^�H;H�H;�H;��H;U�H;��H;��H;��H;O�H;��H;��H;��H;i�H;��H;��H;��H;��H;��H;*�H;��H;�H;I�H;��H;��H;��H;��H;�H;��H;��H;��H;��H;M�H;�H;��H;,�H;��H;��H;��H;��H;��H;g�H;��H;��H;��H;O�H;��H;��H;��H;V�H;��H;�H;I�H;]�H;{�H;ȳH;3�H;ެH;�H;v�H;{�H;��H;�H;      �H;O�H;��H;��H;(�H;��H;h�H;��H;^�H;/�H;/�H;%�H;	�H;�H;��H;�H;��H;��H;��H;�H;��H;�H;"�H;��H;r�H;��H;��H;��H;��H;%�H;��H;�H;D�H;��H;��H;��H;��H;��H;��H;��H;C�H;	�H;��H;&�H;��H;��H;��H;��H;o�H;��H; �H;�H;��H;�H;��H;��H;��H;�H;��H;�H;	�H;#�H;/�H;/�H;_�H;��H;h�H;��H;&�H;��H;��H;I�H;      �sH;XtH;�uH;�xH;'|H;��H;��H;y�H;��H;%�H;ʞH;l�H;�H;+�H;�H;˽H;!�H;��H;V�H;8�H;��H;��H;L�H;��H;��H;G�H;��H;��H;��H;��H;�H;��H;��H;J�H;��H;��H;��H;��H;��H;J�H;��H;��H;�H;��H;��H;��H;��H;G�H;��H;��H;I�H;��H;��H;8�H;V�H;��H;!�H;˽H;�H;)�H;�H;m�H;ȞH;%�H;��H;x�H;��H;��H;%|H;�xH;�uH;XtH;      �OH;QPH;�RH;VH;�ZH;�`H;�gH;moH;�wH;7�H;�H;đH;b�H;��H;��H;�H;θH;�H;��H;��H;N�H;@�H;��H;��H;&�H;D�H;�H;��H;��H;��H;��H;"�H;��H; �H;4�H;X�H;m�H;X�H;4�H;�H;��H;#�H;��H;��H;��H;��H;�H;C�H;%�H;��H;��H;@�H;J�H;��H;��H;�H;͸H;�H;��H;��H;b�H;đH;�H;5�H;�wH;moH;�gH;�`H;�ZH;VH;�RH;PPH;      �H;� H;t#H;1(H;�.H;�6H;@H;]JH;iUH;�`H;�lH;FxH;��H;��H;	�H;��H;��H;ƳH;3�H;��H;��H;��H;�H;��H;�H;��H;�H;��H;i�H;��H;��H;��H;%�H;��H;��H;�H;(�H;�H;��H;��H;%�H;��H;��H;��H;k�H;��H;�H;��H;�H;��H;�H;��H;��H;��H;3�H;ȳH;��H;��H;�H;��H;��H;FxH;�lH;�`H;iUH;[JH;@H;�6H;�.H;-(H;q#H;� H;      4�G;��G;��G;��G;��G;��G;QH;H;�(H;8H;�GH;7WH;RfH;�tH;n�H;!�H;�H;��H;-�H;��H;0�H;��H;g�H;>�H;C�H;��H;��H;��H;��H;��H;��H;��H;��H;�H;��H;��H;��H;��H;��H;�H;��H;��H;��H;��H;��H;��H;��H;��H;B�H;?�H;g�H;��H;,�H;��H;-�H;��H;�H;"�H;n�H;�tH;TfH;6WH;�GH;8H;�(H;H;QH;��G;��G;��G;��G;��G;      bvG;yG;�G;��G;ѝG;��G;��G;��G;��G;�H;EH;�,H;�@H;�SH;�eH;�vH;ԅH;��H;�H;�H;��H;	�H;X�H;|�H;��H;��H;��H;��H;�H;�H;��H;��H;��H;y�H;�H;Z�H;[�H;Z�H;�H;y�H;��H;��H;��H;�H;�H;��H;��H;��H;��H;|�H;W�H;�H;��H;�H;�H;��H;҅H;�vH;�eH;�SH;�@H;�,H;EH;�H;��G;��G;��G;��G;ԝG;��G;�G;yG;      ��F;U�F;֮F;��F;��F;�G;{GG;�pG;J�G;]�G;�G;��G;H;2*H;�AH;}WH;^kH;@}H;M�H;{�H;ħH;]�H;��H;\�H;��H;j�H;��H;��H;��H;I�H;E�H;��H;��H;��H;k�H;��H;�H;��H;o�H;��H;��H;��H;E�H;F�H;��H;��H;��H;k�H;��H;Z�H;��H;]�H;��H;{�H;M�H;C}H;^kH;WH;�AH;2*H;H;��G;�G;\�G;J�G;�pG;}GG;�G;��F;��F;خF;N�F;      �mD;�~D;h�D;��D;�\E;�E;�0F;�F;��F;9G;�vG;�G;f�G;w�G;_H;�0H;dJH;�aH;vH;�H;җH;l�H;��H;ʺH;!�H;��H;��H;E�H;�H;-�H;��H;t�H;��H;	�H;��H;�H;`�H;�H;��H;�H;��H;v�H;��H;,�H;�H;H�H;��H;��H;�H;ȺH;�H;m�H;җH;�H;vH;�aH;cJH;�0H;_H;w�G;g�G;�G;�vG;9G;��F;�F;�0F;�E;�\E;��D;g�D;�~D;      ]`?;ӈ?;�?;س@;��A;��B;̚C;�D;WiE; F;=�F;�G;onG;7�G;�G;m H;�!H;E?H;�YH;�pH;y�H;��H;:�H;w�H;úH;]�H;x�H;:�H;��H;��H;��H;��H;��H;�H;��H;k�H;��H;k�H;��H;�H;��H;��H;��H;��H;��H;<�H;x�H;]�H;��H;v�H;:�H;��H;v�H;�pH;�YH;H?H;�!H;m H;�G;7�G;mnG;�G;:�F;�F;WiE;�D;̚C;�B;ƘA;ڳ@;�?;Ȉ?;      [�4;0�4;j�5;�l7;�_9;z�;;��=;'�?;w�A;�C;��D;��E;�F;�)G;��G;*�G;�G;gH;�6H;TH;4mH;��H;ߔH;;�H;�H;��H;Z�H;e�H;�H;��H;L�H; �H;i�H;��H;��H;��H;��H;��H;��H;��H;g�H; �H;L�H;��H;�H;g�H;W�H;��H;�H;:�H;ߔH;��H;.mH;TH;�6H;iH;
�G;*�G;��G;�)G;�F;��E;��D;�C;w�A;&�?;��=;|�;;�_9;�l7;a�5;�4;      e;% ;x";W%;��(;6j-;L2;݄6;ơ:;�0>;�A;_YC;L�D;&F;7�F;�XG;�G;n�G;�H;�1H;!QH;�kH;��H;��H;i�H;`�H;�H;��H;��H;A�H;��H;�H;��H;��H;��H;��H;��H;��H;��H;��H;��H;�H;��H;?�H;��H;��H;�H;b�H;i�H;��H;��H;�kH;QH;�1H;�H;p�G;!�G;�XG;8�F;&F;L�D;`YC;�A;�0>;ȡ:;ۄ6;L2;5j-;�(;V%;w"; ;      ���:�B�:��:nx;��
;�;9�;�}$;>|,;o�3;�_9;M>;'zA;��C;�E;�F;B5G;��G;��G;mH;�/H; QH;2mH;|�H;͗H;ŧH;��H;-�H;��H;J�H;��H;��H;��H;�H;��H;x�H;��H;y�H;��H;�H;��H;��H;��H;H�H;��H;/�H;��H;ŧH;ϗH;y�H;1mH; QH;�/H;oH;��G;��G;@5G;�F;�E;��C;'zA;K>;�_9;m�3;@|,;�}$;9�;�;��
;lx;��:�B�:      �w[:�Bd:r�}:��:p�:��:�:�;�;j ;�+;��3;�:;(�?;��B;�E;dZF;�G;@�G;��G;oH;�1H;TH;�pH;�H;{�H;�H;��H;��H;��H;1�H;��H;��H;U�H;*�H;J�H;��H;J�H;*�H;U�H;��H;��H;3�H;��H;��H;��H;�H;|�H;�H;�pH; TH;�1H;jH;��G;A�G;�G;dZF;�E;��B;(�?;�:;��3;�+;g ;�;�;�:��:x�:��:b�}:�Bd:      ��S���D�Ė�P��� (78�9r�R:"��:J��:$��:�>;�";�P.;8m7; �=;mB;��D;�9F;@G;D�G;�G;�H;�6H;�YH;vH;P�H; �H;/�H;3�H;��H;T�H;��H;M�H;j�H;��H;��H;(�H;��H;��H;j�H;K�H;��H;V�H;��H;0�H;0�H;�H;S�H;vH;�YH;�6H;�H;}�G;G�G;@G;�9F;��D;mB;�=;9m7;�P.;�";�>;$��:P��: ��:n�R:p�9 (7P���Ė���D�      (E^�0X�rF�L}*�D��Q����D� Ϭ�Di:��:I��:>�;��;O�);��4;)�<;%�A;:�D;�9F;�G;��G;m�G;iH;H?H;�aH;C}H;��H;��H;˳H;�H;��H;��H;��H;O�H;��H;V�H;��H;V�H;��H;O�H;��H;��H;��H;�H;ȳH;��H;��H;F}H;�aH;D?H;gH;n�G;��G;�G;�9F;;�D;$�A;)�<;��4;N�);��;>�;I��:��:Li:@Ϭ���D��P��>��L}*�rF�!0X�      ��ﻺ��p�ܻV�ƻu�����FL���ȸ�� ��:�-:�:���:�;�>&;��3;j9<;'�A;��D;iZF;C5G;"�G;�G;�!H;`JH;`kH;҅H;�H;��H;͸H;�H;��H;��H;�H;��H;��H;'�H;��H;��H;�H;��H;��H;�H;̸H;��H;�H;ЅH;akH;`JH;�!H;	�G;$�G;B5G;jZF;��D;)�A;h9<;��3;�>&;�;���:�:6�-: ��ĸ�����FL����t�V�ƻp�ܻ���      {�V��5S��6H���6�N� �^,��?ػHG���D^���� �D�h��9�4�:�:3�;�%;��3;*�<;nB;�E; �F;�XG;*�G;p H;�0H;WH;�vH;�H;��H;�H;ýH;��H;��H;��H;��H;��H;n�H;��H;��H;��H;��H;��H;ýH;�H;��H;!�H;�vH;�WH;�0H;m H;)�G;�XG; �F;�E;nB;-�<;��3;�%;4�;�:�4�:`��9 �D�����D^�IG���?ػ\,�N� ���6��6H��5S�      '��.��RȤ��������J�f���=����N�ܻ�*��jo5�t��� v(7Z�}:�n�:2�;�>&;��4;��=;��B;�E;4�F;��G;�G;ZH;�AH;�eH;k�H;�H;��H;�H;��H;T�H;��H;��H;��H;��H;��H;��H;��H;R�H;��H;�H;��H;�H;m�H;�eH;�AH;]H;�G;��G;5�F;�E;��B;��=;��4;�>&;2�;�n�:Z�}: v(7v���jo5��*��M�ܻ�����=�I�f��������RȤ�.��      �c��8���������Ҽ����������r�SE:�N,�Zߵ��/X���º Ȭ�b�}:	�:�;Q�);8m7;-�?;��C;&F;~)G;7�G;s�G;0*H;�SH;�tH;��H;��H;"�H;޽H;��H;�H;C�H;��H;��H;��H;C�H;�H;��H;߽H;"�H;��H;��H;�tH;�SH;5*H;t�G;4�G;})G;&F;��C;-�?;8m7;R�);�;�:^�}: Ȭ���º�/X�Zߵ�N,�RE:���r�����������Ҽ�������8�      *'K��G���>��0�cy��c����]��� ��b�V�2��&�ƻ�od���º v(7�4�:���:��;�P.;�:;%zA;J�D;�F;onG;c�G;H;�@H;QfH;��H;[�H;�H;�H;�H;�H;��H;��H;m�H;��H;��H; �H;�H;�H;�H;[�H;��H;QfH;�@H;H;g�G;lnG;�F;J�D;'zA;�:;�P.;��;���:�4�: v(7��º�od�&�ƻ2��b�V� ��]�����会c�cy��0���>��G�      ���6Z��Ӑ����}��c���D�9/%��8���Ҽ7c��?�f����&�ƻ�/X�t���`��9�:?�;�";��3;K>;\YC;��E;�G;�G;��G;�,H;0WH;AxH;��H;b�H;�H;A�H;�H;e�H;u�H;d�H;u�H;e�H;�H;>�H;�H;b�H;��H;?xH;0WH;�,H;��G;�G;�G;��E;\YC;O>;��3;�";?�;�:X��9t����/X�&�ƻ���?�f�6c����Ҽ�8�9/%���D��c���}�Ӑ��6Z��      �Pν!�ʽS8���������Ӑ��g�f���;�7�����JȤ�?�f�2��\ߵ�jo5� �D�2�-:E��:�>;�+;�_9;�A;��D;;�F;�vG;�G;BH;�GH;�lH;�H;ĞH;&�H;Z�H;&�H;��H;4�H;X�H;4�H;��H;&�H;W�H;(�H;ĞH;�H;�lH;�GH;?H;�G;�vG;7�F;��D;�A;�_9;�+;�>;G��:*�-:�D�jo5�\ߵ�2��?�f�JȤ����7����;�g�f�Ґ���������S8��"�ʽ      ���j9�][��s��ؽ���t����}��G������7c��b�V�O,��*�����@����:��:g ;l�3;�0>;�C;�F;9G;]�G;�H;8H;�`H;,�H;�H;+�H;v�H;�H;{�H;�H;C�H;�H;{�H;�H;t�H;+�H;�H;,�H;�`H;8H;�H;_�G;9G;�F;�C;�0>;o�3;f ;��:��:`������*��O,�b�V�7c��������G���}�t�������ؽ�s�][�j9�      ��=�ڀ:���0��Q"��������Pν�榽C���G�7����Ҽ ��TE:�L�ܻ�D^�ȸ��<i:H��:�;<|,;��:;t�A;UiE;��F;J�G;��G;�(H;fUH;�wH;��H;W�H;³H;$�H;�H;��H;C�H;��H;�H;$�H;��H;W�H;��H;�wH;cUH;�(H;��G;L�G;��F;RiE;s�A;��:;?|,;�;F��:@i:θ���D^�M�ܻTE:� ����Ҽ7���G�C���榽�Pν�������Q"���0�ڀ:�      6Dx�8�s���f�xS�ڀ:����][��7ս�榽��}���;��8�]�����r����HG�����ά�"��:�;�}$;҄6;#�?; �D;�F;�pG;��G;H;VJH;aoH;k�H;��H;*�H;j�H;��H;��H;W�H;��H;��H;j�H;)�H;��H;k�H;aoH;TJH;H;��G;�pG;�F;��D;#�?;҄6;�}$;�; ��:�ά���HG�������r�]����8���;���}��榽�7ս][����ڀ:�xS���f�8�s�      �*���0��ᥒ�>����k��H��#%�][��Pνt��h�f�8/%���伍�����=��?ػ�FL���D�R�R:�:.�;>2;��=;ƚC;�0F;yGG;��G;IH;@H;�gH;��H;^�H;ڬH;ŸH;��H;�H;��H;�H;��H;ŸH;جH;^�H;��H;�gH;@H;JH;��G;zGG;�0F;ÚC;��=;?2;1�;�:R�R:��D��FL��?ػ��=��������8/%�h�f�t���Pν][��#%��H��k�>���ᥒ��0��      *�þ
���"����R��~쏾9�s��H�����������Ӑ����D��c�����J�f�],�����P���9��:�;*j-;p�;;{�B;�E;�G;��G;��G;�6H;�`H;��H;��H;��H;�H;ӾH;}�H;�H;�H;ӾH;�H;��H;��H;��H;�`H;�6H;��G;��G;�G;�E;w�B;r�;;+j-;�;��:�9�P�����],�J�f������c���D�Ӑ�������������H�9�s�~쏾�R��"���
���      D��3�很Yؾ+�þĪ�~쏾�k�ڀ:�����ؽ�����c�cy���Ҽ���N� �v�B�� (7b�:��
;��(;�_9;��A;�\E;��F;ʝG;��G;�.H;�ZH;|H;�H;t�H;��H;?�H;�H;��H;�H;=�H;��H;q�H;!�H;|H;�ZH;�.H;��G;̝G;��F;�\E;��A;�_9;��(;��
;b�: (7@��w�N� ������Ҽcy��c�������ؽ��ڀ:��k�~쏾Ī�+�þ�Yؾ3��      %��P������AI�+�þ S��=���yS��Q"��s������}��0��켐�����6�U�ƻP}*�x�����:nx;Z%;�l7;س@;��D;��F;��G;��G;,(H;VH;�xH;��H;p�H;ϲH;�H;��H;��H;��H;�H;ϲH;o�H;��H;�xH;VH;)(H;��G;��G;��F;��D;Գ@;�l7;Z%;px;��:x���P}*�V�ƻ��6��������0���}�����s��Q"�yS�=����R��+�þAIᾧ���P��      ���T��;�
������Yؾ"���ᥒ���f���0�][�S8��Ӑ����>�����SȤ��6H�q�ܻ"rF����F�}:Ά�:c";U�5;��?;u�D;ծF;�G;��G;j#H;~RH;�uH;~�H;�H;��H;��H;�H;��H;�H;��H;��H;�H;~�H;�uH;{RH;g#H;��G;�G;ծF;u�D;��?;X�5;c";І�:F�}:���!rF�r�ܻ�6H�SȤ�������>�Ӑ��S8��][���0���f�ᥒ�"����Yؾ����;�
�T��      �� ����T��P��3��
����0��8�s�ڀ:�j9�!�ʽ5Z���G��8�.���5S����0X���D��Bd:�B�: ;�4;È?;�~D;J�F;yG;��G;� H;FPH;CtH;=�H;��H;��H;_�H;��H;b�H;��H;`�H;��H;��H;>�H;CtH;CPH;� H;��G;yG;K�F;�~D;��?;!�4; ;�B�:�Bd:��D�0X���껺5S�.���8��G�5Z��"�ʽj9�ڀ:�8�s��0��
���3��P��T�����      HEb�c]��N���7����u� ���˾��,�j��!,�v���P��Jm�0��?,˼ʪx�b���1��$�����:Q�:�;B�1;0,>;��C;�wF;��G;� H;�>H;�hH;V�H;y�H;B�H;%�H;��H;4�H;��H;4�H;��H;%�H;A�H;{�H;V�H;�hH;�>H;� H;��G;�wF;��C;.,>;D�1;�;Q�:��:$����1��b��ʪx�?,˼0��Jm�P��v����!,�,�j�����˾u� ������7��N�c]�      c]�g�W��TI�v3� E�������Ǿy����f�<)�)��v;���Fi��k���Ǽ�[t�T�	�6Ȅ�6X���:���:��;YJ2;NZ>;F	D;{F;C�G;H;�?H;�iH;�H;�H;z�H;A�H;��H;`�H;��H;`�H;��H;A�H;y�H;�H;�H;�iH;�?H;H;C�G;{F;F	D;JZ>;^J2;��;���:�:6X��6Ȅ�T�	��[t���Ǽ�k��Fi�v;��*��<)��f�y�����Ǿ���� E�v3��TI�g�W�      �N��TI���;�1�'�l��쾃���{󐾸Z��K ��s�D����&^���"����g�����u�!��3<:���: ;fg3;��>;vBD;��F;�G;�H;LBH;ykH;[�H;�H;1�H;޼H;v�H;��H;N�H;��H;u�H;޼H;/�H;�H;[�H;vkH;JBH;�H;�G;��F;xBD;��>;hg3;�
;���:3<:!���u������g��"����&^�D����s潨K ��Z�{󐾃�����l�1�'���;��TI�      ��7�v3�1�'����u� ��{Ծ!���J���|�F�����ӽ���e�L�Nv��뮼[T����PV���=��)i:\��:�z ;�$5;��?;�D;κF;��G;�H;�FH;�nH;��H;��H;t�H;�H;=�H;\�H;��H;\�H;=�H;�H;r�H;��H;��H;�nH;�FH;�H;��G;κF;	�D;��?;�$5;�z ;^��:�)i:��=��PV����[T��뮼Nv�e�L�����ӽ���|�F�J���!����{Ծu� ����1�'�v3�      ��� E�l�u� �Y�ݾm���X͓��f��>/�����'���섽T�6��t�w��g�:�0Tʻ�.�`۷�jt�:�;��$;�Y7;X�@;�	E;�F;9�G;�H;>LH;�rH;��H;ΤH;'�H;&�H;7�H;O�H;��H;O�H;6�H;&�H;%�H;ФH;��H;�rH;<LH;�H;;�G;�F;�	E;S�@;�Y7;��$;�;ft�:`۷��.�1Tʻg�:�w���t�T�6��섽�'������>/��f�X͓�m���Y�ݾu� �l� E�      u� ��������{Ծm���y���^�x��SC��^���޽C���~�e�,��K�Ѽ+G������R����� ݤ8:�Y;P�);��9;��A;��E;�G;�G;i!H;BSH;�wH;x�H;��H;D�H;��H;}�H;��H;��H;��H;}�H;��H;D�H;��H;x�H;�wH;>SH;h!H;�G;�G;��E;��A;��9;P�);�Y;釲: ݤ8����R�����+G��K�Ѽ,��~�e�C�����޽�^��SC�^�x�x���m����{Ծ�쾣���      ��˾��Ǿ����!���X͓�_�x���J��K �s���"������?����뮼5�[�+���"3|��W��x�:j�:�';n/;fg<;�C;mF;�NG;��G;/-H;o[H;�}H;ɗH;ʪH;��H;��H;�H;��H;�H;��H;�H;��H;��H;˪H;ɗH;�}H;m[H;/-H;��G;�NG;iF;�C;dg<;n/;�';d�:x�:�W��$3|�+���5�[��뮼���?����"��s����K ���J�_�x�X͓�"���������Ǿ      ��y���{�J����f��SC��K �sn���Ž����Z��k�'}ռ2X��iy-�7���x.����P�:�+�:��;4;9�>;�D;�wF;5�G;��G;�9H;ZdH;v�H;��H;d�H;r�H;��H;��H;X�H;u�H;X�H;��H;��H;q�H;f�H;��H;u�H;WdH;�9H;��G;5�G;�wF;�D;7�>;4;��;�+�:�P�:���y.�7���iy-�2X��'}ռ�k��Z�����Žsn���K ��SC��f�J���{�y���      ,�j��f��Z�|�F��>/��^�s����ŽJ ���Fi��Q+��t�uT��x�W�����1��6Ⱥ X�9�P�:�Y;��(;
�8;�A;�E;	�F;k�G;�H;�FH;�mH;��H;ġH;C�H;q�H;��H;��H;��H;��H;��H;��H;��H;q�H;D�H;ġH;��H;�mH;�FH;�H;m�G;�F;�E;�A;
�8;��(;�Y;�P�:X�96Ⱥ�1�����x�W�uT���t�Q+��Fi�J ���Žs����^��>/�|�F��Z��f�      �!,�<)��K ���������޽"������Fi��0����鷼��x�����.��_�(�����*i:���:>�;��0;O�<;�C;��E;=G;��G;�$H;hTH;�wH;�H;�H;Q�H;��H;C�H;��H;��H;�H;��H;��H;C�H;��H;R�H;�H;�H;�wH;gTH;�$H; �G;=G;��E;�C;M�<;��0;<�;���: +i:���_�(��.�������x�鷼����0��Fi����"����޽�������K �<)�      v���)��s��ӽ�'��C�������Z��Q+�����"��"G��ɻ0��׻ܕb�JW�� Y�9ҡ�:*`;�*';�Y7;$@;+�D;��F;�G;��G;;8H;bH;�H;\�H;��H;w�H;��H;��H;��H;U�H;A�H;U�H;��H;��H;��H;z�H;��H;[�H;��H;bH;:8H;��G;�G;��F;(�D;$@;�Y7;�*';,`;ء�:�X�9JW��ڕb��׻Ȼ0�"G���"������Q+��Z����C����'���ӽ�s�*��      Q��v;��D�������섽~�e��?��k��t�鷼"G���e7����Ȅ��0���t�,u�:,�:{;�1;X�<;f�B;+�E;�G;��G;dH;wJH;aoH;�H;��H;�H;��H;��H;"�H;��H;�H;��H;�H;��H;$�H;��H;��H;�H;��H;�H;aoH;tJH;eH;��G;�G;(�E;f�B;X�<;�1;{;,�:(u�:��t��0�Ȅ���껌e7�"G��鷼�t��k��?�~�e��섽���D���v;��      Jm��Fi��&^�e�L�T�6�,����'}ռuT����x�Ȼ0�������"���ط��n`:��:�;+�*;>�8;�@;=�D;l�F;�}G;��G;�1H;�[H;s|H;ÕH;�H;��H;��H;��H;��H;��H;��H;{�H;��H;��H;��H;��H;��H;��H;ߨH;��H;s|H;�[H;�1H;��G;�}G;h�F;=�D;�@;>�8;+�*;"�;��:�n`:�ط�"��������Ȼ0���x�uT��'}ռ��,��U�6�e�L��&^��Fi�      0���k��Nv��t�J�Ѽ�뮼2X��w�W������׻Ȅ�!��8��
5<:a��:�Y;�t%;�$5;�Z>;aC;��E;;*G;i�G;H;HH;rlH;��H;
�H;ɯH;׼H;��H;��H;�H;~�H;v�H;6�H;v�H;~�H;�H;��H;��H;׼H;ȯH;�H;��H;plH;HH;H;h�G;5*G;��E;aC;�Z>;�$5;�t%;�Y;a��:5<:0��"��Ȅ� �׻���w�W�2X���뮼I�Ѽ�t�Nv���k�      >,˼��Ǽ�"���뮼w��+G��5�[�jy-�����.��ܕb��0㺸ط�5<:�L�:�\;��!;�J2;�g<;V0B;1CE;0�F;U�G;��G;�4H;�\H;|H;��H;��H;`�H;��H;G�H;��H;W�H;X�H;�H;��H;�H;Z�H;Z�H;��H;H�H;��H;]�H;��H;��H;|H;�\H;�4H;��G;O�G;/�F;/CE;X0B;�g<;�J2;��!;�\;�L�:5<:�ط��0�ڕb��.�����jy-�5�[�+G��w���뮼�"����Ǽ      Ȫx��[t���g�ZT�g�:����(���7����1��]�(�LW����t��n`:a��:�\;{ ;��0;b;;=A;�D;�wF;�cG;[�G;�!H;�MH;�oH;{�H;��H;˯H;��H;m�H;��H;a�H;v�H;�H;��H;-�H;��H;�H;v�H;^�H;��H;m�H;��H;ƯH;��H;x�H;�oH;�MH;�!H;X�G;�cG;�wF;�D;=A;b;;��0;{ ;�\;e��:�n`:@�t�HW��_�(��1��7���'������g�:�YT���g��[t�      a��P�	������/Tʻ�R��3|�w.�4Ⱥ���Y�9*u�:��:�Y;��!;��0;�:;��@;CD;�2F;}8G;��G;�H;p@H;-dH;ʀH;}�H;M�H;P�H;U�H;��H;��H;��H;v�H;��H;�H;��H;�H;��H;w�H;��H;��H;��H;R�H;N�H;M�H;x�H;̀H;,dH;k@H;�H;��G;|8G;�2F;CD;��@;�:;��0;��!;�Y;��:*u�: Y�9���0Ⱥw.�3|��R��.Tʻ�����S�	�      �1��6Ȅ��u��PV��.�����W�����X�9+i:ء�:,�: �;�t%;�J2;_;;��@;sD;F;.G;��G;�H;�5H;�ZH;;xH;E�H;2�H;�H;�H;c�H;u�H;#�H;8�H;2�H;F�H;b�H;��H;b�H;F�H;2�H;5�H;#�H;u�H;a�H;�H;�H;-�H;H�H;;xH;�ZH;�5H;�H;}�G;/G;F;tD;��@;_;;�J2;�t%; �;	,�:ء�: +i: X�9���W������.��PV��u�:Ȅ�      ���0X��� ����=�`۷� ޤ8��:�P�:�P�:���:,`;~;+�*;�$5;�g<;=A;CD;F;�G;��G;n�G;�-H;!SH;_qH;�H;ǝH;��H;�H;B�H;��H;��H;��H;]�H;��H;��H;��H;��H;��H;��H;��H;\�H;��H;��H;��H;?�H;�H;��H;ǝH;�H;[qH;SH;�-H;i�G;��G;�G;F;CD;=A;�g<;�$5;-�*;~;,`;���:�P�:�P�:��:�ޤ80۷���=�� ��0X��      ��:`�:.3<:�)i:lt�:뇲:f�:�+�:�Y;@�;�*';�1;:�8;�Z>;S0B;�D;�2F;+G;��G;#�G;�)H;�NH;zlH;S�H;p�H;��H;��H;8�H;��H;�H;B�H;2�H;<�H;c�H;��H;��H;��H;��H;��H;c�H;:�H;2�H;@�H;�H;��H;6�H;��H;��H;o�H;N�H;wlH;�NH;�)H;"�G;��G;+G;�2F;�D;S0B;�Z>;<�8;�1;�*';>�;�Y;�+�:j�:�:�t�:�)i:.3<:D�:      m�:��:��:V��:�;�Y;�';��;��(;��0;�Y7;T�<;�@;aC;1CE;�wF;8G;��G;l�G;�)H;�LH;jH;<�H;d�H;��H;ٳH;ľH;m�H;.�H;��H;�H;^�H;��H;��H;��H;��H;��H;��H;��H;��H;��H;^�H;�H;��H;+�H;k�H;þH;׳H;��H;_�H;:�H;jH;�LH;�)H;l�G;��G;|8G;�wF;1CE;aC;�@;T�<;�Y7;��0;��(;��;�';�Y;�;Z��:��:���:      �;��;;�z ;��$;\�);{/;(4;�8;R�<;$@;i�B;?�D;��E;2�F;�cG;��G;�H;�-H;�NH;jH;P�H;��H;��H;�H;ɼH;��H;��H;U�H;��H;��H;;�H;U�H;��H;��H;u�H;��H;u�H;��H;��H;R�H;;�H;�H;��H;O�H;��H;��H;ʼH;�H;��H;��H;N�H;jH;�NH;�-H;�H;��G;�cG;3�F;��E;?�D;i�B;$@;R�<;�8;(4;{/;_�);��$;�z ;;��;      J�1;aJ2;kg3;�$5;�Y7;��9;jg<;=�>;�A;�C;-�D;.�E;l�F;;*G;S�G;Y�G;�H;�5H;SH;}lH;=�H;��H;4�H;�H;��H;u�H;k�H;=�H;��H;��H;��H;��H;��H;��H;��H;6�H;��H;6�H;��H;��H;��H;��H;��H;��H;��H;=�H;h�H;u�H;��H;ްH;1�H;��H;7�H;}lH;SH;�5H;�H;X�G;S�G;9*G;l�F;.�E;.�D;�C;A;=�>;jg<;��9;�Y7;�$5;mg3;VJ2;      J,>;dZ>; �>;��?;]�@;��A;�C;�D;�E;��E;��F;G;�}G;j�G;��G;�!H;m@H;�ZH;^qH;S�H;`�H;��H;�H;(�H;��H;��H;V�H;!�H; �H;�H;u�H;E�H;��H;��H;q�H;��H;�H;��H;q�H;��H;��H;E�H;t�H;�H;��H; �H;T�H;��H;��H;#�H;ްH;��H;\�H;Q�H;\qH;�ZH;k@H;�!H;��G;j�G;�}G;G;��F;��E;�E; D;�C;��A;f�@;��?;��>;VZ>;      ��C;T	D;kBD;�D;�	E;ĄE;oF;�wF;	�F;=G;�G;��G;��G;H;�4H;�MH;3dH;>xH;�H;w�H;��H;�H;��H;��H;U�H;�H;��H;��H;��H;��H;��H;��H;��H;h�H;�H;l�H;s�H;k�H;�H;g�H;��H;��H;��H;��H;��H;��H;��H;�H;U�H;��H;��H;�H;��H;v�H;�H;?xH;.dH;�MH;�4H;H;��G;��G;�G;=G;
�F;�wF;oF;ĄE;
E;�D;jBD;S	D;      �wF;�F;��F;ҺF;!�F;�G;�NG;7�G;m�G;��G;��G;fH;�1H;HH;�\H;�oH;̀H;E�H;ÝH;��H;ֳH;ǼH;r�H;��H;�H;}�H;H�H;E�H;��H;��H;B�H;|�H;`�H;#�H;��H;��H;��H;��H;��H;"�H;\�H;|�H;@�H;��H;��H;D�H;F�H;|�H;�H;��H;r�H;ǼH;ҳH;��H;ÝH;E�H;ǀH;�oH;�\H;HH;�1H;hH;��G;��G;o�G;7�G;�NG;�G;(�F;ҺF;��F;�F;      �G;K�G;�G;��G;E�G;(�G;��G;��G;�H;�$H;>8H;{JH;�[H;slH;|H;|�H;}�H;/�H;��H;��H;žH;��H;j�H;Z�H;��H;L�H;,�H;��H;t�H; �H;c�H;;�H;�H;��H;��H;2�H;@�H;2�H;��H;��H;�H;:�H;`�H;�H;r�H;��H;,�H;H�H;��H;W�H;h�H;��H;þH;��H;��H;0�H;|�H;{�H;|H;slH;�[H;{JH;?8H;�$H;�H;��G;��G;&�G;J�G; �G;�G;J�G;      � H;#H;�H;�H;�H;n!H;7-H;�9H;�FH;nTH;	bH;hoH;v|H;��H;��H;��H;L�H;�H;�H;;�H;k�H;��H;@�H;$�H;}�H;E�H;��H;��H;�H;2�H;3�H;�H;��H;�H;F�H;��H;��H;��H;F�H;�H;��H;�H;2�H;.�H;�H;��H;��H;E�H;}�H;#�H;=�H;��H;h�H;9�H;�H;�H;J�H;��H;��H;��H;u|H;hoH;bH;nTH;�FH;�9H;7-H;n!H;�H;�H;�H;/H;      ?H;�?H;RBH;�FH;CLH;GSH;x[H;adH;�mH;�wH;�H;�H;ƕH;
�H;��H;̯H;R�H;�H;A�H;��H;0�H;R�H;��H;�H;��H;��H;o�H;�H;O�H;�H;��H;��H;�H;e�H;��H;��H;��H;��H;��H;e�H;��H;��H;��H;�H;N�H;�H;r�H;��H;��H;�H;��H;Q�H;,�H;��H;A�H;�H;P�H;̯H;��H;
�H;ƕH;�H;�H;�wH;�mH;adH;x[H;ESH;JLH;�FH;RBH;�?H;      iH;�iH;�kH;�nH;�rH;�wH;�}H;~�H;��H;��H;g�H;áH;�H;ӯH;c�H;��H;X�H;^�H;��H;�H;��H;��H;��H;�H;��H;��H;�H;2�H;�H;��H;��H;	�H;Q�H;��H;��H;��H;��H;��H;��H;��H;N�H;�H;��H;��H;�H;/�H;�H;��H;��H;�H;��H;��H;��H;�H;��H;^�H;U�H;��H;c�H;ЯH;�H;��H;i�H;��H;��H;��H;�}H;�wH;�rH;�nH;�kH;�iH;      `�H;�H;m�H;��H;ȏH;{�H;ԗH;��H;ΡH;"�H;��H;'�H;��H;߼H;��H;u�H;��H;u�H;��H;G�H;#�H;��H;��H;x�H;��H;C�H;_�H;4�H;��H;��H;	�H;_�H;��H;��H;��H;�H;�H;�H;��H;��H;��H;a�H;	�H;��H;��H;4�H;`�H;@�H;��H;x�H;��H;��H; �H;G�H;��H;t�H;��H;t�H;��H;޼H;��H;%�H;��H;%�H;ΡH;��H;ԗH;}�H;ŏH;��H;k�H;�H;      ��H;��H;��H;��H;ۤH;��H;ҪH;r�H;K�H;U�H;��H;��H;��H;��H;N�H;��H;�H;#�H;��H;;�H;e�H;=�H;��H;I�H;��H;|�H;:�H;�H;��H;�H;^�H;��H;��H;�H;�H;5�H;Q�H;5�H;�H;�H;��H;��H;^�H;�H;��H;�H;:�H;z�H;��H;I�H;��H;=�H;d�H;;�H;��H;&�H; �H;��H;N�H;��H;��H;��H;��H;V�H;N�H;p�H;ӪH;��H;ڤH;��H;��H;��H;      L�H;��H;?�H;��H;5�H;H�H;ƸH;��H;z�H;��H;��H;��H;��H;��H;��H;g�H;��H;4�H;_�H;A�H;��H;U�H;��H;��H;��H;`�H;�H;��H;�H;W�H;��H;��H;�H;+�H;N�H;D�H;7�H;C�H;M�H;)�H;��H;��H;��H;X�H;�H;��H;�H;^�H;��H;��H;��H;U�H;��H;B�H;_�H;5�H;��H;g�H;��H;��H;��H;��H;��H;��H;{�H;�H;ƸH;M�H;.�H;��H;?�H;��H;      5�H;Q�H;߼H;�H;2�H;��H;��H;��H;��H;I�H;��H;,�H;��H;�H;^�H;��H;}�H;2�H;��H;k�H;��H;��H;��H;��H;c�H; �H;��H;�H;c�H;��H;��H;�H;$�H;7�H;c�H;n�H;N�H;n�H;c�H;6�H;!�H;�H;��H;��H;f�H;�H;��H; �H;d�H;��H;��H;��H;��H;k�H;��H;3�H;{�H;�H;\�H;�H;��H;,�H;��H;I�H;��H;��H;��H;��H;(�H;�H;�H;J�H;      ��H;
�H;��H;I�H;U�H;}�H;�H;��H;��H;��H;��H;��H;��H;��H;`�H;�H;��H;C�H;��H;��H;��H;��H;��H;v�H;�H;��H;��H;F�H;��H;��H;��H;�H;K�H;d�H;G�H;d�H;��H;d�H;G�H;d�H;H�H;�H;��H;��H;��H;F�H;��H;��H;�H;u�H;��H;��H;��H;��H;��H;D�H;��H;�H;`�H;��H;��H;��H;��H;��H;��H;��H;�H;��H;K�H;G�H;��H;�H;      4�H;n�H;��H;f�H;d�H;��H;��H;f�H;
�H;��H;^�H; �H;��H;��H;�H;��H;�H;]�H;��H;��H;��H;w�H;7�H;��H;g�H;��H;/�H;��H;��H;��H;�H;7�H;C�H;r�H;d�H;[�H;k�H;[�H;d�H;p�H;?�H;:�H;�H;��H;��H;��H;/�H;��H;h�H;��H;7�H;w�H;��H;��H;��H;_�H;�H;��H;�H;~�H;��H; �H;]�H;��H;
�H;c�H;��H;��H;Y�H;f�H;��H;e�H;      ��H;��H;c�H;��H;��H;��H;�H;��H;�H;��H;J�H;��H;��H;@�H;��H;7�H;��H;��H;��H;��H;��H;��H;��H;�H;n�H;��H;=�H;��H;��H;��H;�H;V�H;7�H;R�H;~�H;m�H;Y�H;m�H;~�H;R�H;5�H;X�H;�H;��H;��H;��H;=�H;��H;n�H;�H;��H;��H;��H;��H;��H;��H;��H;7�H;��H;@�H;��H;��H;J�H;��H;�H;}�H;�H;��H;��H;��H;c�H;��H;      4�H;n�H;��H;f�H;d�H;��H;��H;f�H;
�H;��H;^�H; �H;��H;��H;�H;��H;�H;]�H;��H;��H;��H;w�H;7�H;��H;h�H;��H;/�H;��H;��H;��H;�H;7�H;A�H;r�H;d�H;[�H;k�H;[�H;d�H;p�H;@�H;:�H;�H;��H;��H;��H;/�H;��H;g�H;��H;7�H;w�H;��H;��H;��H;_�H;�H;��H;�H;~�H;��H; �H;^�H;��H;
�H;c�H;��H;��H;Y�H;f�H;��H;d�H;      ��H;
�H;��H;I�H;U�H;}�H;�H;��H;��H;��H;��H;��H;��H;��H;`�H;�H;��H;C�H;��H;��H;��H;��H;��H;v�H;�H;��H;��H;F�H;��H;��H;��H;�H;K�H;d�H;G�H;d�H;��H;d�H;G�H;d�H;H�H;�H;��H;��H;��H;F�H;��H;��H;�H;t�H;��H;��H;��H;��H;��H;D�H;��H;�H;`�H;��H;��H;��H;��H;��H;��H;��H;�H;��H;K�H;I�H;��H;�H;      7�H;Q�H;߼H;�H;2�H;��H;��H;��H;��H;I�H;��H;,�H;��H;�H;\�H;�H;}�H;2�H;��H;k�H;��H;��H;��H;��H;d�H;"�H;��H;�H;c�H;��H;��H;��H;"�H;6�H;c�H;n�H;N�H;n�H;c�H;7�H;"�H;�H;��H;��H;f�H;�H;��H;"�H;c�H;��H;��H;��H;��H;k�H;��H;3�H;{�H;��H;^�H;�H;��H;,�H;��H;I�H;��H;��H;��H;��H;(�H;�H;�H;J�H;      O�H;��H;@�H;��H;3�H;J�H;ƸH;�H;{�H;��H;��H;��H;��H;��H;��H;g�H;��H;3�H;_�H;A�H;��H;U�H;��H;��H;��H;`�H;�H;��H;�H;W�H;��H;��H;��H;(�H;M�H;C�H;7�H;D�H;N�H;)�H;��H;��H;��H;X�H;�H;��H;�H;^�H;��H;��H;��H;U�H;��H;B�H;_�H;4�H;��H;g�H;��H;��H;��H;��H;��H;��H;z�H;|�H;ŸH;M�H;,�H;��H;?�H;��H;      ��H;��H;��H;��H;ڤH;��H;ժH;q�H;K�H;V�H;��H;��H;��H;��H;N�H;��H;�H;#�H;��H;<�H;h�H;=�H;��H;I�H;��H;{�H;:�H;�H;��H;�H;^�H;��H;��H;�H;�H;5�H;Q�H;5�H;�H;�H;��H;��H;^�H;�H;��H;�H;:�H;{�H;��H;I�H;��H;=�H;d�H;;�H;��H;%�H; �H;��H;N�H;��H;��H;��H;��H;V�H;M�H;p�H;ժH;��H;פH;��H;��H;��H;      `�H;�H;k�H;��H;ȏH;|�H;ԗH;��H;ΡH;#�H;��H;%�H;��H;߼H;��H;u�H;��H;r�H;��H;I�H;%�H;��H;��H;z�H;��H;B�H;`�H;4�H;��H;��H;	�H;_�H;��H;��H;��H;�H;�H;�H;�H;��H;��H;a�H;	�H;��H;��H;4�H;`�H;B�H;��H;x�H;��H;��H; �H;G�H;��H;u�H;��H;u�H;��H;߼H;��H;'�H;��H;#�H;ΡH;��H;ԗH;}�H;ŏH;��H;m�H;�H;      �hH;�iH;�kH;�nH;�rH;�wH;�}H;��H;��H;��H;g�H;��H;�H;ӯH;c�H;��H;V�H;]�H;��H;�H;��H;��H;��H;�H;��H;��H;�H;/�H;�H;��H;��H;	�H;P�H;��H;��H;��H;��H;��H;��H;��H;P�H;�H;��H;��H;�H;2�H;�H;��H;��H;�H;��H;��H;��H;�H;��H;`�H;V�H;��H;c�H;үH;�H;��H;g�H;��H;��H;��H;�}H;�wH;�rH;�nH;�kH;�iH;      ?H;�?H;XBH;�FH;HLH;BSH;{[H;ddH;�mH;�wH;�H;�H;ƕH;
�H;��H;̯H;R�H;�H;A�H;��H;2�H;Q�H;��H;�H;��H;��H;o�H;�H;N�H;�H;��H;��H; �H;e�H;��H;��H;��H;��H;��H;e�H; �H;��H;��H;�H;O�H;�H;r�H;��H;��H;�H;��H;R�H;.�H;��H;A�H;�H;P�H;ͯH;��H;
�H;ƕH;�H;�H;�wH;�mH;bdH;{[H;ESH;ELH;�FH;UBH;�?H;      � H;#H;�H;�H;�H;n!H;7-H;�9H;�FH;nTH;	bH;hoH;u|H;��H;��H;��H;L�H;�H;�H;;�H;n�H;��H;?�H;#�H;}�H;E�H;��H;��H;�H;0�H;2�H;�H;��H;�H;D�H;��H;��H;��H;F�H;�H;��H;�H;3�H;/�H;�H;��H;��H;E�H;}�H;$�H;?�H;��H;h�H;9�H;�H;�H;J�H;��H;��H;��H;v|H;hoH;bH;nTH;�FH;�9H;7-H;k!H;�H;�H;�H;.H;      �G;J�G;�G;��G;@�G;$�G;��G;��G;�H;�$H;?8H;{JH;�[H;slH;|H;|�H;�H;/�H;��H;��H;ȾH;��H;j�H;X�H;��H;J�H;-�H;��H;t�H; �H;`�H;:�H;�H;��H;��H;2�H;@�H;1�H;��H;��H;�H;=�H;c�H;�H;r�H;��H;,�H;J�H;��H;X�H;h�H;��H;þH;��H;��H;0�H;|�H;{�H;|H;slH;�[H;{JH;?8H;�$H;�H;��G;��G;#�G;C�G;��G;�G;?�G;      �wF;�F;��F;ҺF;"�F;�G;�NG;8�G;m�G; �G;��G;fH;�1H;HH;�\H;�oH;ʀH;C�H;ÝH;��H;׳H;ǼH;p�H;��H;�H;|�H;F�H;D�H;��H;��H;@�H;{�H;]�H;"�H;��H;��H;��H;��H;��H;#�H;]�H;~�H;B�H;��H;��H;E�H;H�H;}�H;�H;��H;r�H;ǼH;ӳH;��H;ÝH;F�H;ɀH;�oH;�\H;HH;�1H;fH;��G;��G;m�G;4�G;�NG;�G;&�F;պF;��F;~F;      ��C;T	D;jBD;�D;�	E;ĄE;oF;�wF;
�F;=G;�G;��G;��G;H;�4H;�MH;0dH;<xH;�H;w�H;��H;�H;��H;��H;U�H;�H;��H;��H;��H;��H;��H;��H;��H;g�H;�H;k�H;s�H;l�H;�H;g�H;��H;��H;��H;��H;��H;��H;��H;�H;U�H;��H;��H;�H;��H;w�H;�H;AxH;0dH;�MH;�4H;H;��G;��G;�G;=G;	�F;�wF;oF;ĄE;�	E;�D;jBD;T	D;      O,>;`Z>;�>;��?;X�@;�A;�C; D;�E;��E;��F;G;�}G;j�G;��G;�!H;m@H;�ZH;\qH;Q�H;`�H;��H;߰H;(�H;��H;��H;V�H; �H;��H;
�H;t�H;C�H;��H;��H;n�H;��H;�H;��H;r�H;��H;��H;F�H;u�H;�H;��H;!�H;V�H;��H;��H;&�H;߰H;��H;]�H;S�H;^qH;�ZH;k@H;�!H;��G;j�G;�}G;G;��F;��E;�E;�D;�C;�A;g�@;��?;�>;RZ>;      G�1;nJ2;yg3;�$5;�Y7;��9;ng<;=�>;�A;�C;-�D;.�E;j�F;9*G;S�G;Y�G;�H;�5H;SH;|lH;=�H;��H;3�H;�H;��H;u�H;k�H;=�H;��H;��H;��H;��H;��H;��H;��H;6�H;��H;6�H;��H;��H;��H;��H;��H;��H;��H;=�H;h�H;u�H;��H;߰H;3�H;��H;9�H;}lH;SH;�5H;�H;Y�G;U�G;;*G;j�F;.�E;-�D;�C;A;;�>;pg<;��9;�Y7;�$5;og3;[J2;      �;��;;�z ;��$;^�);{/;(4;�8;R�<;$@;i�B;?�D;��E;2�F;�cG;��G;�H;�-H;�NH;jH;N�H;��H;��H;�H;ɼH;��H;��H;T�H;��H;�H;;�H;S�H;��H;��H;u�H;��H;u�H;��H;��H;S�H;;�H;��H;��H;Q�H;��H;��H;ʼH;�H;��H;��H;P�H;jH;�NH;�-H;�H;��G;�cG;3�F;��E;?�D;j�B;$@;R�<;�8;'4;{/;\�);��$;�z ;;��;      _�:��:��:Z��:�;�Y;�';��;��(;��0;�Y7;T�<;�@;aC;1CE;�wF;}8G;��G;l�G;�)H;�LH;jH;<�H;c�H;��H;׳H;ľH;k�H;.�H;��H;�H;]�H;��H;��H;��H;��H;��H;��H;��H;��H;��H;`�H;�H;��H;+�H;m�H;þH;ٳH;��H;`�H;:�H;jH;�LH;�)H;l�G;��G;}8G;�wF;1CE;aC;�@;T�<;�Y7;��0;��(;��;�';�Y;�;Z��:��:���:      ��:h�:B3<:�)i:rt�::j�:�+�:�Y;?�;�*';�1;:�8;�Z>;S0B;�D;�2F;)G;��G;"�G;�)H;�NH;ylH;S�H;o�H;��H;��H;6�H;��H;�H;@�H;1�H;<�H;c�H;��H;��H;��H;��H;��H;c�H;;�H;4�H;B�H;�H;��H;8�H;��H;��H;p�H;N�H;wlH;�NH;�)H;#�G;��G;,G;�2F;�D;S0B;�Z>;:�8;�1;�*';?�;�Y;�+�:j�:�:|t�:�)i::3<:@�:      ���2X��� ����=�h۷� ޤ8��:�P�:�P�:���:,`;~;-�*;�$5;�g<;=A;CD;F;�G;��G;l�G;�-H;!SH;_qH;�H;ƝH;��H;�H;B�H;��H;��H;��H;]�H;��H;��H;��H;��H;��H;��H;��H;\�H;��H;��H;��H;?�H;�H;��H;ɝH;�H;[qH;SH;�-H;k�G;��G;�G;F;CD;=A;�g<;�$5;+�*;~;,`;���:�P�:�P�:��:�ޤ88۷���=�� ��0X��      �1��6Ȅ��u��PV��.�����W�����X�9 +i:ء�:	,�: �;�t%;�J2;_;;��@;sD;F;.G;��G;�H;�5H;�ZH;;xH;E�H;0�H;�H;�H;c�H;u�H;"�H;7�H;2�H;F�H;b�H;��H;b�H;F�H;2�H;7�H;%�H;u�H;a�H;�H;�H;/�H;H�H;;xH;�ZH;�5H;�H;��G;/G;F;tD;��@;_;;�J2;�t%; �;,�:ء�:+i: X�9���W������.��PV��u�:Ȅ�      a��Q�	������0Tʻ�R��3|�v.�4Ⱥ���Y�9*u�:��:�Y;��!;��0;�:;��@;CD;�2F;8G;��G;�H;p@H;,dH;ʀH;|�H;M�H;P�H;U�H;��H;��H;��H;w�H;��H;�H;��H;�H;��H;w�H;��H;��H;��H;R�H;N�H;M�H;y�H;̀H;-dH;m@H;�H;��G;}8G;�2F;CD;��@;�:;��0;��!;�Y;��:*u�:Y�9���0Ⱥx.�3|��R��/Tʻ�����S�	�      ɪx��[t���g�YT�g�:����'���7����1��^�(�HW��@�t��n`:a��:�\;{ ;��0;a;;=A;�D;�wF;�cG;Y�G;�!H;�MH;�oH;{�H;��H;̯H;��H;m�H;��H;`�H;v�H;�H;��H;-�H;��H;�H;v�H;`�H;��H;m�H;��H;ƯH;��H;x�H;�oH;�MH;�!H;X�G;�cG;�wF;�D;=A;d;;��0;{ ;�\;a��:�n`:��t�LW��^�(��1��8���(������g�:�ZT���g��[t�      >,˼��Ǽ�"���뮼w��+G��5�[�jy-�����.��ܕb��0㺸ط�5<:�L�:�\;��!;�J2;�g<;V0B;1CE;/�F;U�G;��G;�4H;�\H;|H;��H;��H;`�H;��H;G�H;��H;Z�H;Z�H;�H;��H;�H;X�H;X�H;��H;J�H;��H;_�H;��H;��H;|H;�\H;�4H;��G;O�G;0�F;1CE;X0B;�g<;�J2;��!;�\;�L�:5<:�ط��0�ܕb��.�����jy-�5�[�*G��w���뮼�"����Ǽ      0���k��Nv��t�J�Ѽ�뮼2X��w�W������׻Ȅ�"��8��5<:a��:�Y;�t%;�$5;�Z>;aC;��E;9*G;i�G;H;HH;slH;��H;	�H;ɯH;׼H;��H;��H;�H;~�H;v�H;6�H;v�H;~�H;�H;��H;��H;׼H;ɯH;	�H;��H;plH;HH;H;h�G;7*G;��E;aC;�Z>;�$5;�t%;�Y;a��:
5<:8�� ��Ȅ� �׻���w�W�2X���뮼I�Ѽ�t�Nv���k�      Jm��Fi��&^�e�L�U�6�,����'}ռuT����x�Ȼ0�������#���ط��n`:��: �;+�*;<�8;�@;=�D;l�F;�}G;��G;�1H;�[H;s|H;ÕH;ߨH;��H;��H;��H;��H;��H;��H;{�H;��H;��H;��H;��H;��H;��H;ߨH;��H;s|H;�[H;�1H;��G;�}G;h�F;=�D;�@;>�8;+�*;"�;��:�n`:�ط�"��������Ȼ0���x�uT��'}ռ��,��U�6�e�L��&^��Fi�      Q��v;��D�������섽~�e��?��k��t�鷼"G���e7����Ȅ��0㺀�t�*u�:	,�:{;�1;T�<;f�B;+�E;�G;��G;dH;uJH;aoH;�H;��H;�H;��H;��H;%�H;��H;�H;��H;�H;��H;"�H;��H;��H;�H;��H;�H;aoH;uJH;eH;��G;�G;(�E;f�B;X�<;�1;{;,�:(u�: �t��0�Ȅ���껌e7�"G��鷼�t��k��?�~�e��섽���D���v;��      v���)��s��ӽ�'��C�������Z��Q+�����"��"G��Ȼ0��׻ڕb�JW�� Y�9֡�:,`;�*';�Y7;$@;+�D;��F;�G;��G;;8H;bH;�H;\�H;��H;w�H;��H;��H;��H;U�H;A�H;U�H;��H;��H;��H;x�H;��H;\�H;��H;bH;:8H;��G;�G;��F;(�D;$@;�Y7;�*';*`;ء�:�X�9LW��ܕb��׻ɻ0�"G���"������Q+��Z����C����'���ӽ�s�*��      �!,�<)��K ���������޽"������Fi��0����鷼��x�����.��_�(�����*i:���:>�;��0;M�<;�C;��E;=G;��G;�$H;gTH;�wH;�H;�H;Q�H;��H;C�H;��H;��H;�H;��H;��H;C�H;��H;Q�H;�H;�H;�wH;hTH;�$H; �G;=G;��E;�C;O�<;��0;<�;���: +i: ��`�(��.�������x�鷼����0��Fi����"����޽�������K �<)�      ,�j��f��Z�|�F��>/��^�s����ŽJ ���Fi��Q+��t�uT��x�W�����1��4Ⱥ X�9�P�:�Y;��(;
�8;�A;�E;�F;k�G;�H;�FH;�mH;��H;ġH;C�H;r�H;��H;��H;��H;��H;��H;��H;��H;p�H;C�H;ġH;��H;�mH;�FH;�H;m�G;	�F;�E;�A;
�8;��(;�Y;�P�:X�9:Ⱥ�1�����x�W�uT���t�Q+��Fi�J ���Žs����^��>/�|�F��Z��f�      ��y���{�J����f��SC��K �sn���Ž����Z��k�'}ռ2X��iy-�7���w.����P�:�+�:��;4;7�>;�D;�wF;5�G;��G;�9H;ZdH;v�H;��H;d�H;t�H;��H;��H;X�H;u�H;Y�H;��H;��H;q�H;f�H;��H;v�H;WdH;�9H;��G;4�G;�wF;�D;9�>;4;��;�+�:�P�:���z.�8���iy-�2X��'}ռ�k��Z�����Žsn���K ��SC��f�J���{�y���      ��˾��Ǿ����"���X͓�_�x���J��K �s���"������?����뮼5�[�+���"3|��W��x�:f�:�';n/;fg<;�C;iF;�NG;��G;/-H;o[H;�}H;ɗH;ʪH;¸H;��H;�H;��H;�H;��H;�H;��H;��H;ʪH;ɗH;�}H;n[H;/-H;��G;�NG;mF;�C;dg<;n/;�';d�:x�:�W��$3|�,���5�[��뮼���?����"��s����K ���J�_�x�X͓�!���������Ǿ      u� ��������{Ծm���x���^�x��SC��^���޽C���~�e�,��K�Ѽ+G������R����� ݤ8釲:�Y;P�);��9;��A;��E;�G;�G;h!H;BSH;�wH;x�H;��H;F�H;��H;}�H;��H;��H;��H;}�H;��H;C�H;��H;x�H;�wH;>SH;i!H;�G;�G;��E;��A;��9;P�);�Y;뇲: ݤ8����R�����+G��K�Ѽ,��~�e�C�����޽�^��SC�^�x�x���m����{Ծ�쾣���      ��� E�l�u� �Y�ݾm���X͓��f��>/�����'���섽T�6��t�w��g�:�0Tʻ�.�h۷�ft�:�;��$;�Y7;X�@;�	E;�F;9�G;�H;?LH;�rH;��H;ΤH;'�H;&�H;7�H;O�H;��H;O�H;6�H;&�H;%�H;ФH;��H;�rH;<LH;�H;;�G;�F;�	E;U�@;�Y7;��$;�;ft�:`۷��.�1Tʻg�:�w���t�T�6��섽�'������>/��f�X͓�m���Y�ݾu� �l� E�      ��7�v3�1�'����u� ��{Ծ!���J���|�F�����ӽ���e�L�Nv��뮼[T����PV���=��)i:\��:�z ;�$5;��?;	�D;κF;��G;�H;�FH;�nH;��H;��H;t�H;�H;=�H;\�H;��H;\�H;=�H;�H;r�H;��H;��H;�nH;�FH;�H;��G;κF;�D;��?;�$5;�z ;^��:�)i:��=��PV����[T��뮼Nv�e�L�����ӽ���|�F�J���!����{Ծu� ����1�'�v3�      �N��TI���;�1�'�l��쾂���{󐾸Z��K ��s�D����&^���"����g�����u�!��3<:���: ;fg3;��>;xBD;��F;�G;�H;LBH;ykH;[�H;�H;1�H;޼H;v�H;��H;N�H;��H;v�H;޼H;/�H;�H;[�H;vkH;JBH;�H;�G;��F;vBD;��>;hg3; ;���:3<:!���u������g��"����&^�D����s潨K ��Z�{󐾂�����l�1�'���;��TI�      c]�g�W��TI�v3� E�������Ǿy����f�<)�)��v;���Fi��k���Ǽ�[t�T�	�6Ȅ�6X���:���:��;YJ2;NZ>;F	D;{F;C�G;H;�?H;�iH;�H;�H;z�H;A�H;��H;`�H;��H;`�H;��H;A�H;y�H;�H;�H;�iH;�?H;H;B�G;{F;F	D;KZ>;^J2;��;���:�:6X��6Ȅ�T�	��[t���Ǽ�k��Fi�v;��*��<)��f�y�����Ǿ���� E�v3��TI�g�W�      �?��~h��?v��� ��9�X��O/�2y�C�;㰖��+X����ѽ����dn;�c�������B(�⚩�b�� �e9�:�;�Y.;O�<;�WC;![F;��G;'0H;ojH;S�H;s�H;��H;O�H;��H;��H;��H;��H;��H;��H;��H;N�H;��H;s�H;Q�H;ljH;'0H;��G;"[F;�WC;M�<;�Y.;�;�:�e9b��⚩��B(�����c��dn;������ѽ���+X�㰖�C�;2y��O/�9�X�� ��?v��~h��      ~h��1���c�����y�YvS�rM+��v�9ɾ�����T�"]�\ν����}\8�����x��%�V���~��0�9X-�:p�;��.;�<;�nC;�dF;�G;�1H;kH;ŌH;ѤH;�H;��H;��H;��H;��H;��H;��H;��H;��H;��H;�H;ѤH;H;kH;�1H;�G;�dF;�nC;�<;��.;p�;X-�:(�9~��V���	%��x�����}\8�����\ν"]��T�����9ɾ�v�sM+�YvS���y�c���1���      ?v��c���X ��c�h�9E�Z��m���~㼾���nH�ֈ�}�ý�Ȅ��s/��o��#�����,J��2к@
�9Dg�:�l;S0;]=;��C;�F;y�G;D6H;ZmH;F�H;ХH;��H;&�H;n�H;��H;1�H;�H;1�H;��H;o�H;#�H;��H;ХH;A�H;WmH;D6H;y�G;�F;��C;]=;V0;�l;@g�:(
�90к,J������#���o��s/��Ȅ�}�ýֈ��nH���~㼾m���Z��9E�c�h�X ��c���      � ����y�c�h��N��O/����E�߾B���*|��6�s}�䳽oSt�A�!�vrμIF{��_��X��֓���:��:�Z;�2;�O>;�D;g�F;��G;?=H;�pH;��H;u�H;�H;�H;�H;��H;��H;��H;��H;��H;
�H;�H;�H;u�H;��H;�pH;?=H;��G;f�F;�D;�O>;�2;�Z;��:�:֓���X���_�HF{�vrμA�!�oSt�䳽s}��6��*|�B��E�߾����O/��N�c�h���y�      9�X�YvS�9E��O/��S�LW����������OS\��� ���>����Y�~��փ����]�����0�b���Y���Y:��:s`;b�4;�?;_�D;�F;�G;+FH;zuH;ޓH;��H;��H;?�H;��H;O�H;D�H;%�H;D�H;N�H;��H;=�H;��H;��H;ۓH;yuH;,FH;�G;�F;]�D;�?;d�4;s`;��:��Y:��Y�/�b�������]�փ��~���Y�>����彔� �OS\���������LW���S��O/�9E�YvS�      �O/�rM+�Z�����LW��9ɾB���Mw�� :�l��{�ý M��an;�e���yv���E<��˻��-����y�:�^;�%;��7;��@;:5E;�"G;�G;bPH;2{H;��H;��H;��H;��H;$�H;=�H;�H;��H;�H;=�H;$�H;��H;��H;��H;ݗH;.{H;aPH;�G;�"G;85E;}�@;��7;�%;�^;�y�:����-��˻�E<�yv��e���an;� M��{�ýl��� :��Mw�B��9ɾLW�����Z��rM+�      2y��v�m���E�߾����C��A����nH���Gὠu����d�3O�prμN"�����
	����뺐r89�;�:c�;�+;z|:;�7B;�E;2bG;�H;[H;��H;J�H;ƯH;$�H;r�H;r�H;5�H;�H;��H;�H;5�H;t�H;r�H;$�H;ƯH;I�H;��H;[H;�H;4bG;�E;�7B;y|:;�+;d�;�;�:�r89���
	�����N"��prμ3O���d��u��G����nH�A���C������E�߾m����v�      C�;9ɾ~㼾B�������Mw��nH�����Z�䳽͕��v\8�v#������^N�U��
�b�Ix�P5:��:6�;��0;D]=;R�C;�[F;�G;�)H;fH;��H;D�H;j�H;��H;F�H;��H;[�H;��H;��H;��H;[�H;��H;D�H;��H;k�H;D�H;��H;fH;�)H;�G;�[F;P�C;C]=;��0;6�;��:P5:Ix��b�U��^N�����v#��v\8�͕��䳽�Z񽳯��nH��Mw�����B��~㼾9ɾ      㰖��������*|�OS\�� :����Z�o$�������K�y���Oļ����������>&����V/�:�^;��#;�G6;`�?;�D;r�F;��G; @H;�pH;�H;��H;=�H;|�H;W�H;��H;��H;�H;��H;�H;��H;��H;W�H;}�H;=�H;��H;�H;�pH;@H;��G;o�F;�D;_�?;�G6;��#;�^;V/�:���>&������������Oļy���K�����o$���Z���� :�OS\��*|�������      �+X��T��nH��6��� �l��G�䳽�����mR����ټ�����E<��?ݻ<d\����� !:�d�:��;6�,;��:;�7B;��E;�LG;aH;~SH;�{H;��H;�H;@�H;j�H;{�H;:�H;��H;�H;��H; �H;��H;;�H;z�H;m�H;@�H;�H;��H;�{H;}SH;`H;�LG;��E;7B;��:;6�,;��;�d�:!:����;d\��?ݻ�E<�����ټ����mR�����䳽G�l���� ��6��nH��T�      ��"]�ֈ�s}���{�ý�u��͕���K�����o�nv���&R�#��Z^��~�� p>���:nB;Z";z�4;��>;fD;��F;�G;�)H;�dH;��H;=�H;��H;W�H;Z�H;��H;��H;N�H;:�H;��H;:�H;N�H;��H;��H;\�H;W�H;��H;:�H;��H;�dH;�)H;�G;��F;cD;��>;z�4;W";nB;��: t>�|��Z^��#���&R�nv���o�����K�͕���u��{�ý��s}�ֈ�"]�      �ѽ\ν}�ý䳽>��� M����d�v\8�y��ټnv����Y��_����@���[���Y:l��:^m;�r-;!�:;��A;VoE;�"G;y�G;�GH;�sH;�H;��H;�H;V�H;C�H;��H;��H;��H;T�H;�H;T�H;��H;��H;��H;F�H;V�H;�H;��H;�H;�sH;�GH;s�G;�"G;ToE;��A;!�:;�r-;`m;r��:��Y:�[�?������_���Y�nv��ټy��v\8���d� M��>���䳽}�ý\ν      ���������Ȅ�oSt��Y�an;�3O�v#���Oļ�����&R��_������N3�̅Y�4:$�:ޯ;�?&;�G6;�X?;�D;QxF;ܚG;[!H;�^H;��H;�H;��H;k�H;0�H;&�H;��H;<�H;�H;~�H;<�H;~�H;�H;<�H;��H;(�H;0�H;i�H;��H;�H;��H;�^H;X!H;ךG;MxF;�D;�X?;�G6;�?&;�;"�:4:ȅY��N3������_��&R������Oļv#��3O�an;��Y�oSt��Ȅ�����      dn;�|\8��s/�A�!�~��d���orμ��������E<�"������N3�@Hx���9�:�^;b ;B2;��<;�B;˲E;W5G;*�G;YFH;�qH;ʎH;r�H;ߴH;v�H;��H;��H;)�H;��H;F�H;��H;6�H;��H;F�H;��H;(�H;��H;��H;v�H;ݴH;r�H;ȎH;�qH;XFH;'�G;R5G;˲E;�B;��<;B2;d ;�^;�:�98Hx��N3����"���E<��������orμd���~��A�!��s/�|\8�      b������o�vrμփ��yv��N"��^N�����?ݻZ^��C��ЅY���9�:��:��;`�.;�|:;?A;��D;M�F;ֶG;*H;CaH;=�H;��H;�H;c�H;F�H;c�H;��H;$�H;E�H;��H;��H;
�H;��H;��H;F�H;$�H;��H;c�H;D�H;`�H;�H;��H;@�H;@aH;*H;ѶG;K�F;��D;?A;�|:;c�.;��;��:�:��9ЅY�C��Z^���?ݻ���^N�N"��xv��փ��vrμ�o����      �����x���#��GF{���]��E<����U�뻭���:d\�|�뺤[�4:�:���:�[;|�,;��8;7!@;�0D;�[F;C{G;H;jPH;?vH;�H;i�H;&�H;W�H;��H;��H;�H;�H;��H;��H;��H;��H;��H;��H;��H;�H;�H;��H;��H;S�H;$�H;e�H;�H;<vH;ePH;H;B{G;�[F;�0D;7!@;��8;z�,;�[;���:�:4:�[�|��<d\�����T�뻨���E<���]�GF{��#���x��      �B(�%�����_������˻	���b�>&����� h>���Y:"�:�^;��;x�,;&`8;u�?;�C;�F;GG;l�G;@H;OkH;'�H;,�H;�H;~�H;��H;��H;��H;D�H;��H;	�H;��H;��H;��H;��H;��H;�H;��H;D�H;��H;��H;��H;}�H;�H;/�H;'�H;KkH;@H;l�G;GG;�F;�C;y�?;&`8;x�,;��;�^;"�:��Y: l>�����<&��b�	���˻�����_����%�      㚩�V���*J���X��0�b��-����Ix����!:��:j��:�;` ;c�.;��8;x�?;�C;��E;[#G;�G;2H;bH;o�H;��H;��H;ԷH;
�H;��H;A�H;`�H;c�H;�H;B�H;��H;d�H;��H;d�H;��H;B�H;�H;c�H;`�H;@�H;��H;
�H;зH;��H;��H;l�H;bH;2H;	�G;\#G;��E;�C;u�?;��8;c�.;b ;�;l��:��:!:���Ix������-�+�b��X��*J��Z���      R��z��кȓ����Y���� s89P5:\/�:�d�:pB;`m;�?&;D2;�|:;7!@;�C;��E;�G;��G;}(H;![H;�zH;d�H;�H;ɳH;��H;��H;��H;��H;��H;&�H;y�H;Z�H;x�H;(�H;��H;)�H;x�H;Z�H;x�H;&�H;��H;��H;��H;��H;��H;˳H;�H;b�H;�zH;![H;z(H;��G;�G;��E;߳C;7!@;�|:;D2;�?&;am;rB;�d�:b/�:L5: s89�����Y�ʓ��кx��      @�e9��9h
�9�:��Y:�y�:�;�:��:�^;��;X";�r-;�G6;��<;?A;�0D;�F;X#G;��G;%H;�WH;�vH;��H;j�H;p�H;��H;9�H;��H;��H;d�H;�H;��H;��H;V�H;:�H;��H;&�H;��H;:�H;V�H;��H;��H; �H;a�H;��H;��H;7�H;��H;o�H;e�H;��H;�vH;�WH;%H;��G;X#G;�F;�0D;?A;��<;�G6;�r-;X";��;�^;��:�;�:�y�:��Y:�:h
�9��9      �:�-�:Rg�:��:��:�^;i�;6�;��#;:�,;z�4;�:;�X?;�B;��D;�[F;GG;�G;}(H;�WH;�uH;��H;>�H;%�H;N�H;%�H;��H;�H;�H;��H;��H;�H;��H;�H;��H;��H;��H;��H;��H;�H;��H;�H;��H;��H;�H;�H;��H;#�H;K�H; �H;=�H;��H;�uH;�WH;}(H;�G;GG;�[F;��D;�B;�X?;�:;z�4;:�,;��#;6�;i�;�^;��:��:Tg�:`-�:      ;��;m;�Z;w`;�%;�+;��0;�G6;��:;��>;��A;�D;̲E;P�F;B{G;n�G;2H; [H;�vH;��H;w�H;�H;��H;��H;��H;��H;��H;��H;�H;m�H;f�H;��H;��H;��H;��H;	�H;��H;��H;��H;��H;f�H;k�H;�H;��H;��H;��H;��H;��H;�H;�H;u�H;��H;�vH; [H;2H;l�G;B{G;P�F;̲E;�D;��A;��>;��:;�G6;��0;�+;�%;�`;�Z;m;��;      �Y.;��.;X0;�2;`�4;��7;�|:;H]=;d�?;�7B;gD;YoE;QxF;W5G;ֶG;H;@H;bH;�zH;��H;>�H;�H;v�H;��H;��H;��H;��H;&�H;M�H;��H;��H;��H;��H;u�H;�H;N�H;x�H;N�H;�H;v�H;��H;��H;��H;��H;I�H;$�H;��H;��H;��H;��H;u�H;�H;9�H;��H;�zH;bH;@H;H;ֶG;W5G;PxF;YoE;iD;�7B;f�?;H]=;�|:;��7;h�4;�2;X0;��.;      g�<;-�<;,]=;�O>;��?;��@;�7B;T�C;�D;��E;��F;�"G;ۚG;+�G;*H;hPH;MkH;r�H;c�H;i�H;!�H;��H;��H;e�H;a�H;e�H;w�H;��H;Q�H;k�H;+�H;>�H;;�H;�H;q�H;��H;��H;��H;s�H;�H;8�H;@�H;+�H;h�H;M�H;��H;v�H;e�H;a�H;a�H;��H;��H;�H;h�H;b�H;r�H;KkH;hPH;*H;+�G;ٚG;�"G;��F;��E;�D;U�C;�7B;��@; �?;�O>;,]=;�<;      �WC;oC;�C;�D;f�D;A5E;�E;�[F;s�F;�LG;�G;|�G;[!H;_FH;FaH;AvH;0�H;��H;	�H;w�H;Q�H;��H;��H;h�H;%�H;8�H;q�H;��H;�H;��H;
�H;��H;��H;f�H;��H;�H;�H;	�H;��H;e�H;��H;��H;
�H;��H;�H;��H;o�H;7�H;&�H;e�H;��H;��H;N�H;v�H;�H;��H;*�H;?vH;EaH;\FH;[!H;|�G;�G;�LG;v�F;�[F;�E;A5E;h�D;�D;�C;oC;      2[F;�dF;�F;j�F;�F;�"G;7bG;�G;��G;bH;�)H;�GH;�^H;�qH;=�H;�H;.�H;��H;ƳH;��H;"�H;�H;��H;e�H;1�H;\�H;��H;��H;��H;��H;��H;��H;W�H;��H;�H;F�H;F�H;F�H;�H;��H;S�H;��H;��H;��H;��H;��H;��H;Z�H;3�H;d�H;��H;��H;�H;��H;ųH;��H;,�H;�H;=�H;�qH;�^H;�GH;�)H;bH;��G;�G;7bG;�"G;�F;j�F;�F;�dF;      �G;��G;��G;��G;(�G;&�G;�H;*H;$@H;SH;�dH;�sH;��H;ˎH;��H;i�H;�H;ҷH;��H;<�H;��H;��H;��H;}�H;k�H;��H;��H;s�H;��H;��H;��H;+�H;��H;�H;7�H;i�H;��H;i�H;6�H;�H;��H;(�H;��H;��H;��H;q�H;��H;��H;m�H;y�H;��H;��H;��H;:�H;��H;ӷH;�H;h�H;��H;ˎH;��H;�sH;�dH;SH;&@H;*H;�H;#�G;-�G;��G;}�G;��G;      #0H;�1H;R6H;>=H;5FH;hPH;[H;fH;�pH;�{H;��H;�H;�H;v�H;�H;&�H;~�H;�H;��H;��H;�H;��H;&�H;��H;��H;��H;p�H;��H;��H;��H;2�H;��H;��H;A�H;u�H;��H;z�H;��H;u�H;A�H;��H;��H;1�H;��H;��H;��H;p�H;��H;��H;��H;#�H;��H;�H;��H;��H;�H;|�H;&�H;�H;u�H;�H;�H;��H;�{H;�pH;fH;[H;iPH;@FH;?=H;P6H;�1H;      �jH;%kH;^mH;�pH;�uH;5{H;��H;��H;�H;��H;A�H;��H;��H;�H;d�H;X�H;��H;��H;��H;��H;	�H;��H;J�H;T�H;�H;��H;��H;��H;��H; �H;��H;��H;(�H;d�H;��H;��H;��H;��H;��H;d�H;%�H;��H;��H;�H;��H;��H;��H;��H;�H;T�H;H�H;��H;�H;��H;��H;��H;��H;W�H;c�H;�H;��H;��H;@�H;��H;�H;��H;��H;5{H;�uH;�pH;^mH;kH;      e�H;ьH;T�H;��H;�H;�H;T�H;N�H;��H;�H;��H;!�H;s�H;��H;J�H;��H;��H;?�H;��H;h�H;��H;�H;��H;l�H;��H;��H;��H;��H;�H;{�H;��H;.�H;d�H;��H;��H;��H;��H;��H;��H;��H;b�H;/�H;��H;z�H;�H;��H;��H;��H;��H;k�H;��H;�H;��H;g�H;��H;?�H;��H;��H;J�H;�H;s�H;�H;��H;�H;��H;P�H;T�H;�H;�H;��H;O�H;͌H;      |�H;�H;�H;��H;ΩH;��H;ԯH;{�H;I�H;H�H;a�H;d�H;7�H;��H;g�H;��H;��H;a�H;��H;�H;��H;k�H;��H;.�H;�H;��H;��H;5�H;��H;��H;)�H;[�H;��H;��H;��H;��H;��H;��H;��H;��H;��H;\�H;)�H;��H;��H;5�H;��H;��H;�H;.�H;��H;k�H;��H;�H;��H;a�H;��H;��H;g�H;��H;7�H;a�H;a�H;K�H;K�H;{�H;ԯH;��H;˩H;��H;�H;�H;      εH;�H;ŶH;�H;��H;��H;+�H;��H;��H;q�H;e�H;Q�H;/�H;��H;��H;�H;M�H;d�H;*�H;��H;�H;j�H;��H;B�H;��H;��H;(�H;��H;��H;/�H;Y�H;t�H;��H;��H;��H;��H;��H;��H;��H;��H;��H;u�H;Y�H;2�H;��H;��H;*�H;��H;��H;B�H;��H;j�H;�H;��H;*�H;e�H;L�H;�H;��H;��H;-�H;P�H;e�H;q�H;��H;��H;,�H;��H;��H;�H;ĶH;�H;      Y�H;��H;4�H;�H;M�H;��H;w�H;Q�H;a�H;��H;��H;��H;�H;2�H;*�H;�H;��H;�H;|�H;��H;��H;��H;��H;B�H;��H;U�H;��H;��H;+�H;j�H;��H;��H;��H;��H;��H;��H;��H;��H;��H;��H;��H;��H;��H;k�H;,�H;��H;��H;U�H;��H;A�H;��H;��H;��H;��H;|�H;�H;��H;�H;'�H;2�H;�H;��H;��H;��H;b�H;Q�H;w�H;��H;F�H;�H;3�H;��H;      ��H;�H;o�H;�H;�H;"�H;{�H;�H;��H;A�H;��H;��H;B�H;��H;J�H;��H;�H;B�H;\�H;]�H;"�H;��H;u�H;�H;_�H;��H;	�H;A�H;d�H;��H;��H;��H;��H;��H;��H;��H;��H;��H;��H;��H;��H;��H;��H;��H;g�H;A�H;�H;��H;a�H;�H;s�H;��H;!�H;]�H;\�H;C�H;�H;��H;I�H;��H;B�H;��H;��H;A�H;��H;�H;{�H;(�H;��H;�H;o�H;
�H;      ��H;��H;�H;��H;n�H;=�H;B�H;l�H;��H;��H;X�H;��H;�H;P�H;��H;��H;��H;��H;z�H;A�H; �H;��H;�H;w�H;��H;�H;2�H;u�H;��H;��H;��H;��H;��H;��H;��H;��H;��H;��H;��H;��H;��H;��H;��H;��H;��H;u�H;2�H;�H;��H;v�H;�H;��H;��H;A�H;z�H;��H;��H;��H;��H;P�H;�H;��H;W�H;��H;��H;i�H;A�H;A�H;d�H;��H;�H;��H;      ��H;�H;A�H;��H;Z�H;�H;�H;�H;�H;!�H;E�H;a�H;��H;��H;��H;��H;��H;`�H;,�H;��H;��H;��H;N�H;��H;�H;C�H;f�H;��H;��H;��H;��H;��H;��H;��H;��H;��H;��H;��H;��H;��H;��H;��H;��H;��H;��H;��H;f�H;A�H;�H;��H;N�H;��H;��H;��H;,�H;b�H;��H;��H;��H;��H;��H;a�H;D�H;%�H;�H;�H;�H;�H;N�H;��H;A�H; �H;      ��H;��H;#�H;��H;<�H;��H;��H;��H;��H;��H;�H;&�H;C�H;@�H;�H;��H;��H;��H;��H;,�H;��H;�H;w�H;��H;��H;A�H;��H;�H;��H;��H;��H;��H;��H;��H;��H;��H;��H;��H;��H;��H;��H;��H;��H;��H;��H;�H;��H;C�H;��H;��H;w�H;�H;��H;,�H;��H;��H;��H;��H;�H;@�H;C�H;&�H;�H;��H;��H;��H;��H;��H;/�H;��H;#�H;��H;      ��H;�H;A�H;��H;Z�H;�H;�H;�H;�H;!�H;E�H;a�H;��H;��H;��H;��H;��H;`�H;,�H;��H;��H;��H;N�H;��H;�H;C�H;g�H;��H;��H;��H;��H;��H;��H;��H;��H;��H;��H;��H;��H;��H;��H;��H;��H;��H;��H;��H;f�H;A�H;�H;��H;N�H;��H;��H;��H;,�H;b�H;��H;��H;��H;��H;��H;a�H;E�H;"�H;�H;�H;�H;�H;N�H;��H;<�H;��H;      ��H;��H;�H;��H;p�H;=�H;B�H;l�H;��H;��H;W�H;��H;�H;P�H;��H;��H;��H;��H;z�H;A�H;�H;��H;�H;w�H;��H;�H;2�H;u�H;��H;��H;��H;��H;��H;��H;��H;��H;��H;��H;��H;��H;��H;��H;��H;��H;��H;u�H;2�H;�H;��H;t�H;�H;��H;��H;A�H;z�H;��H;��H;��H;��H;P�H;�H;��H;W�H;��H;��H;i�H;B�H;A�H;d�H;��H;�H;��H;      ��H;�H;o�H;�H;�H;"�H;{�H;�H;��H;A�H;��H;��H;B�H;��H;I�H;��H;�H;B�H;\�H;]�H;&�H;��H;s�H;�H;a�H;��H;�H;A�H;d�H;��H;��H;��H;��H;��H;��H;��H;��H;��H;��H;��H;��H;��H;��H;��H;g�H;A�H;�H;��H;_�H;�H;u�H;��H;"�H;]�H;\�H;C�H;�H;��H;L�H;��H;B�H;��H;��H;A�H;��H;�H;{�H;'�H;��H;�H;o�H;
�H;      \�H;��H;6�H;�H;J�H;��H;w�H;Q�H;a�H;��H;��H;��H;�H;2�H;'�H;�H;��H;�H;|�H;��H;��H;��H;��H;A�H;��H;W�H;��H;��H;+�H;j�H;��H;��H;��H;��H;��H;��H;��H;��H;��H;��H;��H;��H;��H;k�H;,�H;��H;��H;U�H;��H;A�H;��H;��H;��H;��H;|�H;�H;��H;�H;*�H;2�H;�H;��H;��H;��H;a�H;N�H;w�H;��H;D�H;�H;3�H;��H;      еH;�H;ǶH;�H;��H;��H;.�H;��H;��H;r�H;e�H;Q�H;-�H;��H;��H;�H;N�H;d�H;*�H;��H;�H;j�H;��H;D�H;��H;��H;(�H;��H;��H;0�H;Y�H;t�H;��H;��H;��H;��H;��H;��H;��H;��H;��H;u�H;Y�H;0�H;��H;��H;*�H;��H;��H;B�H;��H;j�H;�H;��H;*�H;e�H;L�H;�H;��H;��H;/�H;P�H;e�H;r�H;��H;��H;.�H;��H;��H;�H;ǶH;�H;      |�H;�H;�H;��H;ΩH;��H;ԯH;{�H;I�H;I�H;a�H;a�H;7�H;��H;i�H;��H;��H;`�H;��H;�H;��H;k�H;��H;/�H;�H;��H;��H;5�H;��H;��H;)�H;[�H;��H;��H;��H;��H;��H;��H;��H;��H;��H;\�H;)�H;��H;��H;5�H;��H;��H;�H;.�H;��H;k�H;��H;�H;��H;a�H;��H;��H;g�H;��H;7�H;d�H;`�H;I�H;I�H;{�H;ԯH;��H;ʩH;��H;�H;�H;      ^�H;ьH;R�H;��H;�H;�H;V�H;P�H;��H;�H;��H;!�H;r�H;��H;J�H;��H;��H;=�H;��H;h�H;��H;�H;��H;l�H;��H;��H;��H;��H;�H;{�H;��H;.�H;c�H;��H;��H;��H;��H;��H;��H;��H;c�H;/�H;��H;z�H;�H;��H;��H;��H;��H;k�H;��H;�H;��H;h�H;��H;@�H;��H;��H;J�H;�H;r�H;!�H;��H;�H;��H;P�H;V�H;�H;�H;��H;T�H;ЌH;      �jH; kH;dmH;�pH;�uH;1{H;��H;��H;�H;��H;A�H;��H;��H;�H;c�H;W�H;��H;��H;��H;��H;
�H;��H;I�H;T�H;�H;��H;��H;��H;��H;�H;��H;��H;'�H;d�H;��H;��H;��H;��H;��H;d�H;'�H;��H;��H;�H;��H;��H;��H;��H;�H;T�H;I�H;��H;�H;��H;��H;��H;��H;Z�H;d�H;�H;��H;��H;A�H;��H;�H;��H;��H;2{H;�uH;�pH;bmH; kH;      #0H;�1H;P6H;?=H;3FH;iPH;[H;fH;�pH;�{H;��H;�H;�H;v�H;�H;&�H;~�H;�H;��H;��H;�H;��H;$�H;��H;��H;��H;p�H;��H;��H;��H;1�H;��H;��H;@�H;t�H;��H;z�H;��H;u�H;A�H;��H;��H;2�H;��H;��H;��H;p�H;��H;��H;��H;$�H;��H;�H;��H;��H;�H;|�H;'�H;�H;u�H;�H;�H;��H;�{H;�pH;fH;[H;ePH;=FH;>=H;P6H;�1H;      �G;��G;}�G;��G;#�G;"�G;�H;*H;$@H;�SH;�dH;�sH;��H;ˎH;��H;i�H;�H;ҷH;��H;=�H;��H;��H;��H;|�H;m�H;��H;��H;q�H;��H;��H;��H;*�H;��H;�H;6�H;i�H;��H;g�H;7�H;�H;��H;-�H;��H;��H;��H;s�H;��H;��H;k�H;z�H;��H;��H;��H;:�H;��H;ӷH;�H;h�H;��H;ˎH;��H;�sH;�dH;�SH;$@H; *H;�H; �G;(�G;��G;|�G;�G;      9[F;�dF;�F;j�F;�F;�"G;8bG;�G;��G;dH;�)H;�GH;�^H;�qH;<�H;�H;.�H;��H;ųH;��H;#�H;��H;��H;e�H;3�H;Z�H;��H;��H;��H;��H;��H;��H;T�H;��H;�H;F�H;F�H;F�H;�H;��H;T�H;��H;��H;��H;��H;��H;��H;\�H;1�H;d�H;��H;�H;�H;��H;ƳH;��H;,�H;�H;=�H;�qH;�^H;�GH;�)H;bH;��G;�G;9bG;�"G;�F;m�F; �F;�dF;      �WC;oC;�C;�D;f�D;A5E;�E;�[F;v�F;�LG; �G;|�G;[!H;\FH;EaH;@vH;-�H;��H;�H;v�H;Q�H;��H;��H;h�H;&�H;7�H;o�H;��H;�H;��H;
�H;��H;��H;e�H;��H;	�H;�H;�H;��H;e�H;��H;��H;
�H;��H;�H;��H;q�H;8�H;%�H;g�H;��H;��H;O�H;w�H;	�H;��H;,�H;AvH;FaH;]FH;[!H;|�G;�G;�LG;s�F;�[F;�E;A5E;d�D;�D;�C;oC;      k�<;+�<;2]=;�O>;�?;��@;�7B;T�C;�D;��E;��F;�"G;ۚG;+�G;*H;hPH;LkH;o�H;b�H;h�H;!�H;��H;��H;e�H;a�H;e�H;w�H;��H;O�H;k�H;+�H;>�H;:�H;�H;p�H;��H;��H;��H;s�H;�H;:�H;@�H;+�H;h�H;N�H;��H;v�H;e�H;a�H;b�H;��H;��H;�H;i�H;c�H;s�H;LkH;hPH;*H;+�G;ٚG;�"G;��F;��E;�D;T�C;�7B;��@; �?;�O>;5]=;�<;      �Y.;��.;e0;�2;\�4;��7;�|:;H]=;d�?;�7B;iD;YoE;NxF;W5G;ֶG;H;@H;bH;�zH;��H;>�H;�H;u�H;��H;��H;��H;��H;$�H;L�H;��H;��H;��H;��H;v�H;�H;N�H;x�H;N�H;�H;u�H;��H;��H;��H;��H;J�H;&�H;��H;��H;��H;��H;v�H;�H;:�H;��H;�zH;bH;@H;H;׶G;W5G;PxF;XoE;gD;7B;f�?;G]=;�|:;��7;b�4;�2;]0;��.;      ;��;m;�Z;v`;�%;�+;��0;�G6;��:;��>;��A;�D;̲E;N�F;C{G;l�G;2H; [H;�vH;��H;u�H;�H;��H;��H;��H;��H;��H;��H;�H;k�H;f�H;��H;��H;��H;��H;	�H;��H;��H;��H;��H;f�H;m�H;�H;��H;��H;��H;��H;��H;��H;�H;w�H;��H;�vH; [H;2H;l�G;B{G;Q�F;̲E;�D;��A;��>;��:;�G6;��0;�+;�%;�`;�Z;m;��;      �:x-�:Vg�:��:��:�^;k�;8�;��#;:�,;z�4;�:;�X?;�B;��D;�[F;GG;�G;}(H;�WH;�uH;��H;=�H;%�H;K�H;#�H;��H;�H;�H;��H;��H;�H;��H;�H;��H;��H;��H;��H;��H;�H;��H;�H;��H;��H;�H;�H;��H;%�H;N�H;!�H;>�H;��H;�uH;�WH;}(H;�G;GG;�[F;��D;�B;�X?;�:;z�4;6�,;��#;8�;k�;�^;��:��:Zg�:`-�:       �e9��9�
�9�:��Y:�y�:�;�:��:�^;��;X";�r-;�G6;��<;?A;�0D;�F;V#G;��G;%H;�WH;�vH;��H;j�H;o�H;��H;:�H;��H;��H;d�H; �H;��H;��H;V�H;:�H;��H;&�H;��H;:�H;V�H;��H;��H;�H;a�H;��H;��H;7�H;��H;p�H;f�H;��H;�vH;�WH;%H;��G;Y#G;�F;�0D;?A;��<;�G6;�r-;W";��;�^;��:�;�:�y�:��Y:�:p
�9p�9      R��z��кʓ����Y���� s89L5:\/�:�d�:rB;am;�?&;D2;�|:;7!@;�C;��E;�G;��G;~(H;![H;�zH;f�H;�H;ɳH;��H;��H;��H;��H;��H;$�H;{�H;Z�H;x�H;(�H;��H;(�H;x�H;Z�H;x�H;'�H;��H;��H;��H;��H;��H;̳H;�H;`�H;�zH;![H;z(H; �G;�G;��E;߳C;7!@;�|:;D2;�?&;`m;pB;�d�:`/�:L5: s89�����Y�ȓ��кz��      ⚩�V���)J���X��2�b��-����Ix����!:��:j��:�;` ;c�.;��8;v�?;�C;��E;[#G;�G;2H;bH;o�H;��H;��H;ӷH;
�H;��H;A�H;`�H;a�H;�H;B�H;��H;d�H;��H;d�H;��H;B�H;�H;d�H;`�H;@�H;��H;
�H;ҷH;��H;��H;l�H;bH;2H;
�G;[#G;��E;�C;v�?;��8;c�.;` ;�;j��:��:!:���Ix������-�,�b��X��)J��Z���      �B(�%�����_������˻	���b�=&����� h>���Y:"�:�^;��;x�,;(`8;u�?;�C;�F;GG;l�G;@H;OkH;'�H;.�H;�H;}�H;��H;��H;��H;D�H;��H;�H;��H;��H;��H;��H;��H;
�H;��H;F�H;��H;��H;��H;~�H;�H;/�H;'�H;KkH;@H;l�G;GG;�F;�C;x�?;&`8;x�,;��;�^;"�:��Y: h>�����<&�
�b�	���˻�����_����%�      �����x���#��GF{���]��E<����U�뻬���;d\�|�뺠[�4:�:���:�[;|�,;��8;7!@;�0D;�[F;B{G;H;iPH;<vH;�H;h�H;$�H;W�H;��H;��H;�H;�H;��H;��H;��H;��H;��H;��H;��H;�H;�H;��H;��H;S�H;&�H;f�H;�H;?vH;hPH;H;C{G;�[F;�0D;7!@;��8;z�,;�[;���:�:4:�[�|��;d\�����V�뻨���E<���]�GF{��#���x��      b������o�vrμփ��yv��N"��^N�����?ݻZ^��B��ЅY���9�:��:��;`�.;�|:;?A;��D;K�F;׶G;*H;@aH;?�H;��H;�H;e�H;F�H;c�H;��H;&�H;F�H;��H;��H;
�H;��H;��H;F�H;$�H;��H;c�H;D�H;`�H;�H;��H;@�H;CaH;*H;жG;M�F;��D;?A;�|:;c�.;��;��:�:��9ЅY�C��Z^���?ݻ���^N�N"��xv��փ��vrμ�o����      dn;�|\8��s/�A�!�~��d���orμ��������E<�"������N3�@Hx� �9�:�^;b ;B2;��<;�B;˲E;V5G;*�G;XFH;�qH;ʎH;r�H;ߴH;v�H;��H;��H;)�H;��H;F�H;��H;6�H;��H;F�H;��H;(�H;��H;��H;v�H;޴H;r�H;ȎH;�qH;YFH;(�G;S5G;˲E;�B;��<;B2;b ;�^;�:��9@Hx��N3����"���E<��������orμd���~��A�!��s/�|\8�      ���������Ȅ�oSt��Y�an;�3O�v#���Oļ�����&R��_������N3�ȅY�4:$�:�;�?&;�G6;�X?;�D;QxF;ۚG;X!H;�^H;��H;�H;��H;i�H;0�H;(�H;��H;<�H;�H;~�H;<�H;~�H;�H;<�H;��H;(�H;0�H;k�H;��H;�H;��H;�^H;[!H;ؚG;MxF;�D;�X?;�G6;�?&;�;"�:4:̅Y��N3������_��&R������Oļv#��3O�an;��Y�oSt��Ȅ�����      �ѽ\ν|�ý䳽>��� M����d�v\8�y��ټnv����Y��_����?���[���Y:l��:`m;�r-;�:;��A;VoE;�"G;s�G;�GH;�sH;�H;��H;�H;V�H;C�H;��H;��H;��H;V�H;�H;V�H;��H;��H;��H;E�H;V�H;�H;��H;�H;�sH;�GH;y�G;�"G;ToE;��A;!�:;�r-;^m;r��:��Y:�[�@������_���Y�nv��ټy��v\8���d� M��>���䳽}�ý\ν      ��"]�ֈ�r}���{�ý�u��͕���K�����o�nv���&R�#��Z^��|�� p>���:nB;X";x�4;��>;fD;��F;�G;�)H;�dH;��H;=�H;��H;W�H;Z�H;��H;��H;N�H;:�H;��H;:�H;N�H;��H;��H;[�H;W�H;��H;:�H;��H;�dH;�)H;�G;��F;cD;��>;z�4;X";nB;
��: x>����Z^��#���&R�nv���o�����K�͕���u��{�ý��r}�ֈ�"]�      �+X��T��nH��6��� �l��G�䳽�����mR����ټ�����E<��?ݻ;d\����� !:�d�:��;6�,;��:;�7B;��E;�LG;`H;~SH;�{H;��H;�H;@�H;k�H;|�H;;�H;��H;�H;��H; �H;��H;:�H;z�H;j�H;@�H;�H;��H;�{H;}SH;aH;�LG;��E;7B;��:;6�,;��;�d�:!:����=d\��?ݻ�E<�����ټ����mR�����䳽G�l���� ��6��nH��T�      㰖��������*|�OS\�� :����Z�o$�������K�y���Oļ����������>&����V/�:�^;��#;�G6;`�?;�D;o�F;��G; @H;�pH;�H;��H;=�H;|�H;X�H;��H;��H;�H;��H;�H;��H;��H;V�H;|�H;=�H;��H;�H;�pH;@H;��G;r�F;�D;_�?;�G6;��#;�^;V/�:���A&������������Oļy���K�����o$���Z���� :�OS\��*|�������      C�;9ɾ~㼾B�������Mw��nH�����Z�䳽͕��v\8�v#������^N�U��
�b�Ix�P5:��:4�;��0;C]=;Q�C;�[F;�G;�)H;fH;��H;D�H;k�H;��H;F�H;��H;\�H;��H;��H;��H;[�H;��H;D�H;��H;j�H;D�H;��H;fH;�)H;
�G;�[F;P�C;D]=;��0;6�;��:P5:Ix��b�U��^N�����v#��v\8�͕��䳽�Z񽳯��nH��Mw�����B��~㼾9ɾ      2y��v�m���E�߾����C��A����nH���Gὠu����d�3O�prμN"�����
	����뺐r89�;�:c�;�+;z|:;�7B;�E;4bG;�H;[H;��H;J�H;ƯH;"�H;s�H;u�H;5�H;�H;��H;�H;5�H;r�H;p�H;$�H;ƯH;I�H;��H;[H;�H;4bG;�E;�7B;y|:;�+;d�;�;�:�r89���
	�����N"��prμ3O���d��u��G����nH�A���C������E�߾m����v�      �O/�rM+�Z�����LW��9ɾB���Mw�� :�l��{�ý M��an;�e���yv���E<��˻��-����y�:�^;�%;��7;��@;85E;�"G;�G;aPH;2{H;��H;��H;��H;��H;$�H;=�H;�H;��H;�H;=�H;$�H;��H;��H;��H;ݗH;.{H;bPH;�G;�"G;:5E;}�@;��7;�%;�^;�y�:����-��˻�E<�yv��e���an;� M��{�ýl��� :��Mw�B��9ɾLW�����Z��rM+�      9�X�YvS�9E��O/��S�LW����������OS\��� ���>����Y�~��փ����]�����0�b���Y���Y:��:s`;b�4;�?;]�D;�F;�G;,FH;|uH;ޓH;��H;��H;?�H;��H;O�H;D�H;%�H;D�H;M�H;��H;<�H;��H;��H;ۓH;yuH;+FH;�G;�F;_�D;�?;d�4;s`;��:��Y:��Y�/�b�������]�փ��~���Y�>����彔� �OS\���������LW���S��O/�9E�YvS�      � ����y�c�h��N��O/����E�߾B���*|��6�s}�䳽oSt�A�!�vrμHF{��_��X��֓���:��:�Z;�2;�O>;�D;f�F;��G;?=H;�pH;��H;u�H;�H;�H;
�H;��H;��H;��H;��H;��H;�H;�H;�H;u�H;��H;�pH;?=H;��G;g�F;�D;�O>;�2;�Z;��:�:֓���X���_�IF{�vrμA�!�oSt�䳽s}��6��*|�B��E�߾����O/��N�c�h���y�      ?v��c���X ��c�h�9E�Z��m���~㼾���nH�ֈ�}�ý�Ȅ��s/��o��#�����,J��0к(
�9@g�:�l;S0;]=;��C;�F;y�G;D6H;ZmH;D�H;ХH;��H;&�H;o�H;��H;1�H;�H;1�H;��H;n�H;#�H;��H;ХH;C�H;WmH;D6H;y�G;�F;��C;]=;V0;�l;@g�:0
�90к,J������#���o��s/��Ȅ�}�ýֈ��nH���~㼾m���Z��9E�c�h�X ��c���      ~h��1���c�����y�YvS�rM+��v�9ɾ�����T�"]�\ν����}\8�����x��%�V���~��0�9X-�:p�;��.;�<;�nC;�dF;�G;�1H;kH;ŌH;ѤH;�H;��H;��H;��H;��H;��H;��H;��H;��H;��H;�H;ѤH;H;kH;�1H;�G;�dF;�nC;�<;��.;p�;X-�:(�9~��V���	%��x�����}\8�����\ν"]��T�����9ɾ�v�rM+�YvS���y�c���1���      gܿ5�ֿ�aǿ@^��1���[o���7����iþ�(���-=��` �A���_�4]�3p����I�X�ѻ��)���R���::�
;�*;�:;ѣB;>IF;-�G;�lH;2�H;��H;k�H;��H;��H;}�H;��H;6�H;��H;6�H;��H;}�H;��H;��H;k�H;��H;/�H;�lH;-�G;@IF;ѣB;�:;�*;:�
;��:��R���)�X�ѻ��I�3p��4]��_�A���` ��-=��(���iþ����7�[o�1���@^���aǿ5�ֿ      5�ֿFpѿ�¿������bXi�ѕ3��
�XD��Hl��D�9��.���R��%\� �hx��4�E��ͻ�$�@  �ˍ�:H�;��*;2�:;�B;UF;��G;QnH;̡H;۷H;��H;��H;��H;��H;��H;J�H;��H;J�H;��H;��H;��H;��H;��H;ٷH;ʡH;QnH;��G;UF;�B;0�:;��*;H�;ˍ�:P  ��$��ͻ5�E�hx�� �%\��R���.��D�9�Hl��XD���
�ѕ3�bXi��������¿Fpѿ      �aǿ�¿����������"Y��f'�����9o���.}��k/����(ڟ�'<Q�1#�ע��(;�2���6�� E7���:��;�,;��;;�C;>wF; �G;�rH;Y�H;��H;@�H;$�H;"�H;��H;��H;w�H;�H;w�H;��H;��H;"�H;&�H;@�H;��H;W�H;�rH; �G;>wF;�C;��;;�,;��;��: F7�6��2����(;�ע�1#�'<Q�(ڟ�����k/��.}�9o�������f'��"Y�����������¿      ?^������m���[o���@�*�&�޾����=ce�2��¯ڽ����g@������R���O*�LG������E^9$��:;�d.;�<;��C;2�F;��G;�yH;ĥH;6�H;M�H;��H;��H;�H;�H;��H;D�H;��H;�H;�H;��H;��H;M�H;5�H;��H;�yH;��G;2�F;��C;��<;�d.;;(��:�E^9���LG���O*��R������g@�����¯ڽ2��=ce�����&�޾*���@�[o�m�������      1����������\o��!J�M�#��\��XD������}PH�����b��"C��� +���ټ,����￐�����:%��:X�;�Y1;>;�0D;��F;sH;m�H;��H;*�H;��H;��H;4�H;��H;z�H;��H;��H;��H;y�H;��H;2�H;��H;��H;'�H;��H;m�H;tH;��F;�0D;>;�Y1;X�;)��:�:������,����ټ� +�"C���b�����}PH�����XD���\��M�#��!J�\o��������      [o�bXi��"Y���@�M�#��
��о�A���i���(����yr���_��5��ɺ�v�`��<��i�d�L�\�̒X:�P�:�`;��4;Ƨ?;��D;�8G;�0H;ËH;��H;��H;2�H;��H;��H;'�H;��H;:�H;��H;:�H;��H;'�H;��H;��H;2�H;��H;��H;ËH;�0H;�8G;��D;ħ?;��4;�`;�P�:ĒX:L�\�h�d��<��v�`��ɺ��5��_�yr�������(��i��A���о�
�M�#���@��"Y�bXi�      ��7�ѕ3��f'�*��\���о�����.}��-=�}
���Ľ^��/:����������7�#GĻƃ$��N�����:�{;�D&;,8;&JA;�E;�G;�LH;�H;��H;T�H;�H;2�H;��H;��H;L�H;��H;D�H;��H;L�H;��H;��H;4�H;�H;S�H;��H;�H;�LH;�G;�E;#JA;,8;�D&;�{;���:�N��Ã$�$GĻ�7���������/:�^����Ľ}
��-=��.}������о�\��*��f'�ѕ3�      ���
�����&�޾XD���A���.}�+�D�jt���ڽ�!��\����`�ļ�
v�@��ƿ���Iɺ`S�9���:'(;�-;��;;��B;�IF;��G;:fH;ƝH;�H;O�H;��H;��H;��H;��H;��H;�H;��H;�H;��H;��H;��H;��H;��H;O�H;�H;ƝH;9fH;��G;�IF;��B;��;;�-;'(;���:`S�9�Iɺǿ��@���
v�`�ļ���\��!����ڽjt�+�D��.}��A��XD��&�޾�����
�      �iþXD��9o�����������i��-=�kt����R��mys�~ +� ��|񗼘(;�.�ѻ�s@���!�H4j:�P�:��;�D3;]�>;-FD;��F;�	H;[|H;��H;��H;Y�H; �H;"�H;��H;I�H;_�H;��H;�H;��H;`�H;I�H;��H;#�H; �H;W�H;��H;��H;X|H;�	H;��F;*FD;\�>;�D3;��;�P�:H4j:��!��s@�.�ѻ�(;�|� ��~ +�mys��R����kt��-=��i���������9o��XD��      �(��Hl���.}�=ce�}PH���(�~
���ڽ�R���{�F�6�� �0p��c�`�Ϩ��,��.IҺ�L^9���:��;�~(;K�8;JA; |E;:jG;�=H;g�H;��H;O�H;��H;U�H;��H;��H;�H;��H; �H;z�H; �H;��H;�H;��H;��H;U�H;��H;M�H;��H;g�H;�=H;7jG;|E; JA;J�8;�~(;��;���:M^90IҺ�,��Ϩ�c�`�0p��� �F�6��{��R����ڽ~
���(�}PH�=ce��.}�Hl��      �-=�D�9��k/�2��������Ľ�!��mys�F�6�(#��ɺ��vz����A^��f�$�P~�p�r:(��: �;�Y1;I=;QxC;GwF;K�G;.fH;m�H;��H;��H;��H;�H;�H;
�H;��H;��H;��H;��H;��H;��H;��H;	�H;�H;�H;��H;��H;��H;j�H;/fH;G�G;CwF;NxC;I=;�Y1;��;(��:|�r:X~�c�$�A^������vz��ɺ�(#�F�6�mys��!����Ľ����2���k/�D�9�      �` ��.�����¯ڽ�b��yr��^��\�~ +�� ��ɺ�B��O*�Fͻ�5R� ǅ��:I��:��;�);u8;��@;�*E;�8G;m$H;q�H;i�H;!�H;V�H;��H;��H;��H;.�H;��H; �H;�H;Q�H;�H;"�H;��H;-�H;��H;��H;��H;S�H;!�H;f�H;q�H;l$H;�8G;�*E;��@;u8;�);��;M��:�: ǅ��5R�Fͻ�O*�B��ɺ�� �~ +�\�^��yr���b��¯ڽ��.��      A���R��(ڟ�����"C���_�/:���� ��/p���vz��O*��4ֻk������09b�:1;m� ;�D3;c�=;̐C;lF;��G;�\H;ƗH;w�H;.�H;o�H;��H;��H;��H;+�H;;�H;��H;��H;��H;��H;��H;;�H;*�H;�H;��H;��H;m�H;.�H;t�H;ǗH;�\H;��G;lF;̐C;c�=;�D3;l� ;1;^�: �09���k��4ֻ�O*��vz�0p�� �輧��/:��_�#C������(ڟ��R��      �_�$\�&<Q�g@�� +��5�����_�ļ{�b�`����Eͻk��Hɺ {6�a�:Q�:=�;�d.;p�:;A�A;O|E;�NG;m'H;.�H;��H;��H;��H;\�H;z�H;��H;d�H;)�H;��H;@�H;��H;0�H;��H;@�H;��H;)�H;e�H;��H;z�H;Z�H;��H;��H;��H;+�H;k'H;�NG;O|E;A�A;o�:;�d.;@�;Q�:a�: x6��Hɺk�Eͻ���b�`�{�_�ļ�����5�� +�g@�%<Q�$\�      3]� �1#�������ټ�ɺ������
v��(;�Ϩ�A^���5R���� |6����:��:�;<�*;�+8;�!@;|�D;��F;#�G;fH;��H;��H;пH;��H;�H;��H;T�H;��H;��H;��H;��H;[�H;��H;[�H;��H;��H;��H;��H;T�H;��H;�H;��H;ϿH;��H;��H;�eH;�G;��F;{�D;�!@;�+8;>�*;�;��:���: |6�����5R�@^��Ϩ��(;��
v������ɺ���ټ����1#� �      1p��gx��ע��R��+��v�`��7�?��,�ѻ�,��c�$� ǅ���09[�:��:�;�~(;�Z6;��>;��C;IF;�G;EH;w�H;�H;۹H;A�H;]�H;G�H;*�H;�H;��H;��H;C�H;�H;��H;��H;��H;�H;C�H;��H;��H;�H;*�H;C�H;]�H;?�H;޹H;�H;s�H;EH;�G;IF;�C;��>;�Z6;�~(;�;��:a�:��09 ǅ�c�$��,��+�ѻ?���7�t�`�+���R��ע�hx��      ��I�1�E��(;��O*����<��GĻƿ���s@�,IҺ@~��:\�:Q�:�;�~(;+�5;�>;\C;`�E;�cG;h$H;(|H;i�H;O�H;��H;��H;n�H;�H;T�H;��H;��H;��H;��H;u�H; �H;&�H; �H;u�H;��H;��H;��H;��H;Q�H;	�H;n�H;��H;��H;O�H;e�H;#|H;h$H;�cG;a�E;\C;�>;+�5;�~(;�;Q�:\�:�:P~�,IҺ�s@�ƿ��GĻ�<�����O*��(;�4�E�      X�ѻ�ͻ.���IG��￐�q�d�ă$��Iɺ��!� M^9|�r:I��:1;;�;>�*;�Z6;�>;Y�B;��E;9G;�	H;.nH;H�H;w�H;ٽH;��H;��H;�H;�H;4�H;��H;��H;4�H;/�H;��H;9�H;\�H;9�H;��H;0�H;2�H;��H;��H;3�H;|�H;�H;��H;��H;ؽH;t�H;E�H;/nH;�	H;9G;��E;Z�B;�>;�Z6;>�*;<�;1;I��:|�r:M^9��!��Iɺ$�m�d�쿐�IG��.����ͻ      y�)��$�)��������8�\��N��XS�9T4j:���:*��:��;m� ;�d.;�+8;��>;\C;��E;�)G;��G;AdH;��H;ȫH;��H;��H;j�H; �H;�H;��H;��H;��H;|�H;��H;��H;4�H;j�H;��H;j�H;4�H;��H;��H;}�H;��H;��H;��H;�H;��H;k�H;��H;��H;īH;��H;?dH;��G;�)G;��E;ZC;��>;�+8;�d.;m� ;��;.��:���:\4j:XS�9�N���\�������)���$�      �R��� ;7��E^9��:ĒX:���:���:�P�:��; �;�);�D3;k�:;�!@;�C;_�E;
9G;��G;�`H;��H;H�H;P�H;��H;s�H;h�H;��H;��H;��H;�H;��H;@�H; �H;��H;d�H;��H;��H;��H;d�H;��H;�H;B�H;��H;�H;��H;��H;��H;j�H;r�H;��H;L�H;H�H;��H;�`H;��G;9G;_�E;�C;�!@;k�:;�D3;�); �;��;�P�:���:���:ؒX: �:�E^9 <7����      ��:���:�: ��:��:�P�:�{;'(;��;�~(;�Y1;u8;e�=;?�A;|�D;IF;�cG;�	H;@dH;��H;z�H;�H;f�H;)�H;�H;t�H;�H;��H;\�H;�H;��H;��H;��H;�H;|�H;��H;��H;��H;|�H;�H;��H;��H;��H;�H;X�H;��H;}�H;t�H;�H;#�H;c�H;�H;v�H;��H;@dH;�	H;�cG;IF;|�D;A�A;e�=;u8;�Y1;�~(;��;)(;�{;�P�:#��:$��:�:Ӎ�:      E�
;h�;�;;\�;a;�D&;�-;�D3;Q�8;!I=;��@;͐C;R|E;��F;�G;i$H;.nH;��H;K�H;�H;��H;n�H;T�H;��H;��H;�H;��H;��H;?�H;X�H;,�H;��H;V�H;��H;��H;��H;��H;��H;V�H;��H;,�H;X�H;;�H;��H;��H;�H;��H;��H;P�H;j�H;��H;
�H;K�H;��H;/nH;h$H;�G;��F;Q|E;͐C;��@; I=;N�8;�D3;�-;�D&;a;p�;;�;d�;      �*;��*;�,;�d.;�Y1;��4;!,8;��;;b�>;JA;RxC;�*E;lF;�NG;#�G;EH;(|H;I�H;ȫH;P�H;f�H;p�H;��H;/�H;.�H;��H;B�H;!�H;��H;�H;��H;��H;�H;r�H;��H;��H;��H;��H;��H;q�H;�H;��H;��H;	�H;��H; �H;?�H;��H;/�H;,�H;��H;n�H;`�H;P�H;ūH;I�H;$|H;EH;#�G;�NG;lF;�*E;SxC;JA;b�>;��;;!,8;��4;�Y1;�d.;�,;}�*;      4�:;H�:;��;;�<;>;ȧ?;3JA;��B;2FD;$|E;JwF;�8G;��G;n'H;fH;v�H;i�H;z�H;��H;��H;%�H;Q�H;.�H;�H;N�H;��H;��H;k�H;��H;��H;O�H;��H;U�H;��H;��H;��H;��H;��H;��H;��H;P�H;��H;O�H;��H;��H;j�H;��H;��H;P�H;�H;,�H;Q�H;!�H;��H;��H;z�H;f�H;t�H;fH;n'H;��G;�8G;HwF;"|E;2FD;��B;0JA;ɧ?;>;�<;��;;8�:;      ߣB;"�B;�C;ƐC;�0D;��D;"�E;�IF;��F;:jG;L�G;q$H;�\H;2�H;��H;�H;W�H;۽H;��H;y�H;�H;��H;3�H;U�H;��H;��H;2�H;y�H;a�H;.�H;��H;
�H;h�H;��H;��H;��H;��H;��H;��H;��H;d�H;
�H;��H;,�H;\�H;w�H;/�H;��H;��H;S�H;2�H;��H;�H;y�H;��H;ܽH;S�H;�H;��H;0�H;�\H;q$H;L�G;:jG;��F;�IF;"�E;��D;�0D;ƐC;�C;"�B;      OIF;1UF;9wF;6�F;��F;�8G;��G;��G;�	H;�=H;/fH;u�H;ǗH;��H;��H;ٹH;��H;��H;g�H;h�H;q�H;��H;��H;��H;��H;/�H;^�H;B�H;��H;~�H;��H;Y�H;n�H;��H;��H;��H;��H;��H;��H;��H;j�H;Y�H;��H;|�H;��H;@�H;[�H;/�H;��H;��H;��H;��H;m�H;g�H;g�H;��H;��H;عH;��H;��H;ǗH;u�H;1fH;�=H;�	H;��G;��G;�8G;��F;6�F;9wF;&UF;      @�G;��G;&�G;��G;H;�0H;�LH;?fH;`|H;j�H;q�H;o�H;w�H;��H;пH;A�H;��H;��H;��H;��H;��H;�H;B�H;��H;,�H;a�H;4�H;��H;��H;��H;�H;g�H;��H;��H;��H;��H;��H;��H;��H;��H;��H;e�H;�H;��H;��H;��H;2�H;^�H;/�H;��H;?�H;�H;}�H;��H;��H;��H;��H;A�H;пH;��H;w�H;o�H;q�H;j�H;b|H;?fH;�LH;�0H;�H;��G;$�G;��G;      �lH;\nH;�rH;�yH;v�H;ˋH;�H;ҝH;ĥH;�H;��H;)�H;4�H;��H;��H;]�H;m�H;�H;�H;��H;��H;��H;!�H;n�H;s�H;C�H;��H;m�H;��H;!�H;B�H;q�H;��H;��H;��H;��H;��H;��H;��H;��H;��H;o�H;@�H;�H;��H;k�H;��H;C�H;u�H;k�H; �H;��H;��H;��H;�H;�H;k�H;]�H;��H;��H;0�H;+�H;��H;�H;ťH;ԝH;�H;ˋH;��H;�yH;�rH;hnH;      L�H;֡H;\�H;̥H;�H;��H;��H;!�H;��H;T�H;��H;]�H;r�H;]�H;�H;H�H;�H;|�H;��H;��H;[�H;��H;��H;��H;Z�H;��H;��H;��H;�H;H�H;e�H;��H;��H;��H;��H;��H;��H;��H;��H;��H;��H;��H;d�H;E�H;�H;��H;��H;��H;\�H;��H;��H;��H;W�H;��H;��H;}�H;�H;G�H;�H;]�H;r�H;\�H;��H;T�H;��H;#�H;��H;��H;�H;ͥH;\�H;ˡH;      ��H;�H;͸H;<�H;>�H;��H;^�H;X�H;e�H;��H;��H;��H;��H;��H;��H;/�H;U�H;2�H;��H;	�H;�H;;�H;�H;��H;%�H;|�H;��H;"�H;G�H;\�H;{�H;y�H;��H;��H;��H;��H;��H;��H;��H;��H;��H;{�H;{�H;Z�H;E�H;!�H;��H;z�H;'�H;��H;�H;;�H;�H;�H;��H;2�H;S�H;/�H;��H;��H;��H;��H;��H;��H;h�H;[�H;^�H;��H;>�H;?�H;̸H;�H;      u�H;��H;R�H;^�H;��H;4�H;�H;�H;-�H;^�H;��H;��H;��H;��H;X�H;�H;��H;��H;��H;��H;��H;W�H;��H;T�H;��H;��H;�H;D�H;c�H;}�H;��H;��H;v�H;y�H;��H;��H;g�H;��H;��H;y�H;t�H;��H;��H;|�H;d�H;D�H;�H;��H;��H;R�H;��H;W�H;��H;��H;��H;��H;��H;�H;X�H;��H;��H;��H;��H;a�H;-�H;�H;�H;6�H;��H;^�H;P�H;��H;      ��H;��H;2�H;��H;��H;��H;;�H;��H;*�H;��H;�H;��H;�H;n�H;��H;��H;��H;��H;��H;I�H;��H;0�H;��H;��H;�H;Y�H;d�H;r�H;��H;{�H;��H;��H;x�H;q�H;��H;h�H;^�H;g�H;��H;q�H;r�H;��H;��H;|�H;��H;r�H;e�H;W�H;
�H;��H;��H;0�H;��H;I�H;��H;��H;��H;��H;��H;m�H;�H;��H;�H;��H;-�H;��H;<�H;��H;��H;��H;2�H;��H;      ��H;��H;1�H;��H;F�H;��H;��H;��H;��H;��H;�H;<�H;2�H;2�H;�H;��H;��H;1�H;��H;%�H;��H;��H;�H;Y�H;a�H;n�H;��H;��H;��H;��H;y�H;y�H;|�H;{�H;Y�H;W�H;��H;W�H;Y�H;{�H;x�H;{�H;y�H;��H;��H;��H;��H;m�H;c�H;Y�H;�H;��H;��H;'�H;��H;2�H;��H;��H;�H;2�H;1�H;;�H;�H;��H;��H;��H;��H;��H;?�H;��H;1�H;��H;      ��H;��H;��H;�H;��H;'�H;��H;��H;S�H;�H;��H;��H;A�H; �H;��H;N�H;��H;0�H;��H;��H;#�H;W�H;q�H;��H;��H;��H;��H;��H;��H;��H;x�H;r�H;u�H;d�H;S�H;Z�H;^�H;Z�H;S�H;d�H;t�H;u�H;x�H;��H;��H;��H;��H;��H;��H;��H;r�H;V�H;"�H;��H;��H;2�H;��H;M�H;��H; �H;A�H;��H;��H;�H;S�H;��H;��H;+�H;��H;�H;��H;��H;      ��H;��H;��H;-�H;��H;��H;Z�H;��H;m�H;��H;��H;1�H;��H;J�H;��H;)�H;�H;��H;7�H;j�H;��H;��H;��H;��H;��H;��H;��H;��H;��H;��H;��H;��H;W�H;U�H;^�H;U�H;7�H;U�H;^�H;U�H;U�H;��H;��H;��H;��H;��H;��H;��H;��H;��H;��H;��H;��H;j�H;6�H;��H;|�H;(�H;��H;I�H;��H;1�H;��H;��H;m�H;��H;Z�H;��H;��H;,�H;��H;��H;      5�H;[�H;��H;��H;��H;:�H;��H;-�H;��H;%�H;��H;!�H;��H;��H;b�H;��H;
�H;6�H;n�H;��H;��H;��H;��H;��H;��H;��H;��H;��H;��H;��H;��H;m�H;W�H;^�H;U�H;P�H;A�H;P�H;U�H;\�H;V�H;o�H;��H;��H;��H;��H;��H;��H;��H;��H;��H;��H;��H;��H;n�H;7�H;	�H;��H;b�H;��H;��H;!�H;��H;&�H;��H;,�H;��H;?�H;��H;��H;��H;T�H;      ��H;�H;�H;K�H;��H;��H;N�H;��H;�H;}�H;��H;_�H;��H;<�H;��H;��H;-�H;W�H;��H;��H;��H;��H;��H;��H;��H;��H;��H;��H;��H;��H;k�H;e�H;��H;a�H;7�H;A�H;;�H;A�H;7�H;a�H;��H;g�H;k�H;��H;��H;��H;��H;��H;��H;��H;��H;��H;��H;��H;��H;Y�H;,�H;��H;��H;<�H;��H;_�H;��H;��H; �H;��H;N�H;��H;��H;K�H;�H;��H;      5�H;[�H;��H;��H;��H;:�H;��H;-�H;��H;#�H;��H;!�H;��H;��H;b�H;��H;
�H;6�H;n�H;��H;��H;��H;��H;��H;��H;��H;��H;��H;��H;��H;��H;m�H;W�H;^�H;U�H;P�H;A�H;P�H;U�H;\�H;V�H;o�H;��H;��H;��H;��H;��H;��H;��H;��H;��H;��H;��H;��H;n�H;7�H;�H;��H;b�H;��H;��H;!�H;��H;&�H;��H;,�H;��H;?�H;��H;��H;��H;S�H;      ��H;��H;��H;-�H;��H;��H;Z�H;��H;k�H;��H;��H;1�H;��H;J�H;��H;(�H;~�H;��H;6�H;k�H;��H;��H;��H;��H;��H;��H;��H;��H;��H;��H;��H;��H;W�H;U�H;^�H;U�H;7�H;U�H;^�H;U�H;U�H;��H;��H;��H;��H;��H;��H;��H;��H;��H;��H;��H;��H;j�H;7�H;��H;~�H;)�H;��H;J�H;��H;1�H;��H;��H;m�H;��H;Z�H;��H;��H;,�H;��H;��H;      ��H;��H;��H;�H;��H;'�H;��H;��H;Q�H;�H;��H;��H;A�H; �H;��H;M�H;��H;0�H;��H;��H;&�H;V�H;q�H;��H;��H;��H;��H;��H;��H;��H;x�H;r�H;u�H;d�H;S�H;Z�H;^�H;Z�H;S�H;d�H;t�H;u�H;x�H;��H;��H;��H;��H;��H;��H;��H;r�H;W�H;"�H;��H;��H;2�H;��H;N�H;��H; �H;A�H;��H;��H;�H;T�H;��H;��H;+�H;��H;�H;��H;��H;      ��H;��H;3�H;��H;D�H;��H;��H;��H;��H;��H;�H;;�H;1�H;2�H;�H;��H;��H;1�H;��H;%�H;��H;��H;�H;Y�H;c�H;n�H;��H;��H;��H;��H;y�H;y�H;{�H;y�H;Y�H;W�H;��H;W�H;Y�H;y�H;x�H;|�H;y�H;��H;��H;��H;��H;m�H;a�H;W�H;�H;��H;��H;%�H;��H;1�H;��H;��H;�H;2�H;1�H;;�H;�H;��H;��H;��H;��H;��H;=�H;��H;0�H;��H;      ��H;��H;5�H;��H;��H;��H;=�H;��H;*�H;��H;�H;��H;�H;m�H;��H;��H;��H;��H;��H;J�H;��H;0�H;��H;��H;
�H;Y�H;e�H;r�H;��H;{�H;��H;��H;u�H;q�H;��H;g�H;^�H;g�H;��H;q�H;t�H;��H;��H;|�H;��H;r�H;e�H;W�H;�H;��H;��H;0�H;��H;I�H;��H;��H;��H;��H;��H;n�H;�H;��H;�H;��H;,�H;��H;<�H;��H;��H;��H;4�H;��H;      u�H;��H;R�H;^�H;��H;4�H;�H;�H;-�H;`�H;��H;��H;��H;��H;X�H;�H;��H;��H;��H;��H;��H;W�H;��H;T�H;��H;��H;�H;D�H;d�H;}�H;��H;��H;u�H;y�H;��H;��H;g�H;��H;��H;y�H;t�H;��H;��H;|�H;d�H;D�H;�H;��H;��H;R�H;��H;W�H;��H;��H;��H;��H;��H;�H;X�H;��H;��H;��H;��H;`�H;-�H;�H;�H;6�H;��H;^�H;R�H;��H;      ��H;�H;͸H;?�H;;�H;��H;_�H;Z�H;h�H;��H;��H;��H;��H;��H;��H;/�H;T�H;/�H;��H;�H;�H;;�H;�H;��H;'�H;{�H;��H;!�H;G�H;\�H;{�H;y�H;��H;��H;��H;��H;��H;��H;��H;��H;��H;{�H;{�H;Z�H;G�H;"�H;��H;{�H;%�H;��H;�H;;�H;�H;	�H;��H;2�H;T�H;0�H;��H;��H;��H;��H;��H;��H;h�H;Z�H;_�H;��H;;�H;<�H;͸H;�H;      C�H;ҡH;b�H;˥H;�H;��H;��H;$�H;��H;T�H;��H;]�H;r�H;]�H;�H;G�H;�H;|�H;��H;��H;\�H;��H;��H;��H;\�H;��H;��H;��H;�H;G�H;d�H;��H;��H;��H;��H;��H;��H;��H;��H;��H;��H;��H;e�H;E�H;�H;��H;��H;��H;Z�H;��H;��H;��H;X�H;��H;��H;}�H;�H;J�H;�H;]�H;r�H;]�H;��H;R�H;��H;#�H;��H;��H;�H;ȥH;`�H;ԡH;      �lH;[nH;�rH;�yH;t�H;ˋH;�H;՝H;ĥH;�H;��H;+�H;0�H;��H;��H;]�H;m�H;�H;�H;��H;��H;��H; �H;m�H;u�H;C�H;��H;k�H;��H;!�H;@�H;o�H;��H;��H;��H;��H;��H;��H;��H;��H;��H;r�H;B�H;�H;��H;m�H;��H;C�H;s�H;m�H;!�H;��H;��H;��H;�H;�H;k�H;^�H;��H;��H;4�H;+�H;��H;�H;ťH;ҝH;�H;ȋH;��H;�yH;�rH;hnH;      :�G;��G;$�G;��G;zH;�0H;�LH;?fH;`|H;k�H;q�H;o�H;w�H;��H;пH;C�H;��H;��H;��H;��H;��H;�H;A�H;��H;/�H;`�H;4�H;��H;��H;��H;�H;e�H;��H;��H;��H;��H;��H;��H;��H;��H;��H;h�H;�H;��H;��H;��H;2�H;a�H;,�H;��H;A�H;�H;}�H;��H;��H;��H;��H;@�H;пH;��H;w�H;o�H;s�H;k�H;`|H;=fH;�LH;�0H;~H;��G;#�G;��G;      VIF;*UF;AwF;7�F;��F;�8G;�G;��G;�	H;�=H;/fH;t�H;ǗH;��H;��H;ٹH;��H;��H;g�H;g�H;r�H;��H;��H;��H;��H;/�H;]�H;@�H;��H;~�H;��H;W�H;k�H;��H;��H;��H;��H;��H;��H;��H;k�H;Z�H;��H;{�H;��H;B�H;]�H;0�H;��H;��H;��H;��H;m�H;g�H;g�H;��H;��H;ٹH;��H;��H;ǗH;u�H;/fH;�=H;�	H;��G;�G;�8G;��F;9�F;CwF;"UF;      ߣB;"�B;�C;ƐC;�0D;��D;"�E;�IF;��F;;jG;N�G;q$H;�\H;0�H;��H;�H;T�H;ٽH;��H;y�H;�H;��H;2�H;U�H;��H;��H;0�H;w�H;a�H;.�H;��H;
�H;e�H;��H;��H;��H;��H;��H;��H;��H;g�H;�H;��H;,�H;^�H;y�H;0�H;��H;��H;T�H;2�H;��H;�H;z�H;��H;޽H;S�H;�H;��H;1�H;�\H;q$H;L�G;8jG;��F;�IF;"�E;��D;�0D;ƐC;�C;"�B;      7�:;E�:;��;;�<;>;ͧ?;-JA;��B;4FD;%|E;KwF;�8G;��G;p'H;fH;t�H;g�H;w�H;��H;��H;%�H;Q�H;.�H;�H;P�H;��H;��H;j�H;��H;��H;O�H;��H;R�H;��H;��H;��H;��H;��H;��H;��H;S�H;��H;O�H;��H;��H;k�H;��H;��H;N�H;�H;,�H;Q�H;"�H;��H;��H;{�H;g�H;v�H;fH;p'H;��G;�8G;HwF;$|E;4FD;��B;/JA;ͧ?;>;�<;��;;7�:;      �*;��*;�,;�d.;�Y1;��4;%,8;��;;b�>;JA;SxC;�*E;lF;�NG;#�G;EH;'|H;F�H;ūH;O�H;f�H;n�H;��H;/�H;/�H;��H;B�H; �H;��H;�H;��H;��H;�H;q�H;��H;��H;��H;��H;��H;r�H;�H;��H;��H;	�H;��H;!�H;?�H;��H;.�H;,�H;��H;p�H;b�H;Q�H;ȫH;I�H;'|H;EH;$�G;�NG;lF;�*E;RxC; JA;b�>;��;;%,8; �4;�Y1;�d.;�,;��*;      E�
;j�;�;;X�;a;�D&;�-;�D3;N�8;!I=;��@;͐C;Q|E;��F;�G;h$H;.nH;��H;J�H;�H;��H;m�H;T�H;��H;��H;�H;��H;��H;?�H;X�H;,�H;��H;V�H;��H;��H;��H;��H;��H;V�H;��H;,�H;X�H;;�H;��H;��H;�H;��H;��H;P�H;k�H;��H;�H;M�H;��H;/nH;h$H;�G;��F;R|E;͐C;��@; I=;Q�8;�D3;�-;�D&;a;n�;;�;b�;      ��:퍨:�:"��:��:�P�:�{;+(;��;�~(;�Y1;u8;e�=;A�A;|�D;IF;�cG;�	H;@dH;��H;y�H;�H;d�H;(�H;�H;t�H;�H;��H;[�H;�H;��H;��H;��H;�H;|�H;��H;��H;��H;|�H;�H;��H;��H;��H;�H;X�H;��H;}�H;t�H;�H;%�H;d�H;�H;w�H;��H;@dH;�	H;�cG;IF;|�D;A�A;e�=;u8;�Y1;�~(;��;*(;�{;�P�:)��:"��:�:Ӎ�:       �R���� 87��E^9 �:̒X:���:���:�P�:��; �;�);�D3;k�:;�!@;�C;_�E;9G;��G;�`H;��H;H�H;O�H;��H;r�H;j�H;��H;��H;��H;�H;��H;@�H; �H;��H;d�H;��H;��H;��H;d�H;��H;�H;B�H;��H;�H;��H;��H;��H;h�H;s�H;��H;M�H;H�H;��H;�`H;��G;9G;_�E;�C;�!@;k�:;�D3;�);��;��;�P�:���:���:ВX:�:�E^9 <7����      y�)��$�)��������0�\��N��XS�9X4j:���:.��:��;m� ;�d.;�+8;��>;\C;��E;�)G;��G;AdH;��H;ȫH;��H;��H;j�H; �H;�H;��H;��H;��H;|�H;��H;��H;4�H;h�H;��H;j�H;4�H;��H;��H;}�H;��H;��H;��H;�H;��H;k�H;��H;��H;īH;��H;?dH;��G;�)G;��E;ZC;��>;�+8;�d.;m� ;��;*��:���:\4j:PS�9�N���\�������)���$�      V�ѻ�ͻ.���IG��𿐻s�d�ă$��Iɺ��!�M^9|�r:I��:1;<�;>�*;�Z6;�>;Y�B;��E;9G;�	H;/nH;H�H;x�H;ؽH;��H;��H;�H;��H;4�H;��H;��H;4�H;0�H;��H;9�H;\�H;9�H;��H;/�H;2�H;��H;��H;3�H;|�H;�H;��H;��H;ٽH;s�H;E�H;.nH;�	H;9G;��E;Y�B;�>;�Z6;>�*;;�;1;I��:|�r: M^9��!��Iɺă$�l�d�쿐�IG��.����ͻ      ��I�1�E��(;��O*����<��GĻſ���s@�,IҺ@~��:\�:Q�:�;�~(;.�5;�>;\C;`�E;�cG;h$H;(|H;i�H;O�H;��H;��H;n�H;�H;S�H;��H;��H;��H;��H;u�H; �H;&�H; �H;u�H;��H;��H;��H;��H;Q�H;�H;n�H;��H;��H;O�H;e�H;#|H;h$H;�cG;a�E;\C;�>;+�5;�~(;�;Q�:\�:�:@~�,IҺ�s@�ƿ��GĻ�<�����O*��(;�3�E�      1p��gx��ע��R��+��u�`��7�@��,�ѻ�,��c�$� ǅ���09]�:��:�;�~(;�Z6;��>;�C;IF;�G;EH;w�H;�H;ܹH;A�H;]�H;G�H;*�H;�H;��H;��H;C�H;�H;��H;��H;��H;�H;C�H;��H;��H;�H;*�H;C�H;]�H;@�H;޹H;�H;t�H;EH;�G;IF;��C;��>;�Z6;�~(;�;��:]�:��09 ǅ�c�$��,��*�ѻ@���7�u�`�+���R��ע�hx��      3]� �1#�������ټ�ɺ������
v��(;�Ϩ�A^���5R���� |6����:��:�;<�*;�+8;�!@;|�D;��F;$�G;fH;��H;��H;ϿH;��H;�H;��H;T�H;��H; �H;��H;��H;[�H;��H;[�H;��H;��H;��H;��H;T�H;��H;�H;��H;ϿH;��H;��H;�eH;�G;��F;{�D;�!@;�+8;>�*;�;��:���: |6�����5R�B^��Ϩ��(;��
v������ɺ���ټ����1#� �      �_�$\�%<Q�g@�� +��5�����_�ļ{�b�`����Fͻk��Hɺ y6�a�:Q�:?�;�d.;l�:;A�A;O|E;�NG;m'H;+�H;��H;��H;��H;\�H;z�H;��H;c�H;+�H;��H;@�H;��H;0�H;��H;@�H;��H;(�H;e�H;��H;z�H;Y�H;��H;��H;��H;.�H;k'H;�NG;O|E;A�A;o�:;�d.;@�;Q�:a�: {6��Hɺk�Eͻ���b�`�{�`�ļ�����5�� +�g@�&<Q�$\�      A���R��(ڟ�����"C���_�/:���� ��0p���vz��O*��4ֻk���� �09b�:1;l� ;�D3;c�=;̐C;lF;��G;�\H;ƗH;w�H;.�H;n�H;��H;��H;��H;*�H;;�H;��H;��H;��H;��H;��H;;�H;*�H;��H;��H;��H;m�H;.�H;t�H;ʗH;�\H;��G;lF;̐C;c�=;�D3;m� ;1;^�:��09���k��4ֻ�O*��vz�/p�� �輧��/:��_�"C������(ڟ��R��      �` ��.�����¯ڽ�b��yr��^��\�~ +�� ��ɺ�B��O*�Fͻ�5R� ǅ��:K��:��;�);u8;��@;�*E;�8G;l$H;q�H;h�H;!�H;U�H;��H;��H;��H;.�H;��H;"�H;�H;Q�H;�H; �H;��H;-�H;��H;��H;��H;U�H;!�H;h�H;q�H;m$H;�8G;�*E;��@;u8;�);��;M��:�:ǅ��5R�Fͻ�O*�B��ɺ�� �~ +�\�^��yr���b��¯ڽ��.��      �-=�D�9��k/�2��������Ľ�!��mys�F�6�(#��ɺ��vz����A^��c�$�P~�x�r:(��: �;�Y1;I=;QxC;GwF;G�G;.fH;l�H;��H;��H;��H;�H;�H;
�H;��H;��H;��H;��H;��H;��H;��H;	�H;�H;�H;��H;��H;��H;l�H;.fH;K�G;DwF;NxC;I=;�Y1;��;(��:|�r:X~�g�$�A^������vz��ɺ�(#�F�6�mys��!����Ľ����2���k/�D�9�      �(��Hl���.}�=ce�}PH���(�~
���ڽ�R���{�F�6�� �0p��c�`�Ϩ��,��.IҺ�L^9���:��;�~(;J�8;JA;!|E;7jG;�=H;g�H;��H;O�H;��H;U�H;��H;��H;�H;��H; �H;z�H; �H;��H;�H;��H;��H;U�H;��H;M�H;��H;f�H;�=H;:jG;|E; JA;K�8;�~(;��;���:M^90IҺ�,��Ϩ�c�`�0p��� �F�6��{��R����ڽ~
���(�}PH�=ce��.}�Hl��      �iþXD��9o�����������i��-=�jt����R��mys�~ +� ��|񗼗(;�.�ѻ�s@���!�H4j:�P�:��;�D3;]�>;-FD;��F;�	H;[|H;��H;��H;W�H; �H;"�H;��H;I�H;`�H;��H;�H;��H;_�H;I�H;��H;"�H; �H;W�H;��H;��H;X|H;�	H;��F;+FD;\�>;�D3;��;�P�:H4j:��!��s@�.�ѻ�(;�|� ��~ +�mys��R����kt��-=��i���������9o��XD��      ���
�����&�޾XD���A���.}�+�D�jt���ڽ�!��\����`�ļ�
v�@��ƿ���Iɺ`S�9���:&(;�-;��;;��B;�IF;��G;:fH;ƝH;�H;O�H;��H;��H;��H;��H;��H;�H;��H;�H;��H;��H;��H;��H;��H;O�H;�H;ƝH;9fH;��G;�IF;��B;��;;�-;)(;���:`S�9�Iɺȿ��@���
v�`�ļ���\��!����ڽjt�+�D��.}��A��XD��&�޾�����
�      ��7�ѕ3��f'�*��\���о�����.}��-=�}
���Ľ^��/:����������7�"GĻă$��N�����:�{;�D&;,8;(JA;�E;�G;�LH;�H;��H;T�H;�H;2�H;��H;��H;L�H;��H;D�H;��H;L�H;��H;��H;2�H;�H;S�H;��H;�H;�LH;�G;�E;%JA;,8;�D&;�{;���:�N��ă$�$GĻ�7���������/:�^����Ľ}
��-=��.}������о�\��*��f'�ѕ3�      [o�bXi��"Y���@�M�#��
��о�A���i���(����yr���_��5��ɺ�v�`��<��h�d�L�\�ĒX:�P�:�`;�4;Ƨ?;��D;�8G;�0H;ËH;��H;��H;2�H;��H;��H;'�H;��H;:�H;��H;<�H;��H;'�H;��H;��H;2�H;��H;��H;ËH;�0H;�8G;��D;ħ?;��4;�`;�P�:ĒX:L�\�h�d��<��v�`��ɺ��5��_�yr�������(��i��A���о�
�M�#���@��"Y�bXi�      1����������\o��!J�M�#��\��XD������}PH�����b��"C��� +���ټ,����￐�����:%��:X�;�Y1;>;�0D;��F;sH;m�H;��H;*�H;��H;��H;4�H;��H;z�H;��H;��H;��H;y�H;��H;2�H;��H;��H;'�H;��H;m�H;tH;��F;�0D;>;�Y1;X�;)��:�:���￐���,����ټ� +�"C���b�����}PH�����XD���\��M�#��!J�\o��������      ?^������m���[o���@�*�&�޾����=ce�2��¯ڽ����g@������R���O*�LG������E^9"��:;�d.;�<;��C;2�F;��G;�yH;ĥH;7�H;M�H;��H;��H;�H;�H;��H;D�H;��H;�H;�H;��H;��H;M�H;5�H;��H;�yH;��G;2�F;��C;��<;�d.;;(��:�E^9���LG���O*��R������g@�����¯ڽ2��=ce�����&�޾*���@�[o�m�������      �aǿ�¿����������"Y��f'�����9o���.}��k/����(ڟ�'<Q�1#�ע��(;�2���6�� F7���:��;�,;��;;�C;>wF; �G;�rH;Y�H;��H;@�H;&�H;#�H;��H;��H;w�H;�H;w�H;��H;��H; �H;$�H;@�H;��H;W�H;�rH; �G;>wF;�C;��;;�,;��;��: F7�7��2����(;�ע�1#�'<Q�(ڟ�����k/��.}�9o�������f'��"Y�����������¿      5�ֿFpѿ�¿������bXi�ѕ3��
�XD��Hl��D�9��.���R��%\� �hx��4�E��ͻ�$�@  �ˍ�:H�;��*;2�:;�B;UF;��G;QnH;̡H;۷H;��H;��H;��H;��H;��H;J�H;��H;J�H;��H;��H;��H;��H;��H;ٷH;ʡH;QnH;��G;UF;�B;0�:;��*;H�;ˍ�:P  ��$��ͻ5�E�hx�� �%\��R���.��D�9�Hl��XD���
�ѕ3�bXi��������¿Fpѿ      ��"$������꿱�ſ�ޞ�(3s��2�A����� j���}Hͽȸ����'�F<ͼt�n�h���@Q^�d-.�h��:zW;�S%;ao8;��A;`DF;�H;��H;��H;��H;Q�H;G�H;S�H;��H;��H;��H;8�H;��H;��H;��H;R�H;H�H;Q�H;��H;��H;��H;�H;`DF;��A;`o8;�S%;zW;l��:l-.�@Q^�g���u�n�F<ͼ��'�ȸ��}Hͽ�� j���A����2�(3s��ޞ���ſ������"$�      "$�������忊�����"cm�X�-�����Sh��Yde�$-�۪ɽ�v��+�$���ɼ|mj�;���X�����ņ:ux;A�%;/�8;mB;mRF;H;0�H;V�H;�H;u�H;K�H;D�H;��H;��H;��H;3�H;��H;��H;��H;B�H;K�H;u�H;�H;T�H;0�H;H;mRF;mB;-�8;G�%;wx;�ņ:���X�:���|mj���ɼ+�$��v��۪ɽ$-�Yde�Sh������X�-�"cm��������忞����      ��������� �ԿNw�����=�\�"����m��\0X�����;����w����������]�#���F�����ɒ:��;9�';��9;!pB;�zF;�!H;��H;:�H;!�H;��H;Q�H;H�H;��H;��H;��H;�H;��H;��H;��H;G�H;Q�H;��H;�H;7�H;��H;�!H;�zF;!pB;��9;<�';��;�ɒ:����F�"�黯�]����������w��;�����\0X�m�����"�=�\����Nw�� �Կ��𿞏�      ����� �Կp���ޞ�bF�j�C�.E�%�;�I���D���!"��k�c���֯���J��ѻɢ)��}K� ��:�
;�M*;s�:;�C;�F;�8H;V�H;��H;x�H;��H;J�H;G�H;��H;��H;��H;
�H;��H;��H;��H;G�H;J�H;��H;w�H;��H;Y�H;�8H;�F;�C;p�:;�M*;�
;$��:�}K�ɢ)��ѻ��J��֯��k�c�!"�����D��I��%�;.E�j�C�bF��ޞ�p�� �Կ��      ��ſ���Nw���ޞ�����A�W�7�%�����jɰ��|x�h{+�ձ� ���J��  �ж��[�1�*���+��"
9 �:��;�-;��<;��C;�G;�TH;P�H; �H;��H;��H;`�H;>�H;��H;��H;��H;��H;��H;��H;��H;=�H;b�H;��H;��H;��H;P�H;�TH;�G;��C;��<;�-;��; �:P"
9+�*���\�1�ж���  ��J� ��ձ�h{+��|x�jɰ�����7�%�A�W������ޞ�Nw�����      �ޞ�������bF�A�W�Y�-����BKɾ�G����O����ƽɸ��҄-���ۼㄼ44�ǐ��ζ��]:��:�;��1;�c>;o�D;�\G;FsH;��H;n�H;i�H;+�H;~�H;6�H;x�H;��H;��H;��H;��H;��H;y�H;6�H;��H;+�H;f�H;j�H;��H;DsH;�\G;m�D;�c>;��1;�;	��:�]:�ζ�ǐ�54�ㄼ��ۼ҄-�ɸ��ƽ�����O��G��BKɾ���Y�-�A�W�bF�������      (3s�!cm�=�\�j�C�7�%�����TҾl�� j��C(����aP����[�~������Y�8��aX�0�<���k:M��:�� ;�5;GR@;fuE;�G;5�H;J�H;��H;�H;N�H;w�H;2�H;q�H;�H;d�H;��H;d�H;�H;q�H;2�H;x�H;N�H;�H;��H;K�H;4�H;�G;cuE;CR@; �5;�� ;Q��:��k:0�<�^X�8����Y����~���[�aP����콭C(� j�l���TҾ���7�%�j�C�=�\�!cm�      �2�W�-�"�.E�����BKɾl����s�;�5���y㻽�v��z0��;��+���*����+6��=S��M�:]�	;��(;�9;�/B;yDF;TH;ԫH;��H;��H;��H;{�H;��H;�H;@�H;N�H;K�H;j�H;K�H;N�H;@�H;�H;��H;{�H;��H;��H;��H;ҫH;TH;vDF;�/B;�9;��(;_�	;�M�:�=S�*6�����*��+���;�z0��v��y㻽��;�5���s�l��BKɾ����.E�"�W�-�      A����������%�;jɰ��G�� j�;�5��	�Ҫɽ[����J�u���沼��]�����	x�<	��`n:ͤ�:�v;��/;�-=;��C;G�F;IH;��H;'�H;��H;'�H;��H;��H;��H;�H;�H;#�H;4�H;#�H;�H;�H;��H;��H;��H;&�H;��H;'�H;��H; IH;D�F;��C;�-=;��/;�v;ˤ�:dn::	���	x������]��沼u���J�[���Ҫɽ�	�;�5� j��G��jɰ�%�;��徹���      ��Sh��m���I���|x���O��C(���Ӫɽ����VDX�K��*<ͼㄼ�X!��s���W��tK�F��:�y;�#;I6;6R@;�PE;��G;��H;��H;6�H;��H;��H;��H;��H;��H;��H;��H;��H;��H;��H;��H;��H;��H;��H;��H;��H;��H;5�H;��H;��H;��G;�PE;5R@;I6;�#;�y;F��:�tK��W��s���X!�ㄼ*<ͼK��VDX�����Ӫɽ���C(���O��|x��I��m��Sh��       j�Yde�\0X��D�h{+�������y㻽\���VDX������ۼ;����;�E>ۻX��y�(?":޽�:��;ڷ-;��;;��B;�zF;�H;��H;�H;)�H;��H;��H;��H;{�H;��H;��H;��H;��H;��H;��H;��H;��H;��H;~�H;��H;��H;��H;(�H;~�H;��H;�H;�zF;��B;��;;ٷ-;��;޽�:8?":�y�X�E>ۻ��;�;����ۼ���VDX�[���y㻽��콄��h{+��D�\0X�Yde�      ��$-������ձ�ƽaP���v���J�J����ۼ��d�J������+��rrѺ�)
9�M�:��;� $;�5;�?;��D;d\G;fH;��H;��H;��H;��H;(�H;��H;c�H;�H;m�H;f�H;r�H;K�H;t�H;i�H;n�H;�H;d�H;��H;(�H;��H;��H;��H;��H;fH;b\G;��D;��?;�5;� $;��;�M�:p)
9prѺ�+������d�J�����ۼJ���J��v��aP��ƽձ轅����$-�      }Hͽ۪ɽ�;�� "�� ��ɸ����[�z0�u��*<ͼ;��e�J�����j��m*�����:[b�:V�;��/;�L<;C;1mF;��G;�H;�H;�H;�H;P�H;a�H;��H;7�H;C�H;/�H;)�H;�H;�H;�H;)�H;/�H;C�H;7�H;��H;a�H;M�H;�H;�H;�H;�H;��G;-mF;C;�L<;��/;V�;ab�:��:��m*��j�����d�J�;��*<ͼu��z0���[�ɸ�� �� "���;��۪ɽ      ȸ���v����w�j�c��J�ф-�~��;缈沼
ㄼ��;������j���5���H?Q:s��:gi;�M*;��8;��@;�PE;�uG;EiH;��H;��H;�H;0�H;��H;��H;��H;	�H;��H;��H;��H;��H;��H;��H;��H;��H;��H;�H;��H;��H;��H;/�H;�H;��H;��H;BiH;�uG;�PE;��@;��8;�M*;ji;o��:H?Q:п깙5��j��������;�
ㄼ�沼�;�~�ф-��J�j�c���w��v��      ��'�*�$����~��  ���ۼ����+����]��X!�F>ۻ�+��p*����>:���:�;:�%;�5;��>;�(D;�F;�!H;?�H;_�H;��H;��H;��H;��H;~�H;��H;��H;��H;��H;~�H;c�H;��H;e�H;��H;��H;��H;��H;��H;{�H;��H;��H;��H; �H;]�H;9�H;�!H;�F;�(D;��>;�5;>�%;�;���:�>:��p*��+��D>ۻ�X!���]��+�������ۼ�  �~����+�$�      E<ͼ��ɼ�����֯�϶��ㄼ��Y��*�����s��X�prѺ��H?Q:���:��
;V�#;j�3;�c=;$C;/DF;�G;�H;��H;�H;H�H;	�H;i�H;6�H;z�H;��H;w�H;M�H;f�H;!�H; �H;�H; �H;!�H;f�H;L�H;x�H;��H;x�H;2�H;i�H;�H;I�H;�H;��H;�H;�G;,DF;$C;�c=;l�3;T�#;��
;���:L?Q:��prѺX��s������*���Y�ㄼж���֯�������ɼ      s�n�xmj���]���J�[�1�34�2������	x��W��y��)
9��:m��:�;Q�#;`�2;�<;upB;3�E;��G;�eH;�H;C�H;��H;�H;��H;��H;Q�H;_�H;N�H;&�H;�H;��H;��H;��H;��H;��H;��H;��H;�H;'�H;N�H;\�H;M�H;��H;��H;	�H;��H;@�H;��H;�eH;��G;4�E;wpB;�<;`�2;Q�#;�;m��:��:�)
9�y��W��	x����3��34�[�1���J���]�zmj�      h���8������ѻ*���ǐ�\X�+6�4	���tK�8?":�M�:Yb�:fi;<�%;g�3;�<;M0B;��E;�\G;�HH;U�H;��H;m�H;�H;I�H;Q�H;��H;.�H;1�H;��H;��H;��H;w�H;k�H;i�H;H�H;i�H;k�H;y�H;��H;��H;��H;/�H;*�H;��H;P�H;K�H;�H;j�H;��H;U�H;�HH;�\G;��E;P0B;�<;i�3;<�%;ii;_b�:�M�:8?":�tK�4	��+6�\X�ǐ�&����ѻ��<���      4Q^�X��F�¢)�+��ζ��<� >S�tn:F��:��:��;V�;�M*;��5;�c=;wpB;��E;�JG;b8H;{�H;��H;%�H;?�H;��H;��H;��H;��H;�H;��H;��H;��H;o�H;�H;�H;�H;��H;�H;�H;�H;n�H;��H;��H;��H;��H;��H;��H;��H;��H;:�H;�H;��H;x�H;c8H;�JG;��E;tpB;�c=;��5;�M*;V�;��;��:F��:|n:�=S��<��ζ�+�¢)��F�X�      D-.�D��x��`}K��"
9�]:��k:�M�:ˤ�:�y;��;� $;��/;��8;��>;$C;3�E;�\G;_8H;֥H;�H;4�H;��H;K�H;��H;i�H;��H;��H;��H;��H;V�H;,�H;��H;��H;��H;��H;��H;��H;��H;��H;��H;-�H;V�H;��H;��H;��H;��H;k�H;��H;D�H;��H;3�H;�H;֥H;_8H;�\G;2�E;$C;��>;��8;��/;� $;��;�y;ˤ�:�M�:��k:�]:P#
9`}K�x��X��      ���:Ɔ:�ɒ:��:��:��:W��:]�	;�v;�#;ڷ-;�5;�L<;��@;�(D;-DF;��G;�HH;|�H;�H;��H;a�H;��H;u�H;8�H;��H;��H;��H;z�H;<�H; �H;��H;��H;|�H;N�H;>�H;A�H;@�H;O�H;}�H;��H;��H; �H;:�H;w�H;��H;��H;��H;8�H;q�H;��H;a�H;��H;�H;{�H;�HH;��G;-DF;�(D;��@;�L<;�5;ٷ-;�#;�v;_�	;S��:��:��: ��: ʒ:�ņ:      �W;�x;�;�
;��;�;� ;��(;��/;I6;��;;�?;C;�PE;�F;�G;�eH;U�H;��H;6�H;`�H;��H;H�H;�H;}�H;��H;��H;��H;�H;��H;��H;c�H;;�H;*�H;��H;��H;��H;��H;��H;*�H;9�H;c�H;��H;��H;�H;��H;��H;��H;~�H;�H;E�H;��H;^�H;6�H;��H;U�H;�eH;�G;�F;�PE;C;�?;��;;I6;��/;��(;� ;�;ȅ;�
;�;�x;      �S%;H�%;=�';�M*;�-;��1;�5;�9;�-=;:R@;��B;��D;2mF;�uG;�!H;�H;�H;��H;#�H;��H;��H;I�H;�H;}�H;��H;��H;V�H;�H;��H;��H;D�H;�H;��H;��H;��H;��H;u�H;��H;��H;��H;��H;�H;B�H;��H;��H;�H;Q�H;��H;��H;z�H;�H;I�H;��H;��H;"�H;��H;�H;�H;�!H;�uG;2mF;��D;��B;9R@;�-=;�9;�5;��1;�-;�M*;=�';;�%;      |o8;C�8;ˏ9;v�:;��<;�c>;RR@;�/B;��C;�PE;�zF;i\G;��G;FiH;=�H;��H;F�H;p�H;>�H;H�H;q�H;�H;}�H;��H;��H;h�H;�H;��H;��H;3�H;��H;��H;��H;Q�H;K�H;@�H;�H;@�H;N�H;Q�H;�H;��H;��H;/�H;��H;��H;�H;h�H;��H;��H;|�H;�H;n�H;H�H;<�H;q�H;B�H;��H;=�H;FiH;��G;h\G;�zF;�PE;��C;�/B;QR@;�c>;��<;v�:;ˏ9;4�8;      ��A;~B;pB;�C;��C;v�D;huE;|DF;J�F;��G;�H;fH;�H;��H;c�H;!�H;��H;�H;��H;��H;;�H;��H;��H;��H;I�H;��H;��H;��H;)�H;��H;��H;g�H;6�H;�H;��H;��H;��H;��H;��H;�H;3�H;g�H;��H;��H;&�H;��H;��H;��H;I�H;��H;��H;��H;8�H;��H;��H;�H;��H; �H;c�H;��H;�H;fH;�H;��G;J�F;zDF;huE;v�D;��C;�C;pB;|B;      nDF;�RF;�zF;�F;�G;�\G;
�G;VH;#IH;��H;��H;��H;�H;��H;��H;F�H;	�H;I�H;��H;h�H;��H;��H;��H;h�H;��H;��H;��H;"�H;��H;��H;D�H;�H;��H;��H;��H;��H;��H;��H;��H;��H;��H;�H;A�H;��H;��H;"�H;��H;��H;��H;d�H;��H;��H;��H;h�H;��H;K�H;�H;F�H;��H;��H;�H;��H;��H;��H;#IH;VH;
�G;�\G;�G;�F;�zF;tRF;      �H;H;�!H;�8H;�TH;NsH;B�H;ثH;��H;��H;��H;��H;�H;�H;��H;	�H;��H;O�H;��H;��H;��H;��H;T�H;
�H;��H;��H;�H;��H;q�H;A�H;��H;��H;��H;s�H;W�H;4�H;G�H;4�H;U�H;q�H;��H;��H;��H;?�H;p�H;��H;�H;��H;��H;�H;S�H;��H;��H;��H;��H;P�H;��H;�H;��H;�H;�H;��H;��H;��H;��H;ثH;@�H;JsH;�TH;�8H;�!H;H;      ��H;;�H;��H;Y�H;X�H;��H;T�H;��H;0�H;=�H;3�H;��H;�H;6�H;��H;k�H;��H;��H;��H;��H;��H;��H;�H;��H;��H;"�H;��H;��H;2�H;��H;��H;t�H;N�H;�H;�H; �H; �H; �H;�H;�H;L�H;t�H;��H;��H;/�H;��H;��H;"�H;��H;��H;�H;��H;��H;��H;��H;��H;��H;i�H;��H;4�H;�H;��H;2�H;=�H;1�H;��H;T�H;��H;c�H;Y�H;��H;F�H;      �H;_�H;<�H;��H;�H;s�H;��H;��H;��H;��H;��H;��H;S�H;��H;��H;8�H;T�H;+�H;�H;��H;}�H;�H;��H;��H;"�H;��H;p�H;3�H;��H;��H;h�H;/�H;��H;��H;��H;��H;��H;��H;��H;��H;��H;1�H;f�H;��H;��H;3�H;n�H;��H;%�H;��H;��H;�H;y�H;��H;�H;+�H;Q�H;6�H;��H;��H;S�H;��H;��H;��H;��H;��H;��H;q�H;�H;��H;<�H;U�H;      	�H;�H;1�H;~�H;�H;q�H;�H;��H;5�H;��H;�H;9�H;i�H;��H;��H;}�H;b�H;-�H;��H;��H;;�H;��H;��H;4�H;��H;��H;=�H;��H;��H;^�H;.�H;��H;��H;��H;��H;}�H;r�H;}�H;��H;��H;��H;��H;.�H;\�H;��H;��H;=�H;��H;��H;2�H;��H;��H;8�H;��H;��H;-�H;a�H;}�H;��H;��H;i�H;9�H;	�H;��H;7�H;��H;�H;r�H;�H;�H;-�H;�H;      Z�H;��H;��H;��H;�H;.�H;\�H;��H;��H;��H;�H;�H;�H;�H;��H;��H;U�H;��H;��H;Z�H;%�H;��H;B�H;��H;��H;D�H;��H;��H;e�H;/�H;��H;��H;��H;r�H;P�H;Z�H;X�H;[�H;Q�H;s�H;��H;��H;��H;.�H;f�H;��H;��H;D�H;��H;��H;@�H;��H;"�H;Z�H;��H;��H;T�H;��H;��H;��H;�H;�H;�H;��H;��H;��H;\�H;/�H; �H;��H;��H;��H;      Y�H;`�H;\�H;Y�H;m�H;��H;��H;��H;��H;��H;��H;q�H;=�H;�H;��H;��H;/�H;��H;��H;4�H;��H;g�H;�H;��H;d�H;�H;��H;v�H;/�H;��H;��H;��H;u�H;B�H;-�H;*�H;.�H;*�H;-�H;B�H;p�H;��H;��H;��H;/�H;v�H;��H;�H;g�H;��H;�H;g�H;��H;4�H;��H;��H;.�H;��H;��H;�H;=�H;p�H;��H;��H;��H;��H;��H;��H;j�H;V�H;\�H;\�H;      Z�H;Y�H;V�H;Y�H;R�H;:�H;9�H;,�H;�H;��H;��H;��H;J�H;��H;��H;T�H;�H;��H;u�H;�H;��H;;�H;��H;��H;/�H;��H;��H;S�H;��H;��H;��H;v�H;0�H;%�H;%�H;��H;��H;��H;%�H;%�H;-�H;w�H;��H;��H;��H;Q�H;��H;��H;0�H;��H;��H;;�H;��H;�H;s�H;��H;�H;T�H;��H;��H;J�H;��H;��H;��H;�H;*�H;:�H;=�H;K�H;Y�H;V�H;S�H;      ��H;��H;��H;��H;��H;y�H;y�H;O�H;�H;��H;��H;z�H;5�H;��H;��H;p�H;��H;z�H; �H;��H;��H;*�H;��H;U�H;�H;��H;o�H;�H;��H;��H;s�H;B�H; �H;�H; �H;��H;��H;��H; �H;�H;�H;F�H;s�H;��H;��H;�H;m�H;��H;�H;T�H;��H;*�H;��H;��H; �H;|�H;��H;q�H;��H;��H;5�H;x�H;��H; �H;�H;P�H;y�H;}�H;��H;��H;��H;��H;      �H;�H;��H;��H;��H;��H;��H;`�H;)�H;��H;��H;z�H;5�H;��H;��H;-�H;��H;k�H;�H;��H;V�H;��H;��H;O�H;��H;��H;U�H;�H;��H;��H;Q�H;0�H;#�H;�H;��H;��H;��H;��H;��H;�H; �H;3�H;Q�H;��H;��H;�H;T�H;��H;��H;N�H;��H;��H;R�H;��H;�H;l�H;��H;-�H;��H;��H;5�H;x�H;��H;��H;)�H;^�H;��H;��H;��H;��H;��H;�H;      ��H;��H;��H;��H;��H;��H;r�H;Z�H;3�H;��H;��H;��H;!�H;��H;j�H;	�H;��H;h�H;�H;��H;G�H;��H;��H;D�H;��H;��H;2�H;�H;��H;~�H;]�H;.�H;��H;��H;��H;��H;��H;��H;��H;��H;��H;1�H;]�H;��H;��H;�H;2�H;��H;��H;C�H;��H;��H;E�H;��H;�H;i�H;��H;	�H;j�H;��H;!�H;��H;��H;��H;4�H;Y�H;r�H;��H;��H;��H;��H;��H;      >�H;C�H;7�H;�H;�H;��H;��H;v�H;@�H;��H;��H;Y�H;	�H;��H;��H;(�H;��H;B�H;��H;��H;B�H;��H;r�H;�H;��H;��H;D�H;�H;��H;v�H;]�H;4�H;��H;��H;��H;��H;��H;��H;��H;��H;��H;5�H;]�H;w�H;��H;�H;D�H;��H;��H;�H;r�H;��H;A�H;��H;��H;C�H;��H;(�H;��H;��H;	�H;Y�H;��H;��H;A�H;u�H;��H;��H;�H;�H;5�H;<�H;      ��H;��H;��H;��H;��H;��H;r�H;Z�H;3�H;��H;��H;��H;!�H;��H;l�H;	�H;��H;h�H;�H;��H;H�H;��H;��H;D�H;��H;��H;4�H;�H;��H;~�H;]�H;.�H;��H;��H;��H;��H;��H;��H;��H;��H;��H;1�H;]�H;��H;��H;�H;2�H;��H;��H;A�H;��H;��H;E�H;��H;�H;i�H;��H;	�H;j�H;��H;!�H;��H;��H;��H;3�H;Y�H;r�H;��H;��H;��H;��H;��H;       �H;�H;��H;��H;��H;��H;��H;`�H;)�H;��H;��H;x�H;5�H;��H;��H;-�H;��H;k�H;�H;��H;W�H;��H;��H;O�H;��H;��H;U�H;�H;��H;��H;Q�H;0�H;#�H;�H;��H;��H;��H;��H;��H;�H; �H;4�H;Q�H;��H;��H;�H;T�H;��H;��H;M�H;��H;��H;R�H;��H;�H;l�H;��H;-�H;��H;��H;5�H;z�H;��H;��H;)�H;^�H;��H;��H;��H;��H;��H;�H;      ��H;��H;��H;��H;��H;y�H;y�H;O�H;�H; �H;��H;x�H;5�H;��H;��H;q�H;��H;z�H; �H;��H;��H;*�H;��H;U�H;�H;��H;m�H;�H;��H;��H;s�H;C�H; �H;�H; �H;��H;��H;��H; �H;�H;�H;F�H;s�H;��H;��H;�H;o�H;��H;�H;T�H;��H;*�H;��H;��H; �H;|�H;��H;p�H;��H;��H;5�H;z�H;��H;��H;�H;O�H;y�H;}�H;��H;��H;��H;��H;      ^�H;Z�H;W�H;Z�H;O�H;9�H;9�H;)�H;�H;��H;��H;��H;J�H;��H;��H;T�H;�H;��H;s�H;�H;��H;;�H;��H;��H;0�H;��H;��H;Q�H;��H;��H;��H;v�H;.�H;#�H;%�H;��H;��H;��H;%�H;#�H;-�H;y�H;��H;��H;��H;S�H;��H;��H;/�H;��H;��H;;�H;��H;�H;u�H;��H;�H;T�H;��H;��H;H�H;��H;��H;��H;�H;)�H;7�H;;�H;H�H;Y�H;U�H;Y�H;      Y�H;`�H;_�H;V�H;j�H;��H;��H;��H;��H;��H;��H;q�H;=�H;�H;��H;��H;/�H;��H;��H;5�H;��H;g�H;�H;��H;g�H;�H;��H;v�H;.�H;��H;��H;��H;s�H;B�H;-�H;*�H;.�H;*�H;-�H;B�H;p�H;��H;��H;��H;1�H;v�H;��H;�H;d�H;��H;�H;g�H;��H;4�H;��H;��H;.�H;��H;��H;�H;=�H;p�H;��H;��H;��H;��H;��H;��H;i�H;V�H;_�H;]�H;      Z�H;��H;��H;��H;�H;/�H;\�H;��H;��H;��H;�H;�H;�H;�H;��H;��H;T�H;��H;��H;Z�H;&�H;��H;B�H;��H;��H;F�H;��H;��H;e�H;/�H;��H;��H;��H;s�H;Q�H;[�H;X�H;Z�H;P�H;r�H;��H;��H;��H;.�H;f�H;��H;��H;C�H;��H;��H;@�H;��H;"�H;Z�H;��H;��H;T�H;��H;��H;�H;�H;�H;��H;��H;��H;��H;\�H;/�H; �H;��H;��H;��H;      �H;�H;.�H;��H;�H;p�H;�H;��H;7�H;��H;	�H;9�H;i�H;��H;��H;}�H;b�H;+�H;��H;��H;>�H;��H;��H;4�H;��H;��H;=�H;��H;��H;^�H;.�H;��H;��H;��H;��H;}�H;r�H;}�H;��H;��H;��H;��H;.�H;\�H;��H;��H;<�H;��H;��H;3�H;��H;��H;:�H;��H;��H;.�H;a�H;~�H;��H;��H;i�H;9�H;�H;��H;7�H;��H;�H;q�H;�H;�H;/�H;�H;      �H;[�H;A�H;��H;
�H;n�H;��H;��H;��H;��H;��H;��H;S�H;��H;��H;6�H;S�H;*�H;�H;��H;~�H;�H;��H;��H;%�H;��H;m�H;3�H;��H;��H;f�H;.�H;��H;��H;��H;��H;��H;��H;��H;��H;��H;1�H;h�H;��H;��H;3�H;q�H;��H;"�H;��H;��H;�H;z�H;��H;�H;-�H;S�H;9�H;��H;��H;S�H;��H;��H;��H;��H;��H;��H;p�H;�H;��H;A�H;[�H;      ��H;:�H;��H;Y�H;W�H;��H;T�H;��H;0�H;=�H;3�H;��H;�H;6�H;��H;i�H;��H;��H;��H;��H;��H;��H;�H;��H;��H;"�H;��H;��H;2�H;��H;��H;t�H;M�H;�H;	�H;��H; �H; �H;	�H;�H;M�H;v�H;��H;��H;0�H;��H;��H;"�H;��H;��H;�H;��H;��H;��H;��H;��H;��H;l�H;��H;4�H;�H;��H;2�H;=�H;1�H;��H;T�H;��H;`�H;Y�H;��H;F�H;      �H;H;�!H;�8H;�TH;JsH;?�H;׫H;��H;��H;��H;��H;�H;�H;��H;	�H;��H;O�H;��H;��H;��H;��H;S�H;�H;��H;��H;�H;��H;q�H;@�H;��H;��H;��H;q�H;U�H;4�H;G�H;2�H;W�H;q�H;��H;��H;��H;@�H;p�H;��H;�H;��H;��H;�H;T�H;��H;��H;��H;��H;P�H;��H;�H;��H;�H;�H;��H;��H;��H;��H;ثH;?�H;HsH;�TH;�8H;�!H;H;      uDF;{RF;�zF;�F;�G;�\G;�G;VH;"IH;��H;��H;��H;�H;��H;��H;H�H;�H;I�H;��H;h�H;��H;��H;��H;g�H;��H;��H;��H;"�H;��H;��H;A�H;�H;��H;��H;��H;��H;��H;��H;��H;��H;��H;�H;D�H;��H;��H;"�H;��H;��H;��H;e�H;��H;��H;��H;h�H;��H;K�H;�H;F�H;��H;��H;�H;��H;��H;��H;"IH;TH;�G;�\G;�G;�F;�zF;pRF;      ��A;~B;pB;�C;��C;v�D;huE;zDF;J�F;��G;�H;fH;�H;��H;c�H;!�H;��H;�H;��H;��H;<�H;��H;��H;��H;I�H;��H;��H;��H;)�H;��H;��H;f�H;5�H;�H;��H;��H;��H;��H;��H;�H;5�H;j�H;��H;��H;&�H;��H;��H;��H;I�H;��H;��H;��H;8�H;��H;��H;�H;��H;!�H;c�H;��H;�H;fH;�H;��G;J�F;zDF;huE;v�D;��C;�C;pB;~B;      o8;B�8;ҏ9;s�:;��<;�c>;NR@;�/B;��C;�PE;�zF;i\G;��G;FiH;=�H;��H;D�H;o�H;<�H;H�H;r�H;�H;|�H;��H;��H;g�H;�H;��H;��H;3�H;��H;��H;��H;O�H;J�H;@�H;�H;@�H;M�H;Q�H;��H;��H;��H;0�H;��H;��H;�H;i�H;��H;��H;|�H;�H;n�H;H�H;>�H;q�H;C�H;��H;=�H;FiH;��G;i\G;�zF;�PE;��C;�/B;NR@;�c>;��<;r�:;ԏ9;4�8;      �S%;V�%;K�';�M*;�-;��1;�5;�9;�-=;:R@;��B;��D;1mF;�uG;�!H;�H;�H;��H;"�H;��H;��H;I�H;�H;~�H;��H;��H;T�H;�H;��H;��H;B�H;�H;��H;��H;��H;��H;u�H;��H;��H;��H;��H;�H;D�H;��H;��H;�H;T�H;��H;��H;z�H;�H;I�H;��H;��H;#�H;��H;�H;�H;�!H;�uG;1mF;��D;��B;7R@;�-=;�9;�5;��1;�-;�M*;C�';E�%;      �W;�x;�;�
;��;�;� ;��(;��/;I6;��;;�?;C;�PE;�F;�G;�eH;S�H;��H;4�H;a�H;��H;H�H;�H;~�H;��H;��H;��H;�H;��H;��H;c�H;:�H;*�H;��H;��H;��H;��H;��H;*�H;:�H;c�H;��H;��H;�H;��H;��H;��H;}�H;
�H;E�H;��H;^�H;7�H;��H;V�H;�eH;�G;�F;�PE;C;�?;��;;I6;��/;��(;� ;�;ƅ;�
;�;�x;      t��:Ɔ:ʒ:��:��:��:Y��:b�	;�v;�#;ڷ-;�5;�L<;��@;�(D;-DF;��G;�HH;{�H;�H;��H;a�H;��H;u�H;8�H;��H;��H;��H;|�H;<�H; �H;��H;��H;|�H;O�H;>�H;A�H;>�H;N�H;|�H;��H;��H; �H;:�H;w�H;��H;��H;��H;8�H;q�H;��H;a�H;��H;�H;|�H;�HH;��G;-DF;�(D;��@;�L<;�5;ڷ-;�#;�v;`�	;[��:��:��:��:ʒ:�ņ:      P-.�4��h��`}K��"
9�]:��k:�M�:ˤ�:�y;��;� $;��/;��8;��>;$C;3�E;�\G;_8H;ԥH;�H;3�H;��H;H�H;��H;k�H;��H;��H;��H;��H;V�H;-�H;��H;��H;��H;��H;��H;��H;��H;��H;��H;-�H;V�H;��H;��H;��H;��H;k�H;��H;F�H;��H;4�H;�H;ץH;_8H;�\G;2�E;$C;��>;��8;��/;� $;��;�y;ͤ�:�M�:��k:�]: #
9p}K�x��`��      4Q^�X��F�¢)�+��ζ��<� >S�tn:F��:��:��;V�;�M*;��5;�c=;upB;��E;�JG;b8H;|�H;��H;#�H;>�H;��H;��H;��H;��H;�H;��H;��H;��H;p�H;�H;�H;�H;��H;�H;�H;�H;n�H;��H;��H;��H; �H;��H;��H;��H;��H;;�H; �H;��H;x�H;c8H;�JG;��E;upB;�c=;��5;�M*;V�;��;��:F��:|n: >S��<��ζ�+�¢)��F�X�      f���8������ѻ*���ǐ�\X�.6�4	���tK�8?":�M�:[b�:gi;<�%;i�3;�<;M0B;��E;�\G;�HH;U�H;��H;o�H;�H;I�H;Q�H;��H;.�H;1�H;��H;��H;��H;y�H;k�H;i�H;H�H;i�H;k�H;w�H;��H;��H;��H;/�H;+�H;��H;O�H;L�H;�H;i�H;��H;U�H;�HH;�\G;��E;N0B;�<;g�3;<�%;gi;[b�:�M�:8?":�tK�4	��16�^X�ǐ�'����ѻ��<���      s�n�xmj���]���J�[�1�44�4������	x��W��y��)
9��:m��:�;Q�#;`�2;�<;wpB;3�E;��G;�eH;�H;D�H;��H;�H;��H;��H;P�H;_�H;N�H;'�H;�H;��H;��H;��H;��H;��H;��H;��H;�H;'�H;N�H;^�H;M�H;��H;��H;	�H;��H;?�H;��H;�eH;��G;4�E;upB;�<;`�2;Q�#;�;m��:��:�)
9�y��W��	x����4��34�[�1���J���]�zmj�      E<ͼ��ɼ�����֯�϶��ㄼ��Y��*�����s��X�prѺ��H?Q:���:��
;V�#;j�3;�c=;$C;/DF;�G;�H;��H;�H;H�H;�H;i�H;8�H;x�H;��H;x�H;M�H;f�H;!�H; �H;�H; �H;!�H;f�H;L�H;x�H;��H;z�H;2�H;i�H;�H;J�H;�H;��H;�H;�G;,DF;$C;�c=;l�3;T�#;��
;���:H?Q:��prѺX��s������*���Y�ㄼ϶���֯�������ɼ      ��'�*�$����~��  ���ۼ����+����]��X!�D>ۻ�+��p*����>:���:�;;�%;�5;��>;�(D;�F;�!H;=�H;]�H; �H;��H;��H;��H;}�H;��H;��H;��H;��H;�H;c�H;��H;c�H;~�H;��H;��H;��H;��H;{�H;��H;��H;��H; �H;_�H;;�H;�!H;�F;�(D;��>;�5;<�%;�;���:�>:��p*��+��F>ۻ�X!���]��+�������ۼ�  �~����+�$�      ȸ���v����w�j�c��J�ф-�~��;缈沼
ㄼ��;������j���5�п�H?Q:s��:ii;�M*;��8;��@;�PE;�uG;EiH;��H;��H;�H;/�H;��H;��H;��H;	�H;��H;��H;��H;��H;��H;��H;��H;��H;��H;�H;��H;��H;��H;0�H;�H;��H;��H;BiH;�uG;�PE;��@;��8;�M*;ji;o��:H?Q:�깚5��j��������;�
ㄼ�沼�;�~�ф-��J�j�c���w��v��      }Hͽ۪ɽ�;�� "�� ��ɸ����[�z0�u��*<ͼ;��d�J�����j��m*�����:_b�:V�;��/;�L<;C;1mF;��G;�H;�H;�H;�H;P�H;a�H;��H;6�H;C�H;/�H;)�H;�H;�H;�H;)�H;/�H;A�H;7�H;��H;a�H;M�H;�H;�H;�H;�H;��G;-mF;C;�L<;��/;V�;ab�:��:��m*��j�����e�J�;��*<ͼu��z0���[�ɸ�� �� "���;��۪ɽ      ��$-������ձ�ƽaP���v���J�J����ۼ��d�J������+��prѺ�)
9�M�:��;� $;	�5;��?;��D;d\G;fH;��H;��H;��H;��H;(�H;��H;b�H;��H;p�H;i�H;t�H;K�H;t�H;f�H;m�H;�H;d�H;��H;(�H;��H;��H;��H;��H;fH;b\G;��D;�?;�5;� $;��;�M�:p)
9vrѺ�+������d�J�����ۼJ���J��v��aP��ƽձ轅����$-�       j�Yde�\0X��D�h{+�������y㻽\���VDX������ۼ;����;�E>ۻX��y�0?":޽�:��;׷-;��;;��B;�zF;�H;��H;�H;(�H;��H;��H;��H;{�H;��H;��H;��H;��H;��H;��H;��H;��H;��H;|�H;��H;��H;��H;)�H;~�H;��H;�H;�zF;��B;��;;ٷ-;��;޽�:0?":�y�X�E>ۻ��;�;����ۼ���VDX�[���y㻽��콄��h{+��D�\0X�Yde�      ��Sh��m���I���|x���O��C(���Ӫɽ����VDX�K��*<ͼㄼ�X!��s���W��tK�F��:�y;�#;I6;6R@;�PE;��G;��H;��H;5�H;��H;��H;��H;��H;��H;��H;��H;��H;��H;��H;��H;��H;��H;��H;��H;��H;��H;6�H;��H;��H;��G;�PE;5R@;I6;�#;�y;F��:�tK��W��s���X!�ㄼ*<ͼK��VDX�����Ҫɽ���C(���O��|x��I��m��Sh��      A����������%�;jɰ��G�� j�;�5��	�Ҫɽ[����J�u���沼��]�����	x�<	��dn:ͤ�:�v;��/;�-=;��C;D�F; IH;��H;'�H;��H;&�H;��H;��H;��H;�H;�H;#�H;4�H;#�H;�H;�H;��H;��H;��H;&�H;��H;'�H;��H;IH;G�F;��C;�-=;��/;�v;ˤ�:`n::	���	x������]��沼u���J�[���Ҫɽ�	�;�5� j��G��jɰ�%�;��徹���      �2�W�-�"�.E�����BKɾl����s�;�5���y㻽�v��z0��;��+���*����+6��=S��M�:\�	;��(;�9;�/B;vDF;TH;ԫH;��H;��H;��H;{�H;��H;�H;A�H;O�H;K�H;j�H;L�H;N�H;A�H;�H;��H;{�H;��H;��H;��H;ҫH;SH;yDF;�/B;�9;��(;_�	;�M�:�=S�*6�����*��+���;�z0��v��y㻽��;�5���s�l��BKɾ����.E�"�W�-�      (3s�!cm�=�\�j�C�7�%�����TҾl�� j��C(����aP����[�~������Y�8��_X�0�<���k:K��:�� ;�5;GR@;cuE;�G;5�H;K�H;��H;�H;N�H;x�H;3�H;r�H;�H;d�H;��H;d�H;�H;q�H;0�H;w�H;N�H;�H;��H;J�H;4�H;�G;fuE;DR@; �5;�� ;M��:��k:0�<�^X�8����Y����~���[�aP����콭C(� j�l���TҾ���7�%�j�C�=�\�!cm�      �ޞ�������bF�A�W�Y�-����BKɾ�G����O����ƽɸ��҄-���ۼㄼ44�ǐ��ζ��]:���:�;��1;�c>;m�D;�\G;FsH;��H;n�H;i�H;+�H;�H;7�H;y�H;��H;��H;��H;��H;��H;x�H;4�H;�H;+�H;f�H;j�H;��H;DsH;�\G;o�D;�c>;��1;�;	��:�]:�ζ�ǐ�54�ㄼ��ۼ҄-�ɸ��ƽ�����O��G��BKɾ���Y�-�A�W�bF�������      ��ſ���Nw���ޞ�����A�W�7�%�����jɰ��|x�h{+�ձ� ���J��  �ж��[�1�*���+�P"
9��:��;�-;��<;��C;�G;�TH;P�H;�H;��H;��H;`�H;>�H;��H;��H;��H;��H;��H;��H;��H;=�H;`�H;��H;��H;��H;P�H;�TH;�G;��C;��<;�-;��;�:P"
9+�*���\�1�ж���  ��J� ��ձ�h{+��|x�jɰ�����7�%�A�W������ޞ�Nw�����      ����� �Կp���ޞ�bF�j�C�.E�%�;�I���D���!"��k�c���֯���J��ѻɢ)��}K���:�
;�M*;s�:;�C;�F;�8H;Y�H;��H;z�H;��H;J�H;H�H;��H;��H;��H;
�H;��H;��H;��H;E�H;H�H;��H;w�H;��H;V�H;�8H;�F;�C;o�:;�M*;�
;$��:�}K�ɢ)��ѻ��J��֯��k�c�!"�����D��I��%�;.E�j�C�bF��ޞ�p�� �Կ��      ��������� �ԿNw�����=�\�"����m��\0X�����;����w����������]�"���F�����ɒ:��;9�';��9;!pB;�zF;�!H;��H;:�H;!�H;��H;Q�H;I�H;��H;��H;��H;�H;��H;��H;��H;G�H;O�H;��H;�H;7�H;��H;�!H;�zF;!pB;��9;<�';��;�ɒ:����F�"�黯�]����������w��;�����\0X�m�����"�=�\����Nw�� �Կ��𿞏�      "$�������忊�����"cm�X�-�����Sh��Yde�$-�۪ɽ�v��+�$���ɼ|mj�;���X�����ņ:wx;A�%;/�8;mB;nRF;H;0�H;V�H;�H;u�H;K�H;D�H;��H;��H;��H;3�H;��H;��H;��H;B�H;K�H;u�H;�H;T�H;0�H;H;lRF;mB;.�8;G�%;ux;�ņ:���X�:���|mj���ɼ+�$��v��۪ɽ$-�Yde�Sh������X�-�"cm��������忞����      �>���8���*�O������˿p��G�b�E\�7m־^��T�:��J�+��H�B�@��������,/�������>:�t�:Op ;�J6;EA;�IF;�NH;�H;"I;�I;I;�I;}I;I;� I;��H;9�H;��H;� I;I;|I;�I;I;�I;"I;�H;�NH;�IF;EA;�J6;Rp ;�t�:�>:���,/���������@��H�B�+���J�T�:�^��7m־E\�G�b�p���˿����O���*���8�      ��8��4��g&�7��>����<ƿ򲗿�>]�î�R�Ѿ�p���*7����'W��OR?�}�q8�������������G:� �:�!;�6;"lA;�YF;�TH;t�H;$"I;�I;�I;�I;VI;�I;r I;��H;"�H;��H;s I; I;UI;�I;�I;�I;!"I;t�H;�TH;�YF;"lA;�6;�!;� �:��G:���������r8��}�OR?�'W�����*7��p��R�Ѿî��>]�򲗿�<ƿ>���7���g&��4�      ��*��g&��#�v�V[�sL�������M�s5��>ľ����,��D�뒐��5�5�ݼ���q
��x��tk���b:Ql�:#;Η7;��A;�F;�dH;�I;b"I;I;uI;MI;I;�I;0 I;��H;��H;��H;. I;�I; I;LI;uI;
I;a"I;�I;�dH;�F;��A;ɗ7;#;Ql�:��b:�tk��x��q
���5�ݼ�5�뒐��DὭ�,����>ľs5���M����sL��V[�v��#��g&�      O�7��v����˿B1��:�y�Ŏ6��z �����5�l�+��ͽ%�����&���˼A�k� �����X�`� ����:O�;&;�9;��B;�F;�}H;�	I;n"I;:I;�I;�I;�I;VI;��H;3�H;��H;3�H;��H;VI;�I;�I;�I;9I;k"I;�	I;�}H;�F;��B;�9;&;M�;���:d� ���X� ���A�k���˼��&�%����ͽ+�5�l������z �Ŏ6�:�y�B1���˿���v�7��      ����>���V[忸˿�T���}�R�î��E۾ԗ����M���	������j��3�d����O�9�׻��/���V��:� 
;*;a;;�jC;�'G;�H;�I;"I;�I;�I;�
I;�I;�I;V�H;��H;�H;��H;U�H;�I;�I;�
I;�I;�I;"I;�I;�H;�'G;�jC;\;;*;� 
;X��: ����/�6�׻��O�d���3���j������	���M�ԗ���E۾î�}�R���T���˿V[�>���      �˿�<ƿsL��B1����>]���)�%��ֳ���{���,�u��)��T`I��J���,���3/��+��� �`/69�4�:�;p.;'.=;laD;�G;p�H;�I;H!I;eI;ZI;�	I;�I;� I;��H;!�H;r�H;!�H;��H;� I;�I;�	I;ZI;bI;F!I;�I;n�H;�G;kaD;".=;p.;�;�4�:P/69� ��+���3/��,���J��T`I�)��u�齧�,���{�ֳ�%����)��>]��B1��sL���<ƿ      p��򲗿���:�y�}�R���)�ov��>ľ^���I�Zl����������&�׮Ҽ�}�0B�Ǯ�������!:	+�:=z;�3;`j?;�\E;��G;��H;vI;�I;�I;�I;�I;�I;) I;��H;s�H;��H;s�H;��H;* I;�I;�I;�I;�I;�I;vI;��H;��G;�\E;^j?;�3;=z;+�:�!:����Ʈ��0B��}�׮Ҽ��&��������Zl��I�^���>ľov���)�}�R�:�y����򲗿      G�b��>]���M�Ŏ6�î�%���>ľ%q��|�Z�+�T9ݽ#W����L����#F���G��׻�;��n��Ȋ:�i;P$;ۘ7;p�A;JF;:CH;��H;� I;vI;|I;&I;:I;�I;%�H;��H;��H;!�H;��H;��H;&�H;�I;=I;&I;|I;rI;� I;��H;:CH;JF;l�A;ۘ7;P$;�i;�Ȋ:�n��;��׻�G�#F�������L�#W��T9ݽ+�|�Z�%q���>ľ%��î�Ŏ6���M��>]�      E\�î�s5��z ��E۾ֳ�^��|�Z�N?#����A����j�'��Gϼ�����µ���lۺ:�9�4�:[�;e�,;��;;>�C;�G;T�H;�I;�!I;�I;MI;6I;�I;MI;,�H;�H;��H;3�H;��H;�H;.�H;NI;�I;4I;KI;�I;�!I;�I;U�H;�G;:�C;��;;e�,;\�;�4�::�9�lۺµ�������Gϼ'����j��A�����N?#�|�Z�^��ֳ��E۾�z �s5�î�      7m־R�Ѿ�>ľ����ԗ����{��I�+�����V���{�@�/�(���,��>=�?�һX�@��� ��k:�:b;��3;8j?;r2E;��G;t�H;=I;| I;�I;�I;.	I;I;��H;	�H;��H;��H;i�H;��H;��H;	�H;��H;
I;.	I;�I;�I;| I;<I;t�H;��G;n2E;6j?;��3;b;�:�k:� �Y�@�?�һ>=��,��(��@�/��{��V�����+��I���{�ԗ�������>ľR�Ѿ      ^���p����5�l���M���,�Zl�T9ݽ�A���{���5��J��
;���T[� ?�����,P���P�9��:��;,*;(�9;dkB;ۇF;�NH;��H;& I;�I;�I;*I;I;OI;q�H;��H;��H;��H;}�H;��H;��H;��H;n�H;RI;I;(I;�I;�I;& I;��H;�NH;ׇF;bkB;(�9;+*;��;��:�P�9.P������ ?��T[�
;���J����5��{��A��T9ݽZl���,���M�5�l����p��      T�:��*7���,�+���	�t�齅���#W����j�@�/��J���I���k�j�.��T��h ���Ȋ:eo�:;dr3;)�>;4�D;t�G;V�H;I;:!I;�I;�I;�
I;I;p I;��H;��H;��H;��H;t�H;��H;��H;��H;��H;r I;I;�
I;�I;�I;7!I;I;T�H;q�G;1�D;'�>;dr3;;eo�:�Ȋ:x ��T��.��j��k��I���J��@�/���j�#W������t�齄�	�+���,��*7�      �J�����D��ͽ���)�������L�'��(��
;���k����eI����/�L/���>:J��:�B;k�,;��:;7�B;�xF;�<H;��H;I;�I;�I;RI;�I;�I;��H;��H;I�H;��H;��H;��H;��H;��H;J�H;��H;��H;�I;�I;OI;�I;�I;I;��H;�<H;�xF;7�B;��:;i�,;�B;R��:��>:D/���/�eI������k�
;��(��'����L����)������ͽ�D����      +��'W��뒐�$�����j�S`I���&����Fϼ�,���T[�j�eI��Q;�`nk��:05�:�;&;ߡ6;�!@;B2E;�G;��H;�I;!I;]I; I;I;II;� I;��H;�H;��H;w�H;��H;\�H;��H;u�H;��H;�H;��H;� I;JI;I;I;]I;!I;�I;��H;ݤG;A2E;�!@;�6;&;�;,5�:�:\nk�Q;�eI��j��T[��,��Fϼ�����&�S`I���j�$���꒐�'W��      G�B�NR?��5���&��3��J��֮Ҽ#F����>=� ?�.����/�dnk����9T׳:��;;!;b3;��=;��C;+�F; dH;�H;�I;I;�I;5I;�I;�I;X�H;�H;��H;��H;X�H;��H;O�H;��H;X�H;��H;��H;�H;X�H;�I;�I;5I;�I;!I;�I;�H;dH;+�F;��C;��=;b3;?!;��;T׳:���9dnk���/�.�� ?�?=���#F��֮Ҽ�J���3���&��5�OR?�      ?��}�2�ݼ��˼d���,���}��G����>�һ����T��D/��:\׳:�;vb;��0;�<;��B;�IF;zH;5�H;�I;� I;*I;JI;m
I;�I;5 I;C�H;h�H;!�H;<�H;8�H;��H;R�H;��H;7�H;<�H;!�H;j�H;C�H;4 I;�I;m
I;GI;+I;� I;�I;/�H;zH;�IF;��B;�<;��0;vb;�;\׳:�:H/�R������?�һ����G��}��,��d����˼2�ݼ}�      ����o8����?�k���O��3/�,B��׻����U�@�&P��h ����>:,5�:��;tb;��/;7;;I�A;��E;ѿG;�H;�
I;w I;I;I;�I;�I;�I;��H;R�H;��H;��H;�H;*�H;��H;J�H;��H;*�H;�H;��H;��H;R�H;��H;�I;�I;�I;I;I;s I;�
I;�H;οG;��E;I�A;9;;��/;tb;��;,5�:��>:h ��&P��V�@������׻,B��3/���O�?�k���q8��      ������q
����6�׻�+��Į���;��lۺ� ��P�9�Ȋ:L��:�;=!;��0;8;;˓A;�pE;��G;܎H;��H;�I;II;jI;6I;�I;�I;�H;Y�H;��H;�H;7�H;�H;�H;z�H;S�H;z�H;�H;�H;5�H;�H;��H;W�H;�H;�I;�I;7I;iI;EI;�I;��H;َH;��G;�pE;͓A;7;;��0;=!;�;P��:�Ȋ:�P�9�� ��lۺ�;�Į���+��4�׻����q
���      &/�������x���X���/� � ������n�H:�9�k:��:ko�:�B;&;d3;�<;K�A;�pE;otG;	}H;<�H;;I;�I;WI; I;�
I;I;h I;g�H;;�H;��H;��H;��H;��H;�H;��H;��H;��H;�H;��H;��H;��H;��H;8�H;d�H;h I;	I;�
I; I;QI;I;:I;7�H;
}H;ptG;�pE;H�A;�<;f3;&;�B;ko�:��:�k:P:�9�n������� ���/���X���x����      쯕�Z���dtk�T� � ��`/69�!:�Ȋ:�4�:�:��;;i�,;ۡ6;��=;��B;��E;��G;}H;��H;�I;' I;�I;nI;�I;?I;�I;_�H;�H;U�H;��H;*�H;��H;��H;�H;��H;��H;��H;
�H;��H;��H;,�H;��H;R�H;��H;_�H;�I;?I;�I;jI;�I;& I;�I;��H;}H;��G;��E;��B;��=;ۡ6;i�,;;��;�:�4�:�Ȋ:�!:�/69���T� �dtk�j���      �>:��G:��b:���:L��:�4�:+�:�i;\�;b;,*;br3;��:;�!@;��C;�IF;ѿG;ێH;<�H;�I;/ I;WI;OI;�I;)I;tI;7�H;��H;��H;��H;d�H;��H;��H;��H;/�H;��H;��H;��H;/�H;��H;��H;��H;d�H;��H;��H;��H;5�H;uI;)I;�I;OI;WI;- I;�I;:�H;ގH;пG;�IF;��C;�!@;��:;br3;+*;b;]�;�i;+�:�4�:L��:���:�b:��G:      �t�:� �:{l�:I�;� 
;��;Jz;(P$;n�,;��3;/�9;+�>;:�B;D2E;.�F;zH;�H;��H;;I;) I;VI;�I;NI;�I;I;��H;;�H;g�H;��H;��H;��H;��H;��H;��H;Q�H;�H;��H;�H;Q�H;��H;��H;��H;��H;��H;��H;g�H;:�H;��H;I;�I;LI;�I;TI;* I;:I;��H;�H;yH;/�F;D2E;:�B;+�>;-�9;��3;l�,;*P$;Jz;��;� 
;I�;}l�:� �:      Yp ;�!;#;&;*;p.;�3;ޘ7;��;;<j?;gkB;8�D;�xF;�G; dH;2�H;�
I;�I;�I;�I;OI;PI;�I;nI;K�H;��H;��H;A�H;�H;/�H;��H;��H;��H;�H;p�H;6�H;#�H;6�H;p�H;�H;��H;��H;��H;,�H; �H;A�H;��H;��H;L�H;kI;�I;PI;KI;�I;�I;�I;�
I;1�H; dH;�G;�xF;8�D;ikB;:j?;��;;��7;�3;	p.;*;&;#;�!;      �J6;(�6;ٗ7;�9;f;;(.=;lj?;p�A;C�C;u2E;އF;x�G;�<H;��H;�H;�I;w I;KI;VI;mI;�I;�I;nI;d�H;��H;��H;{�H;I�H;V�H;��H;��H;��H;��H;D�H;��H;��H;g�H;��H;��H;F�H;��H;��H;��H;��H;T�H;I�H;z�H;��H;��H;`�H;mI;�I;�I;mI;VI;LI;v I;�I;�H;��H;�<H;x�G;݇F;t2E;C�C;s�A;jj?;*.=;m;;�9;ٗ7;�6;      EA;0lA;p�A;��B;kC;raD;�\E;JF;�G;��G;�NH;[�H; �H; I;�I;� I;I;kI;I;�I;,I;I;R�H;��H;�H;��H;Q�H;f�H;��H;��H;��H;��H;��H;|�H;�H;��H;��H;��H;�H;z�H;��H;��H;��H;��H;��H;f�H;O�H;��H;�H;��H;O�H;I;*I;�I;I;nI;I;� I;�I;�I;��H;[�H;�NH;��G;�G;JF;�\E;saD;kC;��B;q�A;0lA;      �IF;�YF;�F;�F;�'G;�G;��G;=CH;[�H;x�H;��H;I;I;!I;I;(I;
I;4I;
I;<I;rI;��H;��H;��H;��H;z�H;��H;��H;��H;��H;��H;��H;S�H;��H;n�H;P�H;@�H;P�H;o�H;��H;O�H;��H;��H;��H;��H;��H;�H;z�H;��H;��H;��H;��H;mI;<I;
I;4I;I;(I;I;!I;I;I;��H;u�H;Y�H;;CH;��G;�G;�'G;�F;�F;�YF;      �NH;�TH;�dH;�}H;��H;x�H;��H;��H;�I;@I;, I;@!I;�I;`I;�I;JI;�I;�I;I;�I;9�H;=�H;��H;~�H;L�H;��H;��H;��H;��H;��H;��H;�H;��H;(�H;��H;��H;��H;��H;��H;&�H;��H;�H;��H;��H;��H;��H;��H;��H;M�H;|�H;��H;;�H;3�H;�I;I;�I;�I;II;�I;`I;�I;@!I;, I;@I;�I;��H;��H;u�H;��H;�}H;�dH;�TH;      	�H;}�H;�I;�	I;I;�I;~I;� I;�!I;� I;�I;�I;�I;$I;7I;n
I;�I;�I;g I;b�H;��H;g�H;C�H;J�H;b�H;��H;��H;��H;}�H;��H;�H;j�H;�H;��H;j�H;:�H;2�H;:�H;j�H;��H;�H;j�H;�H;��H;{�H;��H;��H;��H;c�H;J�H;A�H;g�H;��H;a�H;e I;�I;�I;m
I;6I;"I;�I;�I;�I;� I;�!I;� I;~I;�I;I;�	I;�I;��H;      !"I;+"I;c"I;x"I;"I;M!I;�I;|I;�I;�I;�I;�I;UI;I;�I;�I;�I;�H;g�H;�H;��H;��H;��H;Y�H;��H;��H;��H;}�H;��H;�H;^�H;��H;{�H;,�H;��H;��H;��H;��H;��H;,�H;x�H;��H;^�H;�H;��H;}�H;��H;��H;��H;Y�H;��H;��H;��H;��H;d�H;�H;�I;�I;�I;I;TI;�I;�I;�I;�I;}I;�I;K!I;"I;x"I;e"I;""I;      �I;�I;I;>I;I;oI;�I;�I;YI;�I;5I;�
I;�I;UI;�I;8 I;��H;U�H;8�H;V�H;��H;��H;)�H;��H;��H;��H;��H;��H;�H;P�H;��H;w�H;��H;��H;��H;~�H;l�H;~�H;��H;��H;��H;x�H;��H;N�H;�H;��H;��H;��H;��H;��H;(�H;��H;��H;V�H;8�H;V�H;��H;8 I;�I;SI;�I;�
I;6I;�I;[I;�I;�I;oI;I;@I;I;�I;      'I;I;�I;�I;�I;]I;�I;5I;BI;8	I;)I;I;�I;� I;]�H;J�H;[�H;��H;��H;�H;h�H;��H;��H;��H;��H;��H;��H;�H;^�H;��H;[�H;��H;��H;p�H;=�H; �H;�H; �H;=�H;p�H;��H;��H;Y�H;��H;^�H;�H;��H;��H;��H;��H;��H;��H;e�H;�H;��H;��H;X�H;J�H;]�H;� I;�I;I;)I;;	I;BI;5I;�I;^I;�I;�I;�I;I;      �I;�I;WI;�I;�
I;�	I;�I;II;�I;I;[I;~ I;��H;��H;�H;s�H;��H;�H;��H;4�H;��H;��H;��H;��H;��H;��H;�H;m�H;��H;w�H;��H;��H;U�H;.�H;��H;��H;��H;��H;��H;.�H;S�H;��H;��H;x�H;��H;m�H;�H;��H;��H;��H;��H;��H;��H;3�H;��H;�H;��H;s�H;�H;��H;��H;} I;[I;I;�I;HI;�I;�	I;�
I;�I;WI;�I;      �I;mI;I;�I;�I;�I;�I;�I;[I;��H;{�H;��H;��H; �H;��H;(�H;��H;5�H;��H;��H;��H;��H;��H;��H;��H;S�H;��H;�H;~�H;��H;��H;W�H;�H;��H;��H;��H;��H;��H;��H;��H;�H;X�H;��H;�H;�H;�H;��H;P�H;��H;��H;��H;��H;��H;��H;��H;7�H;��H;)�H;��H; �H;��H;��H;{�H;��H;[I;�I;�I;�I;�I;�I;I;eI;      !I;I;�I;cI;�I;� I;1 I;6�H;6�H;�H;��H;��H;Q�H;��H;��H;F�H;�H;�H;��H;��H;��H;��H;�H;G�H;v�H;��H;#�H;��H;+�H;��H;o�H;.�H;��H;��H;��H;��H;n�H;��H;��H;��H;��H;1�H;o�H;��H;.�H;��H;#�H;��H;v�H;F�H;�H;��H;��H;��H;��H;�H;�H;F�H;��H;��H;P�H;��H;��H;�H;7�H;7�H;1 I;� I;�I;cI;�I;I;      � I;� I;A I;��H;u�H;��H;��H;�H;"�H;��H;��H;��H;��H;~�H;^�H;B�H;6�H;�H;�H;�H;6�H;R�H;m�H;��H;�H;m�H;��H;k�H;��H;��H;=�H;��H;��H;��H;h�H;]�H;^�H;]�H;h�H;��H;��H;��H;=�H;��H;��H;k�H;��H;m�H;�H;��H;o�H;R�H;3�H;�H;�H;�H;4�H;B�H;_�H;~�H;��H;��H;��H; �H;#�H;�H;��H;��H;k�H;��H;? I;� I;      ��H;��H;��H;=�H;��H;!�H;~�H;��H;��H;��H;��H;��H;��H;��H;��H;��H;��H;w�H;��H;��H;��H;	�H;6�H;��H;��H;N�H;��H;<�H;��H;}�H;!�H;��H;��H;��H;]�H;B�H;B�H;B�H;]�H;��H;��H;��H;!�H;~�H;��H;<�H;��H;L�H;��H;��H;6�H;	�H;��H;��H;��H;x�H;��H;��H;��H;��H;��H;��H;��H;��H;��H;��H;~�H;&�H;��H;:�H;��H;��H;      =�H;2�H;�H;��H;&�H;s�H;��H;-�H;=�H;l�H;��H;��H;��H;f�H;T�H;\�H;R�H;N�H;��H;��H;��H;��H; �H;h�H;��H;=�H;��H;7�H;��H;o�H;�H;��H;��H;p�H;^�H;C�H;?�H;C�H;^�H;p�H;��H;��H;�H;p�H;��H;7�H;��H;>�H;��H;e�H; �H;��H;��H;��H;��H;P�H;Q�H;\�H;T�H;f�H;��H;��H;��H;o�H;?�H;,�H;��H;w�H;�H;��H;�H;)�H;      ��H;��H;��H;:�H;��H;!�H;~�H;��H;��H;��H;��H;��H;��H;��H;��H;��H;��H;w�H;��H;��H;��H;	�H;6�H;��H;��H;N�H;��H;<�H;��H;}�H;!�H;��H;��H;��H;]�H;B�H;B�H;B�H;]�H;��H;��H;��H;!�H;~�H;��H;<�H;��H;L�H;��H;��H;6�H;	�H;��H;��H;��H;x�H;��H;��H;��H;��H;��H;��H;��H;��H;��H;��H;~�H;&�H;��H;=�H;��H;��H;      ~ I;� I;? I;��H;u�H;��H;��H;�H;#�H;��H;��H;��H;��H;~�H;_�H;B�H;6�H;�H;�H;�H;7�H;R�H;o�H;��H;�H;k�H;��H;k�H;��H;��H;=�H;��H;��H;��H;h�H;]�H;^�H;]�H;h�H;��H;��H;��H;=�H;��H;��H;k�H;��H;m�H;�H;��H;m�H;R�H;3�H;�H;�H;�H;4�H;B�H;_�H;~�H;��H;��H;��H;��H;"�H;�H;��H;��H;k�H;��H;> I;� I;      "I;I;�I;cI;�I;� I;1 I;6�H;6�H;�H;��H;��H;P�H;��H;��H;F�H;�H;�H;��H;��H;��H;��H;�H;G�H;v�H;��H;#�H;��H;,�H;��H;o�H;.�H;��H;��H;��H;��H;n�H;��H;��H;��H;��H;1�H;o�H;��H;.�H;��H;#�H;��H;v�H;F�H;�H;��H;��H;��H;��H;�H;�H;F�H;��H;��H;Q�H;��H;��H;�H;7�H;6�H;1 I;� I;�I;cI;�I;I;      �I;mI;I;�I;�I;�I;�I;�I;[I;��H;{�H;��H;��H; �H;��H;)�H;��H;5�H;��H;��H;��H;��H;��H;��H;��H;Q�H;��H;�H;~�H;��H;��H;W�H;�H;��H;��H;��H;��H;��H;��H;��H;�H;Z�H;��H;�H;�H;�H;��H;Q�H;��H;��H;��H;��H;��H;��H;��H;5�H;��H;(�H;��H; �H;��H;��H;{�H;��H;[I;�I;�I;�I;�I;�I;I;kI;      �I;�I;ZI;�I;�
I;�	I;�I;HI;�I;I;[I;~ I;��H;��H;�H;s�H;��H;�H;��H;4�H;��H;��H;��H;��H;��H;��H;�H;m�H;��H;w�H;��H;��H;T�H;.�H;��H;��H;��H;��H;��H;.�H;S�H;��H;��H;x�H;��H;m�H;�H;��H;��H;��H;��H;��H;��H;4�H;��H; �H;��H;s�H;�H;��H;��H;} I;[I;I;�I;GI;�I;�	I;�
I;�I;ZI;�I;      'I;I;�I;�I;�I;]I;�I;4I;BI;9	I;)I;I;�I;� I;]�H;L�H;Y�H;��H;��H;�H;j�H;��H;��H;��H;��H;��H;��H;�H;]�H;��H;Y�H;��H;��H;p�H;=�H; �H;�H; �H;=�H;p�H;��H;��H;[�H;��H;`�H;�H;��H;��H;��H;��H;��H;��H;e�H;�H;��H;��H;X�H;J�H;]�H;� I;�I;I;&I;9	I;BI;5I;�I;^I;�I;�I;�I;I;      �I;�I;I;@I;I;lI;�I;�I;\I;�I;6I;�
I;�I;TI;�I;8 I;��H;U�H;8�H;Y�H;��H;��H;)�H;��H;��H;��H;��H;��H;�H;O�H;��H;w�H;��H;��H;��H;~�H;l�H;~�H;��H;��H;��H;x�H;��H;O�H;�H;��H;��H;��H;��H;��H;(�H;��H;��H;V�H;8�H;V�H;��H;: I;�I;TI;�I;�
I;5I;�I;\I;�I;�I;nI;I;>I;I;�I;      "I;'"I;i"I;u"I;"I;H!I;�I;I;�I;�I;�I;�I;TI;I;�I;�I;�I;�H;d�H;�H;��H;��H;��H;Y�H;��H;��H;��H;}�H;��H;�H;^�H;��H;z�H;,�H;��H;��H;��H;��H;��H;,�H;z�H;��H;^�H;�H;��H;}�H;��H;��H;��H;Y�H;��H;��H;��H;�H;g�H;�H;�I;�I;�I;I;UI;�I;�I;�I;�I;I;�I;J!I;"I;s"I;k"I;("I;      	�H;{�H;�I;�	I;I;�I;~I;� I;�!I;� I;�I;�I;�I;$I;7I;m
I;�I;�I;e I;a�H;��H;g�H;C�H;J�H;c�H;��H;��H;��H;}�H;��H;�H;j�H;�H;��H;i�H;:�H;2�H;:�H;j�H;��H;�H;k�H;�H;��H;{�H;��H;��H;��H;b�H;J�H;A�H;g�H;��H;b�H;g I;�I;�I;p
I;7I;"I;�I;�I;�I;� I;�!I;� I;~I;�I;I;�	I;�I;��H;      �NH;�TH;�dH;�}H;��H;t�H;��H;��H;�I;BI;, I;@!I;�I;_I;�I;JI;�I;�I;I;�I;:�H;;�H;��H;~�H;M�H;��H;��H;��H;��H;��H;��H;�H;��H;&�H;��H;��H;��H;��H;��H;&�H;��H;�H;��H;��H;��H;��H;��H;��H;L�H;|�H;��H;=�H;5�H;�I;I;�I;�I;II;�I;`I;�I;@!I;, I;BI;�I;��H;��H;r�H;��H;�}H;�dH;�TH;      �IF;�YF;�F;�F;�'G;�G;��G;;CH;X�H;w�H;��H;I;I;!I;I;(I;
I;3I;
I;<I;tI;��H;��H;��H;��H;z�H;�H;��H;��H;��H;��H;��H;Q�H;��H;m�H;P�H;@�H;P�H;o�H;��H;O�H;��H;��H;��H;��H;��H;�H;z�H;��H;��H;��H;��H;mI;<I;
I;6I;I;(I;I;!I;I;I;��H;u�H;Y�H;;CH;��G;�G;�'G;�F;�F;�YF;      EA;0lA;p�A;��B; kC;raD;�\E;JF;�G;��G;�NH;[�H;��H;�I;�I;� I;I;kI;I;�I;-I;I;P�H;��H;�H;��H;P�H;f�H;��H;��H;��H;��H;��H;z�H;�H;��H;��H;��H;�H;z�H;��H;��H;��H;��H;��H;f�H;P�H;��H;�H;��H;P�H;I;*I;�I;I;nI;I;� I;�I;�I; �H;[�H;�NH;��G;�G;JF;�\E;raD;�jC;��B;q�A;1lA;      �J6;%�6;��7;�9;_;;..=;ij?;q�A;D�C;v2E;އF;x�G;�<H;��H;�H;�I;w I;KI;VI;mI;�I;�I;nI;d�H;��H;��H;{�H;I�H;X�H;��H;��H;��H;��H;D�H;��H;��H;g�H;��H;��H;D�H;��H;��H;��H;��H;T�H;I�H;z�H;��H;��H;d�H;mI;�I;�I;mI;VI;LI;v I;�I;�H;��H;�<H;x�G;݇F;t2E;D�C;q�A;ij?;..=;m;;�9;�7;�6;      Tp ;�!;#;&;*;p.;�3;ޘ7;��;;<j?;ikB;8�D;�xF;�G; dH;2�H;�
I;�I;�I;�I;RI;PI;�I;nI;L�H;��H;��H;A�H;�H;/�H;��H;��H;��H;�H;p�H;6�H;#�H;6�H;p�H;�H;��H;��H;��H;,�H; �H;A�H;��H;��H;K�H;kI;�I;PI;KI;�I;�I;�I;�
I;2�H;"dH;�G;�xF;8�D;ikB;9j?;��;;ޘ7;�3;p.;*;&;#;�!;      �t�:� �:{l�:I�;� 
;��;Jz;)P$;l�,;��3;/�9;+�>;:�B;D2E;.�F;zH;�H;��H;:I;) I;XI;�I;NI;�I;I;��H;;�H;g�H;��H;��H;��H;��H;��H;��H;Q�H;�H;��H;�H;Q�H;��H;��H;��H;��H;��H;��H;g�H;9�H;��H;I;�I;LI;�I;TI;* I;;I;��H;�H;zH;/�F;D2E;:�B;-�>;-�9;��3;n�,;(P$;Jz;��;� 
;I�;}l�:� �:      ��>:��G:�b:���:J��:�4�:+�:�i;\�;b;,*;br3;��:;�!@;��C;�IF;ѿG;܎H;:�H;�I;/ I;WI;OI;�I;)I;uI;6�H;��H;��H;��H;d�H;��H;��H;��H;/�H;��H;��H;��H;/�H;��H;��H;��H;d�H;��H;��H;��H;6�H;tI;)I;�I;NI;WI;- I;�I;<�H;ގH;пG;�IF;��C;�!@;��:;br3;.*;b;_�;�i;+�:�4�:V��:���:�b:��G:      ����V���Xtk�\� ����`/69�!:�Ȋ:�4�:�:��;;h�,;ۡ6;��=;��B;��E;��G;}H;��H;�I;& I;�I;pI;�I;?I;�I;_�H;�H;U�H;��H;*�H;��H;��H;
�H;��H;��H;��H;�H;��H;��H;,�H;��H;R�H;��H;_�H;�I;?I;�I;jI;�I;' I;�I;��H;}H;��G;��E;��B;��=;ۡ6;i�,;;��;�:�4�:�Ȋ:�!:�/69���\� �dtk�j���      &/�������x���X���/� � ������n�H:�9�k:��:ko�:�B;&;d3;�<;K�A;�pE;ptG;	}H;<�H;:I;�I;VI; I;�
I;I;h I;g�H;;�H;��H;��H;��H;��H;�H;��H;��H;��H;�H;��H;��H;��H;��H;8�H;b�H;h I;I;�
I; I;SI;�I;;I;9�H;
}H;otG;�pE;H�A;�<;f3;&;�B;ko�:��:�k:P:�9�n������� ���/���X���x����      ������q
����8�׻ ,��Ʈ���;��lۺ�� ��P�9�Ȋ:P��:�;=!;��0;8;;˓A;�pE;��G;܎H;��H;�I;II;iI;7I;�I;�I;�H;Y�H;��H;�H;7�H;�H;�H;z�H;S�H;z�H;�H;�H;5�H;�H;��H;W�H;�H;�I;�I;7I;jI;EI;�I;��H;؎H;��G;�pE;͓A;7;;��0;=!;�;L��:�Ȋ:�P�9� ��lۺ�;�Ʈ���+��6�׻����q
���      ����o8����@�k���O��3/�-B��׻����V�@�&P��h ����>:,5�:��;tb;��/;7;;I�A;��E;пG;�H;�
I;w I;I;
I;�I;�I;�I;��H;R�H;��H;��H;�H;*�H;�H;J�H;��H;*�H;�H;��H;��H;R�H;��H;�I;�I;�I;I;I;s I;�
I;�H;οG;��E;I�A;9;;��/;tb;��;,5�:��>:h ��&P��V�@������׻-B��3/���O�?�k���p8��      ?��}�2�ݼ��˼d���,���}��G����?�һ����R��H/��:Z׳:�;xb;��0;�<;��B;�IF;zH;2�H;�I;� I;*I;JI;m
I;�I;4 I;C�H;i�H;"�H;<�H;7�H;��H;R�H;��H;8�H;<�H;�H;j�H;C�H;5 I;�I;m
I;GI;+I;� I;�I;1�H;zH;�IF;��B;�<;��0;ub;�;Z׳:�:D/�T������>�һ����G��}��,��d����˼2�ݼ}�      G�B�NR?��5���&��3��J��֮Ҽ#F����?=� ?�.����/�dnk����9T׳:��;<!;b3;��=;��C;+�F; dH;�H;�I;!I;�I;5I;�I;�I;X�H;�H;��H;��H;X�H;��H;O�H;��H;X�H;��H;��H;�H;X�H;�I;�I;5I;�I;I;�I;�H;dH;+�F;��C;��=;b3;=!;��;T׳:���9dnk���/�.�� ?�>=���#F��׮Ҽ�J���3���&��5�OR?�      +��'W��뒐�$�����j�S`I���&����Fϼ�,���T[�j�eI��Q;�\nk��:05�:�;&;ޡ6;�!@;A2E;�G;��H;�I;!I;_I;I;I;JI;� I;��H;�H;��H;u�H;��H;\�H;��H;w�H;��H;�H;��H;� I;II;I; I;]I;!I;�I;��H;ޤG;B2E;�!@;ޡ6;&;�;.5�:�:`nk�Q;�eI��j��T[��,��Fϼ�����&�S`I���j�$���뒐�'W��      �J�����D��ͽ���)�������L�'��(��
;���k����eI����/�H/���>:P��:�B;i�,;��:;7�B;�xF;�<H;��H;I;�I;�I;QI;�I;�I;��H;��H;J�H;��H;��H;��H;��H;��H;I�H;��H;��H;�I;�I;OI;�I;�I;I;��H;�<H;�xF;7�B;��:;i�,;�B;R��:��>:L/���/�eI������k�
;��(��'����L����)������ͽ�D����      T�:��*7���,�+���	�t�齅���#W����j�@�/��J���I���k�j�.��T��p ���Ȋ:eo�:;ar3;'�>;4�D;t�G;T�H;I;9!I;�I;�I;�
I;I;o I;��H;��H;��H;��H;t�H;��H;��H;��H;��H;r I;I;�
I;�I;�I;9!I;I;V�H;q�G;1�D;)�>;dr3;;eo�:�Ȋ:p ��U��.��j��k��I���J��@�/���j�#W������t�齄�	�+���,��*7�      ^���p����5�l���M���,�Zl�T9ݽ�A���{���5��J��
;���T[� ?�����,P���P�9��:��;**;(�9;ckB;ۇF;�NH;��H;& I;�I;�I;(I;I;NI;p�H;��H;��H;��H;}�H;��H;��H;��H;p�H;QI;I;*I;�I;�I;& I;��H;�NH;ׇF;bkB;(�9;**;��;��:�P�9.P������ ?��T[�
;���J����5��{��A��T9ݽZl���,���M�5�l����p��      7m־R�Ѿ�>ľ����ԗ����{��I�+�����V���{�@�/�(���,��?=�?�һX�@��� ��k:�:b;��3;8j?;q2E;��G;t�H;=I;| I;�I;�I;.	I;I;��H;	�H;��H;��H;i�H;��H;��H;	�H;��H;I;.	I;�I;�I;| I;<I;t�H;��G;o2E;6j?;��3;b;�:�k:� �Y�@�@�һ?=��,��(��@�/��{��V�����+��I���{�ԗ�������>ľR�Ѿ      E\�î�s5��z ��E۾ֳ�^��|�Z�N?#����A����j�'��Gϼ�����µ���lۺ:�9�4�:Y�;e�,;��;;=�C;�G;U�H;�I;�!I;�I;KI;4I;�I;PI;.�H;�H;��H;3�H;��H;�H;,�H;LI;�I;6I;KI;�I;�!I;�I;T�H;�G;<�C;��;;e�,;\�;�4�::�9�lۺĵ�������Gϼ'����j��A�����N?#�|�Z�^��ֳ��E۾�z �s5�î�      G�b��>]���M�Ŏ6�î�%���>ľ%q��|�Z�+�T9ݽ#W����L����#F���G��׻�;��n��Ȋ:�i;P$;ۘ7;o�A;JF;:CH;��H;� I;uI;|I;&I;;I;�I;(�H;��H;��H;!�H;��H;��H;&�H;�I;:I;&I;|I;sI;� I;��H;9CH;JF;l�A;ۘ7;P$;�i;�Ȋ:�n��;��׻�G�#F�������L�#W��T9ݽ+�|�Z�%q���>ľ%��î�Ŏ6���M��>]�      p��򲗿���:�y�}�R���)�ov��>ľ^���I�Zl����������&�׮Ҽ�}�/B�Ʈ�������!:+�:=z;�3;bj?;�\E;��G;��H;vI;�I;�I;�I;�I;�I;, I;��H;s�H;��H;s�H;��H;) I;�I;�I;�I;�I;�I;vI;��H;��G;�\E;_j?;�3;=z;+�:�!:����Ʈ��0B��}�׮Ҽ��&��������Zl��I�^���>ľov���)�}�R�:�y����򲗿      �˿�<ƿsL��B1����>]���)�%��ֳ���{���,�u��)��T`I��J���,���3/��+��� �0/69�4�:�;p.;'.=;kaD;�G;p�H;�I;J!I;gI;ZI;�	I;�I;� I;��H;!�H;r�H;#�H;��H;� I;�I;�	I;ZI;bI;D!I;�I;n�H;�G;laD;".=;p.;�;�4�:0/69� ��+���3/��,���J��T`I�)��u�齧�,���{�ֳ�%����)��>]��B1��sL���<ƿ      ����>���V[忸˿�T���}�R�î��E۾ԗ����M���	������j��3�d����O�8�׻��/� ��R��:� 
;*;a;;�jC;�'G;�H;�I;"I;�I;�I;�
I;�I;�I;V�H;��H;�H;��H;U�H;�I;�I;�
I;�I;�I;"I;�I;�H;�'G;�jC;^;;*;� 
;X��: ����/�8�׻��O�d���3���j������	���M�ԗ���E۾î�}�R���T���˿V[�>���      O�7��v����˿B1��:�y�Ŏ6��z �����5�l�+��ͽ%�����&���˼A�k� �����X�`� ����:M�;&;�9;��B;�F;�}H;�	I;n"I;;I;�I;�I;�I;VI;��H;3�H;��H;3�H;��H;VI;�I;�I;�I;9I;k"I;�	I;�}H;�F;��B;�9;&;O�;���:d� ���X� ���B�k���˼��&�%����ͽ+�5�l������z �Ŏ6�:�y�B1���˿���v�7��      ��*��g&��#�v�V[�sL�������M�s5��>ľ����,��D�뒐��5�5�ݼ���q
��x��tk���b:Ql�:#;Η7;��A;�F;�dH;�I;c"I;I;uI;MI;I;�I;0 I;��H;��H;��H;0 I;�I; I;LI;uI;
I;_"I;�I;�dH;�F;��A;ɗ7;#;Ql�:��b:�tk��x��q
���5�ݼ�5�뒐��DὭ�,����>ľs5���M����sL��V[�v��#��g&�      ��8��4��g&�7��>����<ƿ򲗿�>]�î�R�Ѿ�p���*7����'W��OR?�}�q8�������������G:� �:�!;�6;"lA;�YF;�TH;t�H;$"I;�I;�I;�I;VI; I;r I;��H;"�H;��H;s I;�I;UI;�I;�I;�I;!"I;t�H;�TH;�YF;"lA;�6;�!;� �:��G:���������r8��}�OR?�'W�����*7��p��R�Ѿî��>]�򲗿�<ƿ>���7���g&��4�      �Aq���i���U�H:�@�����>���w���}A�f5�� ���^Z�����A���]�����d��J",��5��^�Ѻ���9��:^�;bY4;r�@;�VF;��H;�GI;�bI;9OI;J:I;*I;NI;�I;�I;�I;�I;�I;�I;�I;MI;*I;J:I;7OI;�bI;�GI;��H;�VF;r�@;^Y4;a�;��:���9b�Ѻ�5��I",��d������]��A������^Z�� ��f5�}A�w���>�������@�H:���U���i�      ��i���b�\�O�.5�2i�������������q<���� f��c
V�IE	�!���IY�k9�D�����(��R����Ⱥx�:{��: �;H�4;l�@;khF;×H;9II;�bI;�NI;�9I;�)I;I;�I;�I;�I;�I;�I;�I;�I;I;�)I;�9I;�NI;�bI;9II;×H;khF;l�@;D�4;$�;{��:|�:��Ⱥ�R����(�E���k9��IY�!��IE	�c
V� f������q<������������2i�.5�\�O���b�      ��U�\�O�J-?�/�'���O�ῶ欿d�{�ga/���뾟���I����f���ZN�`5������;H�\ �������":��:��;��5;�`A;ܛF;^�H;?MI;"bI;�MI;�8I;)I;qI;I;oI;5I;7I;5I;nI;I;pI;)I;�8I;�MI;bI;AMI;_�H;ܛF;�`A;��5;��;��:��":���\ ��:H�����`5���ZN�f������I�������ga/�d�{��欿O����/�'�J-?�\�O�      H:�.5�/�'��������lȿ���n$_���Y�Ҿݕ���6�����*���`=�?�漮)��FG�6��d��T�Q:��:0";�7;�&B;�F;��H;SI;�`I;�KI;L7I;�'I;kI;II;�I;�I;�
I;�I;�I;JI;kI;�'I;L7I;�KI;�`I;SI;��H;�F;�&B;�7;0";��:\�Q:f��6��FG��)��>���`=��*������6�ݕ��Y�Ҿ��n$_����lȿ�������/�'�.5�      @�2i�������K�ѿl������q<��:��a����q����Wн齅���'�Wb̼�zl��.��;�X�����:��;�&;٫9;RC;zMG;�H;cYI;�^I;�HI;5I;	&I;I;9I;�I;�
I;�	I;�
I;�I;9I;I;&I;5I;�HI;�^I;cYI;�H;xMG;PC;ի9;�&;��;�:���;�X��.���zl�Wb̼��'�齅��Wн����q��a���:��q<���l���K�ѿ������2i�      �������O��lȿl���������O���~]׾|����I�����A��A�d�o�֮�RH��jλ=�$�0&����:bN;ǆ+;�<;'4D;�G;�I;�^I;�[I;EI;Q2I;�#I;pI;�I;�I;�	I;�I;�	I;�I;�I;pI;�#I;Q2I;EI;�[I;�^I;�I;�G;&4D;�<;ǆ+;bN;���:@&�=�$��jλRH�֮�o�A�d��A������I�|���~]׾����O�����l���lȿO�Ῥ��      >��������欿�������O��x����� ���l���"��ܽ���`=����v���k"�&R��ۺ ��9�?�:xL;��0;͟>;�ME;#H;�%I;�aI;3WI;�@I;#/I;p!I;kI;3I;@I;}I;�I;}I;@I;4I;kI;q!I;#/I;�@I;0WI;�aI;�%I;�#H;�ME;ɟ>;��0;xL;�?�:�9ۺ$R���k"�v������`=����ܽ��"��l�� ����뾂x���O�������欿����      w�������c�{�n$_��q<������~��	w���6�����!���h����㷾�� d�w.���^e��H[�t�Z:���:�, ;��5;�A;�VF;҄H;AI;�bI;�QI;<I;o+I;�I;<I;jI;�	I;I;`I;I;�	I;iI;;I;�I;o+I;<I;�QI;�bI;AI;ЄH;�VF;�A;��5;�, ;���:l�Z:�H[��^e�x.��� d�㷾�����h�!�������6�	w��~��������q<�n$_�c�{�����      }A��q<�ga/����:�~]׾� ��	w��>�EE	�����۽����3�b�꼚���",��W��I���Q�ʰ�:�M
;�f);ޅ:;I@C; @G;��H;oTI;�_I;XKI;7I;}'I;�I;�I;nI;I;�I;�I;�I;I;oI;�I;�I;}'I;7I;UKI;�_I;mTI;��H;@G;F@C;ޅ:;�f);�M
;İ�:�Q�H���W��",�����b�꼚�3�۽������EE	�>�	w��� ��~]׾�:���ga/��q<�      f5�������Y�Ҿ�a��|����l��6�EE	���Ƚk���aG����e֮��W����W�k����$d,:���:�;��1;o�>;bE;T�G;KI;Q_I;rZI;hDI;�1I;a#I;sI;*I;5
I;=I;I;PI;I;?I;6
I;'I;sI;`#I;�1I;eDI;pZI;P_I;LI;Q�G;_E;l�>;��1;�;���:$d,:���X�k�����W�e֮�����aG�k����ȽEE	��6��l�|����a��Y�Ҿ������      � �� f�����ݕ����q��I���"���������k���ZN�\�"¼P�y��$��Q��p� � X��:D0;K�&;x8;� B;��F;�H;�@I;#bI;�RI;J=I;B,I;I;I;�I;I;kI;MI;�I;MI;kI;I;�I;I;I;A,I;G=I;�RI; bI;�@I;�H;��F;� B;x8;I�&;D0;�: �W�r� ��Q���$�P�y�"¼\��ZN�k������������"��I���q�ݕ����� f��      �^Z�c
V��I��6�������ܽ!��۽���aG�\��ȼ�)��z�(�^��6G5�@���Z:\�:8S;0'1;��=;ӠD;Y�G;�H;�XI;G^I;�II;(6I;�&I;�I;�I;�
I;�I;�I;� I;��H;� I;�I;�I;�
I;�I;�I;�&I;%6I;�II;G^I;�XI;�H;T�G;ѠD;��=;0'1;6S;\�:�Z:L��6G5�_��z�(��)���ȼ\��aG�۽��!���ܽ������6��I�c
V�      ���HE	��������Wн�A�����h���3����"¼�)��/x/��һ\�X�B#����9���:�>;^f);�`9;�&B;��F;�}H;7I;�aI;�UI;�@I;	/I;-!I;zI;YI;I;�I;� I;��H;0�H;��H;� I;�I;I;[I;{I;.!I;/I;�@I;�UI;�aI;7I;�}H;ۊF;�&B;�`9;]f);�>;���:��9>#��\�X��һ/x/��)��"¼�����3��h��󑽤A���Wн��콻��IE	�      �A��!��e���*��轅�@�d��`=����a��e֮�N�y�z�(��һ�]e�����@�f9챩:T�;l1";H�4;�m?;E;��G;��H;�WI;�^I;;KI;�7I;&(I;�I;[I;�
I;UI;PI;��H;�H;r�H;	�H;��H;PI;UI;�
I;YI;�I;%(I;�7I;:KI;�^I;�WI;��H;��G;E;�m?;H�4;l1";W�;豩: �f9�����]e��һz�(�N�y�e֮�a�꼙���`=�@�d�轅��*��e��!��      �]��IY��ZN��`=���'�o����㷾������W��$�_��\�X�����9���:���:��;̸0;�<;�C;OG;*�H;�?I;\aI;UI;o@I;D/I;�!I;�I;DI;�I;�I;�H;��H;A�H;��H;A�H;��H;�H;�I;�I;DI;�I;�!I;D/I;n@I;UI;[aI;�?I;%�H;OG;}�C;
�<;̸0;��;���:���:9����\�X�_���$��W�����㷾����n���'��`=��ZN��IY�      ���j9�]5��=��Vb̼~֮�u��� d�	",�����Q��4G5�B#��@�f9���:��:5�;��-;��:;
LB;gVF;EKH;I;
]I;U\I;�HI;96I;R'I;OI;�I;N
I;uI;1 I;��H;��H;��H;!�H;��H;��H;��H;. I;vI;N
I;�I;KI;S'I;76I;�HI;S\I;]I;I;EKH;eVF;
LB;��:;��-;2�;��:���:@�f9B#��4G5��Q�����
",�� d�u��~֮�Vb̼=��]5��j9�      �d��B��������)���zl�	RH��k"�t.���W��Q�k�m� �<����9챩:���:1�;�-;�9;paA;�E;V�G;��H;3SI;H`I;PI;�<I;�,I;�I;hI;DI;�I;�I;��H;��H;�H;��H;��H;��H;�H;��H;��H;�I;�I;CI;eI;�I;�,I;�<I;PI;B`I;/SI;��H;T�G;�E;paA;��9;�-;1�;���:챩:��9<��n� �S�k��W��t.���k"�RH��zl��)������D���      J",���(�8H�DG��.���jλ#R���^e�D����� �W��Z:���:T�;��;��-;�9;�A;dE;R�G;��H;�GI;(aI;�UI;tBI;�1I; $I;�I;"I;�I;)I;��H;��H;�H;A�H;K�H;�H;M�H;A�H;�H;��H;��H;)I;�I;I;�I;$I;�1I;uBI;�UI;$aI;�GI;��H;S�G;dE;�A;�9;��-;��;U�;���:�Z: �W����E���^e�#R���jλ�.��DG�8H���(�      �5���R��U ��6��;�X�3�$�ۺ�H[��Q�0d,:�:d�:�>;o1";ϸ0;��:;qaA;dE;%�G;��H;�=I;``I;�YI;#GI;6I;�'I;#I;�I;0I;�I; I;;�H;W�H;-�H;��H;��H;v�H;��H;��H;-�H;U�H;<�H;  I;�I;/I;�I;I;�'I;6I;GI;�YI;_`I;�=I;��H;%�G;dE;oaA;��:;Ѹ0;o1";�>;b�:�:0d,: Q��H[�ۺ/�$�5�X�6��U ���R��      T�Ѻ��Ⱥ
���^�����0&����9l�Z:ʰ�:���:F0;8S;]f);D�4;�<;LB;�E;P�G;��H;�:I;�_I;�[I;UJI;89I;�*I;�I;+I;6I;�I;GI;!�H;��H;H�H;e�H;0�H;j�H;�H;k�H;1�H;f�H;H�H;��H; �H;CI;�I;6I;*I;�I;�*I;59I;RJI;�[I;�_I;�:I;��H;R�G;�E;LB;�<;D�4;]f);8S;F0;���:Ȱ�:t�Z: ��9�%����`��
�����Ⱥ      ���9ĺ:ī":H�Q:�:���:�?�:���:�M
;�;L�&;0'1;�`9;�m?;��C;fVF;W�G;��H;�=I;�_I;E\I;�KI;I;I;-I;!I;(I;�I;I;�I;�H;n�H;��H;p�H;��H;��H;�H;��H;�H;��H;��H;o�H;��H;n�H;�H;~I;I;�I;&I;!I; -I;H;I;�KI;B\I;�_I;�=I;��H;T�G;fVF;�C;�m?;�`9;0'1;K�&;�;�M
;���:�?�:���:�:H�Q:ī":��:      ��:���:��:��:��;nN;�L;�, ;�f);��1;x8;��=;�&B;E;QG;DKH;��H;�GI;``I;�[I;�KI;�;I;!.I;f"I;lI;JI;Q	I;�I;��H;%�H;�H;��H;��H;U�H;x�H;��H;��H;��H;x�H;U�H;��H;��H;�H;!�H;��H;�I;N	I;MI;lI;`"I;.I;�;I;�KI;�[I;``I;�GI;��H;CKH;RG;E;�&B;��=;x8;��1;�f);�, ;�L;pN;��;��:��:���:      h�;$�;��;0";�&;ˆ+;��0;��5;�:;r�>;� B;٠D;��F;��G;*�H;I;3SI;)aI;�YI;VJI;I;I;%.I;�"I;5I;�I;3
I;dI;��H;��H;��H;��H;��H;3�H;�H;*�H;��H;��H;��H;,�H;�H;2�H;��H;��H;��H;��H;�H;aI;6
I;�I;1I;�"I;$.I;E;I;WJI;�YI;+aI;1SI;I;*�H;��G;��F;ؠD;� B;p�>;�:;��5;��0;̆+;
�&;0";��;�;      zY4;Y�4;��5;�7;ݫ9;�<;ן>;�A;N@C;gE;��F;]�G;�}H;��H;�?I;]I;H`I;�UI;"GI;59I;-I;d"I;5I;XI;�
I;�I;# I; �H;��H;!�H;��H;/�H;��H;��H;��H;��H;��H;��H;��H;��H;��H;/�H;��H;�H;��H;�H;" I;�I;�
I;UI;4I;f"I;�,I;59I;"GI;�UI;E`I;]I;�?I;��H;�}H;Z�G;��F;dE;L@C;�A;ן>;�<;�9;�7;��5;K�4;      ~�@;x�@;�`A;�&B;XC;-4D;�ME;�VF;#@G;S�G;	�H;#�H;7I;�WI;_aI;V\I;"PI;uBI;6I;�*I;!I;pI;�I;�
I;$I;T I;k�H;�H;[�H;�H;:�H;��H;��H;��H;�H;��H;��H;��H;�H;��H;��H;��H;:�H;�H;X�H;�H;h�H;T I;&I;�
I;�I;pI;!I;�*I;6I;xBI; PI;U\I;_aI;�WI;7I;!�H;	�H;S�G;#@G;�VF;�ME;.4D;XC;�&B;�`A;x�@;      �VF;hF;қF;�F;MG;�G;�#H;҄H;��H;OI;�@I;�XI;�aI;�^I;UI;�HI;�<I;�1I;�'I;�I;%I;JI;0
I;�I;M I;��H;P�H;��H;&�H;3�H;��H;��H;x�H;��H;?�H;��H;��H;��H;@�H;��H;u�H;��H;��H;2�H;%�H;��H;M�H;��H;O I;�I;0
I;JI;!I;�I;�'I;�1I;�<I;�HI;UI;�^I;�aI;�XI;�@I;LI;��H;҄H;�#H;�G;�MG;�F;ӛF;thF;      ��H;ȗH;_�H;��H;�H;�I;&I;AI;vTI;U_I;&bI;N^I;�UI;<KI;r@I;:6I;�,I;$I;#I;-I;�I;Q	I;bI;% I;d�H;Q�H;��H;J�H;c�H;��H;d�H;H�H;v�H;��H;r�H;�H;�H;�H;p�H;��H;q�H;G�H;d�H;��H;b�H;J�H;��H;Q�H;e�H;# I;aI;Q	I;�I;-I;#I;$I;�,I;76I;r@I;<KI;�UI;M^I;&bI;T_I;wTI;AI;�%I;�I;�H;��H;_�H;ɗH;      �GI;AII;IMI;SI;jYI;�^I;bI;�bI; `I;yZI;�RI;�II;�@I;�7I;G/I;S'I;�I;�I;�I;8I;I;�I;�H;"�H;�H;��H;I�H;@�H;��H;e�H;?�H;D�H;��H;�H;��H;y�H;q�H;y�H;��H;�H;��H;D�H;=�H;a�H;��H;@�H;H�H;��H;�H; �H;}�H;�I;I;8I;�I;�I;�I;S'I;G/I;�7I;�@I;�II;�RI;yZI; `I;�bI;bI;�^I;uYI;SI;KMI;MII;      cI;�bI;"bI;�`I;�^I;�[I;:WI;�QI;]KI;lDI;N=I;06I;/I;'(I;�!I;OI;jI;I;2I;�I;�I;��H;��H;��H;T�H;'�H;`�H;��H;Y�H;:�H;2�H;u�H;��H;d�H;�H;��H;��H;��H;�H;d�H;��H;v�H;2�H;9�H;V�H;��H;b�H;'�H;V�H;��H;��H;��H;I;�I;2I; I;hI;OI;�!I;'(I;
/I;/6I;M=I;lDI;]KI;�QI;:WI;�[I;�^I;�`I;"bI;�bI;      HOI;�NI;�MI;�KI;�HI;EI;�@I;"<I;7I;�1I;M,I;�&I;6!I;�I;�I;�I;II;�I;�I;II;�H;"�H;��H; �H;�H;0�H;��H;c�H;9�H;;�H;d�H;��H;0�H;��H;|�H;[�H;V�H;\�H;|�H;��H;-�H;��H;d�H;9�H;7�H;d�H;��H;0�H;�H; �H;��H;!�H;�H;GI;�I;�I;FI;�I;�I;�I;6!I;�&I;M,I;�1I;7I;&<I;�@I;EI;�HI;�KI;�MI;�NI;      T:I;�9I;�8I;^7I;&5I;T2I;0/I;|+I;�'I;j#I;I;�I;�I;cI;JI;V
I;�I;,I; I;&�H;t�H;�H;��H;��H;5�H;��H;c�H;?�H;/�H;e�H;��H;)�H;��H;K�H;�H;��H;��H;��H;�H;K�H;��H;*�H;��H;d�H;1�H;?�H;`�H;��H;6�H;��H;��H;�H;p�H;&�H; I;,I;�I;V
I;KI;bI;�I;�I;I;m#I;�'I;|+I;//I;U2I;#5I;^7I;�8I;�9I;      *I;�)I;)I;�'I;&I;�#I;w!I;�I;�I;zI;!I;�I;_I;�
I;�I;~I;�I;��H;A�H;��H;��H;��H;��H;2�H;��H;��H;G�H;D�H;r�H;��H;(�H;��H;)�H;��H;��H;��H;s�H;��H;��H;��H;'�H;��H;)�H;��H;s�H;D�H;G�H;�H;��H;2�H;��H;��H;��H;��H;A�H;��H;�I;}I;�I;�
I;_I;�I;!I;zI;�I;�I;w!I;�#I;&I;�'I;)I;�)I;      UI;+I;~I;|I;"I;tI;qI;FI;�I;.I;�I;�
I;I;^I;�I;7 I;��H;�H;[�H;L�H;v�H;��H;2�H;��H;��H;z�H;t�H;��H;��H;3�H;��H;,�H;��H;��H;G�H;=�H;J�H;=�H;G�H;��H;��H;.�H;��H;4�H;��H;��H;q�H;w�H;��H;��H;0�H;��H;t�H;N�H;[�H;��H;��H;7 I;�I;\I;I;�
I;�I;0I;�I;GI;qI;vI;I;|I;}I;$I;      �I;�I;I;WI;GI;�I;;I;wI;wI;:
I;I;�I;�I;ZI;�H; �H;��H;�H;2�H;l�H;��H;V�H;�H;��H;��H;��H;��H;�H;c�H;��H;H�H;��H;��H;W�H;�H;�H;��H;�H;�H;W�H;��H;��H;H�H;��H;e�H;�H;��H;��H;��H;��H;�H;V�H;��H;l�H;2�H;�H;��H; �H;�H;ZI;�I;�I;I;<
I;wI;xI;;I;�I;;I;WI;I;�I;      �I;�I;}I;�I;�I;�I;HI;�	I;I;DI;vI;�I;� I;��H;��H;��H;�H;@�H;��H;8�H;��H;}�H;,�H;�H;�H;=�H;n�H;��H;�H;|�H;�H;��H;G�H;�H;�H;��H;��H;��H;�H;�H;D�H;��H;�H;~�H;
�H;��H;l�H;=�H;�H; �H;)�H;{�H;��H;7�H;��H;@�H;�H;��H;��H;��H;� I;�I;vI;FI;I;�	I;HI;�I;�I;�I;}I;�I;      �I;�I;CI;�I;�
I;�	I;�I;)I;�I;I;YI;� I;��H;�H;H�H;��H;��H;J�H;��H;r�H;�H;��H;��H;��H;��H;��H;�H;y�H;��H;[�H;��H;��H;=�H;�H;��H;��H;��H;��H;��H;�H;<�H;��H;��H;\�H;��H;y�H;�H;��H;��H;��H;��H;��H;�H;r�H;��H;K�H;��H;��H;H�H;�H;��H;� I;VI;I;�I;)I;�I;�	I;�
I;�I;BI;�I;      �I;�I;KI;�
I;�	I;�I;�I;jI;�I;SI;�I;��H;7�H;|�H;��H;*�H;��H;�H;z�H;&�H;��H;��H;��H;��H;��H;��H;�H;t�H;��H;Y�H;��H;x�H;L�H;��H;��H;��H;��H;��H;��H;��H;I�H;z�H;��H;\�H;��H;t�H; �H;��H;��H;��H;��H;��H;��H;&�H;z�H;�H;��H;*�H;��H;|�H;7�H;��H;�I;VI;�I;iI;�I;�I;�	I;�
I;KI;�I;      �I;�I;CI;�I;�
I;�	I;�I;)I;�I;I;YI;� I;��H;�H;H�H;��H;��H;J�H;��H;r�H;�H;��H;��H;��H;��H;��H;�H;y�H;��H;[�H;��H;��H;=�H;�H;��H;��H;��H;��H;��H;�H;<�H;��H;��H;\�H;��H;y�H;�H;��H;��H;��H;��H;��H;�H;r�H;��H;K�H;��H;��H;H�H;�H;��H;� I;XI;
I;�I;)I;�I;�	I;�
I;�I;?I;�I;      �I;�I;}I;�I;�I;�I;HI;�	I;I;FI;vI;�I;� I;��H;��H;��H;�H;@�H;��H;7�H;��H;{�H;*�H;�H;�H;=�H;o�H;��H;	�H;|�H;�H;��H;G�H;�H;�H;��H;��H;��H;�H;�H;D�H;��H;�H;~�H;
�H;��H;l�H;=�H;�H;��H;*�H;}�H;��H;8�H;��H;@�H;�H;��H;��H;��H;� I;�I;uI;FI;I;�	I;HI;�I;�I;�I;|I;�I;      �I;�I;I;WI;GI;�I;;I;wI;vI;<
I;I;�I;�I;ZI;�H; �H;��H;�H;2�H;l�H;��H;V�H;�H;��H;��H;��H;��H;�H;c�H;��H;H�H;��H;��H;W�H;�H;�H;��H;�H;�H;W�H;��H;��H;H�H;��H;e�H;�H;��H;��H;��H;��H;�H;V�H;��H;l�H;2�H;�H;��H; �H;�H;ZI;�I;�I;I;:
I;yI;wI;;I;�I;;I;WI;I;�I;      XI;,I;I;}I;!I;sI;oI;DI;�I;.I;�I;�
I;I;\I;�I;7 I;��H;�H;[�H;L�H;w�H;��H;3�H;��H;��H;x�H;t�H;��H;��H;3�H;��H;,�H;��H;��H;G�H;=�H;J�H;=�H;G�H;��H;��H;/�H;��H;4�H;��H;��H;p�H;x�H;��H;��H;0�H;��H;s�H;N�H;[�H;�H;��H;7 I;�I;^I;I;�
I;�I;0I;�I;DI;qI;vI;I;}I;}I;)I;      *I;�)I;)I;�'I;&I;�#I;x!I;�I;�I;zI;!I;�I;_I;�
I;�I;}I;�I;��H;A�H;��H;��H;��H;��H;2�H;��H;��H;G�H;D�H;s�H;��H;)�H;��H;)�H;��H;��H;��H;s�H;��H;��H;��H;'�H;��H;(�H;��H;s�H;D�H;F�H;��H;��H;2�H;��H;��H;��H;��H;A�H;��H;�I;~I;�I;�
I;_I;�I;!I;|I;�I;�I;z!I;�#I;&I;�'I;)I;�)I;      T:I;�9I;�8I;^7I;$5I;T2I;//I;{+I;�'I;k#I;I;�I;�I;cI;KI;X
I;�I;*I; I;$�H;t�H;�H;��H;��H;6�H;��H;`�H;?�H;/�H;e�H;��H;*�H;��H;K�H;�H;��H;��H;��H;�H;K�H;��H;*�H;��H;d�H;1�H;?�H;a�H;��H;5�H;��H;��H;�H;p�H;'�H; I;,I;�I;V
I;KI;cI;�I;�I;I;k#I;�'I;|+I;0/I;U2I;#5I;^7I;�8I;�9I;      >OI;�NI;�MI;�KI;�HI;EI;�@I;#<I;7I;�1I;M,I;�&I;6!I;�I;�I;�I;GI;�I;�I;II;�H;!�H;��H; �H;�H;2�H;��H;c�H;:�H;;�H;d�H;��H;/�H;��H;|�H;[�H;V�H;\�H;|�H;��H;/�H;��H;d�H;9�H;9�H;c�H;��H;0�H;�H; �H;��H;"�H;�H;II;�I;�I;FI;�I;�I;�I;5!I;�&I;M,I;�1I;7I;%<I;�@I;EI;�HI;�KI;�MI;�NI;      �bI;�bI;(bI;�`I;�^I;�[I;<WI;�QI;]KI;lDI;P=I;06I;
/I;'(I;�!I;OI;jI;I;2I;�I;�I;��H;��H;��H;V�H;'�H;_�H;��H;W�H;:�H;2�H;s�H;��H;d�H;�H;��H;��H;��H;�H;d�H;��H;v�H;2�H;9�H;W�H;��H;`�H;'�H;T�H;��H;��H;��H;~I;�I;2I; I;hI;PI;�!I;)(I;/I;06I;N=I;kDI;]KI;�QI;<WI;�[I;�^I;�`I;(bI;�bI;      �GI;@II;KMI;SI;hYI;�^I;bI;�bI;�_I;yZI;�RI;�II;�@I;�7I;G/I;S'I;�I;�I;�I;8I; I;�I;�H; �H;�H;��H;H�H;@�H;��H;c�H;=�H;D�H;��H;�H;��H;y�H;q�H;y�H;��H;�H;��H;F�H;?�H;c�H;��H;@�H;H�H;��H;�H;#�H;�H;�I;I;8I;�I;�I;�I;U'I;G/I;�7I;�@I;�II;�RI;yZI; `I;�bI;bI;�^I;sYI;SI;KMI;OII;      ��H;ƗH;d�H;��H;	�H;�I;�%I;AI;vTI;U_I;&bI;M^I;�UI;<KI;r@I;96I;�,I;$I;#I;.I;�I;Q	I;bI;% I;e�H;Q�H;��H;J�H;c�H;��H;d�H;G�H;t�H;��H;p�H;�H;�H;�H;r�H;��H;t�H;J�H;d�H;��H;b�H;J�H;��H;S�H;d�H;% I;aI;Q	I;�I;-I;#I;$I;�,I;96I;r@I;>KI;�UI;N^I;'bI;U_I;tTI;AI;�%I;�I;�H;��H;a�H;��H;      �VF;{hF;ܛF;�F;MG;�G;�#H;҄H;��H;OI;�@I;�XI;�aI;�^I;UI;�HI;�<I;�1I;�'I;�I;&I;JI;0
I;�I;O I;��H;N�H;��H;'�H;3�H;��H;��H;w�H;��H;?�H;��H;��H;��H;@�H;��H;u�H;��H;��H;0�H;%�H;��H;M�H;��H;M I;�I;2
I;JI;!I;�I;�'I;�1I;�<I;�HI;UI;�^I;�aI;�XI;�@I;LI;��H;҄H;�#H;�G;�MG;�F;ݛF;qhF;      ~�@;z�@;�`A;�&B;XC;-4D;�ME;�VF;%@G;T�G;�H;!�H;7I;�WI;_aI;V\I;!PI;uBI;6I;�*I;!I;pI;�I;�
I;&I;T I;i�H;�H;[�H;�H;:�H;��H;��H;��H;�H;��H;��H;��H;�H;��H;��H;��H;:�H;�H;X�H;�H;h�H;T I;$I;�
I;�I;pI;!I;�*I;6I;xBI; PI;V\I;_aI;�WI;7I;#�H;	�H;Q�G;#@G;�VF;�ME;-4D;VC;�&B;�`A;z�@;      |Y4;Y�4;��5;�7;֫9;<;ԟ>;�A;N@C;gE;��F;[�G;�}H;��H;�?I;]I;H`I;�UI;"GI;59I;-I;f"I;5I;XI;�
I;�I;# I;�H;��H;!�H;��H;/�H;��H;��H;��H;��H;��H;��H;��H;��H;��H;0�H;��H;�H;��H; �H;" I;�I;�
I;WI;4I;d"I;�,I;59I;"GI;�UI;G`I;]I;�?I;��H;�}H;]�G;��F;eE;O@C;�A;ԟ>;<;�9;�7;��5;L�4;      d�;2�;��;0"; �&;φ+;��0;��5;�:;r�>;� B;ؠD;ߊF;��G;*�H;I;3SI;(aI;�YI;VJI;K;I;$.I;�"I;5I;�I;5
I;dI;�H;��H;��H;��H;��H;3�H;�H;,�H;��H;��H;��H;*�H;�H;2�H;��H;��H;��H;��H;��H;aI;6
I;�I;4I;�"I;%.I;E;I;WJI;�YI;+aI;3SI;I;,�H;��G;��F;ؠD;� B;o�>;�:;��5;��0;ц+;�&;0";��; �;      ��:���:��:��:��;nN;�L;�, ;�f);��1;x8;��=;�&B;E;OG;DKH;��H;�GI;``I;�[I;�KI;�;I;!.I;d"I;lI;LI;P	I;�I;��H;%�H;�H;��H;��H;U�H;x�H;��H;��H;��H;x�H;U�H;��H;��H;�H;!�H;��H;�I;M	I;MI;lI;c"I;.I;�;I;�KI;�[I;``I;�GI;��H;DKH;RG;E;�&B; �=;x8;��1;�f);�, ;�L;nN;��;��:��:���:      ���9��:ث":L�Q:�:���:�?�:���:�M
;�;L�&;0'1;�`9;�m?;�C;fVF;V�G;��H;�=I;�_I;E\I;�KI;I;I;-I;!I;&I;�I;I;�I;�H;n�H;��H;p�H;��H;��H;�H;��H;�H;��H;��H;p�H;��H;n�H;�H;~I;I;�I;(I;!I; -I;H;I;�KI;B\I;�_I;�=I;��H;T�G;fVF;��C;�m?;�`9;0'1;N�&;�;�M
;���:�?�:���:�:L�Q:ܫ":��:      Z�Ѻ��Ⱥ���`�����&� ��9l�Z:ʰ�:���:H0;6S;]f);D�4;�<;LB;�E;P�G;��H;�:I;�_I;�[I;UJI;99I;�*I;�I;+I;6I;�I;FI; �H;��H;I�H;f�H;1�H;k�H;�H;k�H;0�H;e�H;G�H;��H;!�H;CI;�I;6I;(I;�I;�*I;49I;RJI;�[I;�_I;�:I;��H;R�G;�E;LB;�<;E�4;]f);6S;D0;���:ʰ�:x�Z: ��9 &����`��
�����Ⱥ      �5���R��U ��6��<�X�4�$�ۺ�H[� Q�0d,:�:b�:�>;o1";ϸ0;��:;qaA;dE;%�G;��H;�=I;_`I;�YI;#GI;6I;�'I;"I;�I;2I;�I;  I;;�H;W�H;-�H;��H;��H;v�H;��H;��H;-�H;U�H;<�H; I;�I;-I;�I; I;�'I;6I;GI;�YI;``I;�=I;��H;%�G;dE;paA;��:;Ѹ0;o1";�>;d�:�:0d,:�Q��H[�ۺ/�$�7�X�6��U ���R��      I",���(�8H�DG��.���jλ$R���^e�E����� �W��Z:���:T�;��;��-;�9;�A;dE;R�G;��H;�GI;(aI;�UI;uBI;�1I;$I;�I;#I;�I;)I;��H;��H;�H;A�H;K�H;�H;K�H;A�H;�H;��H;��H;)I;�I;I;�I;$I;�1I;tBI;�UI;%aI;�GI;��H;S�G;dE;�A;�9;��-;��;T�;���:�Z: �W����E���^e�$R���jλ�.��DG�8H���(�      �d��B��������)���zl�
RH��k"�t.���W��S�k�m� �<����9챩:���:1�;�-;�9;paA;�E;V�G;��H;4SI;G`I;PI;�<I;�,I;�I;iI;DI;�I;�I;��H;��H;�H;��H;��H;��H;�H;��H;��H;�I;�I;CI;eI;�I;�,I;�<I;PI;D`I;-SI;��H;T�G;�E;paA;��9;�-;1�;���:챩:��9<��m� �S�k��W��t.���k"�	RH��zl��)������D���      ���j9�]5��=��Vb̼~֮�u��� d�
",�����Q��4G5�B#��@�f9���:��:5�;��-;��:;
LB;gVF;EKH;
I;
]I;S\I;�HI;:6I;S'I;OI;�I;N
I;uI;0 I;��H;��H;��H;!�H;��H;��H;��H;0 I;vI;N
I;�I;KI;R'I;76I;�HI;U\I;]I;	I;EKH;eVF;
LB;��:;��-;4�;��:���:@�f9B#��4G5��Q�����	",�� d�u��~֮�Vb̼=��]5��j9�      �]��IY��ZN��`=���'�o����㷾������W��$�_��\�X����� 9���:���:��;̸0;�<;}�C;OG;*�H;�?I;[aI;UI;o@I;D/I;�!I;�I;DI;�I;�I;�H;��H;A�H;��H;A�H;��H;�H;�I;�I;DI;�I;�!I;D/I;o@I;UI;\aI;�?I;%�H;OG;}�C;	�<;̸0;��;���:���:9����\�X�_���$��W�����㷾����n���'��`=��ZN��IY�      �A��!��e���*��轅�@�d��`=����a��e֮�N�y�z�(��һ�]e����� �f9챩:U�;l1";G�4;�m?;E;��G;��H;�WI;�^I;:KI;�7I;'(I;�I;YI;�
I;WI;QI;��H;�H;r�H;�H;��H;NI;TI;�
I;[I;�I;%(I;�7I;:KI;�^I;�WI;��H;��G;E;�m?;G�4;l1";W�;豩:@�f9�����]e��һz�(�N�y�e֮�`�꼙���`=�@�d�轅��*��e��!��      ���HE	��������Wн�A�����h���3����"¼�)��/x/��һ\�X�B#����9���:�>;]f);�`9;�&B;ߊF;�}H;7I;�aI;�UI;�@I;
/I;.!I;{I;YI;I;�I;� I;��H;0�H;��H;� I;�I;I;YI;zI;-!I;/I;�@I;�UI;�aI;7I;�}H;܊F;�&B;�`9;]f);�>;���:��9B#��\�X��һ/x/��)��"¼�����3��h��󑽤A���Wн��콻��IE	�      �^Z�c
V��I��6�������ܽ!��۽���aG�\��ȼ�)��{�(�_��6G5�@���Z:\�:6S;.'1;��=;ӠD;W�G;�H;�XI;G^I;�II;(6I;�&I;�I;�I;�
I;�I;�I;� I;��H;� I;�I;�I;�
I;�I;�I;�&I;'6I;�II;F^I;�XI;�H;T�G;ѠD;��=;0'1;6S;\�:�Z:D��7G5�_��z�(��)���ȼ\��aG�۽��!���ܽ������6��I�c
V�      � �� f�����ݕ����q��I���"���������k���ZN�\�"¼P�y��$��Q��p� � �W��:D0;H�&;x8;� B;��F;�H;�@I;"bI;�RI;J=I;A,I;I;I;�I;I;kI;MI;�I;MI;kI;I;�I;I;I;B,I;G=I;�RI;"bI;�@I;�H;��F;� B;x8;I�&;D0;�: �W�q� ��Q���$�P�y�"¼\��ZN�k������������"��I���q�ݕ����� f��      f5�������Y�Ҿ�a��|����l��6�EE	���Ƚk���aG����e֮��W����W�k���$d,:���:�;��1;m�>;bE;Q�G;LI;Q_I;pZI;hDI;�1I;`#I;sI;)I;6
I;=I;I;PI;I;=I;5
I;)I;rI;a#I;�1I;eDI;rZI;P_I;KI;T�G;_E;m�>;��1;�;���:$d,:���W�k�����W�e֮�����aG�k����ȽEE	��6��l�|����a��Y�Ҿ������      }A��q<�ga/����:�~]׾� ��	w��>�EE	�����۽����3�b�꼚���",��W��I���Q�Ȱ�:�M
;�f);ޅ:;I@C;@G;��H;pTI;�_I;XKI;7I;}'I;�I;�I;oI;I;�I;�I;�I;I;nI;�I;�I;}'I;7I;UKI;�_I;mTI;��H; @G;F@C;ޅ:;�f);�M
;Ȱ�:�Q�H���W��",�����b�꼚�3�۽������EE	�>�	w��� ��~]׾�:���ga/��q<�      w�������c�{�n$_��q<������~��	w���6�����!���h����㷾�� d�v.���^e��H[�t�Z:���:�, ;��5;�A;�VF;҄H;AI;�bI;�QI;<I;o+I;�I;<I;jI;�	I;I;`I;I;�	I;kI;;I;�I;o+I;<I;�QI;�bI;
AI;ЄH;�VF;�A;��5;�, ;���:l�Z:�H[��^e�x.��� d�㷾�����h�!�������6�	w��~��������q<�n$_�c�{�����      >��������欿�������O��x����� ���l���"��ܽ���`=����v���k"�%R��ۺ���9�?�:xL;��0;͟>;�ME;�#H;�%I;�aI;5WI;�@I;#/I;p!I;mI;5I;@I;}I;�I;}I;@I;3I;jI;p!I;#/I;�@I;2WI;�aI;�%I;�#H;�ME;ʟ>;��0;xL;�?�:�9ۺ$R���k"�v������`=����ܽ��"��l�� ����뾂x���O�������欿����      �������O��lȿl���������O���~]׾|����I�����A��A�d�o�֮�RH��jλ=�$�@&����:bN;ņ+;�<;&4D;�G;�I;�^I;�[I;EI;Q2I;�#I;qI;�I;�I;�	I;�I;�	I;�I;�I;oI;�#I;Q2I;EI;�[I;�^I;�I;�G;'4D;�<;ǆ+;bN;���:@&�=�$��jλRH�֮�o�A�d��A������I�|���~]׾����O�����l���lȿO�Ῥ��      @�2i�������K�ѿl������q<��:��a����q����Wн齅���'�Wb̼�zl��.��;�X�����:��;�&;٫9;PC;zMG;�H;cYI;�^I;�HI;5I;	&I;I;9I;�I;�
I;�	I;�
I;�I;9I;I;&I;5I;�HI;�^I;cYI;�H;xMG;RC;֫9;�&;��;
�:���;�X��.���zl�Wb̼��'�齅��Wн����q��a���:��q<���l���K�ѿ������2i�      H:�.5�/�'��������lȿ���n$_���Y�Ҿݕ���6�����*���`=�>�漮)��FG�6��d��T�Q:��:0";�7;�&B;�F;��H;SI;�`I;�KI;N7I;�'I;lI;JI;�I;�I;�
I;�I;�I;II;iI;�'I;L7I;�KI;�`I;SI;��H;�F;�&B;�7;0";��:X�Q:f��6��FG��)��?���`=��*������6�ݕ��Y�Ҿ��n$_����lȿ�������/�'�.5�      ��U�\�O�J-?�/�'���O�ῶ欿d�{�ga/���뾟���I����f���ZN�`5������:H�\ �������":��:��;��5;�`A;ܛF;_�H;AMI;"bI;�MI;�8I;)I;qI;I;oI;5I;7I;5I;oI;I;pI;)I;�8I;�MI;bI;?MI;^�H;ڛF;�`A;��5;��;��:��":���\ ��:H�����`5���ZN�f������I�������ga/�d�{��欿O����/�'�J-?�\�O�      ��i���b�\�O�.5�2i�������������q<���� f��c
V�IE	�!���IY�k9�D�����(��R����Ⱥ|�:{��: �;H�4;l�@;khF;×H;9II;�bI;�NI;�9I;�)I;I;�I;�I;�I;�I;�I;�I;�I;I;�)I;�9I;�NI;�bI;9II;H;khF;l�@;E�4;$�;{��:x�:��Ⱥ�R����(�E���k9��IY�!��IE	�c
V� f������q<������������2i�.5�\�O���b�      ᶕ�T���Ҭ��0�_���7�|�!}߿����,b��V�/l¾Kx�e.���Ž��t�*��e����?�N����� �x9���:��;��2;]@@;�fF;J�H;��I;��I;@|I;�[I;�CI;62I;�%I;�I;�I;aI;�I;�I;�%I;52I;�CI;�[I;?|I;��I;��I;J�H;�fF;]@@;��2;��;���:@�x9���N����?�e��*����t���Že.�Kx�/l¾�V��,b����!}߿|���7�0�_�Ҭ��T���      T���E���%}��+Y��3�����$ڿ&��ƽ\����(���s��3�8����p�d�T���<<�1��Z���ȗ�9z��:�;Z%3;rp@;zF;��H;&�I;!�I;�{I;|[I;�CI;�1I;�%I;UI;�I;4I;�I;WI;�%I;�1I;�CI;|[I;�{I;�I;&�I;��H;zF;rp@;W%3;�;z��:ȗ�9\���1���<<�T��d��p�8����3��s�(�����ƽ\�&���$ڿ����3��+Y�%}�F���      Ҭ��%}�?tf��lG�آ%��p�0�ʿ\����>M����W�����d�ʤ�̷�1�d��
��I���1�\����� ��9���:V;�U4;��@;�F;I�H;	�I;�I;�yI;�YI;qBI;1I;�$I;�I;I;�I;I;�I;�$I;1I;pBI;�YI;�yI;�I;	�I;I�H;�F;��@;�U4;X;���: ��9��\����1��I���
�1�d�̷�ʤ���d�W�������>M�\���0�ʿ�p�آ%��lG�?tf�%}�      0�_��+Y��lG�!f.�|���꿴���O䂿��5���󾏰��Q�N�X��T��#�Q����{����h!�~g��񳺨	:�
�:%�;l16;��A;|G;I;a�I;��I;�vI;{WI;�@I;�/I;�#I;�I;;I;�I;;I;�I;�#I;�/I;�@I;{WI;�vI;��I;c�I;I;|G;��A;h16;(�;�
�:�	: �~g���h!�|������#�Q�T��X��Q�N���������5�O䂿�������|�!f.��lG��+Y�      ��7��3�آ%�|��<����ſ
���Ž\�=����Ͼ����b�3��载z��~�9�`�Ἑ���z��7}��ct�h�^:�+�:գ#;��8;��B;KsG;�%I;ٙI;�I;.rI;ATI;>I;�-I;A"I;~I;I;�I;I;|I;A"I;�-I;>I;BTI;+rI;�I;ۙI;�%I;JsG;��B;��8;أ#;�+�:p�^:�ct��7}��z����`���9��z����b�3�������Ͼ=��Ž\�
�����ſ�<��|�آ%��3�      |�����p������ſ&���Ps���1�4r���d���d�~I�ЈŽ��}�`*�KC���^��B�c�D��E๼ �:��;�);77;;WD;p�G;uHI;؝I;؏I;�lI; PI;�:I;E+I;J I;�I;�I;]I;�I;�I;L I;E+I;�:I; PI;�lI;ԏI;؝I;tHI;o�G;VD;37;;�);��;� �:�E�c�D��B��^�LC��`*���}�ЈŽ~I��d��d��4r����1��Ps�&����ſ��꿄p����      !}߿�$ڿ0�ʿ����
����Ps�SX:����'l¾�ǆ���7����:5���Q�����t���75�b������ �8ʼ:��;��.;��=;�EE;�YH;�hI;O�I;�I;OfI;KKI;V7I;r(I;I;!I;�I;�I;�I;!I;I;r(I;W7I;KKI;NfI;�I;O�I;�hI;�YH;�EE;��=;��.;��;ʼ:` �8���a���75��t������Q�:5�������7��ǆ�'l¾���SX:��Ps�
�������0�ʿ�$ڿ      ���&��\���O䂿Ľ\���1�����J˾Ꝓ�F�N�z��K������X�'�e�Ҽ��|��z��n��x��\�&:�P�:Ш;�W4;�@;TgF;��H;9�I;K�I;c�I;E_I;FI;73I;P%I;vI;�I;I;�I;I;�I;uI;N%I;73I;FI;E_I;`�I;K�I;9�I;��H;RgF;�@;�W4;Ш;�P�:P�&:x���n���z���|�e�ҼX�'����K���z��F�N�Ꝓ��J˾�����1�Ľ\�O䂿\���&��      �,b�ƽ\��>M���5�=��4r��'l¾Ꝓ�%&W��3�;Sؽ�z��\G����{I����?���̻v�-��	��`��:��;��&;M|9;�C;�dG;�I;j�I;~�I;�vI;�WI;Z@I;�.I;�!I;�I;�I;I;�I;I;�I;�I;�!I;�.I;Z@I;�WI;~vI;~�I;h�I;�I;�dG;�C;M|9;��&;��;^��:�	��t�-���̻��?�{I�����\G��z��;Sؽ�3�%&W�Ꝓ�'l¾4r��=����5��>M�ƽ\�      �V������������Ͼ�d���ǆ�F�N��3��c�[����\�4��*C���o���	��눻𳺐��9b��:�h;w�/;e�=;lE;(3H;�WI;�I;(�I;�kI;�OI;T:I;*I;QI;�I;#I;�I;�I;�I;#I;�I;OI;*I;T:I;�OI;�kI;(�I;�I;�WI;%3H;hE;e�=;v�/;�h;`��:���9��눻��	��o�*C��4����\�[���cི3�F�N��ǆ��d����Ͼ���������      /l¾(��V������������d���7�z��;Sؽ[���d�D*�dkּ+\����'�"���R�h}����:�Z;��#;a=7;X�A;@�F;��H;��I;�I;�I;aI;�GI;"4I;U%I;�I;�I;�I;|
I;	I;|
I;�I;�I;�I;W%I;"4I;�GI;aI;�I;�I;��I;��H;<�F;U�A;a=7;��#;�Z;��:`}���R�"����'�+\��dkּD*��d�[��;Sؽz����7��d���������V���(��      Kx��s���d�P�N�b�3�~I����K����z����\�D*��ݼH���-<<���ڻ��V��ct���&:���:iC;�</;xD=;�D;��G;$9I;��I;ӔI;CtI;\VI;�?I;�-I;� I;�I;�I;�
I;*I;EI;*I;�
I;�I;�I;� I;�-I;�?I;\VI;CtI;ӔI;��I;9I;��G;�D;xD=;�</;hC;���:��&:�ct���V���ڻ-<<�H����ݼD*���\��z��K������~I�b�3�P�N���d��s�      e.��3�ʤ�X����ЈŽ:5�����[G�3��dkּH����xC��>�P6}�଼� �x9���:.	;]�&;�;8;��A;ΟF;޹H;eyI;��I;$�I;bfI;�KI;}7I;�'I;�I;�I;�I;FI;�I;�I;�I;EI;�I;�I;�I;�'I;}7I;�KI;bfI;#�I;I;dyI;ڹH;ʟF;��A;�;8;[�&;.	;���:��x9ެ��P6}��>��xC�H���dkּ3��[G����:5��ЈŽ��X��ʤ��3�      ��Ž7���̷�S���z����}��Q�X�'����*C��+\��,<<��>�zn������x��:u��:7�;�'3;��>;�E;�H;�<I;�I;ԕI;�vI;�XI;�AI;�/I;�!I;I;!I;�	I;�I;VI;�I;VI;�I;�	I;"I;I;�!I;�/I;�AI;�XI;�vI;ԕI; �I;�<I;�H;�E;��>;�'3;7�;w��:t��:����xn���>�,<<�+\��*C�����X�'��Q���}��z��S��̷�7���      ��t��p�0�d�"�Q�~�9�`*����e�Ҽ{I���o���'���ڻN6}��ຠ7���:�m�:��;�.;E<;�oC;k7G;��H;�I;
�I;�I;OfI;pLI;,8I;(I;I;�I;�I;|I;�I;� I;� I;� I;�I;I;�I;�I;I;(I;)8I;rLI;NfI;	�I;	�I;��I;��H;k7G;�oC;F<;�.;��;�m�:��:�7���P6}���ڻ��'��o�{I��e�Ҽ���`*�~�9�"�Q�0�d��p�      *��c��
����_��KC���t����|���?���	� ���V�ެ������:�:�h;D�+;�9;��A;�fF;��H;�_I;��I;ɑI;5sI;�VI;�@I;/I; !I;�I;?I;I;�I;� I;��H;<�H;��H;� I;�I;I;@I;�I; !I;/I;�@I;�VI;6sI;ǑI;��I;�_I;��H;�fF;��A;�9;E�+;�h;�:��:��ެ���V� ����	���?���|��t��JC��_������
�d�      d��R���I��{�������^��75��z���̻�눻�R��ct� �x9z��:�m�:�h;��*; �8;�@;�E;g(H;�8I;��I;H�I;�~I;�`I;�HI;�5I;�&I;�I;lI;/
I;�I;� I;%�H;��H;�H;��H;'�H;� I;�I;/
I;jI;�I;�&I;�5I;�HI;�`I;�~I;B�I;�I;�8I;e(H;�E;�@;�8;��*;�h;�m�:z��:��x9�ct��R��눻��̻�z��75��^����{����I��S��      ��?��<<� �1��h!��z��B�`���n��p�-��@}����&:���:u��:��;A�+;�8;f�@;^E;��G;uI;�I;��I;e�I;�iI;nPI;<<I;�+I;�I;�I;�I;`I;�I;�H;��H;��H;�H;��H;��H;�H;�I;bI;�I;�I;�I;�+I;;<I;nPI;�iI;a�I;}�I;�I;rI;��G;^E;h�@;��8;A�+;��;u��:���:��&:H}���p�-��n��`���B黴z��h!� �1��<<�      N��.��U���{g���7}�Z�D�z��x��p	�����9��:���:4	;;�;�.;�9;�@;^E;��G;qI;�I;8�I;�I;�pI;�VI;�AI;�0I;�"I;�I;"I;&I;�I;��H;��H;��H;��H;�H;��H;��H;��H;��H;�I;&I;I;�I;�"I;�0I;�AI;�VI;�pI;z�I;8�I;	�I;qI;��G;^E;�@;�9;�.;;�;4	;���:��:���9p	��x��{��U�D�7}�{g��U���.��      ���0��� ����ct��E๠ �8P�&:d��:h��:�Z;kC;[�&;�'3;C<;��A;�E;��G;oI;�|I;��I;ӐI;�uI;�[I;@FI;�4I;c&I;�I;�I;
I;)I;n�H;��H;l�H;��H;��H;U�H;��H;��H;l�H;��H;o�H;)I;
I;~I;�I;`&I;�4I;@FI;�[I;�uI;ӐI;�I;�|I;oI;��G;�E;��A;C<;�'3;[�&;iC;�Z;b��:`��:\�&:� �8�E๼ct����@���      ��x9X��9`��9�	:X�^:� �:!ʼ:�P�:��;�h;��#;�</;�;8;��>;�oC;�fF;i(H;wI;�I;��I;�I;1xI;�^I;oII;�7I;@)I;@I;�I;�I;�I;� I;~�H;��H;n�H;��H;��H;��H;��H;��H;o�H;��H;��H;� I;I;�I;�I;@I;B)I;�7I;jII;�^I;0xI;ߑI;��I;�I;xI;g(H;�fF;�oC;��>;�;8;�</;��#;�h;��;�P�:ʼ:� �:\�^:�	:`��9ȗ�9      ���:���:���:�
�:�+�:��;��;٨;��&;{�/;h=7;|D=;��A;�E;n7G;��H;�8I;�I;8�I;ӐI;0xI;�_I;KI;�9I;-+I;4I;oI;sI;�I;vI;9�H;��H;R�H;s�H;�H;E�H;�H;E�H;�H;t�H;P�H;��H;9�H;qI;�I;sI;lI;6I;/+I;�9I;KI;�_I;+xI;ԐI;8�I;�I;�8I;��H;n7G;�E;��A;|D=;g=7;z�/;��&;ڨ;��;��;�+�:�
�:���:���:      ��;�;Z;"�;ѣ#;�);��.;�W4;T|9;i�=;Z�A;�D;џF;�H;��H;�_I;�I;��I;��I;�uI;�^I;KI;[:I;V,I;p I;�I;�I;�I;[I;��H;<�H;k�H;B�H;��H;��H;��H;��H;��H;��H;��H;@�H;k�H;<�H;��H;XI;�I;�I;�I;r I;S,I;Y:I;KI;�^I;�uI;��I;��I;�I;�_I;��H;�H;ϟF;	�D;\�A;h�=;S|9;�W4;��.;�);٣#;"�;[;�;      Ǽ2;l%3;�U4;p16;8;97;;��=;�@;�C;oE;C�F;��G;ܹH;�<I;�I;��I;H�I;h�I;�pI;�[I;lII;�9I;T,I;� I;SI;YI;�I;I;��H;��H;��H;c�H;x�H;�H;$�H;��H;;�H;��H;&�H;�H;u�H;e�H;��H;��H;~�H;I;�I;YI;UI;� I;S,I;�9I;iII;�[I;�pI;j�I;F�I;��I;�I;�<I;ܹH;��G;B�F;lE;�C;�@;��=;:7;;ɍ8;r16;�U4;a%3;      m@@;�p@;��@;��A;��B;]D;�EE;SgF;�dG;&3H;��H;(9I;gyI;�I;�I;͑I;�~I;�iI;�VI;FFI;�7I;2+I;v I;ZI;�I;�I;vI;��H;�H;��H;X�H;Z�H;��H;��H;��H;W�H;6�H;W�H;��H;��H;��H;\�H;X�H;��H;�H;��H;uI;�I;�I;VI;u I;2+I;�7I;GFI;�VI;�iI;�~I;ʑI;�I;�I;dyI;%9I;��H;&3H;�dG;SgF;�EE;^D;��B;��A;��@;�p@;      �fF;zF;�F;G;NsG;j�G;�YH;��H;�I;�WI;��I; �I;I;֕I;	�I;5sI;�`I;lPI;�AI;�4I;=)I;3I;�I;VI;�I;�I;%�H;:�H;�H;��H;m�H;��H;P�H;g�H;��H;G�H;M�H;G�H;��H;g�H;M�H;��H;k�H;��H; �H;:�H;#�H;�I;�I;VI;�I;3I;9)I;�4I;�AI;oPI;�`I;4sI;	�I;֕I;I; �I;��I;�WI;�I;��H;�YH;j�G;RsG;�G;�F;zF;      Y�H;��H;K�H;#I;�%I;|HI;�hI;:�I;n�I;�I;�I;ڔI;&�I;�vI;QfI;�VI;�HI;;<I;�0I;c&I;DI;pI;�I;�I;rI;(�H;@�H;"�H;��H;o�H;��H;.�H;�H;D�H;��H;L�H;L�H;L�H;��H;D�H;�H;.�H;��H;n�H;��H;"�H;;�H;&�H;uI;�I;�I;pI;?I;c&I;�0I;<<I;�HI;�VI;QfI;�vI;&�I;ؔI;�I;�I;o�I;<�I;�hI;zHI;�%I;#I;K�H;��H;      ��I;2�I;�I;e�I;ߙI;ޝI;V�I;U�I;��I;-�I;�I;MtI;ffI;YI;uLI;�@I;�5I;�+I;�"I;�I;�I;sI;�I;I;��H;;�H; �H;��H;��H;��H;"�H;��H;��H;;�H;��H;z�H;a�H;z�H;��H;;�H;��H;��H;"�H;��H;�H;��H; �H;;�H;��H;I;�I;sI;�I;�I;�"I;�+I;�5I;�@I;uLI;YI;bfI;JtI;�I;,�I;��I;W�I;V�I;ޝI;�I;d�I;�I;<�I;      ��I;%�I;�I;��I; �I;ڏI;�I;g�I;�vI;�kI;aI;dVI;�KI;�AI;.8I;/I;�&I;�I;�I;�I;�I;�I;YI;��H;
�H;�H;��H;��H;��H;�H;��H;��H;��H;`�H;�H;��H;��H;��H;�H;`�H;��H;��H;��H;�H;��H;��H;��H;�H;�H;��H;XI;�I;�I;�I;�I;�I;�&I;/I;.8I;�AI;�KI;cVI;aI;�kI;�vI;i�I;�I;ڏI;'�I;��I;�I;�I;      P|I;�{I;�yI;�vI;BrI;�lI;YfI;N_I;�WI;�OI;�GI;�?I;�7I;�/I;(I;$!I;�I;�I;!I;
I;�I;sI;��H;��H;��H;��H;m�H;��H;�H;��H;��H;��H;8�H;��H;E�H;�H;��H;�H;E�H;��H;5�H;��H;��H;��H;�H;��H;k�H;��H;��H;��H;��H;sI;�I;
I;!I;�I;�I;$!I;(I;�/I;�7I;�?I;�GI;�OI;�WI;P_I;YfI;�lI;>rI;�vI;�yI;�{I;      \I;�[I;�YI;�WI;STI;"PI;VKI;FI;h@I;]:I;.4I;�-I;�'I;�!I;I;�I;tI;�I;*I;.I;� I;9�H;<�H;��H;U�H;m�H;��H;"�H;��H;��H;��H;�H;��H;�H;��H;��H;��H;��H;��H;�H;��H;�H;��H;��H;��H;"�H;��H;k�H;U�H;��H;9�H;9�H;� I;.I;)I;�I;sI;�I;I;�!I;�'I;�-I;-4I;_:I;h@I;FI;UKI;#PI;PTI;�WI;�YI;�[I;      �CI;�CI;zBI;�@I;>I; ;I;]7I;B3I;�.I; *I;^%I;� I;�I;I;�I;GI;:
I;bI;�I;v�H;��H;��H;m�H;f�H;W�H;��H;-�H;��H;��H;��H;�H;}�H;��H;��H;N�H;�H;�H;�H;N�H;��H;��H;��H;�H;��H;��H;��H;-�H;��H;Z�H;e�H;k�H;��H;��H;v�H;�I;cI;9
I;GI;�I;I;�I;� I;^%I; *I;�.I;B3I;\7I;;I;>I;�@I;{BI;�CI;      =2I;�1I;1I;�/I;�-I;H+I;v(I;W%I;�!I;TI;�I;�I;I;)I;�I;I;�I;�I;��H;��H;��H;S�H;D�H;{�H;��H;P�H;�H;��H;��H;;�H;��H;��H;m�H;'�H;��H;��H;��H;��H;��H;'�H;i�H;��H;��H;<�H;��H;��H;�H;O�H;��H;{�H;B�H;R�H;��H; �H;��H;�I;�I;I;�I;)I; I;�I;�I;UI;�!I;X%I;v(I;K+I;�-I;�/I;1I;�1I;      �%I;�%I;�$I;�#I;O"I;I I;I;�I;�I;�I;�I;�I;�I;�	I;�I;�I;� I;�H;��H;s�H;y�H;w�H;��H;	�H;��H;e�H;A�H;8�H;^�H;��H;�H;��H;"�H;��H;��H;w�H;\�H;w�H;��H;��H;!�H;��H;�H;��H;a�H;9�H;@�H;d�H;��H;�H;��H;w�H;u�H;t�H;��H;�H;� I;�I;�I;�	I;�I;�I;�I;�I;�I;�I;I;M I;D"I;�#I;�$I;�%I;      �I;lI;�I;�I;�I;�I;(I;�I;�I;)I;�I;�
I;MI;�I;�I;� I;0�H;��H;��H;��H;��H;�H;��H;'�H;��H;��H;��H;��H;�H;G�H;��H;R�H;��H;��H;N�H;B�H;J�H;B�H;N�H;��H;��H;U�H;��H;H�H;�H;��H;��H;��H;��H;'�H;��H;�H;��H;��H;��H;��H;/�H;� I;�I;�I;OI;�
I;�I;*I;�I;�I;(I;�I;�I;�I;�I;cI;      �I;�I;I;DI;)I;�I;�I;I;I;�I;�
I;8I;�I;aI;I;��H;��H;��H;��H;��H;��H;H�H;��H;��H;S�H;D�H;L�H;z�H;��H;�H;��H; �H;��H;}�H;C�H;+�H;&�H;+�H;C�H;z�H;��H;"�H;��H;�H;��H;z�H;I�H;C�H;U�H;��H;��H;H�H;��H;��H;��H;��H;��H;��H;I;`I;�I;8I;�
I;�I;I;I;�I;�I; I;BI;I;�I;      aI;AI;�I;�I;�I;]I;�I;�I;�I;�I;�	I;SI;�I;�I;� I;D�H;"�H;�H;�H;\�H;��H;#�H;��H;<�H;2�H;H�H;I�H;e�H;��H;�H;��H;�H;��H;c�H;L�H;'�H;�H;'�H;L�H;c�H;��H;�H;��H;�H;��H;e�H;F�H;J�H;2�H;:�H;��H;#�H;��H;\�H;�H;�H; �H;D�H;� I;�I;�I;SI;�	I;�I;�I;�I;�I;aI;�I;�I;�I;9I;      �I;�I;I;BI;)I;�I;�I;I;I;�I;�
I;8I;�I;aI;I;��H;��H;��H;��H;��H;��H;H�H;��H;��H;U�H;D�H;L�H;z�H;��H;�H;��H; �H;��H;}�H;C�H;+�H;&�H;+�H;C�H;z�H;��H;"�H;��H;�H;��H;z�H;I�H;C�H;S�H;��H;��H;H�H;��H;��H;��H;��H;��H;��H;I;`I;�I;8I;�
I;�I;I;I;�I;�I;I;DI;I;�I;      �I;lI;�I;�I;�I;�I;(I;�I;�I;)I;�I;�
I;OI;�I;�I;� I;0�H;��H;��H;��H;��H;�H;��H;(�H;��H;��H;��H;��H;�H;G�H;��H;R�H;��H;��H;N�H;B�H;J�H;B�H;N�H;��H;��H;V�H;��H;H�H;�H;��H;��H;��H;��H;$�H;��H;�H;��H;��H;��H;��H;/�H;� I;�I;�I;MI;�
I;�I;*I;�I;�I;(I;�I;�I;�I;�I;cI;      �%I;�%I;�$I;�#I;N"I;I I;I;�I;�I;�I;�I;�I;�I;�	I;�I;�I;� I;�H;��H;s�H;{�H;w�H;��H;	�H;��H;e�H;@�H;9�H;^�H;��H;�H;��H;"�H;��H;��H;w�H;\�H;w�H;��H;��H;!�H;��H;�H;��H;a�H;8�H;@�H;e�H;��H;�H;��H;w�H;v�H;t�H;��H;�H;� I;�I;�I;�	I;�I;�I;�I;�I;�I;�I;I;M I;D"I;�#I;�$I;�%I;      @2I;�1I;1I;�/I;�-I;G+I;u(I;U%I;�!I;TI;�I;�I; I;)I;�I;I;�I;�I;��H;��H;��H;R�H;C�H;{�H;��H;P�H;�H;��H;��H;;�H;��H;��H;j�H;%�H;��H;��H;��H;��H;��H;%�H;j�H;��H;��H;<�H;��H;��H;�H;O�H;��H;y�H;C�H;S�H;��H; �H;��H;�I;�I;I;�I;)I; I;�I;�I;UI;�!I;U%I;v(I;I+I;�-I;�/I;1I;�1I;      �CI;�CI;~BI;�@I;>I;�:I;^7I;A3I;�.I; *I;^%I;� I;�I;I;�I;GI;:
I;cI;�I;x�H;��H;��H;m�H;e�H;Z�H;��H;-�H;��H;��H;��H;�H;�H;��H;��H;N�H;�H;�H;�H;N�H;��H;��H;�H;�H;��H;��H;��H;-�H;��H;W�H;f�H;k�H;��H;��H;v�H;�I;cI;9
I;GI;�I;I;�I;� I;^%I;!*I;�.I;A3I;^7I;;I;>I;�@I;~BI;�CI;      \I;�[I;�YI;�WI;STI;"PI;UKI;FI;h@I;]:I;-4I;�-I;�'I;�!I;I;�I;sI;�I;)I;.I;� I;9�H;<�H;��H;U�H;m�H;��H;"�H;��H;��H;��H;�H;��H;�H;��H;��H;��H;��H;��H;�H;��H;�H;��H;��H;��H;"�H;��H;k�H;U�H;��H;9�H;9�H;� I;.I;*I;�I;sI;�I;I;�!I;�'I;�-I;-4I;_:I;g@I;FI;VKI;#PI;PTI;�WI;�YI;�[I;      F|I;�{I;�yI;�vI;<rI;�lI;YfI;N_I;�WI;�OI;�GI;�?I;�7I;�/I;(I;$!I;�I;�I;!I;
I;�I;sI;��H;��H;��H;��H;m�H;��H;�H;��H;��H;��H;7�H;��H;E�H;�H;��H;�H;E�H;��H;7�H;��H;��H;��H;�H;��H;k�H;��H;��H;��H;��H;sI;�I;
I;!I;�I;�I;&!I;(I;�/I;�7I;�?I;�GI;�OI;�WI;O_I;YfI;�lI;>rI;�vI;�yI;�{I;      ��I;!�I;�I;��I;%�I;ՏI;��I;i�I;�vI;�kI;aI;dVI;�KI;�AI;.8I;/I;�&I;�I;�I;�I;�I;�I;YI;��H;�H;�H;��H;��H;��H;�H;��H;��H;��H;`�H;�H;��H;��H;��H;�H;`�H;��H;��H;��H;�H;��H;��H;��H;�H;
�H;��H;XI;�I;�I;�I;�I;�I;�&I;/I;.8I;�AI;�KI;dVI;aI;�kI;�vI;j�I;��I;؏I;!�I;��I;�I;!�I;      ��I;/�I;�I;d�I;ޙI;ޝI;V�I;U�I;��I;,�I;�I;JtI;bfI;YI;uLI;�@I;�5I;�+I;�"I;�I;�I;sI;�I;I;��H;;�H; �H;��H;��H;��H;"�H;��H;��H;9�H;��H;z�H;a�H;z�H;��H;;�H;��H;��H;"�H;��H;�H;��H; �H;;�H;��H;I;�I;sI;�I;�I;�"I;�+I;�5I;�@I;uLI;YI;ffI;MtI;�I;-�I;��I;X�I;V�I;۝I;�I;e�I;�I;=�I;      T�H;��H;N�H;I;�%I;xHI;�hI;:�I;o�I;�I;�I;ؔI;&�I;�vI;QfI;�VI;�HI;;<I;�0I;d&I;FI;pI;�I;�I;uI;(�H;>�H;"�H;��H;o�H;��H;.�H;�H;D�H;��H;L�H;L�H;J�H;��H;C�H;�H;0�H;��H;n�H;��H;"�H;;�H;(�H;rI;�I;�I;pI;@I;d&I;�0I;<<I;�HI;�VI;QfI;�vI;&�I;ڔI;�I;�I;n�I;:�I;�hI;xHI;�%I;I;L�H;��H;      �fF;zF;�F;�G;OsG;l�G;�YH;��H;�I;�WI;��I;��I;I;֕I;�I;5sI;�`I;nPI;�AI;�4I;@)I;3I;�I;VI;�I;�I;%�H;:�H;�H;��H;k�H;��H;O�H;g�H;��H;G�H;M�H;G�H;��H;g�H;M�H;��H;m�H;��H; �H;:�H;#�H;�I;�I;VI;�I;3I;9)I;�4I;�AI;nPI;�`I;5sI;	�I;וI;ÝI; �I;��I;�WI;�I;��H;�YH;l�G;RsG;�G;�F;zF;      m@@;�p@;��@;��A;��B;]D;�EE;SgF;�dG;(3H;��H;%9I;dyI;�I;�I;ˑI;�~I;�iI;�VI;GFI;�7I;2+I;v I;YI;�I;�I;vI;��H;�H;��H;X�H;Z�H;��H;��H;��H;W�H;6�H;W�H;��H;��H;��H;]�H;X�H;��H;�H;��H;uI;�I;�I;YI;u I;2+I;�7I;GFI;�VI;�iI;�~I;͑I;�I;�I;gyI;(9I;��H;%3H;�dG;SgF;�EE;]D;��B;��A;��@;�p@;      ʼ2;l%3;�U4;n16;��8;=7;;��=;�@;�C;oE;B�F;��G;޹H;�<I;�I;��I;H�I;g�I;�pI;�[I;mII;�9I;T,I;� I;UI;YI;�I;I;��H;��H;��H;c�H;v�H;�H;#�H;��H;;�H;��H;&�H;�H;v�H;e�H;��H;��H;~�H;I;�I;YI;SI;� I;S,I;�9I;hII;�[I;�pI;k�I;F�I;��I;�I;�<I;ܹH;��G;B�F;mE;�C;�@;��=;=7;;ˍ8;n16;�U4;_%3;      ��;�;k;$�;ϣ#;�);��.;�W4;T|9;i�=;Z�A;	�D;ΟF;�H;��H;�_I;�I;��I;��I;�uI;�^I;KI;[:I;V,I;r I;�I;�I;�I;[I;��H;<�H;k�H;B�H;��H;��H;��H;��H;��H;��H;��H;@�H;k�H;<�H;��H;XI;�I;�I;�I;p I;S,I;Y:I;KI;�^I;�uI;��I;��I;�I;�_I;��H;�H;ϟF;�D;\�A;g�=;S|9;�W4;��.;�);գ#;$�;a;�;      ���:���:���:�
�:�+�:��;��;٨;��&;z�/;h=7;|D=;��A;�E;l7G;��H;�8I;�I;8�I;ӐI;0xI;�_I;KI;�9I;/+I;4I;mI;sI;�I;vI;9�H;��H;R�H;t�H;�H;E�H;�H;E�H;�H;s�H;P�H;��H;9�H;qI;�I;sI;jI;6I;-+I;�9I;KI;�_I;-xI;ԐI;8�I;�I;�8I;��H;o7G;�E;��A;~D=;g=7;{�/;��&;ڨ;��;��;�+�:�
�:���:���:      p�x90��9���9�	:X�^:� �:#ʼ:�P�:��;�h;��#;�</;�;8;��>;�oC;�fF;h(H;wI;�I;��I;�I;0xI;�^I;oII;�7I;B)I;@I;�I;�I;�I;� I;~�H;��H;n�H;��H;��H;��H;��H;��H;n�H;��H;��H;� I;I;�I;�I;?I;B)I;�7I;jII;�^I;1xI;ݑI;��I;�I;xI;h(H;�fF;�oC;��>;�;8;�</;��#;�h;��;�P�:'ʼ:� �:p�^:�	:���9ؗ�9      ���*��������ct��E๠ �8T�&:d��:d��:�Z;iC;[�&;�'3;C<;��A;�E;��G;oI;�|I;��I;ӐI;�uI;�[I;@FI;�4I;c&I;�I;�I;
I;)I;n�H;��H;l�H;��H;��H;U�H;��H;��H;l�H;��H;o�H;)I;
I;I;�I;`&I;�4I;@FI;�[I;�uI;ӐI;�I;�|I;oI;��G;�E;��A;C<;�'3;[�&;iC;�Z;b��:d��:\�&:� �8�E��ct�� ��@���      N��.��T���{g���7}�[�D�{��x��x	�����9��:���:4	;;�;�.;�9;�@;^E;��G;oI;�I;8�I;�I;�pI;�VI;�AI;�0I;�"I;�I;!I;&I;�I;��H;��H;��H;��H;�H;��H;��H;��H;��H;�I;&I;I;�I;�"I;�0I;�AI;�VI;�pI;z�I;8�I;�I;rI;��G;^E;�@;�9;�.;;�;4	;���:��:���9p	��x��z��U�D�7}�{g��T���.��      ��?��<<� �1��h!��z��B�`���n��p�-��@}����&:���:q��:��;A�+; �8;f�@;^E;��G;uI;�I;��I;e�I;�iI;lPI;<<I;�+I;�I;�I;�I;`I;�I;�H;��H;��H;�H;��H;��H;�H;�I;bI;�I;�I;�I;�+I;:<I;oPI;�iI;a�I;}�I;�I;qI;��G;^E;h�@; �8;A�+;��;u��:���:��&:@}���p�-��n��`���B黴z��h!� �1��<<�      d��R���I��{�������^��75��z���̻�눻�R��ct���x9z��:�m�:�h;��*; �8;�@;�E;g(H;�8I;�I;F�I;�~I;�`I;�HI;�5I;�&I;�I;jI;/
I;�I;� I;'�H;��H;�H;��H;%�H;� I;�I;0
I;lI;�I;�&I;�5I;�HI;�`I;�~I;D�I;�I;�8I;e(H;�E;�@;�8;��*;�h;�m�:z��: �x9�ct��R��눻��̻�z��75��^����{����I��S��      *��c��
����_��KC���t����|���?���	� ���V�ެ������:�:�h;D�+;�9;��A;�fF;��H;�_I;��I;ǑI;6sI;�VI;�@I;/I; !I;�I;?I;I;�I;� I;��H;<�H;��H;� I;�I;I;@I;�I; !I;/I;�@I;�VI;6sI;ɑI;��I;�_I;��H;�fF;��A;�9;E�+;�h;�:��:��ެ���V� ����	���?���|��t��JC��_������
�d�      ��t��p�0�d�"�Q�~�9�`*����e�Ҽ{I���o���'���ڻP6}��ະ7���:�m�:��;�.;E<;�oC;k7G;��H;�I;	�I;�I;OfI;rLI;-8I;(I;I;�I;�I;I;�I;� I;� I;� I;�I;~I;�I;�I;I;(I;)8I;pLI;NfI;	�I;
�I;��I;��H;k7G;�oC;F<;�.;��;�m�:��:�7���N6}���ڻ��'��o�{I��e�Ҽ���`*�~�9�"�Q�0�d��p�      ��Ž7���̷�S���z����}��Q�X�'����*C��+\��,<<��>�zn������x��:u��:7�;�'3;��>;�E;�H;�<I; �I;ԕI;�vI;�XI;�AI;�/I;�!I;I;"I;�	I;�I;VI;�I;VI;�I;�	I;I;I;�!I;�/I;�AI;�XI;�vI;֕I;�I;�<I;�H;�E;��>;�'3;7�;y��:t��:����zn���>�,<<�+\��*C�����X�'��Q���}��z��S��̷�7���      e.��3�ʤ�X����ЈŽ:5�����[G�3��dkּH����xC��>�P6}�଼���x9���:.	;[�&;�;8;��A;ΟF;޹H;dyI;I;#�I;bfI;�KI;}7I;�'I;�I;�I;�I;EI;�I;�I;�I;FI;�I;�I;�I;�'I;}7I;�KI;bfI;!�I;ÝI;eyI;عH;ʟF;��A;�;8;[�&;.	;���:��x9଼�P6}��>��xC�H���dkּ3��[G����:5��ЈŽ��X��ʤ��3�      Kx��s���d�P�N�b�3�~I����K����z����\�D*��ݼH���-<<���ڻ��V��ct���&:���:hC;�</;xD=;�D;��G;9I;��I;ԔI;CtI;]VI;�?I;�-I;� I;�I;�I;�
I;,I;EI;,I;�
I;�I;�I;� I;�-I;�?I;[VI;CtI;ӔI;��I;$9I;��G;�D;xD=;�</;hC;���:��&:�ct���V���ڻ-<<�H����ݼD*���\��z��K������~I�b�3�P�N���d��s�      /l¾(��V������������d���7�z��;Sؽ[���d�D*�dkּ,\����'�"���R�h}����:�Z;��#;a=7;X�A;@�F;��H;��I;�I;�I;aI;�GI;"4I;T%I;�I;�I;�I;|
I;	I;|
I;�I;�I;�I;W%I;"4I;�GI;aI;�I;�I;��I;��H;;�F;U�A;a=7;��#;�Z;��:X}���R�#����'�+\��dkּD*��d�[��;Sؽz����7��d���������V���(��      �V������������Ͼ�d���ǆ�F�N��3��c�[����\�4��*C���o���	��눻𳺐��9b��:�h;v�/;e�=;jE;%3H;�WI;�I;(�I;�kI;�OI;T:I;*I;QI;�I;#I;�I;�I;�I;#I;�I;OI;*I;T:I;�OI;�kI;(�I;�I;�WI;(3H;iE;d�=;w�/;�h;`��:���9��눻��	��o�*C��4����\�[���cི3�F�N��ǆ��d����Ͼ���������      �,b�ƽ\��>M���5�=��4r��'l¾Ꝓ�%&W��3�;Sؽ�z��\G����{I����?���̻v�-��	��`��:��;��&;M|9;�C;�dG;�I;j�I;~�I;�vI;�WI;Z@I;�.I;�!I;�I;�I;I;�I;I;�I;�I;�!I;�.I;Z@I;�WI;~vI;~�I;g�I;�I;�dG;�C;L|9;��&;��;^��:�	��t�-���̻��?�{I�����\G��z��;Sؽ�3�%&W�Ꝓ�'l¾4r��=����5��>M�ƽ\�      ���&��\���O䂿Ľ\���1�����J˾Ꝓ�F�N�z��K������X�'�e�Ҽ��|��z��n��x��P�&:�P�:Ш;�W4;�@;RgF;��H;:�I;K�I;d�I;E_I;FI;73I;N%I;vI;�I;I;�I;I;�I;xI;N%I;63I;FI;E_I;`�I;K�I;9�I;��H;TgF;�@;�W4;Ш;�P�:P�&:x���n���z���|�e�ҼX�'����K���z��F�N�Ꝓ��J˾�����1�Ľ\�O䂿\���&��      !}߿�$ڿ0�ʿ����
����Ps�SX:����'l¾�ǆ���7����:5���Q�����t���75�b������ �8ʼ:��;��.;��=;�EE;�YH;�hI;O�I;�I;OfI;KKI;V7I;s(I;I;!I;�I;�I;�I;!I;I;p(I;V7I;KKI;NfI;�I;O�I;�hI;�YH;�EE;��=;��.;��;ʼ:  �8���a���75��t������Q�:5�������7��ǆ�'l¾���SX:��Ps�
�������0�ʿ�$ڿ      |�����p������ſ&���Ps���1�4r���d���d�~I�ЈŽ��}�`*�LC���^��B�c�D��E๸ �:��;�);77;;VD;p�G;uHI;؝I;؏I;�lI; PI;�:I;G+I;L I;�I;�I;]I;�I;�I;J I;D+I;�:I; PI;�lI;ԏI;؝I;tHI;o�G;WD;37;;�);��;� �:�E�c�D��B��^�LC��`*���}�ЈŽ~I��d��d��4r����1��Ps�&����ſ��꿄p����      ��7��3�آ%�|��<����ſ
���Ľ\�=����Ͼ����b�3��载z��~�9�`�Ἑ���z��7}��ct�d�^:�+�:գ#;��8;��B;KsG;�%I;ۙI; �I;.rI;BTI;>I;�-I;A"I;~I;I;�I;I;|I;A"I;�-I;>I;ATI;+rI;�I;ٙI;�%I;JsG;��B;��8;أ#;�+�:h�^:�ct��7}��z����`���9��z����b�3�������Ͼ=��Ľ\�
�����ſ�<��|�آ%��3�      0�_��+Y��lG�!f.�|���꿴���O䂿��5���󾏰��Q�N�X��T��#�Q����|����h!�~g��񳺤	:�
�:%�;l16;��A;|G;I;c�I;��I;�vI;{WI;�@I;�/I;�#I;�I;;I;�I;;I;�I;�#I;�/I;�@I;{WI;�vI;��I;a�I;I;|G;��A;h16;(�;�
�:�	: �~g���h!�|������#�Q�T��X��Q�N���������5�O䂿�������|�!f.��lG��+Y�      Ҭ��%}�?tf��lG�آ%��p�0�ʿ\����>M����W�����d�ʤ�̷�1�d��
��I���1�\�������9���:V;�U4;��@;�F;I�H;	�I;�I;�yI;�YI;qBI;1I;�$I;�I;I;�I;I;�I;�$I;1I;pBI;�YI;�yI;�I;	�I;I�H;�F;��@;�U4;X;���: ��9��\����1��I���
�1�d�̷�ʤ���d�W�������>M�\���0�ʿ�p�آ%��lG�?tf�%}�      T���E���%}��+Y��3�����$ڿ&��ƽ\����(���s��3�8����p�d�T���<<�1��X���ȗ�9z��:�;Z%3;rp@;zF;��H;&�I;!�I;�{I;|[I;�CI;�1I;�%I;UI;�I;4I;�I;WI;�%I;�1I;�CI;|[I;�{I;�I;&�I;��H;zF;rp@;X%3;�;z��:ȗ�9\���1���<<�T��d��p�8����3��s�(�����ƽ\�&���$ڿ����3��+Y�%}�E���      ����,������U���L�Q�Ǚ$�6�����>�}�J(�B�׾�T���L+���սl����L���iO���ͻe��@%m8�o�:��;d�1;��?;vF;} I;��I;��I;��I;�vI;�WI;�AI;"2I;(I;"I;  I;"I;(I;"2I;�AI;�WI;�vI;��I;��I;��I;{ I;vF;��?;`�1;��;�o�:�%m8f����ͻ�iO� L����l����ս�L+��T��B�׾J(�>�}���6���Ǚ$�L�Q�U��������,��      �,��b��$P���{���K��x �����r�����w��$���Ҿh��� (���ѽӷ��(����ޔK�:ɻ�����8���:��;��1;@;��F;8I;
�I;C�I;ϞI;�uI;]WI;�AI;�1I;�'I;�!I;�I;�!I;�'I;�1I;�AI;^WI;�uI;͞I;A�I;�I;8I;��F;@;��1;��;���:���8��:ɻޔK����(�ӷ����ѽ (�h�����Ҿ�$���w�r��������x ���K��{�$P��b��      ����$P�������d���;�$���㿴���#f�f�� ž��z���?�ƽ'0v�V5�0����o@�z���Qi�bu9tK�:L];�73;P�@;(�F;cI;��I;��I;{�I;tI;�UI;r@I;1I;'I;=!I;aI;=!I;'I;1I;p@I;�UI;tI;y�I;��I;��I;aI;(�F;P�@;�73;O];tK�: bu9Si�{����o@�0���V5�'0v�?�ƽ����z� žf��#f�������$����;���d����$P��      U����{���d��F�Ǚ$�;����ɿ0蒿��K�R���j��Zb�H�4���t�a����>�����.��d���غ���9�Y�:dX;�25;R�A;�!G;f7I;��I;|�I;v�I;�pI;�SI;�>I;�/I;�%I;T I;cI;T I;�%I;�/I;�>I;�SI;�pI;u�I;z�I;��I;f7I;�!G;P�A;�25;gX;�Y�:���9 �غ�d����.�>������t�a�4���H�Zb��j��R����K�0蒿��ɿ;��Ǚ$��F���d��{�      L�Q���K���;�Ǚ$��;
��޿�����w�t,���澟���)�D������I��&�G�����N�������������9:���:�n!;��7;�B;��G;ZI;Z�I;��I;�I;�lI;�PI;F<I;�-I;E$I;�I;�I;�I;C$I;�-I;F<I;�PI;�lI;�I;��I;Z�I;ZI;��G;�B;��7;�n!;���:��9:����������N�����&�G��I������)�D��������t,���w�����޿�;
�Ǚ$���;���K�      Ǚ$��x �$��;���޿q���˅���F��
��~����z��$���ս���B2+���ϼPp�����3�]�x�*�R��:;�;9';Ō:;*�C;:H;�}I;M�I;��I; �I;�gI;�LI;M9I;j+I;X"I;'I;\I;'I;X"I;j+I;M9I;�LI;�gI;��I;��I;N�I;�}I;9H;'�C;��:;9';;�;V��:��*�3�]�����Pp���ϼB2+������ս�$���z��~���
��F�˅��q����޿;��$���x �      6��������㿌�ɿ���˅����P�e��>�׾�`��V�H����@��T�a���̡���D��ɻ� ��ҭ�X�:�;�I-;W|=;TCE;ՅH;6�I;�I;��I;�I;�aI;THI;�5I;�(I; I;I;�I;I; I;�(I;�5I;THI;�aI;�I;��I;�I;4�I;ՅH;QCE;R|=;�I-;�;X�:`ӭ�� ��ɻ�D�̡����T�a��@����V�H��`��>�׾e����P�˅�������ɿ�㿵���      ��r�������0蒿��w��F�e��Ͱ�"����Yb�+����ѽ�%��D4�ڟ�X������G���潺(��9�r�: ;:3;JQ@;�vF;G�H;6�I;��I;��I;�zI;�ZI;ECI;�1I;�%I;vI;�I;VI;�I;vI;�%I;�1I;GCI;�ZI;�zI;��I;��I;4�I;G�H;�vF;FQ@;:3; ;�r�: ��9�潺�G�����X��ڟ�D4��%����ѽ+���Yb�"���Ͱ�e���F���w�0蒿����r���      >�}���w�#f���K�s,��
�>�׾"�����k���'�hz꽟I���;V�=M�����iO�^G�SoE�<�����:h� ;Ͽ$;ݴ8;��B;.�G;gKI;A�I;F�I;u�I;6qI;�SI;�=I;�-I;:"I;�I;JI;�I;JI;�I;:"I;�-I;�=I;�SI;6qI;q�I;F�I;@�I;eKI;+�G;�B;۴8;ο$;h� ;���:<��QoE�^G໧iO����=M��;V��I��iz���'���k�"���>�׾�
�t,���K�#f���w�      J(��$�f��R������~���`���Yb���'��U�J$��F�m�&����ϼ�/��9������^�غp9�9���:G;H.;C|=;pE;�\H;R�I;��I;��I;,�I;2gI;3LI;8I;;)I;�I;�I;�I;\I;�I;�I;�I;9)I;8I;3LI;2gI;)�I;��I;��I;R�I;�\H;mE;B|=;H.;G;���:p9�9Z�غ����9���/����ϼ&��F�m�J$���U���'��Yb��`���~�����R��f���$�      B�׾��Ҿ ž�j��������z�V�H�+��iz�J$���/v�2+�ސ�����5��ɻ4�@'�����:���:do!;:P6;8lA;�F;��H;÷I;��I;�I;}I;�\I;�DI;92I;�$I;�I;�I;�I;�I;�I;�I;�I;�$I;<2I;�DI;�\I;}}I;�I;��I;ķI;��H;�F;5lA;:P6;bo!;���:���:('��4��ɻ��5���ސ�2+��/v�J$��iz�+��V�H���z������j�� ž��Ҿ      �T��h�����z�Zb�)�D��$�����ѽ�I��F�m�2+�������F�K���z�p����Г�9vT�: 0;��-;��<;xzD;�H;�mI;�I;��I;��I;�oI;�RI;�<I;4,I;�I;AI;fI;�I;�I;�I;iI;BI;�I;7,I;�<I;�RI;�oI;ÕI;��I;�I;�mI;�H;vzD;��<;��-;�/;vT�:ؓ�9���|�p���F�K�������2+�F�m��I����ѽ���$�)�D�Zb���z�h���      �L+� (���H�������ս�@���%���;V�&��ݐ�����zMS�H����>D⺀o8Hq�:�;��$;-_7;\�A;��F;*�H;��I;��I;��I;�I;�bI;�HI;B5I;X&I;cI;tI;$I;I;=
I;I;$I;rI;aI;Y&I;B5I;�HI;�bI;�I;��I;��I;��I;$�H;��F;\�A;,_7;��$;�;Nq�:@o8:D���H��zMS�����ݐ�&���;V��%���@����ս����H��� (�      ��ս��ѽ?�ƽ3����I�����S�a�D4�<M���ϼ��F�K�H��?G��=f���o���:*C�:�Y;�1;}l>;E;0H;MqI;5�I;�I;�I;6sI;�UI;"?I;�-I;� I;�I;�I;�
I;II;kI;II;�
I;�I;�I;� I;�-I;#?I;�UI;6sI;�I; �I;2�I;JqI;0H;E;}l>;�1;�Y;.C�:��:��o�=f�>G��H��F�K�����ϼ<M�D4�S�a�����I��3���>�ƽ��ѽ      k��ҷ��&0v�t�a�%�G�A2+���ڟ�����/����5�����?f��׬�t�g:��:2�;DI-;Jg;;.OC;:SG;�I;��I;R�I;2�I;;�I;@cI;�II;�5I;�&I;�I;mI;I;�I;�I;�I;�I;�I;I;mI; I;�&I;�5I;�II;@cI;:�I;5�I;Q�I;��I;�I;:SG;-OC;Kg;;DI-;3�;��:t�g:�׬�?f�������5��/�����ڟ���A2+�%�G�t�a�&0v�ӷ��      ��'�U5���������ϼʡ��X���iO�8���ɻy�p�:D⺰�o���g:C`�:pG;�*;�9;��A;�uF;N�H;��I;��I;ܻI;|�I;�pI;kTI;�>I;Q-I;�I;�I;/I;�I;�I;�I;I;�I;�I;�I;.I;�I;�I;Q-I;�>I;kTI;�pI;}�I;ڻI;��I;�I;O�H;�uF;��A;�9;�*;nG;?`�:��g:��o�:D�|�p��ɻ9���iO�X��ʡ����ϼ������T5�(�      L�����/���=����N��Pp��D����\G�����4�����@o8��:��:nG;0�(;ɶ7;��@;��E;�QH;JmI;��I;,�I;ϢI;\}I;�^I;�FI;4I;%I;�I;�I;(
I;DI;I; I;��H; I;I;FI;'
I;�I;�I;%I;4I;�FI;�^I;\}I;ϢI;)�I;��I;ImI;�QH;��E;��@;˶7;0�(;nG;��:��:@o8 ���4�����[Gໂ���D�Pp��N��=���/������      �iO�ܔK��o@���.���������ɻ�G��JoE�T�غ'��ؓ�9Nq�:,C�:3�;�*;ɶ7;�P@;�\E;#H;JI;��I;��I;?�I;��I;shI;�NI;�:I;t*I;�I;�I;I;NI;DI;e�H;��H;�H;��H;e�H;FI;MI;I;�I;�I;p*I;�:I;�NI;vhI;��I;=�I;��I;��I;�II;#H;�\E;�P@;ƶ7;�*;3�;,C�:Hq�:ؓ�9'��X�غLoE��G���ɻ����~����.��o@�ޔK�      ��ͻ5ɻr����d�����'�]�� ��潺���9�9���:�T�:�;�Y;FI-;�9;��@;�\E;��G;g5I;�I;z�I;�I;��I;�pI;�UI;�@I;k/I;�!I;�I;zI;�I;�I;V�H;��H;O�H;��H;O�H;��H;W�H;�I;�I;zI;�I;�!I;k/I;�@I;�UI;�pI;��I;
�I;z�I;�I;h5I;��G;�\E;��@;�9;HI-;�Y;�;~T�:���:�9�9 ���潺� �$�]�����d��r���6ɻ      ^����Li��غ����x�*��ҭ���9���:���:���: 0;��$;�1;Ig;;��A;��E;"H;e5I;n�I;��I;��I;̗I;�vI;�[I;�EI;�3I;l%I;�I;�I;�	I;�I;��H;��H;]�H;!�H;��H;#�H;]�H;��H;��H;�I;�	I;�I;�I;m%I;�3I;�EI;�[I;�vI;ɗI;��I;��I;o�I;e5I;#H;��E;��A;Ig;;�1;��$; 0;���:���:���:(��9�ҭ�p�*�쓛��غJi����      �(m8 ��8�bu9x��9��9:`��:#X�:�r�:l� ;G;fo!;��-;-_7;~l>;0OC;�uF;�QH;JI;�I;��I;�I;�I;�zI;�_I;{II;�7I;�(I;�I;I;VI;I;` I;��H;��H;:�H;�H;��H;�H;:�H;��H;��H;a I;I;UI;	I;�I;�(I;�7I;{II;�_I;�zI;�I;�I;��I;�I;JI;�QH;�uF;0OC;}l>;-_7;��-;bo!;G;l� ;�r�:!X�:f��:��9:���9�bu9��8      �o�:��:�K�:�Y�:���:H�;�; ;ؿ$;	H.;BP6;��<;]�A;E;;SG;N�H;JmI;��I;{�I;��I;�I;|I;�aI;�KI;�9I;+I;�I;�I;�I;`I;'I;-�H;	�H;��H;(�H;G�H;	�H;G�H;(�H;��H;�H;-�H;'I;]I;�I;�I;�I;+I;�9I;�KI;�aI;|I;�I;��I;{�I;��I;ImI;L�H;=SG;E;\�A;��<;@P6;H.;ٿ$; ;�;I�;̨�:�Y�:�K�:��:      ��;��;U];dX;�n!;9';�I-;:3;�8;I|=;<lA;~zD;��F;0H;�I;��I;��I;��I;�I;͗I;�zI;�aI;�LI;V;I;�,I;k I;]I;/I;tI;I;��H;6�H;��H;��H;A�H;��H;\�H;��H;B�H;��H;��H;6�H;��H;I;qI;0I;[I;n I;�,I;S;I;�LI;�aI;�zI;ЗI;�I;��I;��I;�I;�I;0H;��F;}zD;;lA;F|=;�8;:3;�I-;9';�n!;dX;V];��;      |�1;��1;�73;�25;��7;Ȍ:;b|=;JQ@;��B;tE;�F;�H;'�H;PqI;��I;��I;,�I;B�I;��I;�vI;�_I;�KI;U;I;-I;$!I;SI;I;PI;�I;3�H;��H;��H;_�H;��H;��H;	�H;��H;	�H;��H;��H;\�H;��H;��H;0�H;�I;PI;I;UI;&!I;-I;S;I;�KI;�_I;�vI;��I;D�I;*�I;��I;��I;NqI;&�H;�H;�F;qE;��B;MQ@;a|=;Ɍ:;��7;�25;�73;��1;      ��?;-@;B�@;Z�A;�B;.�C;TCE;�vF;/�G;�\H;��H;�mI;��I;8�I;U�I;ݻI;֢I;��I;�pI;�[I;II;�9I;�,I;*!I;�I;�I;�I;2I;��H;��H;��H;c�H;��H;)�H;(�H;��H;i�H;��H;(�H;)�H;��H;f�H;��H;��H;��H;0I;�I;�I;�I;'!I;�,I;�9I;~II;�[I;�pI;��I;ԢI;ܻI;U�I;6�I;��I;�mI;��H;�\H;/�G;�vF;TCE;/�C;�B;Z�A;A�@;,@;      )vF;ȊF;�F;�!G;��G;8H;مH;G�H;lKI;U�I;ŷI;�I;��I;�I;4�I;z�I;^}I;shI;�UI;�EI;�7I;+I;h I;PI;�I;	I;�I;��H;)�H;�H;b�H;v�H;��H;��H;��H;R�H;#�H;R�H;��H;��H;��H;x�H;b�H;�H;(�H;��H;�I;	I;�I;PI;h I;+I;�7I;�EI;�UI;uhI;\}I;z�I;4�I; �I;��I;�I;ŷI;S�I;kKI;I�H;مH;8H;��G;�!G;�F;��F;      � I;?I;cI;p7I;ZI;�}I;=�I;4�I;G�I;��I;��I;��I;��I;�I;<�I;�pI;�^I;�NI;�@I;�3I;�(I;�I;\I;I;�I;�I;�H;^�H;�H;p�H;`�H;��H;S�H;U�H;��H;@�H;�H;@�H;��H;S�H;Q�H;��H;`�H;o�H;�H;^�H;�H;�I;�I;I;[I;�I;�(I;�3I;�@I;�NI;�^I;�pI;<�I;�I;��I;��I;��I;��I;G�I;6�I;=�I;�}I;ZI;n7I;dI;@I;      ��I;�I;��I;��I;^�I;R�I;�I;��I;N�I;��I;�I;ʕI;�I;;sI;DcI;lTI;�FI;�:I;m/I;o%I;�I;�I;2I;SI;/I;��H;]�H;4�H;}�H;`�H;��H;�H;�H;?�H;��H;;�H;*�H;<�H;��H;?�H;�H;�H;��H;]�H;{�H;5�H;]�H;��H;/I;SI;0I;�I;�I;o%I;k/I;�:I;�FI;lTI;BcI;9sI;�I;ʕI;�I;��I;P�I;��I;�I;R�I;h�I;��I;��I;"�I;      �I;E�I;��I;��I;��I;��I;��I;��I;v�I;-�I;�}I;�oI;�bI;�UI;�II;�>I;4I;q*I;�!I;�I;I;�I;rI;�I;��H;*�H;�H;}�H;g�H;��H;�H;��H;��H;6�H;��H;o�H;g�H;o�H;��H;6�H;��H;��H;�H;��H;g�H;}�H;�H;)�H;��H;�I;qI;�I;
I;�I;�!I;r*I;4I;�>I;�II;�UI;�bI;�oI;}I;-�I;v�I;��I;��I;��I;��I;��I;��I;<�I;      ��I;ڞI;��I;|�I;��I;
�I;�I;�zI;BqI;=gI;�\I;�RI;�HI;,?I;�5I;U-I;%I;�I;�I;�I;WI;_I;I;2�H;��H;�H;m�H;^�H;��H;�H;��H;��H;��H;Z�H;��H;��H;��H;��H;��H;Z�H;��H;��H;��H; �H;��H;^�H;l�H; �H;��H;3�H;�I;_I;VI;�I;�I;�I;%I;U-I;�5I;*?I;�HI;�RI;�\I;;gI;BqI;�zI;�I;�I;�I;}�I;��I;ڞI;      �vI;�uI;tI;�pI;�lI;�gI;�aI;[I;�SI;<LI;�DI;�<I;J5I;�-I;�&I;�I;�I;�I;~I;�	I;'I;*I;��H;��H;��H;c�H;]�H;��H;�H;��H;��H;��H;&�H;��H;G�H;�H;��H;�H;G�H;��H;#�H;��H;��H;��H;�H;��H;]�H;b�H;��H;��H;��H;(I;!I;�	I;~I;�I;�I;�I;�&I;�-I;I5I;�<I;�DI;>LI;�SI;[I;�aI;�gI;�lI;�pI;tI;�uI;      �WI;nWI;VI;�SI;�PI;�LI;XHI;OCI;�=I;8I;A2I;B,I;_&I;� I;	I;�I;�I;I;�I;�I;i I;1�H;9�H;��H;b�H;v�H;��H;�H;��H;��H;��H;"�H;��H;�H;��H;��H;��H;��H;��H;�H;}�H;#�H;��H;��H;��H;�H;��H;u�H;e�H;��H;6�H;1�H;e I;�I;�I;I;�I;�I;	I;� I;]&I;A,I;A2I;8I;�=I;OCI;WHI;�LI;�PI;�SI;VI;jWI;      BI;�AI;|@I;�>I;S<I;P9I;�5I;�1I;�-I;<)I;�$I; I;gI;�I;rI;3I;0
I;KI;�I;��H;��H;	�H;��H;b�H;��H;��H;V�H;�H;��H;��H;'�H;��H;��H;��H;G�H;�H;%�H;�H;G�H;��H;��H;��H;'�H;��H;��H;�H;Q�H;��H;��H;b�H;��H;	�H;��H;��H;�I;MI;.
I;3I;qI;�I;eI;�I;�$I;=)I;�-I;�1I;�5I;Q9I;L<I;�>I;|@I;�AI;      32I;�1I;1I;�/I;�-I;h+I;�(I;�%I;C"I;�I;�I;LI;xI;�I;I;�I;PI;GI;^�H;��H;��H;��H;��H;��H;%�H;��H;P�H;=�H;5�H;X�H;��H;�H;��H;.�H;�H;��H;��H;��H;�H;.�H;��H;�H;��H;Z�H;6�H;=�H;P�H;��H;(�H;��H;��H;��H;��H;��H;^�H;HI;NI;�I;I;�I;xI;LI;�I;�I;D"I;�%I;�(I;m+I;�-I;�/I;1I;�1I;      (I;�'I;"'I;�%I;]$I;U"I; I;~I;�I;�I;�I;vI;+I; I;�I;�I; I;e�H;��H;d�H;C�H;+�H;B�H;��H;!�H;��H;��H;��H;��H;��H;H�H;��H;G�H;�H;��H;��H;��H;��H;��H;�H;D�H;��H;H�H;��H;��H;��H;��H;��H;!�H;��H;A�H;+�H;A�H;d�H;��H;e�H;I;�I;�I; I;+I;vI;�I;�I;�I;~I; I;X"I;S$I;�%I;"'I;�'I;      "I;�!I;I!I;[ I;I;&I;I;�I;YI;�I;�I;�I;I;TI;�I;�I;* I;��H;U�H;(�H;&�H;I�H;��H;�H;��H;P�H;@�H;;�H;r�H;��H;�H;��H;�H;��H;��H;j�H;e�H;j�H;��H;��H;�H;��H;�H;��H;s�H;;�H;?�H;O�H;��H;�H;��H;I�H;%�H;*�H;U�H;��H;' I;�I;�I;SI;I;�I;�I;�I;YI;�I;I;*I;�I;Z I;I!I;�!I;      " I; I;oI;jI;I;ZI;�I;]I;�I;\I;�I;I;A
I;tI;�I;I;��H;�H;��H;��H;��H;�H;\�H;��H;e�H;!�H;�H;.�H;i�H;��H;��H;��H;'�H;��H;��H;f�H;L�H;f�H;��H;��H;"�H;��H;��H;��H;l�H;.�H;�H;"�H;e�H;��H;\�H;�H;��H;��H;��H;�H;��H;I;�I;tI;A
I;I;�I;_I;�I;]I;�I;`I;�I;jI;oI; I;      "I;�!I;I!I;Z I;I;&I;I;�I;[I;�I;�I;�I;I;TI;�I;�I;* I;��H;U�H;(�H;(�H;I�H;��H;�H;��H;P�H;@�H;;�H;r�H;��H;�H;��H;�H;��H;��H;j�H;e�H;j�H;��H;��H;�H;��H;�H;��H;s�H;;�H;=�H;O�H;��H;�H;��H;I�H;%�H;*�H;U�H;��H;' I;�I;�I;SI;I;�I;�I;�I;YI;�I;I;*I;�I;[ I;F!I;�!I;      (I;�'I;!'I;�%I;]$I;U"I; I;~I;�I;�I;�I;vI;+I; I;�I;�I; I;e�H;��H;d�H;E�H;+�H;B�H;��H;!�H;��H;��H;��H;��H;��H;H�H;��H;G�H;�H;��H;��H;��H;��H;��H;�H;D�H;��H;H�H;��H;��H;��H;��H;��H;!�H;��H;A�H;+�H;A�H;d�H;��H;e�H;I;�I;�I; I;+I;vI;�I;�I;�I;~I; I;X"I;S$I;�%I;!'I;�'I;      52I;�1I;1I;�/I;�-I;h+I;�(I;�%I;C"I;�I;�I;LI;xI;�I;I;�I;PI;GI;^�H;��H;��H;��H;��H;��H;(�H;��H;P�H;=�H;5�H;X�H;��H;�H;��H;.�H;�H;��H;��H;��H;�H;.�H;��H;�H;��H;Z�H;8�H;=�H;P�H;��H;%�H;��H;��H;��H;��H;��H;^�H;HI;NI;�I;I;�I;xI;LI;�I;�I;D"I;�%I;�(I;m+I;�-I;�/I;1I;�1I;      BI;�AI;}@I;�>I;Q<I;N9I;�5I;�1I;�-I;<)I;�$I;�I;eI;�I;qI;3I;0
I;KI;�I;��H;��H;	�H;��H;b�H;��H;��H;T�H;�H;��H;��H;'�H;��H;��H;��H;G�H;�H;%�H;�H;G�H;��H;��H;��H;'�H;��H;��H;�H;Q�H;��H;��H;a�H;��H;	�H;��H;��H;�I;KI;.
I;3I;rI;�I;eI; I;�$I;=)I;�-I;�1I;�5I;Q9I;L<I;�>I;|@I;�AI;      �WI;nWI;	VI;�SI;�PI;�LI;ZHI;OCI;�=I;8I;A2I;A,I;]&I;� I;	I;�I;�I;I;�I;�I;k I;1�H;9�H;��H;e�H;v�H;��H;�H;��H;��H;��H;"�H;�H;�H;��H;��H;��H;��H;��H;�H;}�H;#�H;��H;��H;��H;�H;��H;u�H;b�H;��H;7�H;1�H;g I;�I;�I;I;�I;�I;	I;� I;_&I;B,I;A2I; 8I;�=I;OCI;ZHI;�LI;�PI;�SI;	VI;kWI;      �vI;�uI;tI;�pI;�lI;�gI;�aI; [I;�SI;<LI;�DI;�<I;I5I;�-I;�&I;�I;�I;�I;~I;�	I;'I;(I;��H;��H;��H;c�H;]�H;��H;�H;��H;��H;��H;%�H;��H;G�H;�H;��H;�H;G�H;��H;#�H;��H;��H;��H;�H;��H;]�H;b�H;��H;��H;��H;*I;#I;�	I;~I;�I;�I;�I;�&I;�-I;J5I;�<I;�DI;>LI;�SI;[I;�aI;�gI;�lI;�pI;tI;�uI;      ��I;ڞI;��I;|�I;�I;�I;�I;�zI;CqI;:gI;�\I;�RI;�HI;,?I;�5I;U-I;%I;�I;�I;�I;ZI;_I;I;2�H;��H;�H;m�H;^�H;��H;�H;��H;��H;��H;X�H;��H;��H;��H;��H;��H;Z�H;��H;��H;��H; �H;��H;^�H;l�H; �H;��H;3�H;I;_I;VI;�I;�I;�I;%I;W-I;�5I;,?I;�HI;�RI;�\I;;gI;CqI;�zI;�I;
�I;�I;|�I;��I;ݞI;      ��I;A�I;��I;��I;��I;��I;��I;��I;v�I;-�I;�}I;�oI;�bI;�UI;�II;�>I;4I;r*I;�!I;�I;I;�I;tI;�I;��H;*�H;�H;}�H;g�H;��H;�H;��H;��H;6�H;��H;o�H;g�H;o�H;��H;6�H;��H;��H;�H;��H;g�H;}�H;�H;)�H;��H;�I;qI;�I;
I;�I;�!I;r*I;4I;�>I;�II;�UI;�bI;�oI;�}I;,�I;x�I;¤I;��I;��I;��I;��I;��I;C�I;      ��I;�I;��I;��I;\�I;R�I;�I;��I;N�I;��I;�I;ʕI;�I;:sI;DcI;lTI;�FI;�:I;k/I;o%I;�I;�I;2I;SI;/I;��H;]�H;5�H;}�H;`�H;��H;�H;�H;=�H;��H;;�H;*�H;<�H;��H;?�H;�H;�H;��H;]�H;{�H;4�H;]�H;��H;/I;SI;0I;�I;�I;o%I;m/I;�:I;�FI;nTI;DcI;:sI;�I;˕I;�I;��I;N�I;��I;�I;O�I;j�I;��I;��I;"�I;      � I;=I;fI;j7I;ZI;�}I;;�I;4�I;G�I;��I;��I;��I;��I;�I;<�I;�pI;�^I;�NI;�@I;�3I;�(I;�I;\I;I;�I;�I;�H;^�H;�H;p�H;`�H;��H;S�H;S�H;��H;@�H;�H;?�H;��H;S�H;Q�H;��H;`�H;o�H;�H;^�H;�H;�I;�I;I;[I;�I;�(I;�3I;�@I;�NI;�^I;�pI;<�I;�I;��I;��I;��I;��I;E�I;4�I;;�I;�}I;ZI;j7I;dI;5I;      .vF;ÊF;*�F;�!G;��G;9H;مH;G�H;kKI;U�I;ŷI;�I;��I; �I;2�I;z�I;^}I;uhI;�UI;�EI;�7I;+I;h I;PI;�I;	I;�I;��H;)�H;�H;b�H;v�H;��H;��H;��H;R�H;#�H;R�H;��H;��H;��H;x�H;b�H;�H;(�H;��H;�I;	I;�I;PI;h I;+I;7I;�EI;�UI;uhI;\}I;z�I;4�I; �I;��I;�I;ŷI;R�I;iKI;G�H;܅H;8H;��G;�!G;(�F;��F;      ��?;-@;B�@;Z�A;�B;.�C;TCE;�vF;/�G;�\H;��H;�mI;��I;6�I;U�I;ݻI;բI;��I;�pI;�[I;�II;�9I;�,I;*!I;�I;�I;�I;0I;��H;��H;��H;e�H;��H;)�H;'�H;��H;i�H;��H;(�H;(�H;��H;f�H;��H;��H;��H;2I;�I;�I;�I;(!I;�,I;�9I;}II;�[I;�pI;��I;ԢI;ݻI;U�I;6�I;��I;�mI;��H;�\H;.�G;�vF;TCE;.�C;�B;Z�A;A�@;-@;      ��1;��1;�73;�25;��7;͌:;^|=;KQ@;��B;tE;�F;�H;(�H;NqI;��I;��I;,�I;B�I;��I;�vI;�_I;�KI;V;I;-I;&!I;UI;I;PI;�I;3�H;��H;��H;^�H;��H;��H;	�H;��H;	�H;��H;��H;^�H;��H;��H;0�H;�I;PI;I;SI;$!I;	-I;S;I;�KI;�_I;�vI;��I;D�I;*�I;��I;��I;QqI;'�H;�H;�F;qE;��B;KQ@;^|=;͌:;��7;�25;�73;��1;      ��;��;f];dX;�n!;9';�I-;:3;�8;G|=;;lA;}zD;��F;0H;�I;��I;��I;��I;�I;͗I;�zI;�aI;�LI;V;I;�,I;l I;\I;0I;tI;I;��H;6�H;��H;��H;B�H;��H;\�H;��H;A�H;��H;��H;6�H;��H;I;qI;/I;YI;l I;�,I;S;I;�LI;�aI;�zI;ЗI;�I;��I;��I;��I;�I;0H;��F;}zD;=lA;G|=;�8;:3;�I-;9';�n!;fX;[];��;      �o�:��:�K�:�Y�:���:H�;�; ;ؿ$;H.;BP6;��<;\�A;E;;SG;N�H;ImI;��I;{�I;��I;�I;|I;�aI;�KI;�9I;+I;�I;�I;�I;bI;'I;-�H;�H;��H;(�H;G�H;	�H;G�H;(�H;��H;�H;-�H;'I;]I;�I;�I;�I;+I;�9I;�KI;�aI;|I;�I;��I;{�I;��I;ImI;N�H;=SG;E;]�A;��<;@P6;	H.;ؿ$; ;�;H�;̨�:�Y�:�K�:��:      �&m8@��8�bu9���9��9:R��:'X�:�r�:l� ;G;do!;��-;-_7;}l>;0OC;�uF;�QH;JI;�I;��I;�I;�I;�zI;�_I;{II;�7I;�(I;�I;I;VI;I;` I;��H;��H;:�H;�H;��H;�H;:�H;��H;��H;a I;I;SI;	I;�I;�(I;�7I;{II;�_I;�zI;�I;�I;��I;�I;JI;�QH;�uF;0OC;~l>;-_7;��-;fo!;G;n� ;�r�:'X�:f��:�9:���9�bu9��8      _����Hi��غ����t�*��ҭ� ��9���:���:���: 0;��$;�1;Gg;;��A;��E;"H;e5I;n�I;��I;��I;͗I;�vI;�[I;�EI;�3I;m%I;�I;�I;�	I;�I;��H;��H;]�H;#�H;��H;#�H;]�H;��H;��H;�I;�	I;�I;�I;l%I;�3I;�EI;�[I;�vI;ɗI;��I;��I;o�I;e5I;#H;��E;��A;Ig;;�1;��$; 0;���:���:���:8��9�ҭ�p�*�쓛��غJi����      ��ͻ5ɻr����d�����)�]�� ��潺 ���9�9���:~T�:�;�Y;FI-;�9;��@;�\E;��G;g5I;�I;z�I;�I;��I;�pI;�UI;�@I;k/I;�!I;�I;zI;�I;�I;W�H;��H;O�H;��H;O�H;��H;V�H;�I;�I;zI;�I;�!I;k/I;�@I;�UI;�pI;��I;�I;z�I;�I;h5I;��G;�\E;��@;�9;HI-;�Y;�;�T�:���:�9�9���潺� �"�]�����d��r���6ɻ      �iO�۔K��o@���.���������ɻ�G��LoE�Z�غ'��ؓ�9Hq�:*C�:3�;�*;ɶ7;�P@;�\E;"H; JI;��I;��I;A�I;��I;uhI;�NI;�:I;r*I;�I;�I;I;NI;FI;e�H;��H;�H;��H;e�H;DI;MI;I;�I;�I;q*I;�:I;�NI;vhI;��I;:�I;��I;��I;�II;$H;�\E;�P@;ȶ7;�*;3�;,C�:Nq�:ؓ�9'��T�غLoE��G���ɻ����~����.��o@�ޔK�      L�����/���=����N��Pp��D����\G�����4� ���@o8��:��:nG;1�(;ȶ7;��@;��E;�QH;ImI;��I;-�I;ϢI;[}I;�^I;�FI;4I;%I;�I;�I;(
I;FI;I; I;��H; I;I;FI;'
I;�I;�I;%I;4I;�FI;�^I;^}I;ϢI;'�I;��I;JmI;QH;��E;��@;̶7;0�(;nG;��:��:@o8����4�����[Gໂ���D�Pp��N��=���/������      ��'�U5���������ϼʡ��X���iO�8���ɻ|�p�:D���o���g:?`�:pG;�*;�9;��A;�uF;O�H;��I;��I;ڻI;|�I;�pI;kTI;�>I;Q-I;�I;�I;/I;�I;�I;�I;I;�I;�I;�I;.I;�I;�I;Q-I;�>I;kTI;�pI;}�I;ܻI;��I;�I;N�H;�uF;��A;�9;�*;oG;C`�:��g:��o�:D�y�p��ɻ8���iO�X��ʡ����ϼ������U5�(�      k��ӷ��&0v�t�a�%�G�A2+���ڟ�����/����5�����?f��׬�t�g:��:0�;DI-;Jg;;-OC;:SG;�I;��I;Q�I;4�I;;�I;@cI;�II;�5I;�&I;�I;nI;I;�I;�I;�I;�I;�I;I;mI;I;�&I;�5I;�II;@cI;:�I;4�I;R�I;��I;�I;:SG;-OC;Kg;;DI-;5�;��:t�g:�׬�=f�������5��/�����ڟ���A2+�%�G�t�a�&0v�ӷ��      ��ս��ѽ>�ƽ4����I�����S�a�D4�<M���ϼ��F�K�H��?G��=f���o���:,C�:�Y;�1;{l>;E;0H;NqI;2�I;�I;�I;6sI;�UI;"?I;�-I;� I;�I;�I;�
I;II;kI;II;�
I;�I;�I;� I;�-I;"?I;�UI;6sI;�I;�I;5�I;JqI;0H;E;}l>;�1;�Y;.C�:��:��o�=f�>G��H��F�K�����ϼ<M�D4�S�a�����I��3���>�ƽ��ѽ      �L+� (���H�������ս�@���%���;V�&��ݐ�����zMS�H����>D��o8Lq�:�;��$;+_7;\�A;��F;(�H;��I;��I;��I;�I;�bI;�HI;B5I;X&I;aI;rI;$I;I;=
I;I;$I;tI;aI;X&I;B5I;�HI;�bI;�I;��I;��I;��I;#�H;��F;\�A;,_7;��$;�;Pq�:�o8>D���G��zMS�����ݐ�&���;V��%���@����ս����H��� (�      �T��h�����z�Zb�)�D��$�����ѽ�I��F�m�2+�������F�K���|�p����Г�9vT�:�/;��-;��<;xzD;�H;�mI;�I;��I;ÕI;�oI;�RI;�<I;4,I;�I;DI;iI;�I;�I;�I;fI;AI;�I;5,I;�<I;�RI;�oI;��I;��I;�I;�mI;�H;vzD;��<;��-; 0;vT�:��9���}�p���F�K�������2+�F�m��I����ѽ���$�)�D�Zb���z�h���      B�׾��Ҿ ž�j��������z�V�H�+��iz�J$���/v�2+�ސ�����5��ɻ4�0'�����:���:`o!;:P6;8lA;�F;��H;ķI;��I;�I;}I;�\I;�DI;92I;�$I;�I;�I;�I;�I;�I;�I;�I;�$I;:2I;�DI;�\I;}}I;�I;��I;÷I;��H;	�F;6lA;:P6;bo!;���:���:('��4��ɻ��5���ސ�2+��/v�J$��hz�+��V�H���z������j�� ž��Ҿ      J(��$�f��R������~���`���Yb���'��U�J$��F�m�&����ϼ�/��9������^�غp9�9���:G;H.;C|=;qE;�\H;S�I;��I;��I;,�I;2gI;3LI;8I;;)I;�I;�I;�I;\I;�I;�I;�I;9)I;8I;3LI;2gI;)�I;��I;��I;R�I;�\H;mE;B|=;H.;G;���:p9�9X�غ����9���/����ϼ&��F�m�J$���U���'��Yb��`���~�����R��f���$�      >�}���w�#f���K�s,��
�>�׾"�����k���'�hz꽟I���;V�=M�����iO�^G�QoE�<�����:f� ;ο$;ݴ8;��B;+�G;gKI;B�I;F�I;s�I;5qI;�SI;�=I;�-I;:"I;�I;JI;�I;JI;�I;:"I;�-I;�=I;�SI;5qI;r�I;F�I;@�I;gKI;.�G;��B;۴8;Ͽ$;h� ;���:<��PoE�`G໧iO����=M��;V��I��iz���'���k�"���>�׾�
�t,���K�#f���w�      ��r�������0蒿��w��F�e��Ͱ�"����Yb�+����ѽ�%��D4�ڟ�X������G���潺(��9�r�: ;:3;HQ@;�vF;I�H;6�I;��I;��I;�zI;�ZI;ECI;�1I;�%I;wI;�I;VI;�I;vI;�%I;�1I;DCI;�ZI;�zI;��I;��I;4�I;F�H;�vF;FQ@;:3; ;�r�:��9�潺�G�����X��ڟ�D4��%����ѽ+���Yb�"���Ͱ�e���F���w�0蒿����r���      6��������㿌�ɿ���˅����P�e��>�׾�`��V�H����@��T�a���̡���D��ɻ� �@ӭ�X�:�;�I-;W|=;QCE;ׅH;4�I;�I;��I;�I;�aI;THI;�5I;�(I; I;I;�I;I; I;�(I;�5I;SHI;�aI;�I;��I;�I;4�I;ՅH;TCE;T|=;�I-;�;X�:@ӭ�� ��ɻ�D�̡����T�a��@����V�H��`��>�׾e����P�˅�������ɿ�㿵���      Ǚ$��x �$��;���޿q���˅���F��
��~����z��$���ս���B2+���ϼPp�����3�]���*�N��:;�;
9';Ō:;'�C;:H;�}I;N�I;��I;�I;�gI;�LI;M9I;j+I;X"I;'I;\I;(I;X"I;j+I;L9I;�LI;�gI;��I;��I;M�I;�}I;9H;*�C;��:;9';;�;V��:��*�3�]�����Pp���ϼB2+������ս�$���z��~���
��F�˅��q����޿;��$���x �      L�Q���K���;�Ǚ$��;
��޿�����w�t,���澟���)�D������I��&�G�����N�������������9:���:�n!;��7;�B;��G;ZI;Z�I;��I;�I;�lI;�PI;F<I;�-I;E$I;�I;�I;�I;C$I;�-I;E<I;�PI;�lI;�I;��I;Z�I;ZI;��G;�B;��7;�n!;���:��9:����������N�����&�G��I������)�D��������t,���w�����޿�;
�Ǚ$���;���K�      U����{���d��F�Ǚ$�;����ɿ0蒿��K�R���j��Zb�H�4���t�a����>�����.��d���غ���9�Y�:dX;�25;P�A;�!G;f7I;��I;|�I;w�I;�pI;�SI;�>I;�/I;�%I;T I;cI;T I;�%I;�/I;�>I;�SI;�pI;u�I;z�I;��I;f7I;�!G;R�A;�25;gX;�Y�:���9 �غ�d����.�>������t�a�4���H�Zb��j��R����K�0蒿��ɿ;��Ǚ$��F���d��{�      ����$P�������d���;�$���㿴���#f�f�� ž��z���?�ƽ'0v�V5�0����o@�{���Si��au9tK�:L];�73;P�@;(�F;cI;��I;��I;{�I;tI;�UI;r@I;1I;'I;=!I;aI;=!I;'I;1I;p@I;�UI;tI;y�I;��I;��I;aI;(�F;P�@;�73;O];tK�:bu9Si�z����o@�0���V5�'0v�?�ƽ����z� žf��#f�������$����;���d����$P��      �,��b��$P���{���K��x �����r�����w��$���Ҿh��� (���ѽӷ��(����ޔK�:ɻ�����8���:��;��1;@;��F;8I;�I;C�I;ОI;�uI;]WI;�AI;�1I;�'I;�!I;�I;�!I;�'I;�1I;�AI;^WI;�uI;͞I;A�I;
�I;6I;��F;@;��1;��;���:���8��:ɻޔK����(�ӷ����ѽ (�h�����Ҿ�$���w�r��������x ���K��{�$P��b��      E(��r'���o��O�d��X1��x�Ŀ����3�y���x����4�n��[+���'���ü4yY��kٻ�o&���p�}��:t;��0;��?;�F;� I;-�I;��I;S�I;��I;�dI;�KI;�9I;�.I;�'I;�%I;�'I;�.I;�9I;�KI;�dI;��I;Q�I;��I;-�I; I;�F;��?;��0;v;}��:@�p��o&��kٻ4yY���ü�'�[+��n�ཿ�4��x��y���3����Ŀ�x��X1�d�O��o��r'��      r'���X��g^�������]]���,�Q9�7g��U�����/����o��i1��hܽ���-$�_l���|U�Z�ԻV!� �,���:;�51;��?;|�F;Z'I;��I;H�I;d�I;цI;
dI;oKI;�9I;X.I;�'I;�%I;�'I;X.I;�9I;nKI;dI;цI;b�I;E�I;��I;Z'I;|�F;��?;�51;;��: �,�W!�Z�Ի�|U�_l���-$����hܽi1��o���ྜ�/�U���7g��Q9���,��]]�����g^���X��      �o��g^���ē��4z�6K�i��T��(ﱿV�v��X#���Ѿń�	�&�s�нd̀�`��t���F�I��ǻ�4��#9�:l�;4�2;��@;�F;;I; �I;,�I;ŲI;��I;�bI;.JI;�8I;�-I;�&I;%I;�&I;�-I;�8I;,JI;�bI;��I;²I;+�I; �I;;I;�F;��@;0�2;o�;�:�#9�4��ǻF�I�u���`��d̀�s�н	�&�ń���Ѿ�X#�V�v�(ﱿT��i��6K��4z��ē�g^��      O������4z���V��X1��<�uؿ����RZ��	�*���LUo����`y��/l�[��R��=�7�������Ƴ9:��:�;q�4;�tA;�2G;�XI;��I;��I;3�I;'�I;�_I;,HI;U7I;0,I;�%I;�#I;�%I;0,I;V7I;*HI;�_I;'�I;2�I;��I;��I;�XI;�2G;�tA;l�4;�;:��:�Ƴ9������=�7��R��[�0l�`y�����LUo�*����	��RZ����uؿ�<��X1���V��4z�����      d��]]�6K��X1�[f��pQ��U���]58��A���נ���O���a什�Q����>ߓ��� ��V��*氺p�":��:: ;17;6�B;p�G;|I;�I;��I;�I;l|I;k\I;{EI;N5I;j*I;a$I;]"I;a$I;i*I;P5I;zEI;k\I;l|I;ߧI;��I;�I;|I;n�G;6�B;17;< ;��:t�":,氺�V���� �>ߓ�����Q�a什����O��נ��A��]58�U���pQ���[f��X1�6K��]]�      �X1���,�i���<��7g��f_���U�ς�،Ⱦ
ń�,�-�k��R ��'�2�
?ټ^�{��!��n�p�O��u:Q ;�&;K#:;r�C;1&H;?�I;S�I;��I;�I;�vI;XI; BI;�2I;F(I;t"I;� I;t"I;F(I;�2I; BI;XI;�vI;
�I;��I;S�I;=�I;0&H;o�C;D#:;�&;Q ;�u:t�O��n��!�_�{�
?ټ'�2�R ��k��,�-�
ń�،Ⱦς��U�f_��7g��<�i����,�      �x�Q9�T��uؿpQ��g_��8�_��X#�s���f��<�S�{�����l�C�w���M���Ի��+�P:T���:�e;�\,;0=;�BE;��H;��I;�I;��I;�I;�oI;�RI;F>I;�/I;�%I;% I;xI;% I;�%I;�/I;D>I;�RI;�oI;�I;��I;�I;��I;��H;�BE;0=;�\,;�e;��:p:T���+���Ի�M�w��C�l�����{�<�S��f��s���X#�8�_�g_��pQ��uؿT��Q9�      Ŀ7g��(ﱿ���U����U��X#�w��f���KUo�	�#��hܽ����n<����:����� ��᝻��Ժv�9���:�V;��2;� @;��F;I;)�I;p�I;^�I;��I;3hI;@MI;�9I;",I;�"I;�I;�I;�I;�"I;",I;�9I;BMI;3hI;��I;[�I;p�I;'�I;I;��F;� @;��2;�V;���:�u�9��Ժ�᝻�� �:�������n<�����hܽ	�#�KUo�f���w���X#��U�U������(ﱿ7g��      ���U���V�v��RZ�]58�ς�s��f���ioy�`1�bO��]什�`�O�����kyY���t�T�|�1�<�u:P��:p#;C98;3�B;��G;%mI;>�I;/�I;`�I;��I;`I;6GI;'5I;X(I;�I;�I;@I;�I;�I;Z(I;'5I;4GI;`I;��I;]�I;/�I;;�I;%mI;��G;0�B;A98;p#;P��:4�u:|�1�t�T���kyY����O���`�]什bO��`1�ioy�f���s��ς�]58��RZ�V�v�U���      �3���/��X#��	��A��،Ⱦ�f��KUo�`1�ΰ��~n��ռx��'��>ټ�@���k�����Ҵ�P�39�#�:WR;6e-;�/=;�	E;�xH;��I;@�I;��I;5�I;CvI;�WI;�@I;'0I;W$I;sI;�I;kI;�I;sI;X$I;'0I;�@I;�WI;DvI;2�I;��I;?�I;��I;�xH;�	E;�/=;6e-;WR;�#�:0�39δ𺿼���k��@���>ټ�'�ռx�~n��ΰ��`1�KUo��f��،Ⱦ�A���	��X#���/�      y���྅�Ѿ*����נ�
ń�<�S�	�#�bO��~n��K̀���2����}�>��Իk�B�,#��m:0H�:� ;Ƽ5;�FA;��F;�I;��I;��I;ԾI;��I;�jI;�NI;A:I;+I;. I;I;�I;�I;�I;I;0 I;+I;D:I;�NI;�jI;��I;־I;��I;��I;�I;��F;�FA;ȼ5;� ;,H�:�m:(#�l�B��Ի~�>�������2�K̀�~n��bO��	�#�<�S�
ń��נ�*�����Ѿ��      �x���o��ń�LUo���O�,�-�{��hܽ]什ռx���2�tb��TR��Q|U�N2��*���鰺�v�9�:=D;��,;�h<;�rD;|%H;��I;��I;�I;8�I;>�I;_I;<FI;�3I;�%I;I;�I;�I;lI;�I;�I;I;�%I;�3I;=FI;_I;;�I;8�I;�I;��I;��I;y%H;�rD;�h<;��,;<D;�:�v�9�鰺*��N2��R|U�TR��tb����2�ռx�]什�hܽ{�,�-���O�LUo�ń��o��      ��4�i1��&������k�ཇ�������`��'���TR��@�]�x��V���X��@>o����:��;X#;F�6;�tA;��F;�	I;��I;�I;��I;L�I;qI;�SI;�=I;�,I;� I;�I;�I;xI;sI;zI;�I;�I;� I;�,I;�=I;�SI;qI;L�I;��I;�I;��I;�	I;��F;�tA;F�6;Z#;��;���:�>o��X��V��y��@�]�TR����'��`��������k��������&�i1�      m�ེhܽr�н_y��a什R ��l��n<�N���>ټ��P|U�x������f1�x�����u:�l�:4�;�71;�)>;�	E;@JH;��I;��I;��I;�I;�I;�bI;�HI;^5I;�&I;�I;�I;tI;WI;U
I;WI;tI;�I;�I;�&I;^5I;�HI;�bI;�I;�I;��I;��I;��I;=JH;�	E;�)>;�71;4�;�l�:x�u:����d1�����z��P|U����>ټN���n<�l�R ��a什_y��r�н�hܽ      Z+����d̀�/l��Q�&�2�C��������@��}�>�N2��V��g1�p��$R:���:;�\,;l;;<C;�eG;�9I;��I;i�I;��I;u�I;�qI;�TI;�>I;o-I;b I;�I;�I;I;HI;GI;HI;I;�I;�I;g I;o-I;�>I;�TI;�qI;s�I;�I;h�I;��I;�9I;�eG;<C;l;;�\,;;���:�$R:p��g1�V��N2��}�>��@��������C�&�2��Q�/l�d̀���      �'��-$�`��Z����	?ټw��:���hyY��k��Ի*���X�������$R:��:�R;�);�8;��A;��F;h�H;^�I;��I;��I;�I;=�I;aI;*HI;�4I;�%I;|I;I;�I;�I;GI;~I;II;�I;�I;I;~I;�%I;�4I;%HI;aI;;�I;�I;��I;��I;Z�I;f�H;��F;��A;�8;�);�R;��:�$R:x����X��*���Ի�k�iyY�:���w��?ټ���Z�_���-$�      ��ü\l��t����R��=ߓ�\�{��M��� ��컻���e�B��鰺�=o���u:���:�R;^�';B17;�@;1�E;�lH;d�I;��I;��I;@�I;��I; mI;�QI;a<I;�+I;�I;�I;�I;I;|I;`I;�I;`I;zI;I;�I;�I;�I;�+I;]<I;�QI;�lI;��I;?�I;��I;��I;d�I;�lH;1�E;�@;E17;^�';�R;���:��u:@>o��鰺g�B������컆� ��M�\�{�=ߓ��R��t���^l��      4yY��|U�D�I�;�7��� ��!���Ի�᝻n�T�ƴ�#��v�9���:�l�:;�);B17;[ @;m]E;�$H;�kI;?�I;��I;-�I;d�I;�wI;�ZI;�CI;�1I;�#I;`I;�I;f	I;�I;oI;��H;7�H;��H;oI;�I;f	I;�I;`I;�#I;�1I;�CI;�ZI;�wI;d�I;(�I;��I;?�I;�kI;�$H;k]E;] @;?17;�);;�l�:���:�v�9#�δ�o�T��᝻��Ի�!��� �;�7�D�I��|U�      �kٻV�Իwǻ ����V���n���+���ԺT�1���39�m:�:��;8�;�\,;�8;�@;m]E;�
H;�VI;��I;#�I;'�I;��I;;�I;�bI;�JI;]7I;(I;�I;gI;I;sI;pI;��H;�H;��H;�H;��H;pI;pI;I;gI;�I;
(I;]7I;�JI;�bI;;�I;��I;"�I;"�I;��I;�VI;�
H;n]E;�@;�8;�\,;8�;��;�:�m:��39T�1���Ժ��+��n��V�����wǻV�Ի      �o&�?!��4����$氺l�O� :T��u�9H�u:$�:2H�:=D;X#;�71;j;;��A;.�E;�$H;�VI;F�I;��I;K�I;��I;3�I;GiI;dPI;X<I;0,I;WI;�I;�I;�I;�I;i�H;
�H;��H;@�H;��H;
�H;j�H;�I;�I;�I;�I;SI;0,I;V<I;aPI;GiI;.�I;��I;K�I;��I;F�I;VI;�$H;.�E;��A;i;;�71;X#;<D;2H�:$�:<�u:v�90:T�`�O�氺���4�H!�      ��p� �,��$9�Ƴ9p�":<�u:��:���:X��:[R;� ;��,;H�6;�)>;<C;��F;�lH;�kI;��I;��I;��I;P�I;��I;�mI;�TI;b@I;�/I;\"I;�I;�I;I;�I;��H;��H;��H;��H;�H;��H;��H;��H;��H;�I;I;�I;�I;\"I;�/I;b@I;�TI;�mI;��I;P�I;��I;��I;��I;�kI;�lH;��F;<C;�)>;F�6;��,;� ;XR;X��:���:��:H�u:t�":�Ƴ9�$9 �,�      ���:��:I�:8��:��:"Q ;�e;�V;z#;:e-;ͼ5;�h<;�tA;�	E;�eG;f�H;e�I;?�I;#�I;L�I;O�I;/�I;ApI;�WI;)CI;{2I;�$I;�I;�I;	I;�I;2�H;��H;;�H;��H;g�H;	�H;g�H;��H;;�H;��H;3�H;�I;{	I;�I;�I;�$I;|2I;*CI;WI;<pI;.�I;L�I;N�I;#�I;A�I;c�I;d�H;�eG;�	E;�tA;�h<;˼5;8e-;z#;�V;�e;"Q ;E��:8��:I�:��:      �;;v�;�;6 ;&;�\,;�2;M98;�/=;�FA;�rD;��F;DJH;�9I;]�I;��I;��I;'�I;��I;��I;BpI;�XI;�DI;#4I;�&I;]I;"I;�
I;�I;��H;��H;$�H;�H;q�H;~�H;F�H;~�H;s�H;�H;#�H;��H;��H;�I;�
I;!I;ZI;�&I;&4I;�DI;�XI;BpI;��I;��I;'�I;��I;��I;[�I;�9I;CJH;��F;�rD;�FA;�/=;J98;�2;�\,;&;> ;�;x�;;      �0;�51;B�2;x�4;17;N#:;'0=;� @;8�B;�	E;��F;%H;�	I;��I;��I;��I;��I;/�I;��I;1�I;�mI;�WI;�DI;�4I;y'I;nI;=I;�I;qI;k I;k�H;�H;��H;��H;��H;��H;��H;��H;��H;��H;��H;�H;k�H;i I;pI;�I;;I;lI;{'I;�4I;�DI;�WI;�mI;3�I;��I;1�I;��I;��I;��I;��I;�	I;~%H;��F;�	E;8�B;� @;%0=;N#:;17;x�4;@�2;�51;      ƶ?;��?;��@;�tA;9�B;v�C;�BE;��F;��G;�xH;�I;��I;��I;��I;k�I;��I;G�I;f�I;B�I;LiI;�TI;-CI;)4I;�'I;�I;�I;PI;I;� I;��H;Q�H;��H;��H;�H;��H;b�H;-�H;c�H;�H;�H;��H;��H;S�H;��H;� I;I;OI;�I;�I;|'I;'4I;-CI;�TI;NiI;B�I;i�I;C�I;��I;k�I;��I;��I;��I;�I;�xH;��G;��F;�BE;v�C;9�B;�tA;��@;��?;      �F;��F;	�F;�2G;t�G;0&H;��H;
I;)mI;��I;��I;��I;�I;��I;�I;�I;��I;�wI;�bI;aPI;^@I;z2I;�&I;lI;�I;|I;\I;;I;�H;��H;��H;��H;��H;b�H;��H;
�H;��H;�H;��H;b�H;��H;��H;��H;��H;�H;<I;[I;|I;�I;iI;�&I;z2I;Z@I;aPI;�bI;�wI;��I;ߩI;��I;��I;�I;��I;��I;��I;)mI;I;��H;0&H;w�G;�2G;�F;��F;      � I;a'I;;I;�XI;|I;F�I;��I;'�I;D�I;C�I;��I;�I;��I;�I;w�I;=�I;mI;�ZI;�JI;X<I;�/I;�$I;^I;>I;LI;_I;CI;'�H;��H;��H;��H;��H;�H;��H;R�H;��H;��H;��H;P�H;��H;�H;��H;��H;��H;��H;(�H;BI;]I;PI;=I;\I;�$I;�/I;X<I;�JI;�ZI;mI;<�I;w�I;�I;��I;�I;��I;B�I;E�I;)�I;��I;D�I;|I;�XI;;I;`'I;      '�I;��I;*�I;��I;�I;W�I;�I;y�I;8�I;��I;ݾI;?�I;O�I;�I;�qI;aI;�QI;�CI;]7I;1,I;]"I;�I;%I;�I;I;=I;'�H;��H;��H;��H;��H;��H;��H;��H;�H;��H;��H;��H;�H;��H;��H;��H;��H;��H;��H;��H;'�H;=I;I;�I;$I;�I;["I;3,I;]7I;�CI;�QI;aI;�qI;�I;N�I;?�I;۾I;��I;8�I;}�I;�I;W�I;!�I;��I;)�I;��I;      �I;J�I;+�I;��I;��I;��I;��I;_�I;d�I;6�I;��I;C�I;qI;�bI;�TI;)HI;g<I;�1I;(I;YI;�I;�I;�
I;tI;� I;�H;��H;��H;��H;��H;��H;��H;~�H;��H;$�H;��H;��H;��H;$�H;��H;{�H;��H;��H;��H;��H;��H;��H;�H;� I;vI;�
I;�I;�I;WI;(I;�1I;d<I;)HI;�TI;�bI;qI;B�I;��I;5�I;d�I;_�I;��I;��I;��I;��I;+�I;>�I;      _�I;p�I;ϲI;9�I;�I;�I;�I;��I;��I;NvI;�jI;_I;�SI;�HI;�>I;�4I;�+I;�#I;�I;I;�I;}	I;�I;k I;��H;��H;��H;��H;��H;��H;j�H;Q�H;t�H;��H;M�H;
�H;��H;
�H;M�H;��H;q�H;R�H;k�H;��H;��H;��H;��H;��H;��H;k I;�I;}	I;�I;I;�I;�#I;�+I;�4I;�>I;�HI;�SI;_I;�jI;NvI;��I;��I;�I;�I;�I;:�I;ʲI;m�I;      ��I;�I;��I;5�I;||I;�vI;�oI;:hI;`I;�WI;�NI;JFI;�=I;f5I;v-I;�%I;�I;aI;mI;I;I;�I;��H;l�H;M�H;��H;��H;��H;��H;m�H;J�H;M�H;��H;�H;��H;n�H;0�H;n�H;��H;�H;��H;N�H;J�H;k�H;��H;��H;��H;��H;P�H;n�H;��H;�I;I;I;mI;aI;�I;�%I;v-I;e5I;�=I;HFI;�NI;�WI;`I;;hI;�oI;�vI;y|I;5�I;��I;�I;      �dI;dI;�bI;`I;r\I;
XI;�RI;JMI;=GI;�@I;J:I;�3I;-I;�&I;l I;�I;I;�I;I;�I;�I;7�H;��H;�H;��H;��H;��H;��H;��H;Q�H;J�H;��H;��H;d�H;�H;��H;��H;��H;�H;d�H;��H;��H;L�H;R�H;��H;��H;��H;��H;��H;�H;��H;7�H;�I;�I;I;�I;I;�I;l I;�&I;-I;�3I;J:I;�@I;=GI;JMI;�RI;XI;p\I;`I;�bI;dI;      �KI;�KI;7JI;:HI;�EI;$BI;D>I;�9I;/5I;)0I;+I;�%I;� I;�I;�I;I;�I;c	I;wI;�I;��H;��H;$�H;��H;��H;��H;�H;��H;�H;w�H;��H;��H;N�H;��H;��H;Y�H;g�H;Y�H;��H;��H;K�H;��H;��H;x�H;��H;��H;�H;��H;��H;��H;#�H;��H;��H;�I;wI;e	I;�I;I;�I;�I;� I;�%I;+I;*0I;.5I;�9I;D>I;%BI;EI;:HI;7JI;yKI;      :I;�9I;�8I;a7I;X5I;�2I;�/I;*,I;a(I;[$I;8 I;I;�I;�I;�I;�I;&I;�I;wI;p�H;��H;<�H;�H;��H;
�H;a�H;��H;��H;��H;��H;�H;c�H;��H;w�H;5�H;�H;��H;�H;5�H;w�H;��H;e�H;�H;��H;��H;��H;��H;_�H;�H;��H;�H;<�H;��H;q�H;wI;�I;%I;�I;�I;�I;�I;I;7 I;[$I;b(I;-,I;�/I;�2I;N5I;a7I;�8I;�9I;      �.I;k.I;�-I;<,I;�*I;E(I;�%I;�"I;�I;zI;I;�I;�I;{I;I;�I;�I;lI;��H;�H;��H;��H;s�H;��H;��H;��H;O�H;�H;$�H;M�H;��H;�H;��H;6�H;��H;��H;��H;��H;��H;7�H;��H;�H;��H;O�H;'�H;�H;N�H;��H;��H;��H;q�H;��H;��H;�H;��H;mI;�I;�I;I;{I;�I;�I;I;zI;�I;�"I;�%I;H(I;x*I;<,I;�-I;c.I;      �'I;�'I;�&I;�%I;s$I;r"I;- I;�I;�I;�I;�I;�I;I;cI;OI;PI;kI;��H;$�H;��H;��H;i�H;��H;��H;_�H;�H;��H;��H;��H;�H;n�H;��H;V�H;�H;��H;��H;��H;��H;��H;�H;U�H;��H;n�H;
�H;��H;��H;��H;�H;a�H;��H;��H;i�H;��H;��H;$�H;��H;jI;PI;OI;aI;I;�I;�I;�I;�I;�I;- I;w"I;i$I;�%I;�&I;�'I;      �%I;�%I;%I;�#I;j"I;� I;zI;�I;II;kI;�I;vI;wI;]
I;KI;�I;�I;0�H;��H;F�H;�H;�H;F�H;��H;*�H;��H;��H;��H;��H;��H;4�H;��H;i�H;��H;��H;��H;��H;��H;��H;��H;f�H;��H;4�H;��H;��H;��H;��H;��H;*�H;��H;F�H;�H;�H;F�H;��H;2�H;�I;�I;KI;]
I;wI;vI;�I;nI;II;�I;zI;� I;_"I;�#I;%I;�%I;      �'I;�'I;�&I;�%I;s$I;q"I;- I;�I;�I;�I;�I;�I;I;cI;OI;PI;kI;��H;$�H;��H;��H;i�H;��H;��H;a�H;
�H;��H;��H;��H;�H;n�H;��H;V�H;�H;��H;��H;��H;��H;��H;�H;U�H;��H;n�H;
�H;��H;��H;��H;�H;_�H;��H;��H;i�H;��H;��H;$�H;��H;jI;PI;OI;aI;I;�I;�I;�I;�I;�I;- I;w"I;h$I;�%I;�&I;�'I;      �.I;m.I;�-I;;,I;�*I;E(I;�%I;�"I;�I;yI;I;�I;�I;{I;I;�I;�I;lI;��H;�H;��H;��H;s�H;��H;��H;��H;O�H;�H;&�H;M�H;��H;�H;��H;7�H;��H;��H;��H;��H;��H;6�H;��H;�H;��H;O�H;'�H;�H;N�H;��H;��H;��H;s�H;��H;��H;�H;��H;mI;�I;�I;I;{I;�I;�I;I;zI;�I;�"I;�%I;H(I;x*I;<,I;�-I;c.I;      :I;�9I;�8I;a7I;X5I;�2I;�/I;*,I;a(I;[$I;8 I;I;�I;�I;�I;�I;&I;�I;wI;p�H;��H;<�H;�H;��H;�H;a�H;��H;��H;��H;��H;�H;c�H;��H;w�H;5�H;�H;��H;�H;5�H;w�H;��H;e�H;�H;��H;��H;��H;��H;a�H;
�H;��H;�H;<�H;��H;p�H;wI;�I;%I;�I;�I;�I;�I;I;8 I;[$I;b(I;-,I;�/I;�2I;M5I;a7I;�8I;�9I;      �KI;�KI;9JI;;HI;�EI;"BI;D>I;�9I;/5I;)0I;+I;�%I;� I;�I;�I;I;�I;c	I;wI;�I;��H;��H;$�H;��H;��H;��H;�H;��H;�H;w�H;��H;��H;L�H;��H;��H;X�H;g�H;Y�H;��H;��H;K�H;��H;��H;x�H;��H;��H;�H;��H;��H;��H;#�H;��H;��H;�I;wI;c	I;�I;I;�I;�I;� I;�%I;+I;*0I;/5I;�9I;D>I;$BI;EI;;HI;6JI;KI;      �dI;dI;�bI;`I;r\I;
XI;�RI;JMI;=GI;�@I;J:I;�3I;-I;�&I;l I;�I;I;�I;I;�I;�I;7�H;��H;�H;��H;��H;��H;��H;��H;Q�H;L�H;��H;��H;d�H;�H;��H;��H;��H;�H;d�H;��H;��H;J�H;R�H;��H;��H;��H;��H;��H;�H;��H;7�H;�I;�I;I;�I;I;�I;l I;�&I;-I;�3I;J:I;�@I;>GI;JMI;�RI;XI;o\I;`I;�bI;dI;      ��I;�I;��I;5�I;z|I;�vI;�oI;:hI;`I;�WI;�NI;HFI;�=I;f5I;v-I;�%I;�I;aI;mI;I;I;�I;��H;n�H;P�H;��H;��H;��H;��H;m�H;J�H;M�H;��H;�H;��H;n�H;0�H;n�H;��H;�H;��H;N�H;J�H;k�H;��H;��H;��H;��H;M�H;n�H;��H;�I;I;I;mI;aI;�I;�%I;v-I;h5I;�=I;JFI;�NI;�WI;`I;;hI;�oI;�vI;y|I;5�I;��I;�I;      W�I;p�I;ͲI;9�I;�I;�I;�I;��I;��I;MvI;�jI;_I;�SI;�HI;�>I;�4I;�+I;�#I;�I;I;�I;}	I;�I;k I;��H;��H;��H;��H;��H;��H;k�H;Q�H;s�H;��H;M�H;
�H;��H;
�H;M�H;��H;s�H;R�H;j�H;��H;��H;��H;��H;��H;��H;k I;�I;}	I;�I;I;�I;�#I;�+I;�4I;�>I;�HI;�SI;_I;�jI;MvI;��I;��I;�I;�I;�I;9�I;ͲI;q�I;      
�I;E�I;2�I;��I;��I;��I;��I;_�I;c�I;6�I;��I;B�I;qI;�bI;�TI;)HI;e<I;�1I;(I;YI;�I;�I;�
I;tI;� I;�H;��H;��H;��H;��H;��H;��H;|�H;��H;#�H;��H;��H;��H;$�H;��H;|�H;��H;��H;��H;��H;��H;��H;�H;� I;vI;�
I;�I;�I;YI;(I;�1I;e<I;*HI;�TI;�bI;qI;C�I;��I;6�I;d�I;a�I;��I;��I;��I;��I;1�I;E�I;      '�I;��I;*�I;��I;�I;W�I;�I;z�I;8�I;��I;ݾI;?�I;N�I;�I;�qI;aI;�QI;�CI;]7I;3,I;`"I;�I;%I;�I;I;=I;'�H;��H;��H;��H;��H;��H;��H;��H;�H;��H;��H;��H;�H;��H;��H;��H;��H;��H;��H;��H;'�H;=I;I;�I;$I;�I;["I;3,I;]7I;�CI;�QI;aI;�qI;�I;O�I;A�I;۾I;��I;8�I;|�I;�I;T�I;"�I;��I;)�I;��I;      � I;`'I;;I;�XI;|I;B�I;��I;'�I;E�I;C�I;��I;�I;��I;�I;w�I;=�I;mI;�ZI;�JI;Z<I;�/I;�$I;^I;>I;PI;_I;CI;(�H;��H;��H;��H;��H;�H;��H;P�H;��H;��H;��H;R�H;��H;�H;��H;��H;��H;��H;'�H;BI;_I;LI;=I;\I;�$I;�/I;X<I;�JI;�ZI;mI;<�I;w�I;�I;��I;�I;��I;C�I;D�I;'�I;��I;A�I;|I;�XI;;I;V'I;      �F;��F;�F;�2G;t�G;1&H;��H;I;'mI;��I;��I;��I;�I;��I;��I;�I;��I;�wI;�bI;aPI;`@I;z2I;�&I;iI;�I;}I;\I;<I;�H;��H;��H;��H;��H;b�H;��H;
�H;��H;
�H;��H;b�H;��H;��H;��H;��H;�H;;I;[I;|I;�I;kI;�&I;z2I;Z@I;aPI;�bI;�wI;��I;�I;�I;��I;�I;��I;��I;��I;'mI;I;��H;0&H;x�G;�2G;�F;��F;      ƶ?;��?;��@;�tA;9�B;v�C;�BE;��F;��G;�xH;�I;��I;��I;��I;k�I;��I;D�I;g�I;B�I;MiI;�TI;-CI;)4I;'I;�I;�I;PI;I;� I;��H;S�H;��H;��H;�H;��H;b�H;-�H;c�H;��H;�H;��H;��H;Q�H;��H;� I;I;OI;�I;�I;'I;'4I;-CI;�TI;MiI;B�I;i�I;D�I;��I;k�I;��I;��I;��I;�I;�xH;��G;��F;�BE;u�C;6�B;�tA;��@;��?;      �0;�51;G�2;u�4;
17;T#:;"0=;� @;:�B;�	E;��F;~%H;�	I;��I;��I;��I;��I;/�I;��I;3�I;�mI;�WI;�DI;�4I;{'I;nI;=I;�I;sI;k I;k�H;�H;��H;��H;��H;��H;��H;��H;��H;��H;��H;�H;k�H;h I;pI;�I;;I;nI;y'I;�4I;�DI;�WI;�mI;3�I;��I;0�I;��I;��I;��I;��I;�	I;%H;��F;�	E;:�B;� @;"0=;R#:;17;u�4;D�2;�51;      };(;��;�;6 ;&;�\,; �2;K98;�/=;�FA;�rD;��F;CJH;�9I;]�I;��I;��I;'�I;��I;��I;BpI;�XI;�DI;&4I;�&I;]I;!I;�
I;�I;��H;��H;$�H;�H;s�H;~�H;F�H;~�H;q�H;�H;#�H;��H;��H;�I;�
I;"I;ZI;�&I;#4I;�DI;�XI;BpI;��I;��I;'�I;��I;��I;]�I;�9I;EJH;��F;�rD;�FA;�/=;K98;�2;�\,;	&;: ;�;|�;;      ���:��:I�:8��:��:"Q ;�e;�V;z#;8e-;̼5;�h<;�tA;�	E;�eG;e�H;d�I;@�I;#�I;L�I;O�I;.�I;ApI;�WI;*CI;|2I;�$I;�I;�I;	I;�I;3�H;��H;;�H;��H;g�H;	�H;g�H;��H;;�H;��H;2�H;�I;{	I;�I;�I;�$I;|2I;)CI;�WI;<pI;/�I;N�I;N�I;#�I;A�I;d�I;f�H;�eG;�	E;�tA;�h<;ͼ5;:e-;z#;�V;�e;"Q ;K��:8��:G�:��:      ��p� �,��$9�Ƴ9p�": �u:��:���:X��:XR;� ;��,;F�6;�)>;<C;��F;�lH;�kI;��I;��I;��I;P�I;��I;�mI;�TI;b@I;�/I;\"I;�I;�I;I;�I;��H;��H;��H;��H;�H;��H;��H;��H;��H;�I;I;�I;�I;\"I;�/I;b@I;�TI;�mI;��I;P�I;��I;��I;��I;�kI;�lH;��F;<C;�)>;H�6;��,;� ;YR;\��:���:��:D�u:��":�Ƴ9�$9 �,�      �o&�>!��4����氺l�O� :T��u�9H�u:$�:2H�:<D;X#;�71;i;;��A;.�E;�$H;VI;E�I;��I;K�I;��I;3�I;GiI;bPI;W<I;0,I;WI;�I;�I;�I;�I;j�H;
�H;��H;@�H;��H;
�H;i�H;�I;�I;�I;�I;RI;0,I;T<I;bPI;GiI;.�I;��I;K�I;��I;G�I;�VI;�$H;.�E;��A;j;;�71;X#;<D;0H�:$�:H�u:v�9 :T�`�O�氺���4�I!�      �kٻV�Իwǻ����V���n���+���ԺT�1���39�m:�:��;8�;�\,;�8;�@;m]E;�
H;�VI;��I;"�I;'�I;��I;;�I;�bI;�JI;]7I;(I;�I;gI;I;qI;pI;��H;�H;��H;�H;��H;pI;qI;I;gI;�I;
(I;]7I;�JI;�bI;;�I;��I;"�I;#�I;��I;�VI;�
H;n]E;�@;�8;�\,;8�;��;�:�m:��39T�1���Ժ��+��n��V�� ���wǻV�Ի      4yY��|U�D�I�;�7��� ��!���Ի�᝻n�T�δ�#��v�9���:�l�:;�);B17;[ @;k]E;�$H;�kI;?�I;��I;,�I;d�I;�wI;�ZI;�CI;�1I;�#I;`I;�I;f	I;�I;oI;��H;7�H;��H;oI;�I;e	I;�I;`I;�#I;�1I;�CI;�ZI;�wI;d�I;)�I;��I;?�I;�kI;�$H;m]E;^ @;A17;�);;�l�:���:�v�9#�ƴ�n�T��᝻��Ի�!��� �;�7�D�I��|U�      ��ü\l��t����R��=ߓ�\�{��M��� ��컼���e�B��鰺@>o���u:���:�R;a�';B17;�@;0�E;�lH;d�I;��I;��I;?�I;��I; mI;�QI;`<I;�+I;�I;�I;�I;I;zI;`I;�I;`I;|I;I;�I;�I;�I;�+I;^<I;�QI;�lI;��I;@�I;��I;��I;d�I;�lH;3�E;�@;E17;`�';�R;���:��u:�=o��鰺e�B������컆� ��M�\�{�=ߓ��R��t���^l��      �'��-$�_��Z����	?ټw��:���iyY��k��Ի*���X�������$R:��:�R;�);�8;��A;��F;f�H;]�I;��I;��I;�I;=�I;aI;)HI;�4I;�%I;|I;I;�I;�I;GI;~I;GI;�I;�I;I;~I;�%I;�4I;&HI;aI;;�I;�I;��I;��I;Z�I;h�H;��F;��A;�8;�);�R;��:�$R:x����X��*���Ի�k�hyY�:���w��?ټ���Z�_���-$�      Z+����d̀�/l��Q�&�2�C��������@��}�>�N2��V��g1�p��$R:���:;�\,;j;;<C;�eG;�9I;��I;h�I;��I;t�I;�qI;�TI;�>I;o-I;d I;�I;�I;I;HI;GI;HI;I;�I;�I;e I;o-I;�>I;�TI;�qI;t�I;�I;i�I;��I;�9I;�eG;<C;m;;�\,;;���:�$R:p��g1�V��N2��}�>��@��������C�&�2��Q�/l�d̀���      m�ེhܽr�н_y��a什R ��l��n<�N���>ټ��Q|U�z������f1�������u:�l�:4�;�71;�)>;�	E;AJH;��I;��I;��I;�I;�I;�bI;�HI;^5I;�&I;�I;�I;tI;WI;U
I;WI;tI;�I;�I;�&I;^5I;�HI;�bI;�I;�I;��I;��I;��I;<JH;�	E;�)>;�71;4�;�l�:��u:x���g1�����x��P|U����>ټN���n<�l�R ��a什_y��r�н�hܽ      ��4�i1��&������k�ཇ�������`��'���TR��@�]�y��V���X��@>o����:��;X#;D�6;�tA;��F;�	I;��I;�I;��I;L�I;qI;�SI;�=I;�,I;� I;�I;�I;xI;sI;xI;�I;�I;� I;�,I;�=I;�SI;qI;L�I;��I;�I;��I;�	I;��F;�tA;F�6;Z#;��;���:�>o��X��V��x��@�]�TR����'��`��������k��������&�i1�      �x���o��ń�LUo���O�,�-�{��hܽ]什ռx���2�tb��TR��R|U�N2��*���鰺�v�9�:<D;��,;�h<;�rD;|%H;��I;��I;�I;8�I;<�I;_I;=FI;�3I;�%I;I;�I;�I;lI;�I;�I;I;�%I;�3I;<FI;_I;<�I;8�I;�I;��I;��I;y%H;�rD;�h<;��,;<D;�:�v�9�鰺+��N2��Q|U�TR��tb����2�ռx�]什�hܽ{�,�-���O�LUo�ń��o��      y���྅�Ѿ*����נ�
ń�<�S�	�#�bO��~n��K̀���2����~�>��Իk�B�,#��m:0H�:� ;ȼ5;�FA;��F;�I;��I;��I;־I;��I;�jI;�NI;A:I;+I;0 I;I;�I;�I;�I;I;. I;+I;A:I;�NI;�jI;��I;ԾI;��I;��I;�I;��F;�FA;Ƽ5;� ;,H�:�m: #�l�B���Ի}�>�������2�K̀�~n��bO��	�#�<�S�
ń��נ�*�����Ѿ��      �3���/��X#��	��A��،Ⱦ�f��KUo�`1�ΰ��~n��ռx��'��>ټ�@���k�����Ҵ�0�39�#�:UR;6e-;�/=;�	E;�xH;��I;@�I;��I;5�I;CvI;�WI;�@I;'0I;X$I;sI;�I;kI;�I;sI;W$I;&0I;�@I;�WI;CvI;2�I;��I;?�I;��I;�xH;�	E;�/=;6e-;WR;�#�:P�39δ𺿼���k��@���>ټ�'�ռx�~n��ΰ��`1�KUo��f��،Ⱦ�A���	��X#���/�      ���U���V�v��RZ�]58�ς�s��f���ioy�`1�bO��]什�`�O�����kyY���u�T�|�1�<�u:J��:p#;C98;3�B;��G;&mI;>�I;/�I;`�I;��I;`I;3GI;(5I;Z(I;�I;�I;@I;�I;�I;X(I;&5I;4GI;`I;��I;]�I;/�I;;�I;%mI;��G;/�B;A98;p#;R��:4�u:|�1�r�T���kyY����O���`�]什bO��`1�ioy�f���s��ς�]58��RZ�V�v�U���      Ŀ7g��(ﱿ���U����U��X#�w��f���KUo�	�#��hܽ����n<����:����� ��᝻��Ժ�u�9���:�V;��2;� @;��F;I;)�I;p�I;^�I;��I;3hI;@MI;�9I;#,I;�"I;�I;�I;�I;�"I;#,I;�9I;@MI;3hI;��I;[�I;p�I;'�I;I;��F;� @;��2;�V;���:�u�9��Ժ�᝻�� �:�������n<�����hܽ	�#�KUo�f���w���X#��U�U������(ﱿ7g��      �x�Q9�T��uؿpQ��g_��8�_��X#�s���f��<�S�{�����l�C�w���M���Ի��+�`:T���:�e;�\,;0=;�BE;��H;��I;�I;��I;�I;�oI;�RI;D>I;�/I;�%I;% I;xI;% I;�%I;�/I;D>I;�RI;�oI;�I;��I;�I;��I;��H;�BE;0=;�\,;�e;��:p:T���+���Ի�M�w��C�l�����{�<�S��f��s���X#�8�_�g_��pQ��uؿT��Q9�      �X1���,�i���<��7g��f_���U�ς�،Ⱦ
ń�,�-�k��R ��'�2�
?ټ^�{��!��n�t�O��u:Q ;�&;H#:;o�C;1&H;>�I;S�I;��I;�I;�vI;XI;!BI;�2I;F(I;t"I;� I;u"I;F(I;�2I;BI;XI;�vI;
�I;��I;S�I;>�I;0&H;r�C;F#:;�&;Q ; �u:t�O��n��!�_�{�
?ټ'�2�R ��k��,�-�
ń�،Ⱦς��U�f_��7g��<�i����,�      d��]]�6K��X1�[f��pQ��U���]58��A���נ���O���a什�Q����>ߓ��� ��V��,氺l�":��:: ;17;6�B;p�G;|I;�I;��I;�I;l|I;k\I;{EI;P5I;j*I;a$I;]"I;a$I;i*I;N5I;zEI;k\I;l|I;ߧI;��I;�I;|I;n�G;6�B;	17;< ;��:t�":,氺�V���� �>ߓ�����Q�a什����O��נ��A��]58�U���pQ���[f��X1�6K��]]�      O������4z���V��X1��<�uؿ����RZ��	�*���LUo����`y��/l�[��R��=�7�������Ƴ9:��:�;q�4;�tA;�2G;�XI;��I;��I;4�I;'�I;�_I;,HI;V7I;0,I;�%I;�#I;�%I;0,I;U7I;*HI;�_I;'�I;2�I;��I;��I;�XI;�2G;�tA;n�4;�;:��:�Ƴ9������=�7��R��[�0l�`y�����LUo�*����	��RZ����uؿ�<��X1���V��4z�����      �o��g^���ē��4z�6K�i��T��(ﱿV�v��X#���Ѿń�	�&�s�нd̀�`��t���F�I��ǻ�4��#9�:l�;4�2;��@;�F;;I; �I;,�I;ŲI;��I;�bI;.JI;�8I;�-I;�&I;%I;�&I;�-I;�8I;,JI;�bI;��I;²I;+�I; �I;;I;�F;��@;0�2;o�;�:�#9�4��ǻF�I�u���a��d̀�s�н	�&�ń���Ѿ�X#�V�v�(ﱿT��i��6K��4z��ē�g^��      r'���X��g^�������]]���,�Q9�7g��U�����/����o��i1��hܽ���-$�_l���|U�Z�ԻV!� �,���:;�51;��?;|�F;Z'I;��I;H�I;d�I;цI;
dI;oKI;�9I;V.I;�'I;�%I;�'I;Y.I;�9I;nKI;dI;цI;b�I;E�I;��I;Y'I;|�F;��?;�51;;��: �,�W!�Z�Ի�|U�_l���-$����hܽi1��o���ྜ�/�U���7g��Q9���,��]]�����g^���X��      m����������Ѣ��1�j��5���	��ȿ(8����7�G�꾄S���7�3�L���)���Ƽ��\���ݻ]+��Rɸ��:Wx;��0;Ҥ?;��F;,I;��I;�I;��I;U�I;iI;*OI;�<I;1I;�)I;�'I;�)I;1I;�<I;)OI;iI;U�I;��I;�I;��I;,I;��F;Ҥ?;��0;Zx;��:�Rɸ^+���ݻ��\���Ƽ�)�L��3��7��S��G�꾫�7�(8���ȿ��	��5�1�j�Ѣ����������      ��������B��^�����c�821�&X��ÿjڇ�t�3��s��7��~74�d�?ى���&�Nü%�X���ػ`�%�@�J����:�b;��0;��?;H�F;�2I;�I;u�I;�I;z�I;�hI;�NI;d<I;�0I;�)I;�'I;�)I;�0I;d<I;�NI;�hI;z�I;�I;r�I;�I;�2I;H�F;��?;��0;�b;���:@�J�a�%���ػ$�X�Nü��&�?ى�d�~74��7���s�t�3�jڇ��ÿ&X�821���c�^����B�����      �����B����F��y�P���#�P�������x|��'�[D־�X��q�)� Խ�Ă�J<�8_��y-M���ʻ,���)�8���:�;6K2;Ev@;��F;�FI;��I;=�I;U�I;2�I;�fI;pMI;v;I;�/I;�(I;�&I;�(I;�/I;v;I;oMI;�fI;2�I;Q�I;<�I;��I;�FI;��F;Ev@;0K2;�;���:�)�8/����ʻx-M�8_��J<��Ă� Խq�)��X��[D־�'��x|����P�����#�y�P�F�����B��      Ѣ��^���F���/]��5�O���,ݿ-8��sm_��K��t��Z�s�%>����;�o��3��۩���:�`T�������(�9�f�:�<;�_4;=hA;L8G;�dI;3�I;c�I;��I;��I;]dI;LKI;�9I;.I;�'I;�%I;�'I;.I;�9I;KKI;[dI;��I;��I;`�I;3�I;�dI;G8G;<hA;�_4;�<;�f�:�(�9����`T����:��۩��3�;�o����%>�Z�s��t���K�sm_�-8���,ݿO���5��/]�F��^���      1�j���c�y�P��5���u��J���jڇ�Iv<�*���r���_S��������+T��� �*$���G#�����1��|�:���:i�;L7;��B;��G;�I;F�I;��I;��I;��I;�`I;|HI;�7I;�,I;:&I;3$I;:&I;�,I;�7I;zHI;�`I;��I;�I;��I;F�I;�I;��G;��B;H7;j�;���:��:1�������G#�*$���� �+T���������_S�r��*���Iv<�jڇ�J���u�����5�y�P���c�      �5�821���#�O��u���ÿ�ҕ�Z������̾�X����0�3�1W����5��zܼ;��R��?�s��T\���n:%��:�%;��9;��C;/H;B�I;B�I;<�I;��I;�{I;?\I;EI;�4I;_*I;I$I;K"I;I$I;_*I;�4I;EI;?\I;�{I;��I;8�I;B�I;A�I;/H;��C;��9;�%;%��:��n:�T\�@�s�R��<���zܼ��5�1W��3佁�0��X����̾���Z��ҕ��ÿu��O����#�821�      ��	�&X�P����,ݿJ����ҕ��d��'�B��%���{�W����m���4�o��G��*���Q���ػ߮0���~�0�:��;e,;�=;pBE;ĬH;��I;��I;}�I;�I;�tI;�VI;AI;�1I;�'I;�!I; I;�!I;�'I;�1I;AI;�VI;�tI;�I;z�I;��I;��I;ĬH;kBE;�=;d,;��;0�:��~�߮0���ػ�Q��*���G�4�o�m������{�W�%���B�꾎'��d��ҕ�J����,ݿP���&X�      �ȿ�ÿ���-8��jڇ�Z��'�����n8��Z�s�/�&�Z�1j??��V�琼QG#�P7��0Tܺ��9\W�:��;NL2;x@;�F;0I;��I;��I;��I;q�I;�lI;QI;�<I;/.I;�$I;VI;{I;VI;�$I;/.I;�<I;QI;�lI;q�I;��I;��I;��I;0I;�F;t@;PL2;��;^W�:��92TܺP7��RG#�琼�V�j??�1Z�.�&�Z�s�n8�������'�Z�jڇ�-8������ÿ      (8��jڇ��x|�sm_�Iv<����B��n8��'6~�q74��l��|���9nc�5���^����\��9�%Z�H�=���n:���:"#;�8;��B;��G;�xI;��I;��I;��I;�I;idI;�JI;�7I;M*I;l!I;~I;�I;�I;l!I;M*I;�7I;�JI;idI;�I;��I;��I;��I;�xI;��G;��B;�8;"#;���:��n:H�=�$Z��9���\��^��5��9nc�|����l��q74�'6~�n8��B�꾐��Iv<�sm_��x|�jڇ�      ��7�t�3��'��K�*�����̾%���Z�s�q74����#N��Ї|��)�:zܼ�Y��: �{������pV93��:J�;.-;==;�E;6�H;��I;a�I;��I;ޥI;K{I;�[I;�CI;�2I;H&I;I;_I;�I;_I;I;H&I;�2I;�CI;�[I;L{I;ۥI;��I;_�I;��I;3�H;�E;;=;.-;L�;/��:pV9����|��: ��Y��:zܼ�)�Ї|�#N�����q74�Z�s�%�����̾*����K��'�t�3�      G���s�[D־�t��r���X��{�W�.�&��l��#N���Ă�j�5�����{Q����A�7�ػ��G�x!/��f:^b�:��;��5;�9A;s�F;+I;�I;	�I;>�I;��I;aoI;�RI;�<I;P-I;�!I;{I;5I;�I;6I;|I;�!I;M-I;�<I;�RI;aoI;��I;>�I;�I;	�I;+I;o�F;�9A;��5;ߖ;^b�:�f:l!/���G�7�ػ��A�{Q������j�5��Ă�#N���l��.�&�{�W��X��r���t��[D־�s�      �S���7���X��Z�s��_S���0����Z�|���Ї|�j�5�j���ک�3�X�c �h􃻎3���9c��:�;,�,;�L<;�oD;;.H;��I;��I;��I;��I;��I;jcI;�II;6I; (I;I;�I;�I;�I;�I;�I;I; (I;6I;�II;jcI;��I;��I;��I;��I;��I;8.H;�oD;�L<;.�,;�;_��: �9�3��i�c �3�X��ک�k��j�5�Ї|�|���Zཤ����0��_S�Z�s��X���7��      �7�~74�q�)�%>����3�m���08nc��)������ک�pa��Q�B����M�@�ȸp��:�;�#;��6;2hA;��F;�I;n�I;��I;F�I;��I;�uI;�WI;�@I;=/I;�"I;MI;6I;�I;�I;�I;6I;MI;�"I;>/I;�@I;�WI;�uI;��I;B�I;��I;m�I;�I;��F;3hA;��6;�#;�;r��:`�ȸ�M�C����Q�qa��ک������)�8nc�1m���3����%>�q�)�~74�      3�c�Խ�������0W��3�o�j??�4��9zܼzQ��2�X��Q��6�������Ϲ0�n:�m�:=>;��0;�>;aE;�SH;z�I;��I;��I;t�I;��I;gI;XLI;�7I;�(I;BI;*I;�I;SI;vI;SI;�I;(I;BI;�(I;�7I;XLI;gI;��I;r�I;��I;��I;x�I;�SH;`E;�>;��0;=>;�m�:$�n:��Ϲ����6���Q�2�X�{Q��9zܼ4��j??�3�o�0W���������Խc�      ~L��?ى��Ă�:�o�+T���5��G��V��^���Y����A�c �B������(����J:�l�:f;M,;��:;<5C;AlG;EI;0�I;��I;��I;ŝI;�vI;�XI;zAI;�/I;D"I;I;�I;�I;2	I;�I;1	I;�I;�I;I;G"I;�/I;xAI;�XI;�vI;ÝI;��I;��I;,�I;EI;ClG;95C;��:;M,;f;�l�:��J:(�����C���c ���A��Y���^���V��G���5�+T�:�o��Ă�?ى�      �)���&�I<��3��� ��zܼ�*��琼��\�9 �4�ػh��M���Ϲ��J:�j�:��;��(;�e8;͕A;C�F;�H;S�I;��I;7�I;/�I;��I;�eI;�KI;N7I;�'I;I;GI;I;�I;I;bI;I;�I; I;DI;I;�'I;O7I;�KI;�eI;��I;1�I;6�I;��I;O�I;�H;A�F;̕A;�e8;��(;��;�j�:��J:��Ϲ�M�h�4�ػ9 ���\�琼�*���zܼ�� ��3�I<���&�      ��ƼNü7_���۩�)$��9���Q�OG#��9�x����G��3�� �ȸ0�n:�l�:��;G�';�7;�v@;V�E;FvH;)�I;��I;�I;s�I;��I;�qI;�UI;g?I;.I;� I;HI;�I;	I;zI;"I;[I;"I;zI;	I;�I;HI;� I;.I;d?I;�UI;�qI;��I;s�I;�I;��I;'�I;DvH;W�E;�v@;�7;G�';��;�l�:0�n:@�ȸ�3����G�x���9�OG#��Q�8��)$���۩�7_��Nü      ��\�"�X�v-M���:��G#�S����ػP7��Z�����`!/��9p��:�m�:f;��(;�7;�@;T]E;�-H;gwI;��I;��I;��I;�I;}I;	_I;GI;%4I;�%I;�I;I;
I;tI;XI;a I;��H;a I;XI;tI;~
I;I;�I;�%I;"4I;GI;_I;}I;��I;��I;��I;��I;cwI;�-H;T]E;�@;�7;��(;f;�m�:p��:�9`!/�����Z�P7����ػR���G#���:�v-M�%�X�      �ݻ��ػ��ʻ\T������5�s�Ԯ0�(Tܺ �=��V9�f:m��:�;B>;Q,;�e8;�v@;T]E;bH;7bI;D�I;��I;s�I;ʭI;��I;7gI;7NI;:I;"*I;�I;�I;1I;mI;=I;}�H;��H;��H;��H;}�H;=I;mI;3I;�I;�I;*I;:I;3NI;9gI;��I;ƭI;o�I;��I;B�I;8bI;aH;U]E;�v@;�e8;Q,;B>;�;k��:�f:�V9 �=�*TܺԮ0�1�s�����\T����ʻ��ػ      W+�H�%�(������1���T\�P�~���9��n:9��:fb�:�;�#;��0;��:;ǕA;U�E;�-H;4bI;��I;��I;��I;<�I;�I;�mI;5TI;@?I;k.I;#!I;�I;6I;�I;�I;2�H;��H;A�H;��H;B�H;��H;2�H;�I;�I;6I;�I;!I;k.I;=?I;5TI;�mI;�I;8�I;��I;��I;��I;4bI;�-H;S�E;ǕA;��:;��0;�#;�;bb�:3��:��n:��9P�~��T\��0������(��R�%�       Qɸ��J� +�8�(�9x�:�n::�:bW�:���:P�;�;/�,;��6;�>;=5C;A�F;GvH;gwI;D�I;��I;l�I;��I;��I;�rI;�XI;nCI;$2I;a$I;I;&I;	I;yI;x�H;d�H;�H;��H;��H;��H;�H;d�H;x�H;{I;	I;%I;	I;b$I;!2I;nCI;�XI;�rI;��I;��I;h�I;��I;D�I;iwI;FvH;A�F;<5C;�>;��6;,�,;��;N�;���:^W�:8�:�n:��:�(�9�*�8��J�      �:C��:+��:�f�:���:A��:��;��;+#;1-;��5;�L<;5hA;cE;DlG;�H;)�I;��I;��I;��I;��I;&�I;'uI;�[I;�FI;�4I;�&I;jI;�I;�
I;�I;��H;F�H;��H;��H;��H;��H;��H;��H;��H;C�H;��H;�I;�
I;�I;kI;�&I;�4I;�FI;�[I;$uI;&�I;��I;��I;��I;��I;&�I;�H;ElG;cE;3hA;�L<;��5;1-;*#;��;��;G��:%��:�f�:+��:5��:      bx;�b;�;�<;e�;�%;l,;PL2;�8;A=;�9A;�oD;��F;�SH;EI;R�I;��I;��I;t�I;=�I;��I;*uI;�\I;�GI;�6I;�(I;I;xI;�I;�I;~ I;��H;��H;;�H;��H;�H;��H;�H;��H;=�H;��H;��H;} I;�I;�I;yI;I;�(I;�6I;�GI;�\I;*uI;��I;@�I;t�I;��I;��I;Q�I;EI;�SH;��F;�oD;�9A;?=;�8;PL2;l,;�%;m�;�<;�;�b;      ��0;��0;BK2;�_4;P7;��9;�=;z@;��B;�E;v�F;=.H;�I;|�I;3�I;��I;
�I;�I;ʭI;�I;�rI;�[I;�GI;Y7I;�)I;7I;�I;�I;iI;'I;��H;��H;4�H;*�H;��H;>�H;��H;>�H; �H;+�H;3�H;��H;��H;$I;gI;�I;�I;7I;�)I;V7I;�GI;�[I;�rI;�I;ʭI;�I;�I;��I;2�I;|�I;�I;=.H;u�F;�E;��B;{@;�=;��9;V7;�_4;@K2;��0;      �?;��?;6v@;GhA;��B;��C;pBE;�F;��G;5�H;+I;��I;n�I;�I;��I;9�I;y�I;��I;��I;nI;�XI;�FI;�6I;�)I;�I;I;pI;�I;�I;s�H;��H;�H;��H;d�H;N�H;��H;j�H;��H;N�H;c�H;��H;�H;��H;q�H;�I;�I;oI;I;�I;�)I;�6I;�FI;�XI;nI;��I;��I;v�I;7�I;��I;�I;m�I;��I;+I;3�H;��G;�F;pBE;��C;��B;DhA;5v@;��?;      ��F;a�F;��F;S8G;��G;/H;ƬH;,I;�xI;��I;	�I;��I;��I;��I;��I;/�I;��I; }I;4gI;5TI;mCI;�4I;�(I;5I;I;�I;nI;�I;��H;�H;6�H;��H;�H;��H;��H;1�H;)�H;1�H;��H;��H;�H;��H;6�H;�H;��H;�I;mI;�I;I;3I;�(I;�4I;hCI;5TI;6gI;}I;��I;.�I;��I;��I;��I;��I;	�I;��I;�xI;-I;ƬH;/H;��G;Q8G;��F;V�F;      #,I;�2I;�FI;�dI;�I;K�I;��I;��I;��I;d�I;�I;��I;E�I;u�I;ƝI;��I;�qI;_I;9NI;B?I;%2I;�&I;I;�I;lI;oI;(I;��H;M�H;:�H;��H;��H;s�H;[�H;g�H;��H;��H;��H;e�H;Z�H;q�H;��H;��H;:�H;M�H;��H;%I;oI;oI;�I;I;�&I;"2I;B?I;9NI;	_I;�qI;��I;ɝI;u�I;F�I;��I;�I;b�I;��I;��I;��I;F�I;��I;�dI;�FI;�2I;      ��I;�I;��I;6�I;I�I;E�I;��I;��I;��I;��I;E�I;��I;��I;��I;�vI;�eI;�UI;GI;:I;n.I;b$I;kI;{I;�I;�I;�I;��H;m�H;W�H;��H;��H;9�H;��H;��H;\�H;��H;��H;��H;\�H;��H;��H;;�H;��H;��H;W�H;n�H;��H;�I;�I;�I;yI;kI;`$I;n.I;:I;GI;�UI;�eI;�vI;��I;��I;��I;C�I;��I;��I;��I;��I;E�I;S�I;5�I;��I;(�I;      +�I;v�I;<�I;m�I;��I;9�I;~�I;��I;ĵI;�I;��I;��I;�uI;gI;�XI;�KI;k?I;#4I;$*I;!!I;I;�I;�I;kI;�I;��H;K�H;W�H;��H;��H;�H;��H;��H;��H;v�H;�H;��H;�H;v�H;��H;��H;��H;�H;��H;��H;W�H;N�H;��H;�I;kI;�I;�I;I;#!I;$*I;%4I;j?I;�KI;�XI;gI;�uI;��I;��I;ޥI;ĵI;��I;~�I;;�I;��I;m�I;<�I;i�I;      
�I;"�I;]�I;��I;�I;��I; �I;x�I;�I;U{I;koI;xcI;�WI;bLI;~AI;R7I; .I;%I;�I;�I;'I;�
I;�I;'I;m�H;�H;:�H;��H;��H;$�H;��H;��H;��H;��H;]�H;0�H;1�H;0�H;]�H;��H;��H;��H;��H;#�H;��H;��H;9�H;�H;p�H;'I;�I;�
I;&I;�I;�I;�%I;.I;R7I;AI;aLI;�WI;ycI;joI;U{I;�I;|�I;!�I;��I;�I;��I;Y�I;�I;      [�I;��I;<�I;��I;ʁI;�{I;�tI;�lI;udI;�[I;�RI;�II;�@I;8I;�/I;(I;� I;�I;�I;<I;!	I;�I;� I;��H;��H;7�H;��H;��H;�H;��H;x�H;t�H;��H; �H;��H;��H;h�H;��H;��H; �H;��H;v�H;x�H;��H;�H;��H;��H;6�H;��H;��H;} I;�I;	I;<I;�I;�I;� I;(I;�/I;8I;�@I;�II;�RI;�[I;sdI;�lI;�tI;�{I;ɁI;��I;<�I;��I;      iI;�hI;gI;idI;�`I;B\I;�VI;QI;�JI;�CI;�<I;6I;A/I;�(I;M"I;"I;TI;I;8I;�I;�I;��H;��H;��H;�H;��H;��H;;�H;��H;��H;q�H;��H;��H;q�H;%�H;��H;��H;��H;%�H;q�H;��H;��H;s�H;��H;��H;;�H;��H;��H;�H;��H;��H;��H;�I;�I;8I;I;RI;"I;M"I;�(I;A/I;6I;�<I;�CI;�JI;QI;�VI;E\I;�`I;idI;gI;�hI;      2OI;�NI;xMI;YKI;�HI;EI;AI;�<I;�7I;�2I;T-I;(I;�"I;FI; I;II;�I;z
I;qI;�I;��H;H�H;��H;7�H;��H;�H;t�H;��H;��H;��H;��H; �H;P�H; �H;��H;r�H;g�H;r�H;��H; �H;N�H;�H;��H;��H;��H;��H;q�H;�H;��H;9�H;��H;H�H;�H;�I;qI;{
I;�I;II;I;FI;�"I;(I;T-I;�2I;�7I;�<I;AI;EI;}HI;YKI;xMI;�NI;      �<I;p<I;q;I;�9I;�7I;�4I;�1I;7.I;U*I;M&I;�!I;�I;PI;/I;�I;I;$	I;vI;FI;:�H;n�H;��H;=�H;.�H;`�H;��H;W�H;��H;��H;��H;�H;o�H;��H;��H;H�H;.�H;�H;.�H;H�H;��H;��H;r�H;�H;��H;��H;��H;W�H;��H;a�H;-�H;=�H;��H;l�H;:�H;FI;vI;!	I;I;�I;1I;PI;�I;�!I;M&I;V*I;:.I;�1I;�4I;�7I;�9I;r;I;i<I;      1I;�0I;�/I;�.I;�,I;]*I;�'I;�$I;v!I;I;�I;�I;=I;�I;�I;�I;�I;VI;��H;��H;�H;��H;��H;�H;H�H;��H;c�H;[�H;v�H;]�H;��H;(�H;��H;M�H;��H;��H;��H;��H;��H;M�H;��H;)�H;��H;`�H;x�H;[�H;a�H;��H;H�H;�H;��H;��H;�H;��H;��H;XI;�I;�I;�I;�I;;I;�I;�I;I;v!I;�$I;�'I;b*I;�,I;�.I;�/I;�0I;      �)I;�)I;�(I;�'I;N&I;I$I;�!I;cI;�I;cI;=I;�I;�I;^I;9	I;I;-I;^ I;��H;I�H;��H;��H;�H;A�H;��H;.�H;��H;��H;�H;0�H;��H;��H;r�H;3�H;��H;��H;��H;��H;��H;0�H;q�H;��H;��H;0�H;�H;��H;��H;-�H;��H;A�H;�H;��H;��H;K�H;��H;` I;,I;I;9	I;]I;�I;�I;<I;eI;�I;cI;�!I;M$I;D&I;�'I;�(I;�)I;      �'I;�'I;'I;�%I;>$I;M"I; I;�I;�I;�I;�I;�I;�I;I;�I;hI;cI;��H;��H;��H;��H;��H;��H;��H;h�H;%�H;��H;��H;��H;5�H;m�H;��H;j�H;�H;��H;��H;��H;��H;��H;�H;g�H;��H;m�H;7�H;��H;��H;��H;&�H;h�H;��H;��H;��H;��H;��H;��H;��H;bI;hI;�I;I;�I;�I;�I;�I;�I;�I; I;Q"I;3$I;�%I;'I;�'I;      �)I;�)I;�(I;�'I;N&I;I$I;�!I;cI;�I;bI;=I;�I;�I;^I;9	I;I;-I;^ I;��H;I�H;��H;��H;�H;A�H;��H;.�H;��H;��H;�H;.�H;��H;��H;r�H;3�H;��H;��H;��H;��H;��H;0�H;q�H;��H;��H;1�H;�H;��H;��H;-�H;��H;A�H;�H;��H;��H;K�H;��H;` I;,I;I;9	I;]I;�I;�I;=I;cI;�I;cI;�!I;M$I;D&I;�'I;�(I;�)I;      1I;�0I;�/I;�.I;�,I;]*I;�'I;�$I;v!I;I;�I;�I;;I;�I;�I;�I;�I;VI;��H;��H;�H;��H;��H;�H;H�H;��H;c�H;[�H;w�H;]�H;��H;(�H;��H;M�H;��H;��H;��H;��H;��H;M�H;��H;,�H;��H;`�H;x�H;[�H;a�H;��H;H�H; �H;��H;��H;�H;��H;��H;XI;�I;�I;�I;�I;=I;�I;�I;I;v!I;�$I;�'I;b*I;�,I;�.I;�/I;�0I;      �<I;p<I;q;I;�9I;�7I;�4I;�1I;7.I;U*I;M&I;�!I;�I;PI;/I;�I;I;$	I;tI;FI;:�H;p�H;��H;=�H;.�H;a�H;��H;W�H;��H;��H;��H;�H;o�H;��H;��H;H�H;.�H;�H;.�H;H�H;��H;��H;r�H;�H;��H;��H;��H;W�H;��H;`�H;-�H;=�H;��H;l�H;:�H;FI;wI;!	I;I;�I;1I;PI;�I;�!I;M&I;V*I;:.I;�1I;�4I;�7I;�9I;r;I;i<I;      4OI;�NI;zMI;ZKI;�HI;EI;AI;�<I;�7I;�2I;T-I;(I;�"I;FI;I;II;�I;z
I;qI;�I;��H;H�H;��H;9�H;��H;	�H;t�H;��H;��H;��H;��H; �H;O�H;��H;��H;r�H;g�H;r�H;��H;��H;N�H;�H;��H;��H;��H;��H;q�H;�H;��H;7�H;��H;H�H;�H;�I;qI;z
I;�I;II; I;GI;�"I;(I;S-I;�2I;�7I;�<I;AI;EI;}HI;\KI;wMI;�NI;      iI;�hI;	gI;idI;�`I;B\I;�VI;QI;�JI;�CI;�<I;6I;A/I;�(I;M"I;"I;TI;I;8I;�I;�I;��H;��H;��H;�H;��H;��H;;�H;��H;��H;s�H;��H;��H;q�H;%�H;��H;��H;��H;%�H;q�H;��H;��H;q�H;��H;��H;;�H;��H;��H;�H;��H;��H;��H;�I;�I;8I;I;RI;"I;M"I;�(I;A/I;6I;�<I;�CI;�JI;QI;�VI;C\I;�`I;idI;	gI;�hI;      [�I;��I;<�I;��I;ʁI;�{I;�tI;�lI;udI;�[I;�RI;�II;�@I;8I;�/I;(I;� I;�I;�I;:I;#	I;�I;� I; �H;��H;7�H;��H;��H;�H;��H;x�H;t�H;��H; �H;��H;��H;h�H;��H;��H; �H;��H;v�H;x�H;��H;�H;��H;��H;6�H;��H;��H;} I;�I;	I;<I;�I;�I;� I;(I;�/I;8I;�@I;�II;�RI;�[I;sdI;�lI;�tI;�{I;ɁI;��I;<�I;��I;      �I;"�I;\�I;��I;�I;��I; �I;x�I;�I;S{I;koI;xcI;�WI;bLI;~AI;R7I; .I;%I;�I;�I;*I;�
I;�I;&I;p�H;�H;:�H;��H;��H;$�H;��H;��H;��H;��H;]�H;0�H;1�H;0�H;]�H;��H;��H;��H;��H;#�H;��H;��H;9�H;�H;m�H;(I;�I;�
I;&I;�I;�I;�%I;.I;S7I;~AI;aLI;�WI;xcI;koI;U{I;�I;{�I;!�I;��I;�I;��I;\�I;#�I;      &�I;r�I;C�I;k�I;��I;7�I;�I;��I;µI;ޥI;��I;��I;�uI;gI;�XI;�KI;k?I;#4I;$*I;#!I;I;�I;�I;kI;�I;��H;K�H;W�H;��H;��H;�H;��H;��H;��H;t�H;�H;��H;�H;v�H;��H;��H;��H;�H;��H;��H;W�H;M�H;��H;�I;kI;�I;�I;I;#!I;$*I;%4I;j?I;�KI;�XI;gI;�uI;��I;��I;ߥI;ĵI;��I;��I;8�I;��I;i�I;A�I;r�I;      ��I;�I;��I;5�I;I�I;E�I;��I;��I;��I;��I;E�I;��I;��I;��I;�vI;�eI;�UI;GI;:I;n.I;e$I;kI;{I;�I;�I;�I;��H;n�H;W�H;��H;��H;;�H;��H;��H;[�H;��H;��H;��H;\�H;��H;��H;;�H;��H;��H;V�H;m�H;��H;�I;�I;�I;yI;kI;`$I;n.I;:I;GI;�UI;�eI;�vI;��I;��I;��I;C�I;��I;��I;��I;��I;B�I;T�I;6�I;��I;(�I;      ,I;�2I;�FI;�dI;�I;E�I;��I;��I;��I;d�I;�I;��I;F�I;u�I;ȝI;��I;�qI;_I;9NI;D?I;(2I;�&I;I;�I;oI;rI;'I;��H;N�H;;�H;��H;��H;q�H;Z�H;e�H;��H;��H;��H;g�H;Z�H;s�H;��H;��H;:�H;M�H;��H;'I;oI;lI;�I;I;�&I;!2I;B?I;9NI;	_I;�qI;��I;ƝI;u�I;E�I;��I;�I;d�I;��I;��I;��I;D�I;�I;�dI;�FI;�2I;      ��F;Z�F;��F;S8G;��G;/H;ƬH;-I;�xI;��I;	�I;��I;��I;��I;��I;/�I;��I;}I;6gI;5TI;nCI;�4I;�(I;5I;I;�I;mI;�I;��H;�H;6�H;��H;�H;��H;��H;1�H;)�H;1�H;��H;��H;�H;��H;6�H;�H;��H;�I;kI;�I;I;3I;�(I;�4I;gCI;5TI;4gI;}I;��I;/�I;��I;��I;��I;��I;	�I;��I;�xI;-I;ȬH;/H;��G;S8G;��F;Q�F;      �?;��?;6v@;DhA;��B;��C;pBE;�F;��G;5�H;+I;��I;m�I;�I;��I;9�I;w�I;��I;��I;nI;�XI;�FI;�6I;�)I;�I;I;pI;�I;�I;q�H;��H;�H;��H;c�H;M�H;��H;j�H;��H;N�H;c�H;��H;�H;��H;q�H;�I;�I;oI;I;�I;�)I;�6I;�FI;�XI;nI;��I;��I;v�I;9�I;��I;�I;n�I;��I;+I;3�H;��G;�F;pBE;��C;��B;GhA;5v@;��?;      ��0;��0;DK2;�_4;J7;��9;�=;z@;��B;�E;v�F;=.H;�I;|�I;2�I;��I;
�I;�I;ʭI;�I;�rI;�[I;�GI;Y7I;�)I;7I;�I;�I;iI;&I;��H;��H;3�H;*�H;��H;>�H;��H;>�H; �H;*�H;3�H;��H;��H;$I;fI;�I;�I;7I;�)I;W7I;�GI;�[I;�rI;�I;ʭI;�I;�I;��I;2�I;|�I;�I;=.H;u�F;�E;��B;{@;�=;��9;Z7;�_4;DK2;��0;      _x;�b;�;�<;e�;�%;p,;PL2;�8;A=;�9A;�oD;��F;�SH;EI;R�I;��I;��I;t�I;?�I;��I;*uI;�\I;�GI;�6I;�(I;I;yI;�I;�I;} I;��H;��H;=�H;��H;�H;��H;�H;��H;;�H;��H;��H;~ I;�I;�I;xI;I;�(I;�6I;�GI;�\I;*uI;��I;@�I;t�I;��I;��I;R�I;EI;�SH;��F;�oD;�9A;>=;�8;RL2;o,;�%;j�;�<;�;�b;      �:?��:+��:�f�:���:E��:��;��;*#;1-;��5;�L<;3hA;cE;DlG;�H;'�I;��I;��I;��I;��I;&�I;(uI;�[I;�FI;�4I;�&I;kI;�I;�
I;�I;��H;E�H;��H;��H;��H;��H;��H;��H;��H;E�H;��H;�I;�
I;�I;jI;�&I;�4I;�FI;�[I;$uI;&�I;��I;��I;��I;��I;'�I;�H;ElG;cE;5hA;�L<;��5;1-;+#;��;��;A��:'��:�f�:)��:7��:      �Qɸ��J��+�8�(�9|�:��n:>�:dW�:���:N�;�;,�,;��6;�>;;5C;A�F;GvH;gwI;D�I;��I;k�I;��I;��I;�rI;�XI;nCI;!2I;b$I;I;&I;	I;yI;x�H;b�H;�H;��H;��H;��H;�H;d�H;x�H;{I;	I;#I;	I;a$I;!2I;nCI;�XI;�rI;��I;��I;h�I;��I;D�I;iwI;FvH;A�F;<5C;�>;��6;.�,;�;L�;���:jW�:@�:�n:��:�(�9�+�8��J�      Y+�G�%�"������1���T\�@�~���9��n:5��:fb�:�;�#;��0;��:;ǕA;S�E;�-H;4bI;��I;��I;��I;<�I;�I;�mI;5TI;@?I;k.I;!!I;�I;6I;�I;�I;2�H;��H;B�H;��H;B�H;��H;2�H;�I;�I;6I;�I;!I;k.I;=?I;5TI;�mI;�I;9�I;��I;��I;��I;4bI;�-H;U�E;ǕA;��:;��0;�#;�;bb�:5��:��n: �9@�~��T\��0������&��R�%�      �ݻ��ػ��ʻ\T������5�s�Ԯ0�*Tܺ$�=��V9�f:k��:�;B>;P,;�e8;�v@;U]E;aH;7bI;D�I;��I;s�I;ɭI;��I;7gI;6NI;:I;!*I;�I;�I;1I;mI;=I;}�H;��H;��H;��H;}�H;=I;kI;3I;�I;�I; *I;:I;3NI;9gI;��I;ƭI;o�I;��I;@�I;8bI;bH;W]E;�v@;�e8;S,;B>;�;m��:�f:�V9 �=�*TܺԮ0�1�s�����\T����ʻ��ػ      ��\�"�X�v-M���:��G#�T����ػP7��Z�����`!/��9p��:�m�:f;��(;�7;�@;T]E;�-H;dwI;��I;��I;��I;��I; }I;_I;GI;%4I;�%I;�I;I;~
I;tI;XI;a I;��H;a I;XI;tI;|
I;I;�I;�%I;"4I;GI;_I;}I;�I;��I;��I;��I;cwI;�-H;T]E;�@;�7;��(;f;�m�:p��:�9`!/�����Z�P7����ػR���G#���:�v-M�$�X�      ��ƼNü7_���۩�)$��9���Q�OG#��9�x����G��3��@�ȸ0�n:�l�:��;H�';�7;�v@;V�E;FvH;'�I;��I;�I;s�I;��I;�qI;�UI;g?I;.I;� I;HI;�I;	I;zI;"I;[I;"I;zI;	I;�I;HI;� I;.I;d?I;�UI;�qI;��I;s�I;�I;��I;)�I;DvH;W�E;�v@;�7;G�';��;�l�:0�n: �ȸ�3����G�y���9�OG#��Q�8��)$���۩�7_��Nü      �)���&�I<��3��� ��zܼ�*��琼��\�9 �4�ػh��M���Ϲ��J:�j�:��;��(;�e8;̕A;A�F;�H;R�I;��I;6�I;/�I;��I;�eI;�KI;N7I;�'I;I;EI; I;�I;I;bI;I;�I;I;EI;I;�'I;N7I;�KI;�eI;��I;1�I;9�I;��I;O�I;�H;@�F;͕A;�e8;��(;��;�j�:��J:��Ϲ�M�h�4�ػ9 ���\�琼�*���zܼ�� ��3�I<���&�      ~L��?ى��Ă�:�o�+T���5��G��V��^���Y����A�c �B������(����J:�l�:f;M,;��:;95C;ClG;EI;0�I;��I;��I;ƝI;�vI;�XI;xAI;�/I;D"I;I;�I;�I;1	I;�I;2	I;�I;�I;I;F"I;�/I;xAI;�XI;�vI;ÝI;��I;��I;,�I;EI;AlG;;5C;��:;M,;f;�l�:��J:(�����B���c ���A��Y���^���V��G���5�+T�:�o��Ă�?ى�      3�c�Խ�������0W��3�o�j??�4��9zܼzQ��2�X��Q��6�������Ϲ,�n:�m�:=>;��0;�>;`E;�SH;z�I;��I;��I;t�I;��I;gI;WLI;�7I;�(I;CI;*I;�I;SI;vI;SI;�I;(I;@I;�(I;�7I;XLI;gI;��I;r�I;��I;��I;v�I;�SH;aE;�>;��0;=>;�m�:,�n:��Ϲ����6���Q�2�X�zQ��9zܼ4��j??�3�o�0W���������Խc�      �7�~74�q�)�%>����3�m���08nc��)������ک�qa��Q�C����M�@�ȸp��:�;�#;��6;3hA;��F;�I;m�I;��I;E�I;��I;�uI;�WI;�@I;=/I;�"I;MI;6I;�I;�I;�I;6I;MI;�"I;;/I;�@I;�WI;�uI;��I;D�I;��I;n�I;�I;��F;2hA;��6;�#;�;v��:`�ȸ�M�B����Q�pa��ک������)�8nc�1m���3����%>�q�)�~74�      �S���7���X��Z�s��_S���0����Z�|���Ї|�j�5�k���ک�3�X�c �i􃻎3���9_��:�;)�,;�L<;�oD;;.H;��I;��I;��I;��I;��I;jcI;�II;6I;(I;�I;�I;�I;�I;�I;�I;I;�'I;6I;�II;jcI;��I;��I;��I;��I;��I;8.H;�oD;�L<;,�,;�;c��:0�9�3��i�c �3�X��ک�j��j�5�Ї|�|���Zཤ����0��_S�Z�s��X���7��      G���s�[D־�t��r���X��{�W�.�&��l��#N���Ă�j�5�����{Q����A�7�ػ��G�l!/��f:`b�:ݖ;��5;�9A;s�F;+I;	�I;	�I;>�I;��I;aoI;�RI;�<I;N-I;�!I;|I;6I;�I;5I;{I;�!I;N-I;�<I;�RI;aoI;��I;>�I;�I;�I;+I;o�F;�9A;��5;ߖ;^b�:�f:h!/���G�8�ػ��A�{Q������j�5��Ă�#N���l��.�&�{�W��X��r���t��[D־�s�      ��7�t�3��'��K�*�����̾%���Z�s�q74����#N��Ї|��)�:zܼ�Y��: �z������pV93��:H�;.-;==;�E;3�H;��I;a�I;��I;ޥI;K{I;�[I;�CI;�2I;H&I;I;aI;�I;_I;I;H&I;�2I;�CI;�[I;K{I;ۥI;��I;_�I;��I;6�H;�E;;=;.-;J�;/��:pV9����{��: ��Y��:zܼ�)�Ї|�#N�����q74�Z�s�%�����̾*����K��'�t�3�      (8��jڇ��x|�sm_�Iv<����B��n8��'6~�q74��l��|���9nc�5���^����\��9�%Z�H�=���n:���:"#;�8;��B;��G;�xI;��I;��I;��I;
�I;idI;�JI;�7I;M*I;l!I;�I;�I;~I;l!I;M*I;�7I;�JI;idI;�I;��I;��I;��I;�xI;��G;��B;�8;"#;���:��n:H�=�$Z��9���\��^��5��9nc�|����l��q74�'6~�n8��B�꾐��Iv<�sm_��x|�jڇ�      �ȿ�ÿ���-8��jڇ�Z��'�����n8��Z�s�.�&�Z�1j??��V�琼QG#�R7��2Tܺ��9XW�:��;PL2;w@;�F;0I;��I;��I;��I;q�I;�lI;QI;�<I;0.I;�$I;VI;{I;WI;�$I;0.I;�<I;QI;�lI;q�I;��I;��I;��I;/I;�F;t@;NL2;��;^W�:��90TܺP7��RG#�琼�V�j??�1Z�/�&�Z�s�n8�������'�Z�jڇ�-8������ÿ      ��	�&X�P����,ݿJ����ҕ��d��'�B��%���{�W����m���4�o��G��*���Q���ػ߮0���~�*�:��;e,;�=;kBE;ĬH;��I;��I;}�I;�I;�tI;�VI;AI;�1I;�'I;�!I; I;�!I;�'I;�1I;AI;�VI;�tI;�I;{�I;��I;��I;ĬH;pBE;�=;d,;��;2�:��~�߮0���ػ�Q��*���G�4�o�m������{�W�%���B�꾎'��d��ҕ�J����,ݿP���&X�      �5�821���#�O��u���ÿ�ҕ�Z������̾�X����0�3�1W����5��zܼ;��S��@�s��T\���n:%��:�%;��9;��C;/H;B�I;B�I;<�I;��I;�{I;>\I;EI;�4I;_*I;I$I;K"I;J$I;_*I;�4I;EI;A\I;�{I;��I;8�I;B�I;A�I;/H;��C;��9;�%;%��:��n:�T\�?�s�R��<���zܼ��5�1W��3佁�0��X����̾���Z��ҕ��ÿu��O����#�821�      1�j���c�y�P��5���u��J���jڇ�Iv<�*���r���_S��������+T��� �*$���G#�����1��x�:���:i�;L7;��B;��G;�I;F�I;��I;��I;��I;�`I;|HI;�7I;�,I;<&I;3$I;:&I;�,I;�7I;zHI;�`I;��I;�I;��I;F�I;�I;��G;��B;J7;j�;���:��:1�������G#�*$���� �+T���������_S�r��*���Iv<�jڇ�J���u�����5�y�P���c�      Ѣ��^���F���/]��5�O���,ݿ-8��sm_��K��t��Z�s�%>����;�o��3��۩���:�`T�������(�9�f�:�<;�_4;<hA;G8G;�dI;3�I;c�I;��I;��I;]dI;LKI;�9I;.I;�'I;�%I;�'I;.I;�9I;KKI;ZdI;��I;��I;`�I;3�I;�dI;L8G;=hA;�_4;�<;�f�:�(�9����`T����:��۩��3�;�o����%>�Z�s��t���K�sm_�-8���,ݿO���5��/]�F��^���      �����B����F��y�P���#�P�������x|��'�[D־�X��q�)� Խ�Ă�J<�8_��x-M���ʻ/��@)�8���:�;6K2;Ev@;��F;�FI;��I;=�I;S�I;2�I;�fI;pMI;v;I;�/I;�(I;�&I;�(I;�/I;v;I;oMI;�fI;2�I;R�I;<�I;��I;�FI;��F;Ev@;0K2;�;���:�)�8-����ʻx-M�8_��J<��Ă� Խq�)��X��[D־�'��x|����P�����#�y�P�F�����B��      ��������B��^�����c�821�&X��ÿjڇ�t�3��s��7��~74�d�?ى���&�Nü%�X���ػ`�%�@�J����:�b;��0;��?;H�F;�2I;�I;u�I;�I;z�I;�hI;�NI;d<I;�0I;�)I;�'I;�)I;�0I;d<I;�NI;�hI;z�I;�I;r�I;�I;�2I;H�F;��?;��0;�b;���:@�J�a�%���ػ$�X�Nü��&�?ى�d�~74��7���s�t�3�jڇ��ÿ&X�821���c�^����B�����      E(��s'���o��O�d��X1��x�Ŀ����3�z���x����4�o��[+���'���ü4yY��kٻ�o&���p����:u;��0;��?;�F;� I;/�I;��I;T�I;��I;�dI;�KI;�9I;�.I;�'I;�%I;�'I;�.I;�9I;�KI;�dI;��I;T�I;��I;/�I;� I;�F;��?;��0;x;���:@�p��o&��kٻ4yY���ü�'�[+��o�ཿ�4��x��z���3����Ŀ�x��X1�d�O��o��s'��      s'���X��f^�������]]���,�Q9�8g��V�����/����o��i1��hܽ���-$�_l���|U�Z�ԻT!� �,���:;�51;��?;|�F;\'I;��I;H�I;g�I;҆I;dI;qKI;�9I;V.I;�'I;�%I;�'I;X.I;�9I;oKI;dI;҆I;d�I;E�I;��I;\'I;|�F;��?;�51;;��: �,�T!�Z�Ի�|U�_l���-$����hܽi1��o���ྛ�/�V���8g��Q9���,��]]�����f^���X��      �o��f^���ē��4z�6K�j��T��(ﱿX�v��X#���Ѿń��&�r�нd̀�`��v���H�I��ǻ�4��#9#�:l�;6�2;��@;�F;;I;"�I;/�I;ƲI;��I;�bI;/JI;�8I;�-I;�&I;%I;�&I;�-I;�8I;/JI;�bI;��I;òI;,�I;"�I;;I;�F;��@;0�2;o�;#�:�#9�4��ǻH�I�v���`��d̀�r�н�&�ń���Ѿ�X#�X�v�(ﱿT��j��6K��4z��ē�f^��      O������4z���V��X1��<�wؿ����RZ��	�*���LUo����`y��0l�[��R��=�7�������Ƴ9>��:�;r�4;�tA;�2G;�XI;��I;��I;4�I;'�I;�_I;.HI;U7I;.,I;�%I;�#I;�%I;.,I;V7I;-HI;�_I;'�I;3�I;��I;��I;�XI;�2G;�tA;l�4;�;>��:�Ƴ9������=�7��R��[�0l�`y�����LUo�*����	��RZ����wؿ�<��X1���V��4z�����      d��]]�6K��X1�[f��pQ��V���]58��A���נ���O���b什�Q�	���>ߓ��� ��V��&氺t�":��:: ;17;8�B;q�G;|I;�I;��I;�I;n|I;l\I;}EI;N5I;j*I;a$I;]"I;a$I;i*I;N5I;{EI;l\I;l|I;ߧI;��I;�I;|I;p�G;6�B;17;: ;��:|�":*氺�V���� �>ߓ�	����Q�b什����O��נ��A��]58�V���pQ���[f��X1�6K��]]�      �X1���,�i���<��7g��g_���U�ς�،Ⱦ
ń�,�-�m��Q ��'�2�
?ټ\�{��!��n�l�O��u:Q ; &;K#:;r�C;3&H;A�I;T�I;��I;�I;�vI;XI;!BI;�2I;F(I;t"I;� I;t"I;F(I;�2I;!BI;XI;�vI;�I;��I;T�I;?�I;1&H;q�C;F#:; &;Q ; �u:p�O��n��!�]�{�
?ټ'�2�Q ��l��,�-�
ń�،Ⱦς��U�g_��7g��<�i����,�      �x�Q9�T��wؿpQ��g_��8�_��X#�t���f��<�S�{�����l�C�w���M���Ի��+� :T���:�e;�\,;0=;�BE;��H;��I;�I;��I;�I;�oI;�RI;D>I;�/I;�%I;' I;xI;& I;�%I;�/I;D>I;�RI;�oI;�I;��I;�I;��I;��H;�BE;0=;�\,;�e;��:`:T���+���Ի�M�w��C�l�����{�<�S��f��t���X#�8�_�g_��pQ��wؿT��Q9�      Ŀ8g��(ﱿ���V����U��X#�w��f���KUo�	�#��hܽ����n<����:����� ��᝻��Ժv�9���:�V;�2;� @;��F;I;*�I;r�I;_�I;��I;4hI;BMI;�9I;",I;�"I;�I;�I;�I;�"I;",I;�9I;CMI;4hI;��I;\�I;r�I;'�I;I;��F;� @;��2;�V;���:�u�9��Ժ�᝻�� �:�������n<�����hܽ	�#�KUo�f���w���X#��U�V������(ﱿ8g��      ���V���W�v��RZ�]58�ς�t��f���ioy�`1�bO��^什�`�O�����kyY���t�T�x�1�<�u:R��:p#;G98;4�B;��G;'mI;?�I;2�I;a�I;��I;`I;6GI;'5I;[(I;�I;�I;BI;�I;�I;[(I;'5I;7GI;`I;��I;`�I;1�I;;�I;)mI;��G;0�B;F98;p#;V��:4�u:|�1�r�T���kyY����O���`�^什bO��`1�ioy�f���t��ς�]58��RZ�W�v�V���      �3���/��X#��	��A��،Ⱦ�f��KUo�`1�ΰ��n��ռx��'��>ټ�@���k�����δ�P�39$�:XR;8e-;�/=;�	E;�xH;��I;@�I;��I;6�I;DvI;�WI;�@I;)0I;Z$I;uI;�I;mI;�I;uI;Z$I;'0I;�@I;�WI;FvI;4�I;��I;?�I;��I;�xH;�	E;�/=;8e-;XR;$�:P�39δ𺼼���k��@���>ټ�'�ռx�n��ΰ��`1�KUo��f��،Ⱦ�A���	��X#���/�      z���྅�Ѿ*����נ�
ń�<�S�	�#�bO��n��K̀���2����}�>��Իh�B�(#��m:0H�:� ;ȼ5;�FA;��F;�I;��I;��I;׾I;��I;�jI;�NI;C:I;+I;1 I;I;�I;�I;�I;I;1 I;+I;F:I;�NI;�jI;��I;׾I;��I;��I;�I;��F;�FA;ȼ5;� ;,H�:�m:#�k�B��Ի}�>�������2�K̀�n��bO��	�#�<�S�
ń��נ�*�����Ѿ��      �x���o��ń�LUo���O�,�-�{��hܽ^什ռx���2�tb��TR��Q|U�N2��)���鰺�v�9�:@D;��,;�h<;�rD;~%H;��I;��I;�I;:�I;>�I;_I;?FI;�3I;�%I;I;�I;�I;lI;�I;�I;I;�%I;�3I;?FI;_I;<�I;:�I;�I;��I;��I;{%H;�rD;�h<;��,;=D;�:�v�9�鰺*��N2��Q|U�TR��tb����2�ռx�^什�hܽ{�,�-���O�LUo�ń��o��      ��4�i1��&������l�཈�������`��'���TR��@�]�y��V���X���=o����:��;\#;H�6;�tA;��F;�	I;��I;�I;��I;L�I;qI;�SI;�=I;�,I;� I;�I;�I;xI;tI;zI;�I;�I;� I;�,I;�=I;�SI;qI;L�I;��I;�I;��I;�	I;��F;�tA;H�6;Z#;��;���:�>o��X��V��y��@�]�TR����'��`��������l��������&�i1�      n�ཹhܽq�н_y��b什Q ��l��n<�N���>ټ��P|U�y������f1�x�����u:�l�:4�;�71;�)>;�	E;AJH;��I;��I;��I;�I;�I;�bI;�HI;^5I;�&I;�I;�I;uI;WI;V
I;WI;tI;�I;�I;�&I;a5I;�HI;�bI;�I;�I;��I;��I;��I;=JH;�	E;�)>;�71;5�;�l�:��u:x���d1�����y��Q|U����>ټN���n<�l�Q ��b什_y��q�н�hܽ      Z+����d̀�/l��Q�'�2�C��������@��}�>�N2��V��f1�`��$R:���:;�\,;l;;<C;�eG;�9I;��I;i�I;��I;w�I;�qI;�TI;�>I;o-I;d I;�I;�I;I;II;HI;II;I;�I;�I;e I;p-I;�>I;�TI;�qI;t�I;�I;i�I;��I;�9I;�eG;<C;n;;�\,;;���:�$R:`��g1�V��N2��}�>��@��������C�&�2��Q�/l�d̀���      �'��-$�`��Z����	?ټw��:���hyY��k��Ի)���X��x����$R:��:�R;�);�8;��A;��F;h�H;_�I;��I;��I;�I;?�I;aI;*HI;�4I;�%I;~I;I;�I;�I;JI;}I;JI;�I;�I;I;~I;�%I;�4I;&HI;aI;<�I;�I;��I;��I;[�I;h�H;��F;��A;�8;�);�R;��:�$R:p����X��)���Ի�k�hyY�:���w��?ټ	���Z�_���-$�      ��ü\l��u����R��=ߓ�Z�{��M��� ��컹���d�B��鰺�=o���u:��:�R;`�';D17;�@;4�E;�lH;e�I;��I;��I;A�I;��I;mI;�QI;a<I;�+I;�I;�I;�I;I;|I;bI;�I;bI;|I;I;�I;�I;�I;�+I;^<I;�QI;�lI;��I;A�I;��I;��I;e�I;�lH;4�E;�@;F17;^�';�R;��:��u:�=o��鰺g�B������컅� ��M�Z�{�=ߓ��R��u���^l��      4yY��|U�E�I�:�7��� ��!���Ի�᝻n�T�ʴ�#��v�9���:�l�:;�);B17;^ @;m]E;�$H;�kI;@�I;��I;/�I;f�I;�wI;�ZI;�CI;�1I;�#I;aI;�I;h	I;�I;oI;��H;7�H;��H;oI;�I;f	I;�I;aI;�#I;�1I;�CI;�ZI;�wI;f�I;*�I;��I;@�I;�kI;�$H;m]E;^ @;A17;�);;�l�:���:�v�9#�ʴ�n�T��᝻��Ի�!��� �:�7�F�I��|U�      �kٻU�Իwǻ ����V���n���+��ԺP�1���39�m:�:��;9�;�\,;�8;�@;p]E;�
H;�VI;��I;#�I;)�I;��I;<�I;�bI;�JI;^7I;(I;�I;gI;I;sI;pI;��H;�H;��H;�H;��H;pI;qI;I;iI;�I;(I;]7I;�JI;�bI;<�I;��I;#�I;"�I;��I;�VI;�
H;q]E;�@;�8;�\,;9�;��;�:�m:��39P�1��Ժ��+��n��V�� ���wǻV�Ի      �o&�<!��4����$氺d�O� :T��u�9H�u:	$�:8H�:@D;Z#;�71;m;;��A;1�E;�$H;�VI;G�I;��I;K�I;��I;4�I;FiI;ePI;X<I;1,I;YI;�I;�I;�I;�I;j�H;�H;��H;A�H;��H;�H;j�H;�I;�I;�I;�I;UI;1,I;V<I;bPI;FiI;.�I;��I;K�I;��I;G�I;�VI;�$H;1�E;��A;l;;�71;Z#;=D;2H�:$�:@�u:v�9 :T�`�O�氺���4�F!�      ��p� �,��$9�Ƴ9p�":<�u:��:���:^��:\R;� ;��,;H�6;�)>;<C;��F;�lH;�kI;��I;��I;��I;R�I;��I;�mI;�TI;b@I;�/I;]"I;�I;�I;I;�I;��H;��H;��H;��H;�H;��H;��H;��H;��H;�I;I;�I;�I;]"I;�/I;b@I;�TI;�mI;��I;R�I;��I;��I;��I;�kI;�lH;��F;<C;�)>;H�6;��,;� ;[R;\��:���:��:H�u:p�":�Ƴ9�$9 �,�      ���:��:I�::��:��:"Q ;�e;�V;z#;:e-;ϼ5;�h<;�tA;�	E;�eG;h�H;g�I;A�I;#�I;K�I;O�I;/�I;ApI;�WI;*CI;|2I;�$I;�I;�I;	I;�I;3�H;��H;;�H;��H;i�H;�H;i�H;��H;<�H;��H;3�H;�I;}	I;�I;�I;�$I;~2I;,CI;�WI;<pI;/�I;N�I;N�I;#�I;C�I;d�I;e�H;�eG;�	E;�tA;�h<;̼5;:e-;z#;�V;�e;$Q ;E��::��:I�:��:      �; ;x�;�;6 ;&;�\,;�2;O98;�/=;�FA;�rD;��F;EJH;�9I;^�I;��I;��I;)�I;��I;��I;CpI;�XI;�DI;%4I;�&I;^I;$I;�
I;�I;��H;��H;'�H;�H;s�H;��H;F�H;��H;s�H;�H;&�H;��H;��H;�I;�
I;$I;\I;�&I;&4I;�DI;�XI;BpI;��I;��I;)�I;��I;��I;]�I;�9I;DJH;��F;�rD;�FA;�/=;M98;�2;�\,;&;@ ;�;y�;;      �0;�51;B�2;|�4;17;O#:;)0=;� @;;�B;�	E;��F;�%H;�	I;��I;��I;��I;��I;0�I;��I;3�I;�mI;�WI;�DI;�4I;{'I;oI;>I;�I;sI;l I;k�H;�H;��H;��H;��H;��H;��H;��H;��H;��H;��H;�H;l�H;i I;qI;�I;=I;nI;|'I;�4I;�DI;�WI;�mI;3�I;��I;1�I;��I;��I;��I;��I;�	I;�%H;��F;�	E;:�B;� @;'0=;Q#:;17;y�4;@�2;�51;      Ƕ?;��?;��@;�tA;:�B;x�C;�BE;��F;��G;�xH;�I;��I;��I;��I;l�I;��I;H�I;g�I;C�I;LiI;�TI;-CI;*4I;�'I;�I;�I;QI;I;� I;��H;S�H;��H;��H;�H;�H;b�H;/�H;b�H;�H;�H;��H;��H;T�H;��H;� I;I;PI;�I;�I;}'I;'4I;/CI;�TI;MiI;C�I;i�I;D�I;��I;l�I;��I;��I;��I;�I;�xH;��G;��F;�BE;v�C;<�B;�tA;��@;��?;      �F;��F;�F;�2G;s�G;1&H;��H;I;-mI;��I;��I;��I;�I;��I;�I;�I;��I;�wI;�bI;bPI;`@I;{2I;�&I;nI;�I;}I;]I;<I;�H;��H;��H;��H;��H;b�H;��H;
�H;��H;
�H;��H;c�H;��H;��H;��H;��H;�H;=I;\I;}I;�I;kI;�&I;{2I;[@I;bPI;�bI;�wI;��I;�I;��I;��I;�I;��I;��I;��I;,mI;I;��H;1&H;w�G;�2G;�F;��F;      � I;c'I;;I;�XI;|I;I�I;��I;)�I;E�I;D�I;��I;�I;��I; �I;x�I;?�I;mI;�ZI;�JI;Z<I;�/I;�$I;`I;AI;MI;_I;DI;(�H;��H;��H;��H;��H;�H;��H;R�H;��H;��H;��H;P�H;��H;�H;��H;��H;��H;��H;*�H;CI;]I;QI;@I;\I;�$I;�/I;Z<I;�JI;�ZI;mI;=�I;x�I; �I;��I;�I;��I;B�I;F�I;*�I;��I;F�I; |I;�XI;;I;`'I;      &�I;��I;,�I;��I;�I;W�I;�I;|�I;9�I;��I;޾I;A�I;P�I;�I;�qI;aI;�QI;�CI;^7I;3,I;]"I;�I;'I;�I;I;?I;(�H;��H;��H;��H;��H;��H;��H;��H;�H;��H;��H;��H;�H;��H;��H;��H;��H;��H;��H;��H;(�H;?I;I;�I;$I;�I;["I;4,I;^7I;�CI;�QI;aI;�qI;�I;O�I;A�I;ݾI;��I;9�I;}�I;�I;W�I;!�I;��I;*�I;��I;      �I;K�I;,�I;��I;��I;��I;��I;a�I;f�I;9�I;��I;C�I;qI;�bI;�TI;*HI;e<I;�1I;(I;ZI;�I;�I;�
I;vI;� I;�H;��H;��H;��H;��H;��H;��H;|�H;��H;$�H;��H;��H;��H;$�H;��H;{�H;��H;��H;��H;��H;��H;��H;�H;� I;wI;�
I;�I;�I;YI;(I;�1I;d<I;*HI;�TI;�bI;qI;B�I;��I;8�I;f�I;a�I;��I;��I;��I;��I;+�I;=�I;      b�I;q�I;вI;;�I;�I;�I;�I;��I;��I;NvI;�jI;_I;�SI;�HI;�>I;�4I;�+I;�#I;�I;I;�I;~	I;�I;l I;��H;��H;��H;��H;��H;��H;j�H;O�H;s�H;��H;M�H;
�H;��H;
�H;M�H;��H;q�H;Q�H;j�H;��H;��H;��H;��H;��H;��H;l I;�I;~	I;�I;I;�I;�#I;�+I;�4I;�>I;�HI;�SI;_I;�jI;NvI;��I;��I;�I;�I;�I;:�I;ʲI;n�I;      ��I;�I;��I;6�I;z|I;�vI;�oI;:hI;`I;�WI;�NI;JFI;�=I;h5I;w-I;�%I;�I;bI;nI;I;I;�I;��H;n�H;N�H;��H;��H;��H;��H;m�H;J�H;M�H;��H;�H;��H;n�H;0�H;n�H;��H;�H;��H;N�H;J�H;k�H;��H;��H;��H;��H;Q�H;n�H;��H;�I;I;I;nI;bI;�I;�%I;v-I;f5I;�=I;HFI;�NI;�WI;`I;;hI;�oI;�vI;w|I;5�I;��I;�I;      �dI;dI;�bI;`I;p\I;
XI;�RI;JMI;=GI;�@I;J:I;�3I;-I;�&I;n I;�I;I;�I;I;�I;�I;7�H;��H; �H;��H;��H;��H;��H;��H;Q�H;L�H;��H;��H;e�H;�H;��H;��H;��H;�H;e�H;��H;��H;L�H;R�H;��H;��H;��H;��H;��H; �H;��H;9�H;�I;�I;I;�I;I;�I;n I;�&I;-I;�3I;J:I;�@I;=GI;JMI;�RI;XI;o\I;`I;�bI;dI;      �KI;�KI;9JI;:HI;�EI;"BI;D>I;�9I;/5I;*0I;+I;�%I;� I;�I;�I;I;�I;c	I;wI;�I;��H;��H;&�H;��H;��H;��H;�H;��H;�H;w�H;��H;��H;P�H;��H;��H;[�H;j�H;[�H;��H;��H;N�H;��H;��H;x�H;��H;��H;�H;��H;��H;��H;$�H;��H;��H;�I;wI;e	I;�I;I;�I;�I;� I;�%I;+I;*0I;.5I;�9I;D>I;%BI;EI;:HI;:JI;{KI;      :I;�9I;�8I;c7I;Z5I;�2I;�/I;-,I;b(I;^$I;: I;I;�I;�I;�I;�I;'I;�I;xI;q�H;��H;=�H;	�H;��H;�H;a�H;��H;��H;��H;��H;�H;d�H;��H;x�H;5�H;�H;��H;�H;5�H;x�H;��H;g�H;�H;��H;��H;��H;��H;_�H;�H;��H;�H;=�H;��H;q�H;xI;�I;&I;�I;�I;�I;�I;I;7 I;]$I;d(I;-,I;�/I;�2I;P5I;c7I;�8I;�9I;      �.I;m.I;�-I;<,I;�*I;F(I;�%I;�"I;�I;zI;I;�I;�I;|I;I;�I;�I;mI;��H;�H;��H;��H;t�H;��H;��H;��H;O�H;�H;$�H;M�H;��H;�H;��H;9�H;��H;��H;��H;��H;��H;9�H;��H;�H;��H;P�H;'�H;�H;N�H;��H;��H;��H;s�H;��H;��H;�H;��H;oI;�I;�I;I;~I;�I;�I;I;|I;�I;�"I;�%I;I(I;z*I;<,I;�-I;d.I;      �'I;�'I;�&I;�%I;u$I;t"I;. I;�I;�I;�I;�I;�I;�I;dI;PI;QI;mI;��H;$�H;��H;��H;j�H;��H;��H;_�H;�H;��H;��H;��H;�H;o�H;��H;X�H;�H;��H;��H;��H;��H;��H;�H;X�H;��H;o�H;
�H;��H;��H;��H;�H;a�H;��H;��H;j�H;��H;��H;$�H;��H;kI;QI;PI;cI;�I;�I;�I;�I;�I;�I;. I;x"I;k$I;�%I;�&I;�'I;      �%I;�%I;%I;�#I;j"I;� I;{I;�I;II;mI;�I;uI;xI;_
I;LI;�I;�I;2�H;��H;G�H;�H;�H;H�H;��H;+�H;��H;��H;��H;��H;��H;6�H;��H;j�H;��H;��H;��H;��H;��H;��H;��H;i�H;��H;6�H;��H;��H;��H;��H;��H;+�H;��H;H�H;�H;�H;G�H;��H;3�H;�I;�I;LI;_
I;xI;uI;�I;pI;JI;�I;{I;� I;`"I;�#I;%I;�%I;      �'I;�'I;�&I;�%I;u$I;t"I;. I;�I;�I;�I;�I;�I;�I;dI;PI;QI;mI;��H;$�H;��H;��H;j�H;��H;��H;a�H;�H;��H;��H;��H;�H;o�H;��H;X�H;�H;��H;��H;��H;��H;��H;�H;X�H;��H;o�H;
�H;��H;��H;��H;�H;_�H;��H;��H;j�H;��H;��H;$�H;��H;kI;QI;PI;cI;�I;�I;�I;�I;�I;�I;. I;x"I;k$I;�%I;�&I;�'I;      �.I;m.I;�-I;<,I;�*I;F(I;�%I;�"I;�I;zI;I;�I;�I;|I;I;�I;�I;mI;��H;�H;��H;��H;t�H;��H;��H;��H;O�H;�H;&�H;M�H;��H;�H;��H;9�H;��H;��H;��H;��H;��H;9�H;��H;�H;��H;O�H;'�H;�H;N�H;��H;��H;��H;s�H;��H;��H;�H;��H;oI;�I;�I;I;~I;�I;�I;I;|I;�I;�"I;�%I;J(I;z*I;<,I;�-I;d.I;      :I;�9I;�8I;c7I;X5I;�2I;�/I;,,I;b(I;]$I;8 I;I;�I;�I;�I;�I;'I;�I;xI;q�H;��H;=�H;	�H;��H;�H;b�H;��H;��H;��H;��H;�H;d�H;��H;x�H;5�H;�H;��H;�H;5�H;x�H;��H;g�H;�H;��H;��H;��H;��H;a�H;�H;��H;�H;=�H;��H;q�H;xI;�I;&I;�I;�I;�I;�I;I;: I;^$I;e(I;.,I;�/I;�2I;N5I;c7I;�8I;�9I;      �KI;�KI;<JI;<HI;�EI;"BI;D>I;�9I;/5I;)0I;+I;�%I;� I;�I;�I;I;�I;e	I;wI;�I;��H;��H;&�H;��H;��H;��H;�H;��H;�H;w�H;��H;��H;O�H;��H;��H;[�H;j�H;[�H;��H;��H;N�H;��H;��H;x�H;��H;��H;�H;��H;��H;��H;$�H;��H;��H;�I;wI;c	I;�I;I;�I;�I;� I;�%I;+I;,0I;/5I;�9I;D>I;$BI;EI;;HI;9JI;�KI;      �dI;dI;�bI; `I;r\I;
XI;�RI;JMI;=GI;�@I;J:I;�3I;-I;�&I;n I;�I;I;�I;I;�I;�I;9�H;��H; �H;��H;��H;��H;��H;��H;Q�H;L�H;��H;��H;e�H;�H;��H;��H;��H;�H;e�H;��H;��H;L�H;R�H;��H;��H;��H;��H;��H; �H;��H;7�H;�I;�I;I;�I;I;�I;n I;�&I;-I;�3I;J:I;�@I;>GI;JMI;�RI;XI;o\I; `I;�bI;dI;      ��I;�I;��I;5�I;z|I;�vI;�oI;:hI;`I;�WI;�NI;HFI;�=I;h5I;v-I;�%I;�I;aI;nI;I;I;�I;��H;o�H;Q�H;��H;��H;��H;��H;m�H;J�H;M�H;��H;�H;��H;n�H;0�H;n�H;��H;�H;��H;M�H;J�H;k�H;��H;��H;��H;��H;N�H;o�H;��H;�I;I;I;nI;dI;�I;�%I;w-I;i5I;�=I;JFI;�NI;�WI;`I;;hI;�oI;�vI;y|I;6�I;��I;�I;      [�I;p�I;ϲI;:�I;�I;�I;�I;��I;��I;MvI;�jI;_I;�SI;�HI;�>I;�4I;�+I;�#I;�I;I;�I;~	I;�I;l I;��H;��H;��H;��H;��H;��H;j�H;O�H;s�H;��H;M�H;
�H;��H;
�H;M�H;��H;s�H;Q�H;j�H;��H;��H;��H;��H;��H;��H;l I;�I;~	I;�I;I;�I;�#I;�+I;�4I;�>I;�HI;�SI;_I;�jI;NvI;��I;��I;�I;�I;�I;:�I;ϲI;r�I;      	�I;G�I;1�I;��I;��I;��I;��I;a�I;f�I;8�I;��I;C�I;qI;�bI;�TI;*HI;e<I;�1I;(I;ZI;�I;�I;�
I;vI;� I;�H;��H;��H;��H;��H;��H;��H;{�H;��H;#�H;��H;��H;��H;$�H;��H;{�H;��H;��H;��H;��H;��H;��H;�H;� I;wI;�
I;�I;�I;ZI;(I;�1I;d<I;,HI;�TI;�bI;qI;C�I;��I;9�I;f�I;c�I;��I;��I;��I;��I;1�I;G�I;      &�I;��I;,�I;��I;�I;W�I;�I;z�I;9�I;��I;޾I;A�I;O�I;�I;�qI;aI;�QI;�CI;^7I;4,I;`"I;�I;'I;�I;I;?I;(�H;��H;��H;��H;��H;��H;��H;��H;�H;��H;��H;��H;�H;��H;��H;��H;��H;��H;��H;��H;(�H;?I;I;�I;$I;�I;["I;4,I;^7I;�CI;�QI;aI;�qI;�I;P�I;A�I;ݾI;��I;:�I;~�I;�I;T�I;#�I;��I;*�I;��I;      � I;a'I;;I;�XI;|I;E�I;��I;)�I;E�I;C�I;��I;�I;��I; �I;x�I;?�I;mI;�ZI;�JI;[<I;�/I;�$I;^I;@I;QI;`I;DI;*�H;��H;��H;��H;��H;�H;��H;P�H;��H;��H;��H;R�H;��H;�H;��H;��H;��H;��H;(�H;CI;_I;MI;>I;]I;�$I;�/I;Z<I;�JI;�ZI;mI;=�I;x�I; �I;��I;�I;��I;C�I;E�I;*�I;��I;D�I;|I;�XI;;I;V'I;      �F;��F;�F;�2G;s�G;3&H;��H;I;,mI;��I;��I;��I;�I;��I;��I;�I;��I;�wI;�bI;bPI;a@I;{2I;�&I;lI;�I;}I;]I;=I;�H;��H;��H;��H;��H;c�H;��H;
�H;��H;
�H;��H;b�H;��H;��H;��H;��H;�H;<I;\I;}I;�I;kI;�&I;{2I;[@I;bPI;�bI;�wI;��I;�I;�I;��I;�I;��I;��I;��I;*mI;I;��H;1&H;x�G;�2G;�F;��F;      Ƕ?;��?;��@;�tA;:�B;x�C;�BE;��F;��G;�xH;�I;��I;��I;��I;l�I;��I;F�I;g�I;C�I;MiI;�TI;/CI;*4I;�'I;�I;�I;QI;I;� I;��H;T�H;��H;��H;�H;�H;b�H;/�H;b�H;�H;�H;��H;��H;S�H;��H;� I;I;PI;�I;�I;'I;'4I;-CI;�TI;MiI;C�I;j�I;F�I;��I;l�I;��I;��I;��I;�I;�xH;��G;��F;�BE;x�C;9�B;�tA;��@;��?;      �0;�51;E�2;v�4;17;U#:;#0=;� @;=�B;�	E;��F;�%H;�	I;��I;��I;��I;��I;0�I;��I;3�I;�mI;�WI;�DI;�4I;|'I;oI;>I;�I;tI;l I;l�H;�H;��H;��H;��H;��H;��H;��H;��H;��H;��H;�H;k�H;i I;qI;�I;=I;oI;{'I;�4I;�DI;�WI;�mI;4�I;��I;1�I;��I;��I;��I;��I;�	I;�%H;��F;�	E;;�B;� @;#0=;U#:;17;y�4;E�2;�51;      ;*;��;�;6 ;&;�\,;�2;N98;�/=;�FA;�rD;��F;DJH;�9I;^�I;��I;��I;)�I;��I;��I;BpI;�XI;�DI;&4I;�&I;^I;$I;�
I;�I;��H;��H;'�H;�H;s�H;��H;F�H;��H;s�H;�H;&�H;��H;��H;�I;�
I;$I;\I;�&I;%4I;�DI;�XI;CpI;��I;��I;)�I;��I;��I;^�I;�9I;EJH;��F;�rD;�FA;�/=;N98;�2;�\,;
&;< ;�;|�;;      ���:��:I�::��:��:"Q ;�e;�V;z#;:e-;ͼ5;�h<;�tA;�	E;�eG;f�H;d�I;A�I;#�I;L�I;P�I;/�I;ApI;�WI;,CI;~2I;�$I;�I;�I;	I;�I;3�H;��H;<�H;��H;i�H;�H;i�H;��H;;�H;��H;3�H;�I;{	I;�I;�I;�$I;~2I;*CI;�WI;>pI;/�I;N�I;N�I;#�I;C�I;e�I;h�H;�eG;�	E;�tA;�h<;ͼ5;:e-;z#;�V;�e;"Q ;K��::��:I�:��:      ��p� �,� %9�Ƴ9l�":(�u:��:���:\��:[R;� ;��,;H�6;�)>;<C;��F;�lH;�kI;��I;��I;��I;R�I;��I;�mI;�TI;d@I;�/I;]"I;�I;�I;I;�I;��H;��H;��H;��H;�H;��H;��H;��H;��H;�I;I;�I;�I;]"I;�/I;b@I;�TI;�mI;��I;R�I;��I;��I;��I;�kI;�lH;��F;<C;�)>;H�6;��,;� ;YR;^��:���:��:H�u:��":�Ƴ9�$9 �,�      �o&�<!��4����氺d�O� :T�v�9L�u:	$�:2H�:=D;Z#;�71;l;;��A;1�E;�$H;�VI;F�I;��I;K�I;��I;3�I;FiI;dPI;X<I;1,I;YI;�I;�I;�I;�I;j�H;�H;��H;A�H;��H;�H;j�H;�I;�I;�I;�I;SI;1,I;V<I;dPI;FiI;.�I;��I;K�I;��I;I�I;�VI;�$H;1�E;��A;m;;�71;Z#;=D;6H�:$�:L�u: v�9 :T�X�O�氺���4�H!�      �kٻU�Իxǻ ����V���n���+��ԺT�1���39�m:�:��;9�;�\,;�8;�@;p]E;�
H;�VI;��I;"�I;)�I;��I;<�I;�bI;�JI;]7I;(I;�I;iI;I;sI;pI;��H;�H;��H;�H;��H;pI;qI;I;gI;�I;(I;^7I;�JI;�bI;<�I;��I;#�I;#�I;��I;�VI;�
H;q]E;�@;�8;�\,;9�;��;�:�m:��39P�1��Ժ��+��n��V�� ���wǻV�Ի      3yY��|U�E�I�;�7��� ��!���Ի�᝻n�T�̴�#��v�9���:�l�:;�);D17;] @;m]E;�$H;�kI;@�I;��I;-�I;f�I;�wI;�ZI;�CI;�1I;�#I;aI;�I;h	I;�I;oI;��H;7�H;��H;oI;�I;f	I;�I;aI;�#I;�1I;�CI;�ZI;�wI;f�I;)�I;��I;@�I;�kI;�$H;m]E;` @;B17;�);;�l�:���:�v�9#�ʴ�n�T��᝻��Ի�!��� �:�7�F�I��|U�      ��ü\l��u����R��=ߓ�Z�{��M��� ��컹���e�B��鰺�=o���u:��:�R;`�';D17;�@;3�E;�lH;e�I;��I;��I;@�I;��I;mI;�QI;a<I;�+I;�I;�I;�I;I;|I;bI;�I;bI;|I;I;�I;�I;�I;�+I;^<I;�QI;�lI;��I;A�I;��I;��I;e�I;�lH;5�E;�@;F17;`�';�R;��:��u:�=o��鰺d�B������컅� ��M�Z�{�=ߓ��R��u���^l��      �'��-$�`��Z����	?ټw��:���hyY��k��Ի)���X��x����$R:��:�R;�);�8;��A;��F;h�H;^�I;��I;��I;�I;?�I;aI;*HI;�4I;�%I;|I;I;�I;�I;JI;}I;JI;�I;�I;I;I;�%I;�4I;&HI;aI;;�I;�I;��I;��I;[�I;h�H;��F;��A;�8;�);�R;��:�$R:x����X��)���Ի�k�hyY�:���w��?ټ���Z�`���-$�      Z+����d̀�/l��Q�'�2�C��������@��}�>�N2��V��g1�`��$R:���:;�\,;m;;<C;�eG;�9I;��I;i�I;�I;u�I;�qI;�TI;�>I;p-I;b I;�I;�I;I;II;HI;II;I;�I;�I;g I;o-I;�>I;�TI;�qI;u�I;�I;i�I;��I;�9I;�eG;<C;m;;�\,;;���:�$R:`��f1�V��N2��}�>��@��������C�&�2��Q�/l�d̀���      n�ཹhܽq�н_y��b什Q ��l��n<�N���>ټ��Q|U�y������d1�x�����u:�l�:5�;�71;�)>;�	E;AJH;��I;��I;��I;�I;�I;�bI;�HI;a5I;�&I;�I;�I;tI;WI;V
I;WI;uI;�I;�I;�&I;^5I;�HI;�bI;�I;�I;��I;��I;��I;=JH;�	E;�)>;�71;4�;�l�:��u:x���f1�����y��P|U����>ټN���n<�l�Q ��b什_y��q�н�hܽ      ��4�i1��&������l�཈�������`��'���TR��@�]�y��V���X���=o����:��;Z#;F�6;�tA;��F;�	I;��I;�I;��I;L�I;qI;�SI;�=I;�,I;� I;�I;�I;zI;tI;xI;�I;�I;� I;�,I;�=I;�SI;qI;L�I;��I;�I;��I;�	I;��F;�tA;H�6;Z#;��;���:@>o��X��V��y��@�]�TR����'��`��������l��������&�i1�      �x���o��ń�LUo���O�,�-�{��hܽ^什ռx���2�tb��TR��Q|U�N2��*���鰺�v�9�:=D;��,;�h<;�rD;~%H;��I;��I;�I;:�I;>�I;_I;?FI;�3I;�%I;
I;�I;�I;lI;�I;�I;I;�%I;�3I;?FI;_I;<�I;:�I;�I;��I;��I;{%H;�rD;�h<;��,;?D;�:�v�9�鰺*��N2��Q|U�TR��tb����2�ռx�^什�hܽ{�,�-���O�LUo�ń��o��      z���྅�Ѿ*����נ�
ń�<�S�	�#�bO��n��K̀���2����}�>��Իh�B� #��m:2H�:� ;ȼ5;�FA;��F;�I;��I;��I;׾I;��I;�jI;�NI;C:I;+I;1 I;I;�I;�I;�I;I;1 I;+I;D:I;�NI;�jI;��I;׾I;��I;��I;�I;��F;�FA;ȼ5;� ;0H�:�m:#�j�B��Ի}�>�������2�K̀�n��bO��	�#�<�S�
ń��נ�*�����Ѿ��      �3���/��X#��	��A��،Ⱦ�f��KUo�`1�ΰ��n��ռx��'��>ټ�@���k�����Ҵ�P�39$�:WR;8e-;�/=;�	E;�xH;��I;@�I;��I;6�I;DvI;�WI;�@I;'0I;Z$I;uI;�I;mI;�I;uI;Z$I;'0I;�@I;�WI;DvI;4�I;��I;?�I;��I;�xH;�	E;�/=;8e-;XR;$�:P�39ʴ𺼼���k��@���>ټ�'�ռx�n��ΰ��`1�KUo��f��،Ⱦ�A���	��X#���/�      ���V���W�v��RZ�]58�ς�t��f���ioy�`1�bO��^什�`�O�����kyY���t�T�|�1�<�u:P��:p#;G98;3�B;��G;'mI;?�I;1�I;c�I;��I;`I;6GI;(5I;[(I;�I;�I;BI;�I;�I;[(I;&5I;4GI;`I;��I;`�I;2�I;;�I;'mI;��G;0�B;F98;p#;V��:<�u:x�1�r�T���kyY����O���`�^什bO��`1�ioy�f���t��ς�]58��RZ�W�v�V���      Ŀ8g��(ﱿ���V����U��X#�w��f���KUo�	�#��hܽ����n<����:����� ��᝻��Ժv�9���:�V; �2;� @;��F;I;*�I;r�I;_�I;��I;4hI;BMI;�9I;#,I;�"I;�I;�I;�I;�"I;#,I;�9I;BMI;4hI;��I;\�I;r�I;'�I;I;��F;� @; �2;�V;���:�u�9��Ժ�᝻�� �:�������n<�����hܽ	�#�KUo�f���w���X#��U�V������(ﱿ8g��      �x�Q9�T��wؿpQ��g_��8�_��X#�t���f��<�S�{�����l�C�w���M���Ի��+�P:T���:�e;�\,;0=;�BE;��H;��I;�I;��I;�I;�oI;�RI;F>I;�/I;�%I;& I;xI;' I;�%I;�/I;C>I;�RI;�oI;�I;��I;�I;��I;��H;�BE;0=;�\,;�e;��:P:T���+���Ի�M�w��C�l�����{�<�S��f��t���X#�8�_�g_��pQ��wؿT��Q9�      �X1���,�i���<��7g��g_���U�ς�،Ⱦ
ń�,�-�l��Q ��'�2�
?ټ\�{��!��n�p�O��u:Q ;�&;J#:;q�C;3&H;A�I;T�I;��I;�I;�vI;XI;"BI;�2I;F(I;t"I;� I;u"I;F(I;�2I; BI;XI;�vI;�I;��I;T�I;?�I;1&H;r�C;G#:; &;Q ; �u:p�O��n��!�]�{�
?ټ'�2�Q ��m��,�-�
ń�،Ⱦς��U�g_��7g��<�i����,�      d��]]�6K��X1�[f��pQ��V���]58��A���נ���O���b什�Q�
���>ߓ��� ��V��*氺p�":��:: ;17;6�B;q�G;|I;�I;��I;�I;l|I;k\I;}EI;N5I;j*I;a$I;]"I;a$I;i*I;N5I;{EI;l\I;n|I;�I;��I;�I;|I;p�G;8�B;	17;: ;��:|�":*氺�V���� �>ߓ�	����Q�b什����O��נ��A��]58�V���pQ���[f��X1�6K��]]�      O������4z���V��X1��<�wؿ����RZ��	�*���LUo����`y��0l�[��R��=�7�������Ƴ9>��:�;r�4;�tA;�2G;�XI;��I;��I;6�I;'�I;�_I;.HI;V7I;.,I;�%I;�#I;�%I;.,I;U7I;-HI;�_I;'�I;3�I;��I;��I;�XI;�2G;�tA;l�4;�;>��:�Ƴ9������<�7��R��[�0l�`y�����LUo�*����	��RZ����wؿ�<��X1���V��4z�����      �o��f^���ē��4z�6K�i��T��(ﱿX�v��X#���Ѿń��&�r�нd̀�`��v���H�I��ǻ�4��#9#�:l�;6�2;��@;�F;;I;"�I;/�I;ƲI;��I;�bI;/JI;�8I;�-I;�&I;%I;�&I;�-I;�8I;/JI;�bI;��I;òI;,�I;"�I;;I;�F;��@;0�2;q�;#�:�#9�4��ǻH�I�v���a��d̀�r�н�&�ń���Ѿ�X#�X�v�(ﱿT��i��6K��4z��ē�f^��      s'���X��f^�������]]���,�Q9�8g��V�����/����o��i1��hܽ���-$�_l���|U�Z�ԻT!� �,���:;�51;��?;|�F;\'I;��I;H�I;g�I;҆I;dI;qKI;�9I;V.I;�'I;�%I;�'I;X.I;�9I;oKI;dI;҆I;d�I;E�I;��I;Z'I;|�F;��?;�51;;��: �,�T!�Z�Ի�|U�_l���-$����hܽi1��o���ྛ�/�V���8g��Q9���,��]]�����f^���X��      ����,������U���L�Q�ș$�5�����>�}�J(�D�׾�T���L+���սl���� L���iO���ͻ`���%m8�o�:��;d�1;��?;vF;� I;��I;��I;��I;�vI;�WI;�AI;$2I;(I;"I; I;"I;(I;$2I;�AI;�WI;�vI;��I;��I;��I;� I;vF;��?;b�1;��;�o�: &m8a����ͻ�iO� L����l����ս�L+��T��D�׾J(�>�}���5���ș$�L�Q�U��������,��      �,��b��$P���{���K��x �����s�����w��$���Ҿh��� (���ѽӷ��(������K�<ɻ������8���:��;��1;!@;��F;;I;�I;G�I;ӞI;�uI;^WI;�AI;�1I;�'I;�!I;�I;�!I;�'I;�1I;�AI;`WI;�uI;ОI;D�I;�I;;I;��F;!@;��1;��;���:���8���<ɻߔK����(�ӷ����ѽ (�h�����Ҿ�$���w�s��������x ���K��{�$P��b��      ����$P�������d���;�$���㿴���#f�f�� ž��z���@�ƽ(0v�V5�0����o@�z���Oi�0bu9zK�:O];�73;R�@;+�F;dI;��I;��I;~�I;tI;�UI;r@I;1I;'I;=!I;aI;=!I;'I;1I;p@I;�UI;tI;{�I;��I;��I;dI;+�F;R�@;�73;R];|K�:0bu9Pi�z����o@�1���V5�(0v�@�ƽ����z� žf��#f�������$����;���d����$P��      U����{���d��F�ș$�;����ɿ0蒿��K�R���j��Zb�G�4���u�a����?�����.��d���غ���9�Y�:gX;�25;S�A;�!G;g7I;��I;�I;y�I;�pI;�SI;�>I;�/I;�%I;S I;bI;S I;�%I;�/I;�>I;�SI;�pI;w�I;{�I;��I;g7I;�!G;R�A;�25;jX;�Y�:���9�غ�d����.�?������u�a�4���G�Zb��j��R����K�0蒿��ɿ;��ș$��F���d��{�      L�Q���K���;�ș$��;
��޿�����w�s,���澟���)�D������I��&�G�����N�������������9:���:�n!;��7;�B;��G;ZI;\�I;��I;�I;�lI;�PI;H<I;�-I;E$I;�I;�I;�I;C$I;�-I;F<I;�PI;�lI;�I;��I;Z�I;ZI;��G;�B;��7;�n!;���:�9:�����������N�����&�G��I������)�D��������s,���w�����޿�;
�ș$���;���K�      ș$��x �$��;���޿r���˅���F��
��~����z��$���ս���B2+���ϼPp�����2�]�h�*�V��:=�;9';ƌ:;+�C;=H;�}I;Q�I;��I;�I;�gI;�LI;M9I;k+I;V"I;*I;]I;(I;V"I;k+I;M9I;�LI;�gI;�I;��I;Q�I;�}I;<H;*�C;:;9';=�;X��:l�*�2�]�����Pp���ϼB2+������ս�$���z��~���
��F�˅��r����޿;��$���x �      5��������㿌�ɿ���˅����P�e��?�׾�`��W�H����@��T�a���̡���D��ɻ� ��ҭ�X�:�;�I-;X|=;WCE;مH;7�I;�I;��I;�I;�aI;WHI;�5I;�(I; I;I;�I;I; I;�(I;�5I;WHI;�aI;�I;��I;�I;4�I;مH;TCE;T|=;�I-;�;X�: ӭ�� ��ɻ�D�̡����T�a��@����W�H��`��?�׾e����P�˅�������ɿ�㿵���      ��s�������0蒿��w��F�e��Ͱ�"����Yb�+����ѽ�%��D4�ڟ�X������G��~潺@��9�r�: ;:3;MQ@;�vF;K�H;7�I;��I;��I;�zI;�ZI;GCI;�1I;�%I;wI;�I;WI;�I;wI;�%I;�1I;HCI;�ZI;�zI;��I;��I;3�I;K�H;�vF;HQ@;:3; ;�r�:8��9~潺�G�����X��ڟ�D4��%����ѽ+���Yb�"���Ͱ�e���F���w�0蒿����s���      =�}���w�#f���K�s,��
�?�׾"�����k���'�iz꽟I���;V�=M�����iO�\G�NoE�0�����:l� ;ҿ$;ߴ8;��B;1�G;kKI;D�I;I�I;s�I;;qI;�SI;�=I;�-I;<"I;�I;MI;�I;MI;�I;<"I;�-I;�=I;�SI;8qI;q�I;I�I;A�I;iKI;.�G;��B;۴8;ҿ$;n� ;���:4��MoE�\G໦iO����=M��;V��I��iz���'���k�"���?�׾�
�s,���K�#f���w�      J(��$�f��R������~���`���Yb���'��U�J$��G�m�&����ϼ�/��8������X�غ�9�9���:G;	H.;G|=;qE;�\H;X�I;��I;��I;/�I;4gI;7LI;8I;<)I;�I;�I;�I;]I;�I;�I;�I;;)I;8I;5LI;4gI;*�I;��I;��I;V�I;�\H;pE;D|=;H.;G;���:�9�9T�غ����8���/����ϼ&��G�m�J$���U���'��Yb��`���~�����R��f���$�      C�׾��Ҿ ž�j��������z�W�H�+��iz�J$���/v�2+�ސ�����5��ɻ4�('�����:���:fo!;>P6;<lA;�F;��H;ŷI;��I;�I;�}I;�\I;�DI;92I;�$I;�I;�I;�I;�I;�I;�I;�I;�$I;<2I;�DI;�\I;~}I;�I;��I;ǷI;��H;�F;8lA;>P6;fo!;���:���:'��4��ɻ��5���ސ�2+��/v�J$��iz�+��W�H���z������j�� ž��Ҿ      �T��h�����z�Zb�)�D��$�����ѽ�I��G�m�2+�������H�K���|�p� ���ؓ�9|T�:0;��-;��<;{zD;�H;�mI;�I;��I;ĕI;�oI;�RI;�<I;5,I;�I;EI;hI;�I;�I;�I;iI;DI;�I;8,I;�<I;�RI;�oI;ÕI;��I;�I;�mI;�H;xzD;��<;��-;0;|T�:��9���y�p���H�K�������2+�G�m��I����ѽ���$�)�D�Zb���z�h���      �L+� (���G�������ս�@���%���;V�&��ݐ�����zMS�G����8D� o8Nq�:�;��$;-_7;_�A;��F;+�H;��I;��I;��I;�I;�bI;�HI;D5I;[&I;dI;vI;%I;I;?
I;I;$I;uI;cI;[&I;D5I;�HI;�bI;�I;��I;��I;��I;'�H;��F;`�A;-_7;��$;�;Tq�:@o86D���G��zMS�����ސ�&���;V��%���@����ս����G��� (�      ��ս��ѽ?�ƽ4����I�����S�a�D4�<M���ϼ��H�K�G��>G��<f���o���:.C�:�Y;�1;�l>;E; 0H;NqI;6�I;!�I;�I;7sI;�UI;%?I;�-I;� I;�I;�I;�
I;JI;kI;JI;�
I;�I;�I;� I;�-I;%?I;�UI;7sI;�I;"�I;5�I;LqI;0H;E;�l>;�1;�Y;4C�:��:��o�;f�>G��H��H�K�����ϼ<M�D4�S�a�����I��4���>�ƽ��ѽ      l��ӷ��'0v�t�a�%�G�A2+���ڟ�����/����5�����=f��׬���g:��:3�;EI-;Mg;;1OC;=SG;�I;��I;V�I;6�I;;�I;AcI;�II;�5I;�&I;I;nI;I;�I;�I;�I;�I;�I;I;nI;I;�&I;�5I;�II;AcI;:�I;8�I;U�I;��I;�I;=SG;1OC;Ng;;EI-;6�;��:��g:�׬�=f�������5��/�����ڟ���A2+�%�G�t�a�'0v�ӷ��      ��'�U5���������ϼʡ��X���iO�8���ɻy�p�8D⺰�o���g:E`�:rG;�*;�9;��A;�uF;Q�H;��I;��I;߻I;~�I;�pI;nTI;�>I;T-I;�I;�I;0I;�I;�I;�I;	I;�I;�I;�I;/I;�I;�I;T-I;�>I;lTI;�pI;~�I;ݻI;��I;��I;R�H;�uF;��A;�9;�*;pG;C`�:��g:��o�8D�z�p��ɻ8���iO�X��ʡ����ϼ������U5�(�      L�����0���>����N��Pp��D����XG�����4�����@o8��:��:oG;4�(;̶7;��@;��E;�QH;LmI;��I;/�I;ҢI;^}I;�^I;�FI;4I;%I;�I;�I;)
I;FI;I; I;��H; I;I;GI;(
I;�I;�I;%I;4I;�FI;�^I;_}I;ҢI;)�I;��I;LmI;�QH;��E;��@;Ͷ7;3�(;oG;��:��:@o8����4�����XGແ���D�Pp��N��>���0������      �iO�ݔK��o@���.��������ɻ�G��JoE�R�غ�&����9Nq�:.C�:6�;�*;˶7;�P@;�\E;&H;JI;��I;��I;B�I;��I;whI;�NI;�:I;u*I;�I;�I;I;OI;HI;g�H;��H;�H;��H;g�H;GI;NI;I;�I;�I;r*I;�:I;�NI;vhI;��I;>�I;��I;��I; JI;'H;�\E;�P@;ɶ7;�*;6�;2C�:Nq�:��9�&��T�غHoE��G���ɻ����~����.��o@���K�      ��ͻ8ɻr����d�����'�]�� �v潺���9�9���:�T�:�;�Y;KI-;�9;��@;�\E;��G;i5I;�I;}�I;�I;��I;�pI;�UI;�@I;m/I;�!I;�I;{I;�I;�I;Y�H;��H;P�H;��H;P�H;��H;Y�H;�I;�I;{I;�I;�!I;n/I;�@I;�UI;�pI;��I;�I;}�I;�I;k5I;��G;�\E;��@;�9;LI-;�Y;�;�T�:���:�9�9��x潺� �"�]�����d��r���8ɻ      \����Ji��غ����`�*��ҭ�(��9���:���:���:0;��$;�1;Kg;;��A;��E;$H;g5I;q�I;��I;��I;ϗI;�vI;�[I;�EI;�3I;m%I;�I;�I;�	I;�I;��H;��H;_�H;!�H;��H;#�H;_�H;��H;��H;�I;�	I;�I;�I;m%I;�3I;�EI;�[I;�vI;ʗI;��I;��I;r�I;g5I;$H;��E;��A;Kg;;�1;��$;0;���:���:���:8��9�ҭ�T�*�蓛��غIi���      @)m8 ��8�bu9���9��9:d��:'X�:�r�:p� ;G;jo!;��-;-_7;�l>;3OC;�uF;�QH;JI;�I;��I;�I;�I;�zI;�_I;~II;�7I;�(I;�I;I;YI; I;a I;��H;��H;;�H;�H;��H;�H;;�H;��H;��H;b I;!I;VI;I;�I;�(I;�7I;~II;�_I;�zI;�I;�I;��I;�I;JI;�QH;�uF;1OC;�l>;-_7;��-;ho!;G;p� ;�r�:!X�:j��:��9:���9�bu9��8      �o�:���:�K�:�Y�:���:K�;�;# ;ڿ$;H.;DP6;��<;`�A;E;@SG;O�H;MmI;��I;}�I;��I;�I;|I;�aI;�KI;�9I;+I;�I;�I;�I;cI;*I;.�H;	�H;��H;)�H;G�H;	�H;G�H;)�H;��H;�H;.�H;*I;_I;�I;�I;�I;+I;�9I;�KI;�aI;|I;�I;��I;}�I;��I;JmI;N�H;ASG;E;_�A;��<;BP6;H.;ܿ$;! ;�;L�;̨�:�Y�:�K�:��:      ��;��;X];fX;�n!;9';�I-;:3;�8;I|=;?lA;zD;��F;"0H;�I;��I;��I;��I;�I;ЗI;�zI;�aI;�LI;W;I;�,I;n I;_I;2I;vI;I;��H;6�H;��H;��H;B�H;��H;]�H;��H;B�H;��H;��H;7�H;��H;I;tI;3I;\I;o I;�,I;U;I;�LI;�aI;�zI;ӗI;�I;��I;��I;��I;�I;"0H;��F;zD;<lA;G|=;�8;:3;�I-;9'; o!;fX;Y];��;      ��1;��1;�73;�25;��7;Ɍ:;c|=;NQ@;��B;vE;�F;�H;(�H;QqI;��I;��I;0�I;E�I;��I;�vI;�_I;�KI;V;I;-I;'!I;VI;I;SI;�I;3�H;��H;��H;a�H;��H;��H;�H;��H;�H;��H;��H;^�H;��H;��H;0�H;�I;SI;I;VI;(!I;-I;U;I;�KI;�_I;�vI;��I;F�I;-�I;��I;��I;QqI;(�H;�H;�F;sE;��B;NQ@;b|=;ʌ:;��7;�25;�73;��1;      ��?;/@;B�@;\�A;�B;2�C;WCE;�vF;3�G;�\H;��H;�mI;��I;;�I;Y�I;�I;٢I;��I;�pI;�[I;�II;�9I;�,I;.!I;�I;�I;�I;2I;��H;��H;��H;e�H;��H;,�H;*�H;��H;l�H;��H;+�H;+�H;��H;h�H;��H;��H;��H;3I;�I;�I;�I;*!I;�,I;�9I;II;�[I;�pI;��I;֢I;߻I;X�I;9�I;��I;�mI;��H;�\H;2�G;�vF;WCE;1�C;�B;\�A;B�@;/@;      ,vF;͊F;#�F;�!G;��G;<H;܅H;G�H;nKI;X�I;ǷI;�I;��I;"�I;6�I;}�I;_}I;vhI;�UI;�EI;�7I;+I;k I;UI;�I;	I;�I;��H;*�H;�H;e�H;x�H;��H;��H;��H;U�H;&�H;U�H;��H;��H;��H;{�H;e�H;�H;)�H;��H;�I;	I;�I;SI;k I;+I;�7I;�EI;�UI;whI;^}I;|�I;8�I;"�I;��I;�I;ŷI;U�I;kKI;I�H;܅H;:H;��G;�!G;!�F;F;      � I;@I;gI;q7I;ZI;�}I;>�I;7�I;I�I;��I;��I;��I;��I;�I;>�I;�pI;�^I;�NI;�@I;�3I;�(I;�I;_I;I;�I;�I;�H;^�H;�H;s�H;a�H;��H;V�H;V�H;��H;C�H;	�H;C�H;��H;U�H;S�H;��H;c�H;q�H;�H;`�H;�H;�I;�I;I;]I;�I;�(I;�3I;�@I;�NI;�^I;�pI;>�I;�I;��I;��I;��I;��I;I�I;7�I;>�I;�}I;!ZI;q7I;fI;=I;      ��I;�I;��I;��I;^�I;T�I;�I;��I;Q�I;��I;�I;˕I;�I;=sI;DcI;nTI;�FI;�:I;n/I;q%I;�I;�I;5I;VI;/I;��H;^�H;5�H;�H;a�H;��H;�H;�H;A�H;��H;=�H;+�H;=�H;��H;A�H;�H;�H;��H;`�H;~�H;5�H;^�H;��H;2I;VI;3I;�I;�I;q%I;n/I;�:I;�FI;nTI;DcI;=sI;�I;˕I;�I;��I;Q�I;��I;�I;T�I;h�I;��I;��I;$�I;      �I;J�I;��I;��I;��I;��I;��I;��I;x�I;0�I;�}I;�oI;�bI;�UI;�II;�>I;4I;t*I;�!I;�I;I;�I;uI;�I;��H;,�H;�H;}�H;j�H;��H;
�H;��H;��H;8�H;��H;s�H;i�H;s�H;��H;8�H;��H;��H;
�H;��H;j�H;~�H;�H;*�H;��H;�I;tI;�I;I;�I;�!I;u*I;4I;�>I;�II;�UI;�bI;�oI;�}I;-�I;x�I;��I;��I;��I;��I;��I;��I;=�I;      ��I;ݞI;��I;~�I;��I;�I;�I;�zI;CqI;@gI;�\I;�RI;�HI;/?I;6I;X-I;!%I;�I;�I;�I;ZI;`I;I;5�H;��H;�H;o�H;^�H;��H;�H;��H;��H;��H;[�H;��H;��H;��H;��H;��H;[�H;��H;��H;��H;�H;��H;`�H;o�H; �H;��H;3�H;I;bI;YI;�I;�I;�I; %I;W-I;6I;/?I;�HI;�RI;�\I;>gI;CqI;�zI;�I;�I;�I;}�I;��I;ڞI;      �vI;�uI;tI;�pI;�lI;�gI;�aI; [I;�SI;?LI;�DI;�<I;L5I;�-I;�&I;�I;�I;�I;�I;�	I;'I;*I;��H;��H;��H;e�H;^�H;��H;�H;��H;��H;��H;'�H;��H;I�H;�H;��H;�H;I�H;��H;%�H;��H;��H;��H;�H;��H;^�H;b�H;��H;��H;��H;*I;$I;�	I;�I;�I;�I;�I;�&I;�-I;L5I;�<I;�DI;>LI;�SI;[I;�aI;�gI;�lI;�pI;tI;�uI;      �WI;tWI;	VI;�SI;�PI;�LI;XHI;PCI;�=I; 8I;C2I;B,I;`&I;� I;I;�I;�I;I;�I;�I;i I;2�H;9�H;��H;c�H;v�H;��H;�H;��H;��H;��H; �H;��H;�H;��H;��H;��H;��H;��H;�H;�H;#�H;��H;��H;��H;�H;��H;u�H;h�H;��H;7�H;2�H;h I;�I;�I;I;�I;�I;
I;� I;`&I;B,I;C2I; 8I;�=I;PCI;WHI;�LI;�PI;�SI;VI;nWI;      BI;�AI;}@I;�>I;S<I;Q9I;�5I;�1I;�-I;?)I;�$I; I;hI;�I;rI;5I;0
I;MI;�I;��H;��H;	�H;��H;c�H;��H;��H;V�H;�H;��H;��H;)�H;��H;��H;��H;J�H;�H;'�H;�H;J�H;��H;��H;��H;)�H;��H;��H;�H;S�H;��H;��H;c�H;��H;	�H;��H;��H;�I;NI;/
I;3I;qI;�I;hI;  I;�$I;@)I;�-I;�1I;�5I;S9I;M<I;�>I;}@I;�AI;      62I;�1I;1I;�/I;�-I;j+I;�(I;�%I;D"I;�I;�I;LI;yI;�I; I;�I;QI;GI;^�H;��H;��H;��H;��H;��H;%�H;��H;R�H;?�H;6�H;Z�H;��H;�H;��H;/�H;�H;��H;��H;��H;�H;/�H;��H;�H;��H;[�H;;�H;?�H;R�H;��H;'�H;��H;��H;��H;��H;��H;^�H;HI;PI;�I; I;�I;yI;LI;�I;�I;D"I;�%I;�(I;n+I;�-I;�/I;1I;�1I;      (I;�'I;"'I;�%I;^$I;U"I; I;I;�I;�I;�I;vI;,I;I;�I;�I;!I;e�H;��H;d�H;C�H;+�H;B�H;��H;#�H;��H;��H;��H;��H;��H;H�H;��H;H�H;�H;��H;��H;��H;��H;��H;�H;F�H;��H;I�H;��H;��H;��H;��H;��H;#�H;��H;B�H;+�H;B�H;d�H;��H;g�H; I;�I;�I;I;,I;vI;�I;�I;�I;I; I;Y"I;V$I;�%I;"'I;�'I;      "I;�!I;J!I;[ I;I;'I;I;�I;\I;�I;�I;�I;I;VI;�I;�I;* I;��H;V�H;*�H;&�H;J�H;��H;�H;��H;O�H;@�H;<�H;u�H;��H;�H;��H;�H;��H;��H;m�H;h�H;m�H;��H;��H;�H;��H;�H;��H;w�H;<�H;?�H;N�H;��H;�H;��H;J�H;%�H;*�H;V�H;��H;) I;�I;�I;TI;I;�I;�I;�I;\I;�I;I;-I;�I;[ I;J!I;�!I;      # I; I;rI;jI;I;]I;�I;^I;�I;]I;�I;I;A
I;tI;�I;I;��H;�H;��H;��H;��H;�H;]�H;��H;g�H;�H;�H;.�H;k�H;��H;��H;��H;'�H;��H;��H;i�H;M�H;i�H;��H;��H;%�H;��H;��H;��H;n�H;.�H;�H;!�H;g�H;��H;]�H;�H;��H;��H;��H;�H;��H;I;�I;tI;A
I;I;�I;`I;�I;^I;�I;aI;I;jI;rI; I;      "I;�!I;J!I;[ I;I;(I;I;�I;\I;�I;�I;�I;I;VI;�I;�I;* I;��H;V�H;*�H;(�H;J�H;��H;�H;��H;O�H;@�H;<�H;u�H;��H;�H;��H;�H;��H;��H;m�H;h�H;m�H;��H;��H;�H;��H;�H;��H;w�H;<�H;?�H;N�H;��H;�H;��H;J�H;%�H;*�H;V�H;��H;) I;�I;�I;TI;I;�I;�I;�I;\I;�I;I;+I;�I;[ I;G!I;�!I;      (I;�'I;!'I;�%I;^$I;U"I; I;I;�I;�I;�I;vI;,I;I;�I;�I;!I;e�H;��H;d�H;E�H;+�H;B�H;��H;#�H;��H;��H;��H;��H;��H;I�H;��H;H�H;�H;��H;��H;��H;��H;��H;�H;F�H;��H;H�H;��H;��H;��H;��H;��H;#�H;��H;B�H;+�H;B�H;d�H;��H;g�H; I;�I;�I;I;,I;vI;�I;�I;�I;I; I;Y"I;V$I;�%I;!'I;�'I;      72I;�1I;1I;�/I;�-I;j+I;�(I;�%I;C"I;�I;�I;LI;yI;�I; I;�I;QI;GI;^�H;��H;��H;��H;��H;��H;'�H;��H;R�H;?�H;6�H;Z�H;��H;�H;��H;/�H;�H;��H;��H;��H;�H;/�H;��H;�H;��H;[�H;9�H;?�H;R�H;��H;%�H;��H;��H;��H;��H;��H;^�H;HI;PI;�I; I;�I;yI;LI;�I;�I;F"I;�%I;�(I;n+I;�-I;�/I;1I;�1I;      BI;�AI;~@I;�>I;S<I;Q9I;�5I;�1I;�-I;?)I;�$I;  I;hI;�I;qI;3I;0
I;MI;�I;��H;��H;	�H;��H;c�H;��H;��H;V�H;�H;��H;��H;)�H;��H;��H;��H;J�H;�H;'�H;�H;H�H;��H;��H;��H;)�H;��H;��H;�H;S�H;��H;��H;b�H;��H;	�H;��H;��H;�I;MI;/
I;5I;rI;�I;gI; I;�$I;@)I;�-I;�1I;�5I;S9I;L<I;�>I;|@I;�AI;      �WI;tWI;	VI;�SI;�PI;�LI;ZHI;PCI;�=I; 8I;C2I;B,I;`&I;� I;
I;�I;�I;I;�I;�I;l I;2�H;9�H;��H;h�H;v�H;��H;�H;��H;��H;��H; �H;�H;�H;��H;��H;��H;��H;��H;�H;}�H;"�H;��H;��H;��H;�H;��H;u�H;c�H;��H;7�H;2�H;h I;�I;�I;I;�I;�I;
I;� I;`&I;B,I;C2I;#8I;�=I;PCI;[HI;�LI;�PI;�SI;	VI;oWI;      �vI;�uI;tI;�pI;�lI;�gI;�aI; [I;�SI;<LI;�DI;�<I;L5I;�-I;�&I;�I;�I;�I;�I;�	I;(I;*I;��H;��H;��H;e�H;^�H;��H;�H;��H;��H;��H;&�H;��H;I�H;�H;��H;�H;I�H;��H;%�H;��H;��H;��H;
�H;��H;^�H;b�H;��H;��H;��H;*I;$I;�	I;�I;�I;�I;�I;�&I;�-I;L5I;�<I;�DI;ALI;�SI;[I;�aI;�gI;�lI;�pI;tI;�uI;      ��I;۞I;��I;}�I;�I;�I;�I;�zI;DqI;=gI;�\I;�RI;�HI;/?I;6I;W-I;!%I;�I;�I;�I;\I;bI;I;5�H;��H;�H;p�H;`�H;��H;�H;��H;��H;��H;Z�H;��H;��H;��H;��H;��H;[�H;��H;��H;��H;�H;��H;^�H;m�H; �H;��H;6�H;I;`I;YI;�I;�I;�I; %I;Z-I;6I;/?I;�HI;�RI;�\I;>gI;FqI;�zI;�I;�I;�I;}�I;��I;ݞI;      ��I;E�I;��I;��I;��I;��I;��I;��I;x�I;/�I;�}I;�oI;�bI;�UI;�II;�>I;4I;t*I;�!I;�I;I;�I;uI;�I;��H;,�H;�H;~�H;j�H;��H;
�H;��H;��H;8�H;��H;s�H;i�H;s�H;��H;8�H;��H;��H;
�H;��H;h�H;}�H;�H;*�H;��H;�I;tI;�I;I;�I;�!I;u*I;4I;�>I;�II;�UI;�bI;�oI;�}I;0�I;y�I;¤I;��I;��I;��I;��I;��I;E�I;      ��I;�I;��I;��I;^�I;T�I;�I;��I;Q�I;��I;�I;˕I;�I;=sI;DcI;nTI;�FI;�:I;n/I;q%I;�I;�I;5I;VI;2I;��H;^�H;5�H;�H;c�H;��H;�H;�H;@�H;��H;=�H;+�H;=�H;��H;A�H;�H;�H;��H;`�H;~�H;5�H;^�H;��H;/I;VI;3I;�I;�I;q%I;n/I;�:I;�FI;oTI;DcI;=sI;�I;˕I;�I;��I;S�I;��I;�I;Q�I;k�I;��I;��I;"�I;      � I;@I;fI;k7I;ZI;�}I;=�I;7�I;I�I;��I;��I;��I;��I;�I;<�I;�pI;�^I;�NI;�@I;�3I;�(I;�I;_I;I;�I;�I;�H;`�H;�H;s�H;c�H;��H;T�H;U�H;��H;C�H;	�H;A�H;��H;U�H;T�H;��H;a�H;q�H;�H;^�H;�H;�I;�I;I;]I;�I;�(I;�3I;�@I;�NI;�^I;�pI;<�I;�I;��I;��I;��I;��I;I�I;9�I;=�I;�}I;ZI;k7I;cI;5I;      2vF;ŊF;,�F;�!G;��G;=H;܅H;J�H;kKI;V�I;ǷI;�I;��I;"�I;5�I;}�I;_}I;vhI;�UI;�EI;�7I;+I;k I;UI;�I;	I;�I;��H;*�H;�H;e�H;x�H;��H;��H;��H;U�H;&�H;U�H;��H;��H;��H;y�H;e�H;�H;)�H;��H;�I;	I;�I;RI;k I;+I;�7I;�EI;�UI;whI;^}I;}�I;6�I;"�I;��I;�I;ǷI;V�I;lKI;J�H;ޅH;<H;��G;�!G;*�F;��F;      ��?;/@;B�@;\�A;�B;2�C;WCE;�vF;2�G;�\H;��H;�mI;��I;9�I;X�I;�I;آI;��I;�pI;�[I;�II;�9I;�,I;.!I;�I;�I;�I;3I;��H;��H;��H;f�H;��H;+�H;*�H;��H;l�H;��H;*�H;+�H;��H;h�H;��H;��H;��H;2I;�I;�I;�I;+!I;�,I;�9I;~II;�[I;�pI;��I;֢I;�I;Y�I;9�I;��I;�mI;��H;�\H;2�G;�vF;WCE;2�C;�B;\�A;B�@;-@;      ��1;��1; 83;�25;��7;ό:;^|=;NQ@;��B;vE;�F;�H;+�H;QqI;��I;��I;/�I;E�I;��I;�vI;�_I;�KI;V;I;-I;(!I;VI;I;SI;�I;3�H;��H;��H;^�H;��H;��H;�H;��H;�H;��H;��H;_�H;��H;��H;0�H;�I;SI;I;VI;'!I;-I;U;I;�KI;�_I;�vI;��I;F�I;/�I;��I;��I;QqI;*�H;�H;�F;sE;��B;QQ@;^|=;ό:;��7;�25; 83;��1;      ��;��;f];fX;�n!;9';�I-;:3;�8;I|=;<lA;zD;��F;"0H;�I;��I;��I;��I;�I;їI;�zI;�aI;�LI;W;I;�,I;n I;_I;3I;vI;I;��H;7�H;��H;��H;B�H;��H;]�H;��H;B�H;��H;��H;6�H;��H;I;tI;2I;]I;o I;�,I;U;I;�LI;�aI;�zI;ӗI;�I;��I;��I;��I;�I;"0H;��F;zD;?lA;G|=;�8;:3;�I-;9';�n!;fX;\];��;      �o�:���:�K�:�Y�:���:K�;�;  ;ڿ$;H.;BP6;��<;_�A;E;@SG;O�H;LmI;��I;}�I;��I;�I;|I;�aI;�KI;�9I;+I;�I;�I;�I;cI;*I;.�H;�H;��H;)�H;I�H;	�H;G�H;)�H;��H;	�H;-�H;*I;_I;�I;�I;�I;+I;�9I;�KI;�aI;|I;�I;��I;}�I;��I;LmI;O�H;ASG;E;`�A;��<;BP6;H.;ܿ$;# ;�;K�;Ҩ�:�Y�:�K�:��:      �'m8���8 cu9���9��9:X��:'X�:�r�:p� ;G;ho!;��-;-_7;�l>;1OC;�uF;�QH;JI;�I;��I;�I;�I;�zI;�_I;~II;�7I;�(I;�I;I;YI;!I;a I;��H;��H;;�H;�H;��H;�H;;�H;��H;��H;b I; I;VI;
I;�I;�(I;�7I;~II;�_I;�zI;�I;�I;��I;�I;JI;�QH;�uF;3OC;�l>;-_7;��-;jo!;G;p� ;�r�:)X�:j��:�9:���9cu9 ��8      \����Ei��غ�`�*�`ҭ�8��9���:���:���:0;��$;�1;Kg;;��A;��E;#H;g5I;q�I;��I;��I;ϗI;�vI;�[I;�EI;�3I;m%I;�I;�I;�	I;�I;��H;��H;_�H;$�H;��H;#�H;_�H;��H;��H;�I;�	I;�I;�I;m%I;�3I;�EI;�[I;�vI;ʗI;��I;��I;r�I;g5I;&H;��E;��A;Kg;;�1;��$; 0;���:���:���:H��9`ҭ�T�*�ⓛ��غHi����      ��ͻ8ɻr����d�����'�]�� �x潺���9�9���:�T�:�;�Y;KI-;�9;��@;�\E;��G;k5I;�I;}�I;�I;��I;�pI;�UI;�@I;n/I;�!I;�I;{I;�I;�I;Y�H;��H;P�H;��H;P�H;��H;Y�H;�I;�I;{I;�I;�!I;m/I;�@I;�UI;�pI;��I;�I;}�I;�I;l5I;��G;�\E;��@;�9;LI-;�Y;�;�T�:���:�9�9 ��t潺� �"�]�����d��r���8ɻ      �iO�ݔK��o@���.��������ɻ�G��JoE�X�غ�&����9Nq�:.C�:6�;�*;˶7;�P@;�\E;&H;JI;��I;��I;B�I;��I;uhI;�NI;�:I;u*I;�I;�I;I;OI;GI;g�H;��H;�H;��H;g�H;HI;NI;I;�I;�I;r*I;�:I;�NI;whI;��I;>�I;��I;��I;JI;'H;�\E;�P@;˶7;�*;6�;.C�:Nq�:��9�&��R�غHoE��G���ɻ����~����.��o@�ߔK�      L�����0���>����N��Pp��D����XG�����4�����@o8��:��:oG;4�(;̶7;��@;��E;�QH;LmI;��I;-�I;ҢI;^}I;�^I;�FI;4I;%I;�I;�I;)
I;GI;I; I;��H; I;I;GI;(
I;�I;�I;%I;4I;�FI;�^I;_}I;ҢI;)�I;��I;LmI;�QH;��E;��@;϶7;4�(;oG;��:��:@o8����4�����XGແ���D�Pp��N��>���0������      ��'�U5���������ϼʡ��X���iO�8���ɻz�p�8D⺰�o���g:C`�:rG;�*;�9;��A;�uF;R�H;��I;��I;ݻI;~�I;�pI;lTI;�>I;T-I;�I;�I;0I;�I;�I;�I;	I;�I;�I;�I;/I;�I;�I;T-I;�>I;nTI;�pI;��I;߻I;��I;��I;Q�H;�uF;��A;�9;�*;pG;E`�:��g:��o�8D�y�p��ɻ8���iO�X��ʡ����ϼ������U5�(�      l��ӷ��'0v�t�a�%�G�A2+���ڟ�����/����5�����=f��׬���g:��:3�;EI-;Mg;;0OC;=SG;�I;��I;U�I;6�I;<�I;AcI;�II;�5I;�&I;I;nI;I;�I;�I;�I;�I;�I;I;nI;I;�&I;�5I;�II;AcI;:�I;8�I;V�I;��I;�I;=SG;0OC;Pg;;EI-;6�;��:��g:�׬�=f�������5��/�����ڟ���A2+�%�G�t�a�'0v�ӷ��      ��ս��ѽ?�ƽ4����I�����T�a�D4�<M���ϼ��H�K�H��>G��;f���o���:2C�:�Y;�1;~l>;E; 0H;NqI;5�I;!�I;�I;7sI;�UI;#?I;�-I;� I;�I;�I;�
I;JI;kI;JI;�
I;�I;�I;� I;�-I;&?I;�UI;7sI;�I;"�I;6�I;LqI;0H;E;~l>;�1;�Y;4C�:��:��o�<f�>G��G��H�K�����ϼ<M�D4�S�a�����I��4���?�ƽ��ѽ      �L+� (���G�������ս�@���%���;V�&��ސ�����zMS�G����8D⺀o8Pq�:�;��$;,_7;`�A;��F;+�H;��I;��I;��I;�I;�bI;�HI;D5I;Y&I;cI;uI;$I;I;?
I;I;%I;vI;cI;Y&I;D5I;�HI;�bI;�I;��I;��I;��I;&�H;��F;_�A;-_7;��$;�;Tq�:�o88D���G��zMS�����ݐ�&���;V��%���@����ս����G��� (�      �T��h�����z�Zb�)�D��$�����ѽ�I��G�m�2+�������H�K���y�p�������9|T�:0;��-;��<;}zD;�H;�mI;�I;��I;ÕI;�oI;�RI;�<I;5,I;�I;EI;jI;�I;�I;�I;iI;EI;�I;7,I;�<I;�RI;�oI;ĕI;��I;�I;�mI;�H;xzD;��<;��-;0;|T�: ��9���}�p���H�K�������2+�G�m��I����ѽ���$�)�D�Zb���z�h���      C�׾��Ҿ ž�j��������z�W�H�+��iz�J$���/v�2+�ސ�����5��ɻ4� '�����:���:do!;>P6;<lA;�F;��H;ŷI;��I;�I;�}I;�\I;�DI;92I;�$I;�I;�I;�I;�I;�I;�I;�I;�$I;:2I;�DI;�\I;}I;�I;��I;ǷI;��H;�F;8lA;>P6;fo!;���:���:'��4��ɻ��5���ސ�2+��/v�J$��iz�+��W�H���z������j�� ž��Ҿ      J(��$�f��R������~���`���Yb���'��U�J$��G�m�&����ϼ�/��8������X�غ�9�9���:G;H.;G|=;qE;�\H;V�I;��I;��I;-�I;3gI;5LI;8I;<)I;�I;�I;�I;]I;�I;�I;�I;;)I;8I;7LI;6gI;,�I;��I;��I;X�I;�\H;oE;D|=;	H.;G;���:�9�9T�غ����8���/����ϼ&��G�m�J$���U���'��Yb��`���~�����R��f���$�      >�}���w�#f���K�s,��
�?�׾"�����k���'�iz꽟I���;V�=M�����iO�ZG�NoE�4�����:l� ;ҿ$;޴8;��B;.�G;hKI;D�I;I�I;s�I;6qI;�SI;�=I;�-I;<"I;�I;MI;�I;MI;�I;<"I;�-I;�=I;�SI;9qI;r�I;I�I;A�I;kKI;1�G;��B;ݴ8;ҿ$;n� ;���:0��MoE�\G໦iO����=M��;V��I��iz���'���k�"���?�׾�
�s,���K�#f���w�      ��s�������0蒿��w��F�e��Ͱ�"����Yb�+����ѽ�%��D4�ڟ�X������G��~潺@��9�r�: ;:3;KQ@;�vF;K�H;6�I;��I;��I;�zI;�ZI;GCI;�1I;�%I;xI;�I;WI;�I;wI;�%I;�1I;GCI;�ZI;�zI;��I;��I;6�I;J�H;�vF;HQ@;:3; ;�r�:8��9~潺�G�����X��ڟ�D4��%����ѽ+���Yb�"���Ͱ�e���F���w�0蒿����s���      5��������㿌�ɿ���˅����P�e��?�׾�`��W�H����@��T�a���̡���D��ɻ� ��ҭ�X�:�;�I-;X|=;TCE;مH;7�I;�I;��I;�I;�aI;VHI;�5I;�(I; I;I;�I;I; I;�(I;�5I;WHI;�aI;�I;��I;�I;6�I;مH;WCE;U|=;�I-;�;X�:�ҭ�� ��ɻ�D�̡����T�a��@����W�H��`��?�׾e����P�˅�������ɿ�㿵���      ș$��x �$��;���޿r���˅���F��
��~����z��$���ս���B2+���ϼPp�����2�]�l�*�P��:=�;9';ƌ:;*�C;=H;�}I;Q�I;��I;�I;�gI;�LI;N9I;k+I;V"I;*I;]I;*I;V"I;k+I;L9I;�LI;�gI;�I;��I;Q�I;�}I;<H;+�C;:;9';=�;X��:l�*�2�]�����Pp���ϼB2+������ս�$���z��~���
��F�˅��r����޿;��$���x �      L�Q���K���;�ș$��;
��޿�����w�s,���澟���)�D������I��&�G�����N��������������9:���:�n!;��7;�B;��G;ZI;Z�I;��I;�I;�lI;�PI;H<I;�-I;E$I;�I;�I;�I;C$I;�-I;F<I;�PI;�lI;�I;��I;\�I;ZI;��G;�B;��7;�n!;���:�9:�����������N�����&�G��I������)�D��������s,���w�����޿�;
�ș$���;���K�      U����{���d��F�ș$�;����ɿ0蒿��K�R���j��Zb�G�4���u�a����?�����.��d���غx��9�Y�:gX;�25;R�A;�!G;g7I;��I;~�I;z�I;�pI;�SI;�>I;�/I;�%I;S I;bI;S I;�%I;�/I;�>I;�SI;�pI;w�I;|�I;��I;g7I;�!G;S�A;�25;jX;�Y�:���9�غ�d����.�?������u�a�4���G�Zb��j��R����K�0蒿��ɿ;��ș$��F���d��{�      ����$P�������d���;�$���㿴���#f�f�� ž��z���@�ƽ(0v�V5�0����o@�z���Pi�bu9|K�:O];�73;R�@;+�F;dI;��I;��I;~�I;tI;�UI;r@I;1I;'I;=!I;aI;=!I;'I;1I;p@I;�UI;tI;{�I;��I;��I;dI;+�F;R�@;�73;R];zK�:0bu9Pi�z����o@�1���V5�(0v�@�ƽ����z� žf��#f�������$����;���d����$P��      �,��b��$P���{���K��x �����s�����w��$���Ҿh��� (���ѽӷ��(������K�<ɻ������8���:��;��1;!@;��F;;I;�I;G�I;ӞI;�uI;^WI;�AI;�1I;�'I;�!I;�I;�!I;�'I;�1I;�AI;`WI;�uI;ОI;D�I;�I;9I;��F;!@;��1;��;���:���8���<ɻߔK����(�ӷ����ѽ (�h�����Ҿ�$���w�s��������x ���K��{�$P��b��      ᶕ�T���Ҭ��/�_���7�|�!}߿����,b��V�0l¾Lx�f.���Ž��t�*��e����?�N�����`�x9���:��;��2;b@@;�fF;M�H;��I;��I;E|I;�[I;�CI;62I;�%I;�I;�I;`I;�I;�I;�%I;52I;�CI;�[I;E|I;��I;��I;M�H;�fF;b@@;��2;��;���:��x9���N����?�e��*����t���Žf.�Lx�0l¾�V��,b����!}߿|���7�/�_�Ҭ��T���      T���G���&}��+Y��3�����$ڿ'��ƽ\����(���s��3�8����p�d�T���<<�0��R������9���:�;_%3;up@;zF;��H;,�I;%�I;�{I;[I;�CI;�1I;�%I;TI;�I;4I;�I;WI;�%I;�1I;�CI;[I;�{I;"�I;,�I;��H;zF;up@;[%3;�;���:���9R���0���<<�T��d��p�8����3��s�(�����ƽ\�'���$ڿ����3��+Y�&}�G���      Ҭ��&}�@tf��lG�آ%��p�1�ʿ\����>M����X�����d�ʤ�̷�1�d��
��I���1�Z�����(��9���:W;�U4;��@;�F;L�H;�I;�I;�yI;�YI;rBI;1I;�$I;�I;I;�I;I;�I;�$I;1I;rBI;�YI;�yI;�I;�I;L�H;�F;��@;�U4;Z;���:(��9��Z����1��I���
�1�d�̷�ʤ���d�X�������>M�\���1�ʿ�p�آ%��lG�@tf�&}�      /�_��+Y��lG� f.�|���꿳���O䂿��5���󾎰��R�N�X��U��#�Q����|����h!�}g��񳺴	:�
�:(�;r16;��A;G;I;h�I;��I;�vI;}WI;�@I;�/I;�#I;�I;;I;�I;;I;�I;�#I;�/I;�@I;}WI;�vI;��I;h�I;I;G;��A;n16;+�;�
�:�	:�}g���h!�|������#�Q�U��X��R�N���������5�O䂿�������|� f.��lG��+Y�      ��7��3�آ%�|��<����ſ���Ž\�>����Ͼ����c�3��载z���9�`�Ἑ���z��7}��ct�t�^:�+�:أ#;č8;��B;NsG;�%I;��I; �I;0rI;CTI;>I;�-I;C"I;�I;I;�I;I;I;D"I;�-I;>I;CTI;-rI;�I;��I;�%I;LsG;��B;��8;ڣ#;�+�:x�^:�ct��7}��z����`���9��z����c�3�������Ͼ>��Ž\������ſ�<��|�آ%��3�      |�����p������ſ'���Ps���1�4r���d���d�I�шŽ��}�`*�KC���^��B�c�D��E�� �:��;�);<7;;ZD;s�G;xHI;ޝI;ۏI;�lI;"PI;�:I;G+I;O I;�I;�I;^I;�I;�I;O I;G+I;�:I;"PI;�lI;׏I;ܝI;wHI;q�G;XD;77;;�);��;� �:�E�c�D��B��^�KC��`*���}�шŽI��d��d��4r����1��Ps�'����ſ��꿄p����       }߿�$ڿ0�ʿ��������Ps�RX:����)l¾�ǆ���7����:5���Q�����t���75�`������ �8ʼ:��;��.;��=;�EE;�YH;�hI;U�I;�I;UfI;OKI;W7I;u(I;I;"I;�I;�I;�I;"I;I;u(I;Y7I;LKI;RfI;�I;U�I;�hI;�YH;�EE;��=;��.;��;ʼ:� �8���_���75��t������Q�:5�������7��ǆ�)l¾���RX:��Ps��������0�ʿ�$ڿ      ���'��\���O䂿Ž\���1�����J˾띒�H�N�z��K������W�'�e�Ҽ��|��z��n��x��h�&:�P�:֨;�W4;��@;YgF;��H;=�I;P�I;f�I;I_I;FI;:3I;S%I;vI;�I;I;�I;I;�I;vI;P%I;:3I;FI;I_I;c�I;P�I;:�I;��H;VgF;�@;�W4;֨;�P�:d�&:x���n���z���|�e�ҼW�'����K���z��H�N�띒��J˾�����1�Ž\�O䂿\���'��      �,b�ƽ\��>M���5�>��4r��)l¾띒�%&W��3�;Sؽ�z��\G����|I����?���̻r�-��	��j��:��;��&;Q|9;�C;�dG;�I;l�I;��I;�vI;�WI;^@I;�.I;�!I;�I;�I;I;�I;I;�I;�I;�!I;�.I;^@I;�WI;�vI;�I;j�I;�I;�dG;�C;O|9;��&;��;f��:�	��p�-���̻��?�|I�����\G��z��;Sؽ�3�%&W�띒�)l¾4r��>����5��>M�ƽ\�      �V������������Ͼ�d���ǆ�H�N��3��c�[����\�4��*C���o���	��눻𳺰��9h��:�h;z�/;k�=;oE;+3H;�WI;�I;+�I;�kI;�OI;V:I;*I;RI;�I;%I;�I;�I;�I;%I;�I;QI;*I;V:I;�OI;�kI;+�I;�I;�WI;(3H;lE;h�=;z�/;�h;d��:���9��눻��	��o�*C��3����\�[���cཱི3�H�N��ǆ��d����Ͼ���������      0l¾(��X������������d���7�z��;Sؽ[���d�D*�dkּ+\����'� ���R�H}����:�Z;��#;g=7;_�A;B�F;��H;��I;�I;�I;aI;�GI;&4I;X%I;�I;�I;�I;�
I;�	I;
I;�I;�I;�I;Z%I;&4I;�GI;aI;�I;�I;��I;��H;?�F;Z�A;g=7;��#;�Z;��:0}���R�!����'�+\��dkּD*��d�[��;Sؽz����7��d���������X���(��      Kx��s���d�R�N�b�3�~I����K����z����\�D*��ݼG���,<<���ڻ�V��ct���&:���:oC;�</;~D=;�D;��G;(9I; �I;הI;EtI;bVI;�?I;�-I;� I;�I;�I;�
I;-I;II;-I;�
I;�I;�I;� I;�-I;�?I;_VI;EtI;ԔI; �I;%9I;��G;�D;~D=;�</;nC;���:��&:�ct��V���ڻ,<<�G����ݼD*���\��z��K������~I�c�3�R�N���d��s�      e.��3�ʤ�X����ЈŽ:5�����[G�3��dkּG����xC��>�K6}�ج��@�x9���:4	;b�&;�;8;��A;ԟF;�H;kyI;ƝI;'�I;dfI;�KI;�7I;�'I;�I;�I;�I;HI;�I;�I;�I;HI;�I;�I;�I;�'I;�7I;�KI;dfI;#�I;ȝI;hyI;޹H;ΟF;��A;�;8;`�&;4	;���: �x9Ԭ��K6}��>��xC�G���dkּ3��[G����:5��ЈŽ��X��ʤ��3�      ��Ž7���̷�T���z����}��Q�W�'����*C��+\��,<<��>�xn���� ����:y��:;�;�'3;��>;�E;�H;�<I;�I;ٕI;�vI;YI;�AI;�/I;�!I;I;%I;�	I;�I;WI;�I;WI;�I;�	I;%I;I;�!I;�/I;�AI;YI;�vI;ڕI;�I;�<I;�H;�E;��>;�'3;9�;}��:���: � ��xn���>�,<<�+\��*C�����W�'��Q���}��z��T��̷�7���      ��t��p�0�d�"�Q�~�9�`*����e�Ҽ|I���o���'���ڻK6}��຀7���:�m�:��;�.;J<;�oC;q7G;��H;�I;�I;�I;TfI;vLI;.8I;(I;I;�I;�I;I;�I; I;� I; I;�I;�I;�I;�I;I;(I;,8I;vLI;RfI;�I;�I;�I;��H;q7G;�oC;J<;�.;��;�m�:��:�7���M6}���ڻ��'��o�|I��e�Ҽ���`*�~�9�#�Q�0�d��p�      *��c��
����_��JC���t����|���?���	����V�Ԭ�� ��:�:�h;J�+;"�9;��A;�fF;��H;�_I;��I;ΑI;;sI;�VI;�@I;/I;$!I;�I;AI;I;�I;� I;��H;=�H;��H;� I;�I;I;CI;�I;#!I;/I;�@I;�VI;;sI;͑I;��I;�_I;��H;�fF;��A;"�9;K�+;�h;�:�: �Ԭ���V�����	���?���|��t��JC��_������
�d�      d��R���I��z�������^��75��z���̻�눻�R��ct�@�x9���:�m�:�h;��*;�8;�@;�E;l(H;�8I;��I;L�I;�~I;�`I;�HI;�5I;�&I;�I;oI;2
I;�I;� I;(�H;��H;�H;��H;'�H;� I;�I;3
I;mI;�I;�&I;�5I;�HI;�`I;�~I;E�I;�I;�8I;k(H;�E;�@;�8;��*;�h;�m�:���: �x9�ct��R��눻��̻�z��75��^����{����I��S��      ��?��<<���1��h!��z��B�^���n��m�-�� }����&:���:y��:��;G�+;�8;i�@;^E;��G;yI;�I;��I;j�I;�iI;rPI;><I;�+I;�I;�I;�I;cI;�I;�H;��H;��H;�H;��H;��H;�H;�I;dI;�I;�I;�I;�+I;;<I;sPI;�iI;e�I;��I;�I;wI;��G;^E;i�@;�8;G�+;��;}��:���:��&:(}���l�-��n��^���B黵z��h!���1��<<�      N��,��T���zg���7}�Z�D�y��x��P	�����9��:���:4	;>�;�.;"�9;�@;^E;��G;sI;�I;;�I;��I;�pI;�VI;�AI;�0I;�"I;�I;%I;'I;�I;��H;��H;��H;��H;�H;��H;��H;��H;��H;�I;'I;"I;�I;�"I;�0I;�AI;�VI;�pI;�I;;�I;�I;uI;��G;!^E;�@; �9;�.;>�;4	;���:��:���9X	��x��z��U�D�~7}�zg��T���.��      ��$��������ct��E� !�8\�&:j��:n��:�Z;nC;^�&;�'3;I<;��A;�E;��G;qI;�|I;��I;אI;�uI;�[I;CFI;�4I;g&I;�I;�I;
I;,I;q�H;��H;o�H;��H;��H;X�H;��H;��H;o�H;��H;r�H;,I;
I;�I;�I;c&I;�4I;DFI;�[I;�uI;אI;��I;�|I;qI;��G;�E;��A;H<;�'3;^�&;nC;�Z;h��:j��:d�&: !�8�E��ct�����:���      0�x9���9p��9�	:d�^:� �:#ʼ:�P�:��;�h;��#;�</;�;8;��>;�oC;�fF;l(H;yI;�I;��I;�I;2xI;�^I;sII;�7I;D)I;FI;�I;�I;�I;� I;��H;��H;r�H;��H;��H;��H;��H;��H;q�H;��H;��H;� I;�I;�I;�I;CI;C)I;�7I;oII;�^I;4xI;�I;��I;�I;{I;k(H;�fF;�oC;��>;�;8;�</;��#;�h;��;�P�:#ʼ:� �:h�^:�	:x��9���9      ���:���:���:�
�:�+�:��;��;ި;��&;}�/;l=7;�D=;��A;�E;r7G;��H;�8I; �I;;�I;ِI;1xI;�_I;KI;�9I;0+I;9I;sI;tI;�I;wI;<�H;��H;V�H;w�H;�H;H�H;#�H;G�H;�H;w�H;S�H;��H;=�H;sI;�I;vI;oI;9I;3+I;�9I;KI;�_I;0xI;ڐI;;�I; �I;�8I;��H;s7G;�E;��A;�D=;k=7;}�/;��&;ި;��;��;�+�:�
�:���:���:      ��;�;^;&�;գ#;�);��.;�W4;X|9;n�=;`�A;�D;ԟF;�H;��H;�_I;��I;��I;��I;�uI;�^I;KI;_:I;Z,I;u I;�I;�I;�I;_I;��H;?�H;n�H;F�H;��H;��H;��H;��H;��H;��H;��H;D�H;n�H;?�H;��H;]I;�I;�I;�I;v I;V,I;]:I;KI;�^I;�uI;��I;��I;��I;�_I;��H;�H;ԟF;�D;_�A;l�=;W|9;�W4;��.;�);ݣ#;%�;_;�;      ʼ2;v%3;�U4;z16;ȍ8;>7;;��=;��@;�C;pE;G�F;��G;�H;�<I;�I;��I;K�I;k�I;�pI;�[I;oII;�9I;W,I;� I;WI;\I;�I;I;��H;��H;��H;c�H;y�H;	�H;'�H;��H;<�H;��H;(�H;	�H;v�H;f�H;��H;��H;��H;I;�I;ZI;YI;� I;V,I;�9I;mII;�[I;�pI;l�I;I�I;��I;�I;�<I;�H;��G;E�F;oE;�C;��@;��=;@7;;̍8;v16;�U4;h%3;      n@@;�p@;��@;��A;��B;_D;�EE;VgF;�dG;,3H;��H;)9I;iyI;
�I;�I;БI;�~I;�iI;�VI;JFI;�7I;4+I;y I;]I;�I;�I;|I;��H;�H;��H;[�H;Z�H;��H;��H;��H;Z�H;7�H;Z�H;��H;��H;��H;]�H;\�H;��H;�H;��H;{I;�I;�I;ZI;y I;4+I;�7I;KFI;�VI;�iI;�~I;ΑI;�I;�I;hyI;+9I;��H;)3H;�dG;VgF;�EE;_D;��B;��A;��@;�p@;      �fF;!zF;�F;�G;OsG;q�G;ZH;��H;�I;�WI;��I;�I;ŝI;ڕI;�I;8sI;�`I;rPI;�AI;�4I;B)I;7I;�I;ZI;�I;�I;)�H;>�H;�H;��H;m�H;��H;S�H;h�H;��H;J�H;N�H;J�H;��H;h�H;P�H;��H;n�H;��H;�H;>�H;(�H;�I;�I;YI;�I;7I;=)I;�4I;�AI;rPI;�`I;6sI;�I;ڕI;ŝI;�I;��I;�WI;�I;��H;�YH;p�G;UsG;�G;�F;zF;      `�H;��H;O�H;%I;�%I;�HI;�hI;?�I;s�I;�I;�I;ݔI;'�I;�vI;UfI;�VI;�HI;><I;�0I;g&I;FI;sI;�I;�I;uI;*�H;B�H;%�H;��H;q�H;��H;1�H;!�H;F�H;��H;N�H;N�H;N�H;��H;D�H;�H;1�H;��H;q�H;��H;&�H;A�H;(�H;xI;�I;�I;sI;DI;g&I;�0I;><I;�HI;�VI;TfI;�vI;'�I;۔I;�I;�I;s�I;?�I;�hI;|HI;�%I;%I;N�H;��H;      ��I;3�I;�I;g�I;�I;�I;Z�I;X�I;��I;4�I;�I;NtI;gfI;YI;yLI;�@I;�5I;�+I;�"I;�I;�I;vI;�I;
I;��H;>�H;%�H;��H;��H;��H;#�H;��H;��H;<�H;��H;}�H;d�H;}�H;��H;<�H;��H;��H;#�H;��H;��H;��H;%�H;>�H;��H;	I;�I;vI;�I;�I;�"I;�+I;�5I;�@I;yLI;YI;gfI;NtI;�I;2�I;��I;[�I;Z�I;ߝI;�I;h�I;�I;@�I;      ��I;(�I;�I;��I; �I;ۏI;��I;j�I;�vI;�kI;!aI;fVI;�KI;�AI;08I;/I;�&I;�I;�I;�I;�I;�I;\I;��H;�H;�H;��H;��H;��H;�H;��H;��H;��H;b�H;�H;��H;��H;��H;�H;b�H;��H;��H;��H;�H;��H;��H;��H;�H;�H;��H;[I;�I;�I;�I;�I;�I;�&I;/I;08I;�AI;�KI;dVI; aI;�kI;�vI;j�I;��I;ۏI;'�I;��I;�I;�I;      S|I;�{I;�yI;�vI;ArI;�lI;\fI;R_I;�WI;�OI;�GI;�?I;�7I;�/I;(I;'!I;�I;�I;#I;
I;�I;tI;��H;��H;��H;��H;n�H;��H;�H;��H;��H;��H;:�H;��H;I�H;�H;�H;�H;I�H;��H;8�H;��H;��H;��H;�H;��H;m�H;��H;��H;��H;��H;vI;�I;
I;#I;�I;�I;&!I;(I;�/I;�7I;�?I;�GI;�OI;�WI;S_I;[fI;�lI;>rI;�vI;�yI;�{I;      \I;�[I;�YI;�WI;STI;&PI;YKI;FI;i@I;`:I;04I;�-I;�'I;�!I;I;�I;vI;�I;,I;0I;� I;<�H;?�H;��H;U�H;o�H;��H;&�H;��H;��H;��H;�H;��H;�H;��H;��H;��H;��H;��H;�H;��H;
�H;��H;��H;��H;&�H;��H;m�H;X�H;��H;<�H;<�H;� I;0I;,I;�I;tI;�I;I;�!I;�'I;�-I;.4I;`:I;i@I;FI;WKI;%PI;PTI;�WI;�YI;�[I;      �CI;�CI;~BI;�@I;>I;;I;]7I;B3I;�.I;!*I;a%I;� I;�I;!I;�I;JI;<
I;dI;�I;x�H;��H;��H;o�H;h�H;Y�H;��H;0�H;��H;��H;��H;�H;��H;��H;��H;Q�H;�H;�H;�H;Q�H;��H;��H;��H;�H;��H;��H;��H;0�H;��H;\�H;h�H;n�H;��H;��H;x�H;�I;fI;:
I;JI;�I;!I;�I;� I;a%I;!*I;�.I;B3I;\7I;;I;>I;�@I;|BI;�CI;      ?2I;�1I;1I;�/I;�-I;I+I;w(I;X%I;�!I;VI;�I;�I;I;,I;�I;I;�I;�I;��H;�H;��H;U�H;F�H;|�H;��H;Q�H;"�H;�H;��H;>�H;��H;��H;p�H;)�H;��H;��H;��H;��H;��H;)�H;m�H;��H;��H;?�H;��H;�H;�H;O�H;��H;|�H;D�H;U�H;��H;�H;��H;�I;�I;I;�I;,I;I;�I;�I;XI;�!I;X%I;w(I;K+I;�-I;�/I;1I;�1I;      �%I;�%I;�$I;�#I;Q"I;L I;I;�I;�I;�I;�I;�I;�I;�	I;�I;�I;� I;�H;��H;t�H;y�H;x�H;��H;�H;��H;g�H;C�H;<�H;a�H;��H;�H;��H;$�H;��H;��H;{�H;_�H;{�H;��H;��H;"�H;��H;�H;��H;d�H;<�H;C�H;d�H;��H;�H;��H;w�H;x�H;t�H;��H;�H;� I;�I;�I;�	I;�I;�I;�I;�I;�I;�I;I;O I;G"I;�#I;�$I;�%I;      �I;mI;�I;�I;�I;�I;)I;�I;�I;,I;�I;�
I;OI;�I;�I;� I;2�H;��H;��H;��H;��H;�H;��H;+�H;��H;��H;��H;��H;�H;I�H;��H;T�H;��H;��H;P�H;D�H;M�H;D�H;P�H;��H;��H;V�H;��H;K�H;�H;��H;��H;��H;��H;*�H;��H;�H;��H;��H;��H;��H;0�H;� I;�I;�I;OI;�
I;�I;-I;�I;�I;)I;�I;�I;�I;�I;eI;      �I;�I;I;BI;+I;�I;�I;!I;I;�I;�
I;8I;�I;dI;I;��H;��H;��H;��H;��H;��H;I�H;��H;��H;U�H;F�H;M�H;~�H;��H;�H;��H;!�H;��H;�H;D�H;-�H;(�H;.�H;D�H;}�H;��H;$�H;��H;�H;��H;~�H;L�H;D�H;V�H;��H;��H;I�H;��H;��H;��H;��H;��H;��H;I;cI;�I;:I;�
I;�I;I; I;�I;�I; I;AI;I;�I;      cI;BI;�I;�I;�I;^I;�I;�I;�I;�I;�	I;SI;�I;�I;� I;F�H;"�H;�H;�H;\�H;��H;%�H;��H;?�H;3�H;H�H;L�H;h�H;��H;�H;��H;�H;��H;e�H;M�H;*�H;�H;*�H;M�H;e�H;��H;�H;��H;	�H;��H;h�H;J�H;J�H;3�H;<�H;��H;%�H;��H;\�H;�H;�H; �H;F�H;� I;�I;�I;SI;�	I;�I;�I;�I;�I;cI;�I;�I;�I;:I;      �I;�I;I;AI;+I;�I;�I;!I;I;�I;�
I;:I;�I;cI;I;��H;��H;��H;��H;��H;��H;I�H;��H;��H;V�H;F�H;M�H;~�H;��H;�H;��H;!�H;��H;�H;D�H;-�H;(�H;.�H;D�H;}�H;��H;$�H;��H;�H;��H;~�H;L�H;D�H;U�H;��H;��H;I�H;��H;��H;��H;��H;��H;��H;I;cI;�I;:I;�
I;�I;I; I;�I;�I; I;BI;I;�I;      �I;mI;�I;�I;�I;�I;)I;�I;�I;,I;�I;�
I;PI;�I;�I;� I;0�H;��H;��H;��H;��H;�H;��H;+�H;��H;��H;��H;��H;�H;I�H;��H;T�H;��H;��H;P�H;D�H;M�H;D�H;P�H;��H;��H;X�H;��H;K�H;�H;��H;��H;��H;��H;(�H;��H;�H;��H;��H;��H;��H;0�H;� I;�I;�I;PI;�
I;�I;-I;�I;�I;)I;�I;�I;�I;�I;eI;      �%I;�%I;�$I;�#I;O"I;L I;I;�I;�I;�I;�I;�I;�I;�	I;�I;�I;� I;�H;��H;t�H;{�H;w�H;��H;�H;��H;e�H;C�H;<�H;a�H;��H;�H;��H;$�H;��H;��H;{�H;_�H;{�H;��H;��H;"�H;��H;�H;��H;d�H;<�H;C�H;g�H;��H;�H;��H;x�H;x�H;t�H;��H;�H;� I;�I;�I;�	I;�I;�I;�I;�I;�I;�I;I;P I;D"I;�#I;�$I;�%I;      A2I;�1I;1I;�/I;�-I;I+I;w(I;W%I;�!I;VI;�I;�I;I;*I;�I;I;�I;�I;��H; �H;��H;U�H;F�H;|�H;��H;P�H;"�H;�H;��H;>�H;��H;��H;n�H;(�H;��H;��H;��H;��H;��H;(�H;m�H;��H;��H;?�H;��H;�H;�H;P�H;��H;{�H;D�H;U�H;��H;�H;��H;�I;�I;I;�I;,I;I;�I;�I;XI;�!I;W%I;w(I;K+I;�-I;�/I;1I;�1I;      �CI;�CI;|BI;�@I;>I;;I;`7I;D3I;�.I;!*I;a%I;� I;�I;!I;�I;JI;<
I;dI;�I;y�H;��H;��H;o�H;h�H;\�H;��H;0�H;��H;��H;��H;�H;��H;��H;��H;Q�H;�H;�H;�H;Q�H;��H;��H;��H;�H;��H;��H;��H;0�H;��H;Y�H;h�H;n�H;��H;��H;x�H;�I;fI;:
I;JI;�I;!I;�I;� I;a%I;"*I;�.I;D3I;`7I;;I;>I;�@I;|BI;�CI;      \I;�[I;�YI;�WI;TTI;%PI;WKI;FI;i@I;_:I;04I;�-I;�'I;�!I;I;�I;tI;�I;,I;0I;� I;<�H;?�H;��H;X�H;n�H;��H;&�H;��H;��H;��H;�H;��H;�H;��H;��H;��H;��H;��H;�H;��H;
�H;��H;��H;��H;&�H;��H;m�H;U�H;��H;<�H;<�H;� I;0I;,I;�I;tI;�I;I;�!I;�'I;�-I;.4I;b:I;i@I;FI;YKI;&PI;QTI;�WI;�YI;�[I;      M|I;�{I;�yI;�vI;<rI;�lI;[fI;P_I;�WI;�OI;�GI;�?I;�7I;�/I;(I;&!I;�I;�I;#I; 
I;�I;vI;��H;��H;��H;��H;n�H;��H;�H;��H;��H;��H;:�H;��H;I�H;�H;�H;�H;I�H;��H;:�H;��H;��H;��H;�H;��H;m�H;��H;��H;��H;��H;tI;�I;
I;#I;�I;�I;(!I;(I;�/I;�7I;�?I;�GI;�OI;�WI;V_I;]fI;�lI;>rI;�vI;�yI;�{I;      ��I;$�I;�I;��I;%�I;؏I;�I;j�I;�vI;�kI;!aI;fVI;�KI;�AI;08I;/I;�&I;�I;�I;�I;�I;�I;\I;��H;�H;�H;��H;��H;��H;�H;��H;��H;��H;b�H;�H;��H;��H;��H;�H;b�H;��H;��H;��H;�H;��H;��H;��H;�H;�H;��H;[I;�I;�I;�I;�I;�I;�&I;/I;08I;�AI;�KI;fVI;!aI;�kI;�vI;k�I;�I;ۏI;$�I;��I;�I;%�I;      ��I;6�I;�I;h�I;�I;�I;Z�I;Y�I;��I;2�I;�I;NtI;gfI;YI;yLI;�@I;�5I;�+I;�"I;�I;�I;vI;�I;	I;��H;>�H;%�H;��H;��H;��H;#�H;��H;��H;;�H;��H;}�H;d�H;}�H;��H;<�H;��H;��H;#�H;��H;��H;��H;%�H;>�H;��H;	I;�I;vI;�I;�I;�"I;�+I;�5I;�@I;yLI;YI;gfI;MtI;�I;4�I;��I;\�I;Z�I;ޝI;�I;g�I;�I;>�I;      [�H;��H;L�H;I;�%I;|HI;�hI;?�I;s�I;�I;�I;۔I;'�I;�vI;TfI;�VI;�HI;><I;�0I;i&I;II;sI;�I;�I;xI;*�H;D�H;&�H;��H;r�H;��H;1�H;�H;D�H;��H;N�H;N�H;M�H;��H;D�H;�H;1�H;��H;o�H;��H;%�H;A�H;)�H;uI;�I;�I;sI;CI;g&I;�0I;?<I;�HI;�VI;UfI;�vI;'�I;ݔI; �I;�I;s�I;@�I;�hI;{HI;�%I;I;I�H;��H;      �fF;zF;�F;�G;QsG;q�G;�YH;��H;�I;�WI;��I; �I;ŝI;ڕI;
�I;8sI;�`I;pPI;�AI;�4I;B)I;7I;�I;ZI;�I;�I;)�H;>�H;�H;��H;n�H;��H;Q�H;h�H;��H;K�H;N�H;J�H;��H;h�H;P�H;��H;m�H;��H;�H;>�H;(�H;�I;�I;WI;�I;7I;=)I;�4I;�AI;sPI;�`I;8sI;�I;ڕI;ŝI;�I;��I;�WI;�I;��H;ZH;p�G;UsG;�G;�F;zF;      n@@;�p@;��@;��A;��B;_D;�EE;VgF;�dG;+3H;��H;+9I;hyI;�I;�I;БI;�~I;�iI;�VI;KFI;�7I;4+I;y I;]I;�I;�I;|I;��H;�H;��H;\�H;\�H;��H;��H;��H;Z�H;7�H;Z�H;��H;��H;��H;]�H;[�H;��H;�H;��H;{I;�I;�I;\I;w I;4+I;�7I;KFI;�VI;�iI;�~I;БI;�I;�I;iyI;)9I;��H;+3H;�dG;WgF;�EE;aD;��B;��A;��@;�p@;      ϼ2;r%3;�U4;r16;8;D7;;��=;��@;�C;qE;F�F;��G;�H;�<I;�I;��I;K�I;j�I;�pI;�[I;pII;�9I;W,I;� I;YI;\I;�I;I;��H;��H;��H;e�H;x�H;�H;&�H;��H;<�H;��H;(�H;	�H;x�H;e�H;��H;��H;��H;I;�I;\I;WI;� I;V,I;�9I;lII;�[I;�pI;l�I;I�I;��I;�I;�<I;�H;��G;F�F;oE;�C;��@;��=;C7;;ҍ8;v16;�U4;f%3;      ��;#�;l;%�;ӣ#;�);��.;�W4;X|9;n�=;_�A;�D;ҟF;�H;��H;�_I;��I;��I;��I;�uI;�^I;KI;_:I;Z,I;v I;�I;�I;�I;_I;��H;?�H;n�H;D�H;��H;��H;��H;��H;��H;��H;��H;D�H;n�H;?�H;��H;]I;�I;�I;�I;u I;V,I;_:I;KI;�^I;�uI;��I;��I;��I;�_I;��H;�H;ҟF;�D;`�A;k�=;X|9;�W4;��.;�);٣#;%�;b;�;      ���:���:���:�
�:�+�:��;��;ި;��&;}�/;l=7;�D=;��A;�E;r7G;��H;�8I; �I;;�I;ِI;2xI;�_I;KI;�9I;3+I;9I;sI;vI;�I;wI;=�H;��H;U�H;w�H;�H;H�H;#�H;H�H;�H;w�H;U�H;��H;<�H;sI;�I;tI;oI;9I;0+I;�9I;KI;�_I;0xI;ڐI;;�I;"�I;�8I;��H;s7G;�E;��A;�D=;l=7;}�/;��&;�;��;��;�+�:�
�:���:���:      ��x9H��9���9�	:d�^:� �:'ʼ:�P�:��;�h;��#;�</;�;8;��>;�oC;�fF;l(H;yI;�I;��I;�I;4xI;�^I;sII;�7I;D)I;DI;�I;�I;�I;� I;��H;��H;o�H;��H;��H;��H;��H;��H;r�H;��H;��H;� I;�I;�I;�I;CI;D)I;�7I;mII;�^I;2xI;�I;��I;�I;{I;l(H;�fF;�oC;��>;�;8;�</;��#;�h;��;�P�:)ʼ:� �:x�^:�	:���9���9      ��(��������ct��E�@!�8d�&:l��:j��:�Z;nC;^�&;�'3;H<;��A;�E;��G;qI;�|I;��I;אI;�uI;�[I;DFI;�4I;g&I;�I;�I;
I;,I;q�H;��H;o�H;��H;��H;X�H;��H;��H;o�H;��H;r�H;,I;
I;�I;�I;c&I;�4I;CFI;�[I;�uI;אI;��I;�|I;qI;��G;�E;��A;H<;�'3;^�&;lC;�Z;j��:l��:l�&:@!�8�E๸ct�����>���      N��,��T���zg���7}�Z�D�z��x��h	�����9��:���:4	;>�;�.; �9;�@;^E;��G;sI;�I;;�I;��I;�pI;�VI;�AI;�0I;�"I;�I;%I;'I;�I;��H;��H;��H;��H;�H;��H;��H;��H;��H;�I;'I;"I;�I;�"I;�0I;�AI;�VI;�pI;�I;;�I;�I;uI;��G;!^E;�@;"�9;�.;>�;4	;���:��:���9P	��x��y��V�D�{7}�zg��S���.��      ��?��<<���1��h!��z��B�^���n��m�-��(}����&:���:y��:��;G�+;�8;h�@;^E;��G;yI;�I;��I;j�I;�iI;rPI;><I;�+I;�I;�I;�I;cI;�I;�H;��H;��H;�H;��H;��H;�H;�I;dI;�I;�I;�I;�+I;;<I;sPI;�iI;e�I;��I;�I;wI;��G;^E;k�@;�8;G�+;��;y��:���:��&: }���l�-��n��^���B黵z��h!���1��<<�      d��R���I��{�������^��75��z���̻�눻�R��ct� �x9���:�m�:�h;��*;�8;�@;�E;l(H;�8I;��I;I�I;�~I;�`I;�HI;�5I;�&I;�I;mI;3
I;�I;� I;'�H;��H;�H;��H;)�H;� I;�I;2
I;oI;�I;�&I;�5I;�HI;�`I;�~I;F�I;�I;�8I;k(H;�E;�@;	�8;��*;�h;�m�:���:@�x9�ct��R��눻��̻�z��75��^����{����I��S��      *��c��
����^��KC���t����|���?���	����V�Ԭ��@��:�:�h;J�+;"�9;��A;�fF;��H;�_I;��I;͑I;9sI;�VI;�@I;/I;#!I;�I;AI;I;�I;� I;��H;=�H;��H;� I;�I;I;AI;�I;$!I;/I;�@I;�VI;;sI;ΑI;��I;�_I;��H;�fF;��A;"�9;K�+;�h;�:�: �Ԭ���V�����	���?���|��t��JC��_������
�c�      ��t��p�0�d�"�Q�~�9�`*����e�Ҽ|I���o���'���ڻM6}��຀7���:�m�:��;�.;I<;�oC;q7G;��H;�I;�I;�I;TfI;vLI;08I;(I;I;�I;�I;�I;�I; I;� I; I;�I;�I;�I;�I;I;(I;,8I;vLI;RfI;�I;�I;�I;��H;q7G;�oC;L<;�.;��;�m�:��:�7���K6}���ڻ��'��o�|I��e�Ҽ���`*�~�9�"�Q�0�d��p�      ��Ž7���̷�T���z����}��Q�W�'����*C��+\��,<<��>�xn�� �� ����:}��:9�;�'3;��>;�E;�H;�<I;�I;וI;�vI;YI;�AI;�/I;�!I;I;%I;�	I;�I;WI;�I;WI;�I;�	I;#I;I;�!I;�/I;�AI;YI;�vI;ڕI;�I;�<I;�H;�E;��>;�'3;;�;��:���: ���xn���>�,<<�+\��*C�����W�'��Q���}��z��T��̷�7���      e.��3�ʤ�X����ЈŽ:5�����[G�3��dkּG����xC��>�K6}�ج��@�x9���:4	;`�&;�;8;��A;ҟF;�H;hyI;ƝI;'�I;dfI;�KI;�7I;�'I;�I;�I;�I;HI;�I;�I;�I;HI;�I;�I;�I;�'I;�7I;�KI;dfI;#�I;ɝI;kyI;ܹH;ϟF;��A;�;8;a�&;4	;���: �x9ج��K6}��>��xC�G���dkּ3��[G����:5��ЈŽ��X��ʤ��3�      Kx��s���d�R�N�b�3�~I����K����z����\�D*��ݼG���,<<���ڻ�V��ct���&:���:nC;�</;~D=;�D;��G;%9I;�I;הI;EtI;`VI;�?I;�-I;� I;�I;�I;�
I;.I;II;.I;�
I;�I;�I;� I;�-I;�?I;`VI;EtI;ԔI; �I;(9I;��G;�D;~D=;�</;nC;���:��&:�ct��V���ڻ,<<�G����ݼD*���\��z��K������~I�b�3�R�N���d��s�      0l¾(��X������������d���7�z��;Sؽ[���d�D*�dkּ+\����'�!���R�@}����:�Z;��#;g=7;_�A;B�F;��H;��I;�I;�I;aI;�GI;&4I;U%I;�I;�I;�I;�
I;�	I;�
I;�I;�I;�I;Z%I;&4I;�GI;aI;�I;�I;��I;��H;?�F;Z�A;g=7;��#;�Z;��:0}���R�!����'�+\��dkּD*��d�[��;Sؽz����7��d���������X���(��      �V������������Ͼ�d���ǆ�H�N��3��c�[����\�3��*C���o���	��눻𳺰��9h��:�h;z�/;k�=;oE;(3H;�WI;�I;+�I;�kI;�OI;V:I;*I;RI;�I;%I;�I;�I;�I;%I;�I;QI;*I;V:I;�OI;�kI;+�I;�I;�WI;+3H;lE;i�=;z�/;�h;d��:���9��눻��	��o�*C��4����\�[���cཱི3�H�N��ǆ��d����Ͼ���������      �,b�ƽ\��>M���5�>��4r��)l¾띒�%&W��3�;Sؽ�z��\G����|I����?���̻r�-��	��j��:��;��&;Q|9;�C;�dG;�I;l�I;�I;�vI;�WI;^@I;�.I;�!I;�I;�I;I;�I;I;�I;�I;�!I;�.I;^@I;�WI;�vI;��I;j�I;�I;�dG;�C;O|9;��&;��;f��:�	��o�-���̻��?�|I�����\G��z��;Sؽ�3�%&W�띒�)l¾4r��>����5��>M�ƽ\�      ���'��\���O䂿Ž\���1�����J˾띒�H�N�z��K������W�'�e�Ҽ��|��z��n��x��h�&:�P�:֨;�W4;�@;VgF;��H;<�I;P�I;f�I;I_I;FI;:3I;Q%I;xI;�I;I;�I;I;�I;xI;Q%I;:3I;FI;I_I;c�I;P�I;:�I;��H;YgF;�@;�W4;֨;�P�:d�&:x���n���z���|�e�ҼW�'����K���z��H�N�띒��J˾�����1�Ž\�O䂿\���'��       }߿�$ڿ0�ʿ��������Ps�RX:����)l¾�ǆ���7����:5���Q�����t���75�`����� !�8ʼ:��;��.;��=;�EE;�YH;�hI;U�I;�I;RfI;LKI;W7I;v(I;I;"I;�I;�I;�I;"I;I;s(I;W7I;OKI;TfI;�I;U�I;�hI;�YH;�EE;��=;��.;��;ʼ:� �8���_���75��t������Q�:5�������7��ǆ�)l¾���RX:��Ps��������0�ʿ�$ڿ      |�����p������ſ'���Ps���1�4r���d���d�I�шŽ��}�`*�KC���^��B�c�D��E�� �:��;�);<7;;XD;s�G;xHI;ܝI;ۏI;�lI;"PI;�:I;H+I;O I;�I;�I;^I;�I;�I;O I;E+I;�:I;"PI;�lI;׏I;ޝI;wHI;q�G;ZD;77;;�);��;� �:�E�c�D��B��^�KC��`*���}�шŽI��d��d��4r����1��Ps�'����ſ��꿄p����      ��7��3�آ%�|��<����ſ���Ž\�>����Ͼ����c�3��载z���9�`�Ἑ���z��7}��ct�p�^:�+�:أ#;č8;��B;NsG;�%I;��I;!�I;0rI;CTI;>I;�-I;D"I;�I;I;�I;I;I;C"I;�-I;>I;CTI;.rI;�I;��I;�%I;LsG;��B;��8;ڣ#;�+�:x�^:�ct��7}��z����`���9��z����c�3�������Ͼ>��Ž\������ſ�<��|�آ%��3�      /�_��+Y��lG� f.�|���꿳���O䂿��5���󾎰��R�N�X��U��#�Q����|����h!�}g��񳺰	:�
�:(�;r16;��A;G;I;h�I;��I;�vI;}WI;�@I;�/I;�#I;�I;;I;�I;;I;�I;�#I;�/I;�@I;}WI;�vI;��I;h�I;I;G;��A;n16;+�;�
�:�	:�}g���h!�|������#�Q�U��X��R�N���������5�O䂿�������|� f.��lG��+Y�      Ҭ��&}�@tf��lG�آ%��p�1�ʿ\����>M����X�����d�ʤ�̷�1�d��
��I���1�Z����� ��9���:W;�U4;��@;�F;L�H;�I;�I;�yI;�YI;rBI;1I;�$I;�I;I;�I;I;�I;�$I;1I;rBI;�YI;�yI;�I;�I;L�H;�F;��@;�U4;Z;���:(��9��Z����1��I���
�1�d�̷�ʤ���d�X�������>M�\���1�ʿ�p�آ%��lG�@tf�&}�      T���G���&}��+Y��3�����$ڿ'��ƽ\����(���s��3�8����p�d�T���<<�0��N������9���:�;a%3;up@;zF;��H;,�I;%�I;�{I;[I;�CI;�1I;�%I;TI;�I;4I;�I;WI;�%I;�1I;�CI;[I;�{I;"�I;,�I;��H;zF;up@;]%3;�;���:���9R���0���<<�T��d��p�8����3��s�(�����ƽ\�'���$ڿ����3��+Y�&}�G���      �Aq���i���U�I:�@�����=���x���}A�f5�� ���^Z�����A���]�����d��H",��5��V�Ѻ���9��:b�;fY4;v�@;�VF;��H;�GI;�bI;>OI;N:I;*I;QI;�I;�I;�I;�I;�I;�I;�I;OI;*I;N:I;=OI;�bI;�GI;��H;�VF;v�@;bY4;e�;��:���9Z�Ѻ�5��H",��d������]��A������^Z�� ��f5�}A�x���=�������@�I:���U���i�      ��i���b�\�O�.5�4i�������������q<����f��c
V�IE	�!���IY�k9�D�����(��R����Ⱥ��:���:$�;L�4;p�@;qhF;ƗH;@II;�bI;�NI;�9I;�)I;I;�I;�I;�I;�I;�I;�I;�I;I;�)I;�9I;�NI;�bI;@II;ƗH;qhF;p�@;H�4;*�;���:��:��Ⱥ�R����(�D���k9��IY�!��IE	�c
V�f������q<������������4i�.5�\�O���b�      ��U�\�O�J-?�0�'���O�ῶ欿c�{�ha/���뾟���I����f���ZN�`5������9H�Z �������":��:��;��5;�`A;�F;b�H;FMI;(bI;�MI;�8I;)I;sI;I;rI;8I;9I;8I;qI;I;qI;)I;�8I;�MI;%bI;FMI;b�H;�F;�`A;��5;��;��:��":���Z ��9H�����`5���ZN�f������I�������ha/�c�{��欿O����0�'�J-?�\�O�      I:�.5�0�'� ������lȿ���m$_���Z�Ҿޕ���6�����*���`=�>�漮)��FG�6��X��h�Q:�:0";�7;�&B;�F;��H;SI;�`I;�KI;P7I;�'I;nI;LI;�I;�I;�
I;�I;�I;LI;lI;�'I;P7I;�KI;�`I;SI;��H;�F;�&B;�7;0";�:t�Q:Z��6��EG��)��>���`=��*������6�ޕ��Z�Ҿ��m$_����lȿ���� ��0�'�.5�      @�4i�������K�ѿm������q<��:��a����q����Wн齅���'�Vb̼�zl��.��5�X�����:��;
�&;߫9;VC;�MG;�H;hYI;�^I;�HI;5I;&I;I;;I;�I;�
I;�	I;�
I;�I;;I;I;&I;5I;�HI;�^I;hYI;	�H;~MG;TC;ܫ9;�&;��;�:���5�X��.���zl�Vb̼��'�齅��Wн����q��a���:��q<���m���K�ѿ������4i�      �������O��lȿm���������O���}]׾}����I�����A��A�d�o�~֮�	RH��jλ5�$��%����:hN;̆+; <;,4D;�G;�I;�^I;�[I;EI;U2I;�#I;sI;�I;�I;�	I;�I;�	I;�I;�I;sI;�#I;U2I;EI;�[I;�^I;�I;�G;*4D;�<;̆+;hN;���:�%�5�$��jλ	RH�~֮�o�A�d��A������I�}���}]׾����O�����m���lȿO�Ῥ��      =��������欿�������O��x����� ���l���"��ܽ���`=����v���k"�#R��ۺ(��9�?�:�L;��0;ӟ>;�ME;�#H;�%I;bI;7WI;�@I;&/I;s!I;nI;7I;@I;~I;�I;~I;@I;5I;nI;t!I;&/I;�@I;5WI;bI;�%I;�#H;�ME;Ο>;��0;�L;�?�:��9ۺ"R���k"�v������`=����ܽ��"��l�� ����뾃x���O�������欿����      w�������c�{�m$_��q<������~��
w���6�����!���h����䷾�� d�t.��~^e��H[���Z:���:�, ;��5;�A;WF;لH;AI;�bI;�QI;<I;t+I;�I;?I;kI;�	I;I;bI;I;�	I;kI;=I;�I;r+I;<I;�QI;�bI;AI;ׄH; WF;�A;��5;�, ;���:��Z:�H[�}^e�t.��� d�䷾�����h�!�������6�
w��~��������q<�m$_�c�{�����      }A��q<�ha/����:�}]׾� ��
w��>�FE	�����ܽ����3�`�꼘���
",��W��D���Q�װ�:�M
;�f);�:;N@C;%@G;��H;tTI;�_I;\KI;7I;�'I;�I;�I;rI;I;�I;�I;�I;I;rI;�I;�I;�'I;7I;YKI;�_I;pTI;��H;"@G;K@C;�:;�f);�M
;Ӱ�:�Q�B���W��
",�����`�꼛�3�ܽ������FE	�>�
w��� ��}]׾�:���ha/��q<�      f5�������Z�Ҿ�a��}����l��6�FE	���Ƚk���aG����e֮��W����O�k����<d,:���:!�;��1;t�>;gE;X�G;SI;U_I;vZI;lDI;�1I;g#I;wI;-I;9
I;@I;I;UI;I;@I;9
I;,I;yI;e#I;�1I;iDI;vZI;T_I;SI;W�G;dE;s�>;��1;!�;���:<d,:���Q�k�����W�e֮�����aG�k����ȽFE	��6��l�}����a��Z�Ҿ������      � ��f�����ݕ����q��I���"���������k���ZN�\�"¼M�y��$��Q��k� � �W��:K0;P�&;x8;� B;��F;�H;�@I;&bI;�RI;P=I;F,I;I;I;�I;I;nI;QI;�I;QI;nI;I;�I;I;I;F,I;M=I;�RI;$bI;�@I;	�H;��F;� B;x8;O�&;J0;�: �W�m� ��Q���$�M�y�"¼\��ZN�k������������"��I���q�ݕ�����f��      �^Z�c
V��I��6�������ܽ!��ܽ���aG�\��ȼ�)��z�(�\��2G5�(���Z:f�:>S;6'1;�=;ܠD;]�G;#�H;�XI;M^I;�II;,6I;�&I;�I;�I;�
I;�I;�I;� I;��H;� I;�I;�I;�
I;�I;�I;�&I;+6I;�II;J^I;�XI; �H;Z�G;ؠD;�=;6'1;<S;f�:$�Z:0��2G5�]��z�(��)���ȼ\��aG�ܽ��!���ܽ������6��I�c
V�      ���IE	��������Wн�A�����h���3����"¼�)��-x/��һV�X�6#����9���:�>;df);�`9;�&B;�F;�}H;7I;�aI;�UI;�@I;/I;1!I;I;[I;I;�I;� I;��H;2�H;��H;� I;�I;I;\I;I;1!I;/I;�@I;�UI;�aI;7I;�}H;�F;�&B;�`9;bf);�>;���:��94#��W�X��һ-x/��)��"¼�����3��h��󑽤A���Wн��콼��IE	�      �A��!��e���*��轅�@�d��`=����_��e֮�L�y�y�(��һ�]e�������f9���:[�;p1";N�4;�m?;E;��G;��H;�WI;�^I;?KI;�7I;,(I;�I;_I;�
I;ZI;UI;��H;�H;s�H;�H;��H;SI;XI;�
I;]I;�I;*(I;�7I;>KI;�^I;�WI;��H;��G;E;�m?;N�4;p1";\�;���:��f9�����]e��һy�(�L�y�e֮�^�꼚���`=�@�d�轅��*��e��!��      �]��IY��ZN��`=���'�n����䷾������W��$�]��Y�X�����@9���:���:��;Ҹ0;�<;��C;TG;1�H;�?I;baI;	UI;s@I;H/I;�!I;�I;HI;�I;�I;�H;��H;B�H;��H;B�H;��H;�H;�I;�I;HI;�I;�!I;H/I;r@I;	UI;`aI;�?I;,�H;TG;��C;�<;Ҹ0;��;���:���:@9����Y�X�^���$��W�����䷾����n���'��`=��ZN��IY�      ���j9�]5��=��Vb̼~֮�t��� d�",�����Q��0G5�8#��`�f9���:��:;�;��-;��:;LB;mVF;KKH;I;]I;Z\I;�HI;?6I;W'I;UI;�I;R
I;yI;4 I;��H;��H;��H;$�H;��H;��H;��H;3 I;zI;R
I;�I;PI;W'I;<6I;�HI;Y\I;]I;I;KKH;jVF;LB;��:;��-;8�;��:���:��f98#��2G5��Q�����",�� d�t��}֮�Vb̼=��]5��j9�      �d��B��������)���zl�RH��k"�r.���W��M�k�i� �(����9���:���:8�;�-;��9;vaA;�E;Z�G;��H;:SI;L`I; PI;�<I;�,I;�I;lI;GI;�I;�I;��H;��H;�H;��H;��H;��H;�H;��H;��H;�I;�I;GI;iI;�I;�,I;�<I; PI;G`I;4SI;��H;W�G;�E;vaA;��9;�-;5�;���:���:��9(��j� �N�k��W��r.���k"�RH��zl��)������C���      H",���(�7H�DG��.���jλ"R��~^e�A����� �W��Z:���:[�;��;��-;��9;�A;dE;W�G;��H;�GI;-aI;�UI;xBI;�1I;%$I;I;&I;�I;-I;��H;��H;�H;B�H;N�H;!�H;N�H;B�H;�H;��H;��H;-I;�I;#I;I; $I;�1I;zBI;�UI;+aI;�GI;��H;W�G;dE;�A;��9;��-;��;[�;���:�Z: �W����?���^e�"R���jλ�.��DG�7H���(�      �5���R��S ��6��8�X�.�$��ۺ|H[��Q�@d,:�:l�:�>;s1";ո0;��:;waA;dE;)�G;��H;�=I;c`I;�YI;'GI;6I;�'I;'I;�I;4I;�I; I;>�H;[�H;2�H;��H;��H;y�H;��H;��H;/�H;Z�H;?�H; I;�I;2I;�I;%I;�'I;6I;#GI;�YI;d`I;�=I;��H;)�G;dE;taA;��:;ָ0;s1";�>;l�:�:@d,: Q��H[��ۺ*�$�3�X�6��S ���R��      N�Ѻ��Ⱥ���V������%���9��Z:װ�:���:M0;<S;af);H�4;�<;LB;�E;T�G;��H;�:I;�_I;�[I;ZJI;=9I;�*I;�I;/I;9I;�I;JI;$�H;��H;L�H;i�H;4�H;k�H;"�H;m�H;4�H;i�H;K�H;��H;&�H;GI;�I;9I;-I;�I;�*I;99I;YJI;�[I;�_I;�:I;��H;V�G;�E;LB;�<;J�4;af);<S;K0;���:Ӱ�:��Z:��9�%�|��V�� �����Ⱥ      ���9Ժ:Ы":T�Q:�:���:�?�:���:�M
;#�;R�&;6'1;�`9;�m?;��C;lVF;[�G;��H;�=I;�_I;I\I;�KI;O;I;	-I;	!I;,I;�I;"I;�I;�H;q�H;��H;s�H;��H;��H;�H;��H;�H;��H;��H;q�H;��H;q�H;�H;�I;"I;�I;*I;	!I;-I;N;I;�KI;F\I;�_I;�=I;��H;Z�G;lVF;��C;�m?;�`9;6'1;O�&;!�;�M
;���:�?�:���:�:\�Q:ث":��:      "��:���:��:��:��;tN;�L;�, ;�f);1;x8;�=;�&B;E;WG;JKH;��H;�GI;c`I;�[I;�KI;�;I;%.I;j"I;oI;PI;W	I;�I;��H;)�H;�H;��H;��H;X�H;{�H;��H;��H;��H;{�H;X�H;��H;��H;�H;%�H;��H;�I;S	I;QI;rI;f"I;$.I;�;I;�KI;�[I;c`I;�GI;��H;HKH;XG;E;�&B;�=;x8;Ó1;�f);�, ;�L;tN;��;��:��:���:      h�;*�;��;0";�&;Ά+;��0;��5;�:;w�>;� B;ݠD;�F;��G;0�H;I;7SI;,aI;�YI;\JI;N;I;(.I;�"I;;I;�I;9
I;iI;��H;��H;��H;��H;��H;6�H;�H;.�H;��H;��H;��H;.�H;�H;5�H;��H;��H;��H;��H;��H;gI;:
I;�I;8I;�"I;(.I;K;I;]JI;�YI;-aI;6SI;I;0�H;��G;�F;ݠD;� B;v�>;�:;��5;��0;φ+;�&;0";��; �;      ~Y4;b�4;��5; �7;�9; <;۟>;�A;R@C;hE;��F;`�G;�}H;��H;�?I;]I;L`I;�UI;'GI;;9I;-I;i"I;8I;^I;�
I;�I;) I;%�H;��H;$�H;��H;2�H;��H;��H; �H;��H;��H;��H;�H;��H;��H;5�H;��H;"�H;��H;%�H;' I;�I;�
I;[I;8I;i"I;-I;;9I;'GI;�UI;K`I;]I;�?I;��H;�}H;`�G;��F;gE;P@C;�A;۟>;<;�9;�7;��5;T�4;      ��@;|�@;�`A;�&B;ZC;04D;�ME;WF;)@G;X�G;�H;'�H;7I;�WI;eaI;]\I;(PI;{BI; 6I;�*I;!I;sI;�I;�
I;*I;Z I;o�H;!�H;_�H;�H;?�H;��H;��H;��H;�H;��H;��H;��H;�H;��H;��H;��H;?�H;�H;\�H;!�H;l�H;Z I;+I;�
I;�I;sI;!I;�*I; 6I;~BI;%PI;Z\I;eaI;�WI;7I;'�H;�H;V�G;'@G;WF;�ME;04D;\C;�&B;�`A;|�@;      �VF;�hF;֛F;�F;�MG;�G;�#H;ԄH;��H;UI;�@I;�XI;�aI;�^I;	UI;�HI;�<I;�1I;�'I;�I;)I;OI;6
I;�I;S I;��H;S�H;��H;,�H;9�H;��H;��H;|�H;��H;B�H;��H;��H;��H;D�H;��H;z�H;��H;��H;7�H;*�H;��H;Q�H;��H;T I;�I;6
I;PI;&I;�I;�'I;�1I;�<I;�HI;	UI;�^I;�aI;�XI;�@I;QI;��H;ԄH;�#H;�G;�MG;�F;֛F;vhF;      ��H;ɗH;e�H;��H;�H;�I;&I;AI;zTI;[_I;*bI;Q^I;�UI;BKI;v@I;?6I;�,I;"$I;'I;1I;�I;W	I;hI;, I;h�H;U�H;��H;M�H;g�H;��H;h�H;J�H;w�H;��H;v�H; �H;
�H;"�H;u�H;��H;t�H;K�H;h�H;��H;g�H;O�H;��H;T�H;k�H;) I;gI;W	I;�I;1I;'I;#$I;�,I;=6I;v@I;BKI;�UI;Q^I;*bI;X_I;zTI;AI;&I;�I;�H;��H;d�H;ʗH;      �GI;CII;PMI;SI;kYI;�^I;
bI;�bI;`I;~ZI;�RI;�II;�@I;�7I;I/I;W'I;�I; I;�I;=I;"I;�I;��H;'�H;�H;��H;M�H;C�H;��H;h�H;?�H;F�H;��H;�H;��H;|�H;r�H;|�H;��H;�H;��H;G�H;A�H;e�H;��H;C�H;M�H;��H;�H;'�H;��H;�I;I;<I;�I; I;�I;W'I;I/I;�7I;�@I;�II;�RI;~ZI;`I;�bI;
bI;�^I;vYI;SI;PMI;OII;      cI;�bI;$bI;�`I;�^I;�[I;=WI;�QI;bKI;rDI;S=I;26I;/I;,(I;�!I;SI;mI;#I;4I;�I;�I;��H;��H;��H;X�H;,�H;d�H;��H;Z�H;=�H;4�H;v�H;��H;g�H;
�H;��H;��H;��H;
�H;g�H;��H;w�H;4�H;<�H;Z�H;��H;f�H;*�H;[�H;��H;��H;��H;�I;�I;6I;%I;lI;RI;�!I;-(I;/I;06I;Q=I;oDI;bKI;�QI;<WI;�[I;�^I;�`I;%bI;�bI;      KOI;�NI;�MI;�KI;�HI;EI;�@I;&<I;7I;�1I;Q,I;�&I;8!I;�I;�I;�I;MI;�I;�I;MI;�H;&�H;��H;%�H;�H;5�H;��H;d�H;<�H;<�H;e�H;��H;3�H;��H;�H;_�H;[�H;_�H;�H;��H;0�H;��H;e�H;;�H;:�H;g�H;��H;3�H;�H;$�H;��H;&�H;�H;LI;�I;�I;JI;�I;�I;�I;8!I;�&I;P,I;�1I;7I;*<I;�@I;EI;�HI;�KI;�MI;�NI;      U:I;�9I;�8I;`7I;&5I;X2I;3/I;|+I;�'I;o#I;I;�I;�I;gI;NI;[
I;�I;/I; I;*�H;w�H;�H;��H;��H;9�H;��H;d�H;A�H;2�H;h�H;��H;,�H;��H;M�H;�H;��H;��H;��H;�H;N�H;��H;-�H;��H;g�H;4�H;A�H;d�H;��H;:�H;��H;��H;�H;t�H;(�H; I;-I;�I;X
I;MI;fI;�I;�I;I;o#I;�'I;|+I;3/I;X2I;$5I;`7I;�8I;�9I;      *I;�)I;)I;�'I;&I;�#I;x!I;�I;�I;}I;$I;�I;bI;�
I;�I;�I;�I;��H;E�H;��H;��H;��H;��H;6�H;��H;��H;H�H;G�H;u�H;��H;)�H;��H;,�H;��H;��H;��H;t�H;��H;��H;��H;)�H;��H;,�H;��H;w�H;G�H;H�H;��H;��H;6�H;��H;��H;��H;��H;E�H;��H;�I;~I;�I;�
I;bI;�I;#I;|I;�I;�I;x!I;�#I;&I;�'I;)I;�)I;      XI;/I;�I;}I;#I;vI;rI;II;�I;1I;�I;�
I;I;aI;�I;: I;��H;��H;^�H;O�H;w�H;��H;6�H;��H;��H;{�H;v�H;��H;��H;6�H;��H;/�H;��H;��H;L�H;B�H;N�H;B�H;J�H;��H;��H;0�H;��H;7�H;��H;��H;t�H;z�H;��H;��H;5�H;��H;w�H;P�H;^�H;��H;��H;8 I;�I;aI;I;�
I;�I;3I;�I;II;rI;xI;I;}I;~I;(I;      �I;�I;I;XI;HI;�I;<I;xI;yI;?
I;I;�I;�I;[I;!�H;�H;��H;�H;6�H;o�H;��H;Y�H;�H;��H;��H;��H;��H;�H;e�H;��H;K�H;��H;��H;\�H;!�H;�H;��H;�H;!�H;\�H;��H;��H;K�H;��H;h�H;�H;��H;��H;��H;��H;�H;Y�H;��H;o�H;6�H;�H;��H;�H;�H;[I;�I;�I;I;=
I;|I;xI;<I;�I;>I;XI;I;�I;      �I;�I;�I;�I;�I;�I;II;�	I;I;GI;yI;�I;� I;��H;��H;��H;�H;A�H;��H;:�H;��H;~�H;-�H;�H;�H;?�H;p�H;��H;
�H;�H;�H;��H;L�H;$�H;�H;��H;��H;��H;�H;$�H;I�H;��H;�H;��H;�H;��H;p�H;?�H;�H;�H;-�H;~�H;��H;:�H;��H;D�H;�H;��H;��H;��H;� I;�I;wI;HI;I;�	I;II;�I;�I;�I;�I;�I;      �I;�I;FI;�I;�
I;�	I;�I;,I;�I;I;[I;� I;��H;�H;I�H;��H;��H;K�H;��H;t�H;�H;��H;��H;��H;��H;��H;�H;|�H;��H;_�H;��H;��H;C�H;�H;��H;��H;��H;��H;��H;	�H;B�H;��H;��H;`�H;��H;|�H;�H;��H;��H;��H;��H;��H;�H;t�H;��H;M�H;��H;��H;I�H;�H;��H;� I;YI;I;�I;*I;�I;�	I;�
I;�I;EI;�I;      �I;�I;NI;�
I;�	I;�I;�I;kI;�I;VI;�I;��H;9�H;}�H;��H;+�H;��H;�H;|�H;(�H;��H;��H;��H;��H;��H;��H;�H;x�H;��H;]�H;��H;{�H;N�H;��H;��H;��H;��H;��H;��H;��H;M�H;}�H;��H;_�H;��H;x�H;�H;��H;��H;��H;��H;��H;��H;(�H;|�H;�H;��H;+�H;��H;}�H;9�H;��H;�I;YI;�I;jI;�I;�I;�	I;�
I;LI;�I;      �I;�I;FI;�I;�
I;�	I;�I;,I;�I;I;[I;� I;��H;�H;I�H;��H;��H;K�H;��H;t�H;�H;��H;��H;��H;��H;��H;�H;|�H;��H;_�H;��H;��H;B�H;�H;��H;��H;��H;��H;��H;	�H;B�H;��H;��H;`�H;��H;|�H;�H;��H;��H;��H;��H;��H;�H;t�H;��H;M�H;��H;��H;K�H;�H;��H;� I;[I;I;�I;*I;�I;�	I;�
I;�I;BI;�I;      �I;�I;I;�I;�I;�I;II;�	I;I;GI;wI;�I;� I;��H;��H;��H;�H;B�H;��H;:�H;��H;~�H;-�H;�H;�H;?�H;p�H;��H;�H;�H;�H;��H;L�H;$�H;�H;��H;��H;��H;�H;$�H;I�H;��H;�H;��H;�H;��H;p�H;?�H;�H;�H;-�H;~�H;��H;:�H;��H;D�H;�H;��H;��H;��H;� I;�I;wI;HI;I;�	I;II;�I;�I;�I;}I;�I;      �I;�I;I;XI;GI;�I;<I;xI;zI;=
I;I;�I;�I;[I;!�H;�H;��H;�H;6�H;o�H;��H;Y�H;�H;��H;��H;��H;��H;�H;e�H;��H;K�H;��H;��H;\�H;!�H;�H;��H;�H;!�H;\�H;��H;��H;K�H;��H;h�H;�H;��H;��H;��H;��H;�H;Y�H;��H;o�H;6�H;�H;��H;�H;�H;[I;�I;�I;I;?
I;|I;zI;<I;�I;;I;XI;I;�I;      [I;/I;I;~I;"I;vI;rI;GI;�I;1I;�I;�
I;I;aI;�I;8 I;��H;��H;^�H;O�H;x�H;��H;6�H;��H;��H;{�H;w�H;��H;��H;6�H;��H;/�H;��H;��H;J�H;B�H;N�H;B�H;L�H;��H;��H;2�H;��H;7�H;��H;��H;t�H;z�H;��H;��H;5�H;��H;w�H;P�H;^�H;��H;��H;: I;�I;aI;I;�
I;�I;3I;�I;FI;rI;wI;I;~I;}I;,I;      *I;�)I;)I;�'I;&I;�#I;{!I;�I;�I;|I;$I;�I;bI;�
I;�I;�I;�I;��H;E�H;��H;��H;��H;��H;6�H;��H;��H;H�H;G�H;u�H;��H;,�H;��H;+�H;��H;��H;��H;t�H;��H;��H;��H;)�H;��H;)�H;��H;w�H;G�H;H�H;��H;��H;6�H;��H;��H;��H;��H;E�H;��H;�I;�I;�I;�
I;cI;�I;$I;~I;�I;�I;{!I;�#I;&I;�'I;)I;�)I;      U:I;�9I;�8I;`7I;'5I;X2I;3/I;|+I;�'I;n#I;I;�I;�I;gI;MI;Y
I;�I;,I; I;(�H;x�H;�H;��H;��H;:�H;��H;d�H;A�H;2�H;h�H;��H;,�H;��H;N�H;�H;��H;��H;��H;�H;M�H;��H;-�H;��H;e�H;4�H;A�H;d�H;��H;9�H;��H;��H;�H;t�H;*�H; I;/I;�I;[
I;NI;gI;�I;�I;I;q#I;�'I;}+I;3/I;X2I;$5I;`7I;�8I;�9I;      DOI;�NI;�MI;�KI;�HI;EI;�@I;'<I;!7I;�1I;P,I;�&I;9!I;�I;�I;�I;LI;�I;�I;NI;�H;&�H;��H;$�H;�H;5�H;��H;g�H;<�H;=�H;e�H;��H;2�H;��H;�H;_�H;[�H;_�H;�H;��H;2�H;��H;e�H;;�H;<�H;d�H;��H;3�H;�H;$�H;��H;&�H;�H;MI;�I;�I;LI;�I;�I;�I;9!I;�&I;Q,I;�1I;"7I;*<I;�@I;EI;�HI;�KI;�MI;�NI;      �bI;�bI;(bI;�`I;�^I;�[I;>WI;�QI;`KI;oDI;S=I;26I;/I;,(I;�!I;RI;mI;#I;6I;�I;�I;��H;��H;��H;[�H;,�H;d�H;��H;Z�H;=�H;4�H;u�H;��H;g�H;	�H;��H;��H;��H;
�H;g�H;��H;w�H;4�H;<�H;Z�H;��H;f�H;*�H;X�H;��H;��H;��H;�I;�I;4I;%I;lI;UI;�!I;,(I;/I;26I;S=I;pDI;cKI;�QI;AWI;�[I;�^I;�`I;)bI;�bI;      �GI;FII;PMI;SI;lYI;�^I;
bI;�bI;`I;~ZI;�RI;�II;�@I;�7I;I/I;W'I;�I;�I;�I;=I;%I;�I;��H;'�H;�H;��H;M�H;C�H;��H;j�H;A�H;F�H;��H;�H;��H;|�H;r�H;|�H;��H;�H;��H;G�H;?�H;e�H;��H;C�H;M�H;��H;�H;'�H;��H;�I;I;=I;�I; I;�I;Y'I;I/I;�7I;�@I;�II;�RI;~ZI;`I;�bI;
bI;�^I;yYI;SI;PMI;OII;      ��H;ʗH;d�H;��H;�H;�I;&I;AI;yTI;Z_I;*bI;Q^I;�UI;BKI;v@I;?6I;�,I;"$I;'I;2I;�I;W	I;hI;, I;k�H;U�H;��H;O�H;i�H;��H;h�H;K�H;v�H;��H;u�H;"�H;
�H; �H;v�H;��H;v�H;K�H;h�H;��H;f�H;M�H;��H;U�H;h�H;) I;gI;W	I;�I;1I;'I;#$I;�,I;=6I;v@I;BKI;�UI;Q^I;+bI;Z_I;zTI;AI;&I;�I;�H;��H;_�H;��H;      �VF;|hF;��F;�F;�MG;�G;�#H;քH;��H;RI;�@I;�XI;�aI;�^I;UI;�HI;�<I;�1I;�'I;�I;*I;PI;6
I;�I;T I;��H;S�H;��H;,�H;9�H;��H;��H;{�H;��H;B�H;��H;��H;��H;C�H;��H;z�H;��H;��H;6�H;*�H;��H;Q�H;��H;S I;�I;6
I;OI;%I;�I;�'I;�1I;�<I;�HI;	UI;�^I;�aI;�XI;�@I;SI;��H;քH;�#H;�G;�MG; �F;ޛF;rhF;      ��@;~�@;�`A;�&B;\C;04D;�ME;WF;'@G;W�G;�H;'�H;7I;�WI;eaI;\\I;'PI;{BI; 6I;�*I;!I;sI; I;�
I;+I;Z I;n�H;!�H;_�H;�H;?�H;��H;��H;��H;�H;��H;��H;��H;�H;��H;��H;��H;?�H;�H;\�H;!�H;l�H;Z I;*I;�
I;�I;sI;!I;�*I; 6I;~BI;%PI;]\I;eaI;�WI;7I;'�H;�H;W�G;'@G;WF;�ME;04D;XC;�&B;�`A;|�@;      �Y4;^�4;��5;�7;ݫ9;<;ן>;�A;S@C;iE;��F;`�G;�}H;��H;�?I;]I;L`I;�UI;'GI;;9I;-I;i"I;9I;^I;�
I;�I;) I;%�H;��H;%�H;��H;3�H;��H;��H;��H;��H;��H;��H;�H;��H;��H;3�H;��H;!�H;��H;%�H;' I;�I;�
I;[I;6I;i"I;-I;;9I;'GI;�UI;K`I;]I;�?I;��H;�}H;`�G;��F;gE;S@C;�A;ן>;<;�9;�7;��5;S�4;      e�;8�;��;0";�&;ӆ+;¹0;��5;�:;w�>;� B;ݠD;�F;��G;0�H;I;7SI;+aI;�YI;\JI;O;I;(.I;�"I;;I;�I;9
I;iI;��H;��H;��H;��H;��H;6�H;�H;.�H;��H;��H;��H;.�H;�H;5�H;��H;��H;��H;��H;��H;gI;:
I;�I;6I;�"I;(.I;I;I;]JI;�YI;-aI;7SI;I;1�H;��G;�F;ݠD;� B;t�>;�:;��5;¹0;Ն+;
�&;0";��;(�;      "��:���:��:��:��;tN;�L;�, ;�f);Ó1;x8;�=;�&B;E;WG;JKH;��H;�GI;c`I;�[I;�KI;�;I;'.I;j"I;rI;PI;W	I;�I;��H;)�H;�H;��H;��H;X�H;{�H;��H;��H;��H;{�H;X�H;��H;��H;�H;%�H;��H;�I;S	I;PI;oI;g"I;$.I;�;I;�KI;�[I;c`I;�GI;��H;JKH;XG;E;�&B;�=;x8;1;�f);�, ;�L;tN;��;��:��:���:      ���9��:�":X�Q:�:���:�?�:���:�M
;#�;P�&;6'1;�`9;�m?;��C;lVF;[�G;��H;�=I;�_I;H\I;�KI;O;I;	-I;	!I;,I;�I;"I;�I;�H;q�H;��H;s�H;��H;��H;�H;��H;�H;��H;��H;s�H;��H;q�H;�H;�I;"I;�I;,I;	!I;-I;N;I;�KI;F\I;�_I;�=I;��H;Z�G;lVF;��C;�m?;�`9;7'1;P�&;!�;�M
;���:�?�:���:�:X�Q:�":��:      J�Ѻ��Ⱥ����X������%�(��9��Z:ٰ�:���:K0;<S;af);J�4;�<;LB;�E;T�G;��H;�:I;�_I;�[I;\JI;=9I;�*I;�I;/I;9I;�I;JI;&�H;��H;L�H;i�H;4�H;n�H;"�H;m�H;4�H;i�H;K�H;��H;$�H;GI;�I;9I;-I;�I;�*I;99I;WJI;�[I;�_I;�:I;��H;V�G;�E;LB;�<;H�4;af);<S;K0;���:װ�:��Z:(��9�%�p��X��������Ⱥ      �5���R��S ��6��7�X�.�$��ۺ�H[��Q�@d,:�:l�:�>;s1";ո0;��:;vaA;dE;)�G;��H;�=I;d`I;�YI;'GI;6I;�'I;'I;�I;4I;�I; I;>�H;[�H;/�H;��H;��H;y�H;��H;��H;2�H;Z�H;?�H; I;�I;2I;�I;%I;�'I;6I;#GI;�YI;c`I;�=I;��H;)�G;dE;vaA;��:;ָ0;s1";�>;l�:�:@d,: Q�|H[��ۺ*�$�1�X�6��S ���R��      H",���(�7H�DG��.���jλ!R��^e�A����� �W�$�Z:���:Z�;��;��-;��9;�A;dE;V�G;��H;�GI;-aI;�UI;zBI;�1I;%$I;I;%I;�I;-I;��H;��H;�H;B�H;N�H;!�H;N�H;D�H;�H;��H;��H;-I;�I;#I;I;"$I;�1I;xBI;�UI;+aI;�GI;��H;Y�G;dE;�A;��9;��-;��;[�;���:$�Z: �W����?��~^e�!R���jλ�.��DG�7H���(�      �d��B��������)���zl�RH��k"�r.���W��N�k�i� �(����9���:���:5�;�-;��9;vaA;�E;Y�G;��H;:SI;K`I; PI;�<I;�,I;�I;lI;GI;�I;�I;��H;��H;�H;��H;��H;��H;�H;��H;��H;�I;�I;GI;iI;�I;�,I;�<I; PI;G`I;4SI;��H;Y�G;�E;vaA;��9;�-;8�;���:���:��9(��i� �N�k��W��q.���k"�RH��zl��)������C���      ���j9�]5��=��Vb̼~֮�t��� d�",�����Q��2G5�8#��`�f9���:��:9�;��-;��:;LB;lVF;KKH;I;]I;Y\I;�HI;?6I;W'I;UI;�I;R
I;yI;4 I;��H;��H;��H;$�H;��H;��H;��H;3 I;yI;R
I;�I;PI;W'I;<6I;�HI;Z\I;]I;I;KKH;jVF;LB;��:;��-;9�;��:���:`�f98#��/G5��Q�����",�� d�t��}֮�Vb̼=��]5��j9�      �]��IY��ZN��`=���'�o����䷾������W��$�^��Y�X�����@9���:���:��;Ҹ0;�<;��C;TG;1�H;�?I;`aI;UI;s@I;H/I;�!I;�I;HI;�I;�I;�H;��H;B�H;��H;B�H;��H;�H;�I;�I;HI;�I;�!I;H/I;r@I;
UI;baI;�?I;,�H;TG;��C;�<;Ҹ0;��;���:���:@9����Y�X�]���$��W�����䷾����n���'��`=��ZN��IY�      �A��!��e���*��轅�@�d��`=����^��e֮�L�y�z�(��һ�]e�������f9���:[�;p1";L�4;�m?;E;��G;��H;�WI;�^I;?KI;�7I;,(I;�I;]I;�
I;ZI;TI;��H;�H;s�H;�H;��H;TI;XI;�
I;_I;�I;*(I;�7I;>KI;�^I;�WI;��H;��G;E;�m?;L�4;p1";^�;���:��f9�����]e��һy�(�L�y�e֮�^�꼙���`=�@�d�轅��*��e��!��      ���IE	��������Wн�A�����h���3����"¼�)��-x/��һW�X�6#����9���:�>;bf);�`9;�&B;�F;�}H;7I;�aI;�UI;�@I;/I;1!I;I;[I;I;�I;� I;��H;2�H;��H;� I;�I;I;[I;I;1!I;
/I;�@I;�UI;�aI;7I;�}H;�F;�&B;�`9;bf);�>;���:��96#��V�X��һ-x/��)��"¼�����3��h��󑽤A���Wн��콼��IE	�      �^Z�c
V��I��6�������ܽ!��ܽ���aG�\��ȼ�)��z�(�]��2G5�(���Z:f�:<S;3'1;�=;ܠD;[�G; �H;�XI;M^I;�II;,6I;�&I;�I;�I;�
I;�I;�I;� I;��H;� I;�I;�I;�
I;�I;�I;�&I;+6I;�II;J^I;�XI;#�H;Z�G;ؠD;�=;6'1;>S;f�:$�Z:0��3G5�\��z�(��)���ȼ\��aG�ܽ��!���ܽ������6��I�c
V�      � ��f�����ݕ����q��I���"���������k���ZN�\�"¼N�y��$��Q��k� � �W��:K0;N�&;x8;� B;��F;	�H;�@I;&bI;�RI;P=I;F,I;I;I;�I;I;nI;QI;�I;QI;nI;I;�I;I;I;F,I;M=I;�RI;$bI;�@I;�H;��F;� B;x8;O�&;J0;�: �W�m� ��Q���$�N�y�"¼\��ZN�k������������"��I���q�ݕ�����f��      f5�������Z�Ҿ�a��}����l��6�FE	���Ƚk���aG����e֮��W����O�k����<d,:���: �;��1;t�>;gE;W�G;SI;U_I;vZI;lDI;�1I;e#I;wI;-I;9
I;@I;I;UI;I;@I;9
I;,I;wI;g#I;�1I;iDI;vZI;T_I;SI;X�G;eE;s�>;��1;!�;���:<d,:���Q�k�����W�e֮�����aG�k����ȽFE	��6��l�}����a��Z�Ҿ������      }A��q<�ha/����:�}]׾� ��
w��>�FE	�����ܽ����3�`�꼘���
",��W��D���Q�װ�:�M
;�f);�:;N@C;"@G;��H;sTI;�_I;\KI;7I;�'I;�I;�I;rI;I;�I;�I;�I;I;rI;�I;�I;�'I;7I;YKI;�_I;pTI;��H;%@G;K@C;�:;�f);�M
;Ӱ�:�Q�B���W��
",�����`�꼛�3�ܽ������FE	�>�
w��� ��}]׾�:���ha/��q<�      w�������c�{�m$_��q<������~��
w���6�����!���h����䷾�� d�t.��~^e��H[���Z:���:�, ;��5;�A; WF;ׄH;AI;�bI;�QI;<I;r+I;�I;?I;mI;�	I;I;bI;I;�	I;mI;=I;�I;t+I;<I;�QI;�bI;AI;քH;WF;�A;��5;�, ;���:��Z:�H[�}^e�t.��� d�䷾�����h�!�������6�
w��~��������q<�m$_�c�{�����      =��������欿�������O��x����� ���l���"��ܽ���`=����v���k"�"R��ۺ(��9�?�:�L;��0;ӟ>;�ME;�#H;�%I;bI;7WI;�@I;&/I;s!I;oI;7I;@I;~I;�I;~I;@I;7I;mI;s!I;&/I;�@I;7WI;bI;�%I;�#H;�ME;П>;��0;�L;�?�:��9ۺ"R���k"�v������`=����ܽ��"��l�� ����뾃x���O�������欿����      �������O��lȿl���������O���}]׾}����I�����A��A�d�o�~֮�	RH��jλ5�$��%����:hN;̆+;<;*4D;�G;�I;�^I;�[I;EI;U2I;�#I;tI;�I;�I;�	I;�I;�	I;�I;�I;qI;�#I;U2I;EI;�[I;�^I;�I;�G;,4D;�<;̆+;hN;���:�%�5�$��jλ
RH�~֮�o�A�d��A������I�}���}]׾����O�����m���lȿO�Ῥ��      @�4i�������K�ѿm������q<��:��a����q����Wн齅���'�Vb̼�zl��.��5�X�����:��;
�&;߫9;TC;�MG;�H;hYI;�^I;�HI;5I;&I;I;;I;�I;�
I;�	I;�
I;�I;;I;I;&I;5I;�HI;�^I;hYI;	�H;MG;VC;ܫ9;�&;��;�:���5�X��.���zl�Vb̼��'�齅��Wн����q��a���:��q<���m���K�ѿ������4i�      I:�.5�0�'� ������lȿ���m$_���Z�Ҿޕ���6�����*���`=�>�漭)��FG�6��X��h�Q:�:0";�7;�&B;�F;��H;SI;�`I;�KI;P7I;�'I;nI;LI;�I;�I;�
I;�I;�I;LI;lI;�'I;P7I;�KI;�`I;SI;��H;�F;�&B;�7;0";�:p�Q:Z��6��EG��)��>���`=��*������6�ޕ��Z�Ҿ��m$_����lȿ���� ��0�'�.5�      ��U�\�O�J-?�0�'���O�ῶ欿c�{�ha/���뾟���I����f���ZN�`5������9H�Z �������":��:��;��5;�`A;�F;b�H;FMI;&bI;�MI;�8I;)I;sI;I;rI;8I;9I;8I;rI;I;qI;)I;�8I;�MI;%bI;FMI;b�H;��F;�`A;��5;��;��:��":���Z ��9H�����`5���ZN�f������I�������ha/�c�{��欿O����0�'�J-?�\�O�      ��i���b�\�O�.5�4i�������������q<����f��c
V�IE	�!���IY�k9�D�����(��R����Ⱥ��:���:$�;L�4;p�@;qhF;ƗH;@II;�bI;�NI;�9I;�)I;I;�I;�I;�I;�I;�I;�I;�I;I;�)I;�9I;�NI;�bI;@II;ŗH;qhF;p�@;I�4;*�;���:��:��Ⱥ�R����(�D���k9��IY�!��IE	�c
V�f������q<������������4i�.5�\�O���b�      �>���8���*�O������˿p��H�b�E\�7m־^��T�:��J�+��I�B�?��������'/��쯕��>:�t�:Vp ;�J6;EA;�IF;�NH;�H;"I;�I;#I;�I;�I;I;� I;��H;:�H;��H;� I;I;I;�I;#I;�I;"I;�H;�NH;�IF;EA;�J6;Yp ;�t�:�>:�'/���������@��I�B�+���J�T�:�^��7m־E\�H�b�p���˿����O���*���8�      ��8��4��g&�7��>����<ƿ򲗿�>]�î�S�Ѿ�p���*7����'W��PR?�}�p8�������p�����G:� �:�!;�6;&lA;�YF;�TH;{�H;)"I;�I;�I;�I;YI;I;s I;��H;"�H;��H;u I;I;WI;�I;�I;�I;'"I;{�H;�TH;�YF;&lA;�6;�!;� �:��G:r��������p8��}�PR?�'W�����*7��p��S�Ѿî��>]�򲗿�<ƿ>���7���g&��4�      ��*��g&��#�v�X[�rL�������M�t5��>ľ����,��D�뒐��5�4�ݼ���q
��x�`tk��b:_l�:#;ӗ7;��A;�F;�dH;�I;i"I;I;{I;QI;I;�I;3 I;��H;��H;��H;1 I;�I;I;QI;{I;I;f"I;�I;�dH;��F;��A;З7;#;_l�:�b:`tk��x��q
���4�ݼ�5�뒐��DὬ�,����>ľs5���M����rL��X[�v��#��g&�      O�7��v����˿B1��9�y�Ŏ6��z �����5�l�+��ͽ&�����&���˼?�k������X�D� ����:T�;&;�9;��B;�F;�}H;�	I;u"I;@I;�I;�I;�I;[I;��H;6�H;��H;6�H;��H;[I;�I;�I;�I;>I;r"I;�	I;�}H;�F;��B;�9; &;T�;���:D� ���X����@�k���˼��&�&����ͽ+�5�l������z �Ŏ6�9�y�B1���˿���v�7��      ����>���X[忸˿�T���~�R�î��E۾՗����M���	� �����j��3�d����O�4�׻��/����d��:� 
;*;f;;�jC;�'G;��H;I;"I;I;�I;�
I;�I;�I;W�H;��H;�H;��H;W�H;�I;�I;�
I;�I;�I;"I;I;��H;�'G;�jC;e;;*;� 
;f��:�����/�4�׻��O�d���3���j� �����	���M�՗���E۾î�~�R���T���˿X[�>���      �˿�<ƿrL��B1����>]���)�%��ֳ���{���,�u��)��T`I��J���,���3/��+���� ��/69�4�:�;p.;,.=;raD;��G;r�H;�I;O!I;kI;^I;�	I;�I;� I;��H;&�H;v�H;&�H;��H;� I;�I;�	I;`I;hI;K!I;�I;q�H;��G;qaD;*.=;p.;�;�4�:�/69�� ��+���3/��,���J��T`I�)��u�齦�,���{�ֳ�%����)��>]��B1��rL���<ƿ      p��򲗿���9�y�~�R���)�ov��>ľ^���I�Zl����������&�֮Ҽ�}�.B�Į������<�!:+�:Dz;�3;ij?;�\E;��G;��H;}I;�I;�I;�I;�I;�I;. I;��H;v�H;��H;v�H;��H;. I;�I;�I;�I;�I;�I;}I;��H;��G;�\E;ej?;�3;Dz;+�:0�!:����®��.B��}�֮Ҽ��&��������Zl��I�^���>ľov���)�~�R�9�y����򲗿      G�b��>]���M�Ŏ6�î�%���>ľ$q��|�Z�+�U9ݽ#W����L����#F���G��׻�;�Xn��Ȋ:�i;(P$;�7;x�A;JF;BCH;��H;� I;zI;�I;+I;@I;�I;,�H;��H;��H;#�H;��H;��H;,�H;�I;AI;+I;�I;xI;� I;��H;ACH;JF;t�A;�7;&P$;�i;�Ȋ:`n��;��׻�G�#F�������L�#W��U9ݽ+�|�Z�$q���>ľ%��î�Ŏ6���M��>]�      E\�î�s5��z ��E۾ֳ�^��|�Z�N?#����A����j�'��Fϼ����������lۺX:�9�4�:`�;n�,;��;;D�C;�G;]�H;�I;�!I;�I;RI;;I;�I;SI;0�H;�H;��H;6�H;��H;�H;0�H;SI;�I;:I;QI;�I;�!I;�I;\�H;�G;C�C;��;;l�,;b�;�4�:h:�9�lۺ���������Fϼ'����j��A�����N?#�|�Z�^��ֳ��E۾�z �s5�î�      7m־S�Ѿ�>ľ����՗����{��I�+�����V���{�A�/�(���,��==�>�һR�@�ؖ �$�k:!�:b;��3;@j?;x2E;��G;|�H;CI;� I;�I;�I;4	I;I;��H;�H;��H;��H;m�H;��H;��H;�H;��H;I;4	I;�I;�I;� I;BI;|�H;��G;u2E;?j?;��3;b;�:$�k:Ԗ �S�@�>�һ==��,��(��A�/��{��V�����+��I���{�՗�������>ľS�Ѿ      ^���p����4�l���M���,�Zl�T9ݽ�A���{� �5��J��
;���T[�?�����P���P�9��:��;5*;0�9;kkB;�F;�NH;��H;/ I;�I;�I;/I;"I;UI;w�H;��H;��H;��H;��H;��H;��H;��H;u�H;XI;!I;/I;�I;�I;, I;��H;�NH;݇F;ikB;0�9;3*;��;��: Q�9 P������?��T[�
;���J�� �5��{��A��U9ݽZl���,���M�4�l����p��      T�:��*7���,�+���	�u�齅���#W����j�@�/��J���I���k�i�.��N��0 ��Ɋ:so�:";kr3;0�>;<�D;|�G;]�H;I;>!I;�I;�I;�
I;I;v I;��H;��H;��H;��H;y�H;��H;��H;��H;��H;y I;I;�
I;�I;�I;=!I;I;Z�H;x�G;:�D;.�>;kr3; ;so�:
Ɋ:8 ��N��.��j��k��I���J��@�/���j�#W������u�齄�	�+���,��*7�      �J�����D��ͽ ���)�������L�'��(��
;���k����cI����/�0/���>:Y��:�B;r�,;��:;?�B;�xF;�<H;�H;I;�I;�I;XI;�I;�I;��H;��H;N�H;��H;��H;��H;��H;��H;N�H;��H;��H;�I;�I;VI;�I;�I;I;�H;�<H;�xF;>�B;��:;r�,;�B;]��:��>:,/���/�cI������k�
;��'��'����L����)�� ����ͽ�D����      +��'W��뒐�%�����j�S`I���&����Fϼ�,���T[�h�cI��M;�@nk��:<5�:�;&;�6;�!@;H2E;�G;��H;I;!I;dI;%I;I;NI;� I;��H;�H;��H;z�H;��H;a�H;��H;z�H;��H;�H;��H;� I;PI;I;%I;cI;!I; I;��H;�G;H2E;�!@;�6;&;�;:5�:�:<nk�L;�cI��i��T[��,��Fϼ�����&�S`I���j�%���뒐�'W��      H�B�OR?��5���&��3��J��֮Ҽ#F����>=�?�.����/�Lnk�Ю�9b׳:��;B!;h3;�=;��C;2�F;'dH;�H;�I;&I;�I;:I;�I;�I;\�H;�H;��H;��H;[�H;��H;S�H;��H;\�H;��H;��H;�H;\�H;�I;�I;:I;�I;&I;�I;�H;"dH;1�F;��C;�=;h3;D!;��;b׳:Ю�9Lnk���/�.��?�==���#F��֮Ҽ�J���3���&��5�PR?�      >��}�2�ݼ��˼d���,���}��G����>�һ����M��0/��:j׳:�;|b;£0;�<;��B;�IF;�H;<�H;�I;� I;1I;PI;r
I;�I;8 I;H�H;l�H;%�H;@�H;;�H;��H;U�H;��H;;�H;?�H;#�H;m�H;H�H;: I;�I;r
I;MI;1I;� I;�I;6�H;�H;�IF;��B;�<;ģ0;zb;�;j׳:�:0/�N������>�һ����G��}��,��d����˼2�ݼ}�      ����o8����>�k���O��3/�,B��׻����Q�@�P��0 ����>::5�:��;xb;��/;>;;O�A;��E;ԿG;	�H;�
I;~ I;I;I;�I;�I;�I;��H;X�H;��H;��H;�H;/�H;��H;M�H;��H;/�H;�H;��H;��H;X�H;��H;�I;�I;�I;I;I;y I;�
I;	�H;ҿG;��E;O�A;@;;��/;xb;��;:5�:��>:0 ��P��Q�@������׻,B��3/���O�>�k���p8��      ������q
����4�׻�+��®���;��lۺؖ �Q�9Ɋ:Y��:�;D!;��0;?;;ѓA;�pE;��G;�H;��H;�I;OI;pI;;I;�I;�I;�H;^�H;��H; �H;<�H;�H;�H;~�H;W�H;~�H;�H;�H;;�H;!�H;��H;]�H;�H;�I;�I;;I;pI;KI;�I;��H;ߎH;��G;�pE;ғA;>;;��0;C!;�;Y��:Ɋ:Q�9Ԗ ��lۺ�;�®���+��2�׻����q
���      "/�������x���X���/��� �����Xn칀:�9$�k:��:yo�:�B;&;l3;�<;O�A;�pE;ttG;}H;C�H;?I;�I;]I;I;�
I;I;n I;l�H;@�H;��H;��H;��H;��H;�H;��H;��H;��H;�H;��H;��H;��H;��H;=�H;h�H;n I;I;�
I;I;XI;�I;AI;>�H;}H;ttG;�pE;N�A;�<;l3;&;�B;yo�:��: �k:�:�9`n������� ���/���X���x����      毕�N���Ltk�@� �����/690�!:�Ȋ:�4�:!�:��; ;r�,;�6; �=;��B;��E;��G;}H;��H;�I;+ I;�I;tI;�I;FI;�I;e�H;�H;Z�H;�H;/�H;��H;��H;�H;��H;��H;��H;�H;��H;��H;0�H;�H;W�H;�H;e�H;�I;DI;�I;pI;�I;+ I;�I;��H;}H;��G;��E;��B; �=;�6;r�,;;��;!�:�4�:�Ȋ:0�!:�/69���@� �Dtk�b���      (�>:��G:�b:���:V��:�4�:+�:�i;b�;b;6*;ir3;��:;�!@;��C;�IF;׿G;�H;A�H;�I;5 I;]I;UI;�I;0I;{I;=�H;��H;��H;��H;h�H;��H;��H;��H;2�H;��H;��H;��H;2�H;��H;��H;��H;h�H;��H;��H;��H;:�H;{I;0I;�I;SI;]I;2 I;�I;C�H;�H;տG;�IF;��C;�!@;��:;kr3;3*;b;c�;�i;+�:�4�:X��:���: �b:��G:      �t�:� �:}l�:L�;� 
;��;Mz;0P$;r�,;��3;6�9;2�>;A�B;K2E;5�F;�H;�H;��H;AI;- I;[I;�I;TI;�I;I;��H;A�H;l�H;��H;��H;�H;��H;��H;��H;U�H;�H;��H;�H;U�H;��H;��H;��H;�H;��H;��H;l�H;>�H;��H;I;�I;SI;�I;ZI;. I;AI;��H;
�H;�H;6�F;K2E;A�B;2�>;4�9;��3;s�,;/P$;Nz;�;� 
;M�;�l�:� �:      Zp ;�!;#;&;*;p.;�3;�7;��;;Bj?;pkB;?�D;�xF;�G;'dH;9�H;�
I;�I;�I;�I;UI;UI;�I;uI;R�H;��H;��H;G�H;�H;5�H;��H;��H;��H;�H;v�H;;�H;&�H;;�H;v�H;	�H;��H;��H;��H;2�H;�H;H�H;��H;��H;S�H;rI;�I;WI;RI;�I;�I;�I;�
I;8�H;'dH;�G;�xF;?�D;mkB;@j?;��;;�7;�3;p.;*;&;#;�!;      �J6;/�6;ܗ7;�9;i;;+.=;sj?;w�A;H�C;y2E;�F;��G;�<H;��H;�H;�I;| I;PI;[I;tI;�I;�I;tI;j�H;��H;��H;��H;O�H;]�H;��H;��H;��H;��H;I�H;��H;��H;k�H;��H;��H;I�H;��H;��H;��H;��H;[�H;O�H;��H;��H;��H;g�H;rI;�I;�I;tI;]I;RI;| I;�I;�H;��H;�<H;��G;�F;x2E;H�C;x�A;qj?;,.=;p;;�9;ݗ7;�6;      EA;4lA;q�A;��B;kC;vaD;�\E;JF;�G;��G;�NH;`�H;�H;I;�I;� I;I;rI;I;�I;3I;I;V�H;��H;�H;��H;W�H;k�H;��H;��H;��H;��H;��H;��H;�H;��H;��H;��H;�H;��H;��H;��H;��H;��H;��H;k�H;T�H;��H;�H;��H;V�H;I;2I;�I;I;uI;I;� I;�I;I;�H;a�H;�NH;��G;�G;JF;�\E;vaD;kC;��B;r�A;4lA;      �IF;�YF;�F;�F;�'G;�G;��G;=CH;]�H;|�H;��H;I;I;!I;%I;/I;I;:I;�
I;CI;xI;��H;��H;��H;��H;��H;��H;��H;��H;��H;��H;��H;W�H;��H;t�H;V�H;G�H;V�H;u�H;��H;T�H;��H;��H;��H;��H;��H;��H;��H;��H;��H;��H;��H;tI;CI;�
I;;I;I;-I;%I;!I;I;I;��H;{�H;]�H;=CH;��G;�G;�'G;�F;�F;�YF;      �NH;�TH;�dH;�}H;��H;z�H;��H;��H;�I;GI;2 I;D!I;�I;gI;�I;PI;�I;�I;I;�I;=�H;A�H;��H;��H;Q�H;��H;��H;��H;��H;��H;��H;�H;��H;,�H;��H;��H;��H;��H;��H;*�H;��H;�H;��H;��H;��H;��H;��H;��H;T�H;��H;��H;B�H;<�H;�I;I;�I;�I;NI;�I;fI;�I;D!I;0 I;DI;�I;��H;��H;u�H;��H;�}H;�dH;�TH;      	�H;}�H;�I;�	I;I;�I;�I;� I;�!I;� I;�I;�I;�I;)I;<I;t
I;�I;�I;l I;h�H;��H;l�H;G�H;P�H;f�H;��H;��H;��H;��H;��H;�H;o�H;
�H;��H;p�H;@�H;7�H;@�H;p�H;��H;	�H;o�H;�H;��H;��H;��H;��H;��H;i�H;P�H;G�H;l�H;��H;h�H;l I;�I;�I;r
I;<I;(I;�I;�I;�I;� I;�!I;� I;�I;�I;I;�	I;�I;��H;      $"I;/"I;e"I;{"I;"I;O!I;�I;�I;�I;�I;�I;�I;[I;I;�I;�I;�I;�H;k�H;�H;��H;��H;�H;_�H;��H;��H;��H;��H;��H;
�H;d�H;��H;��H;0�H;��H;��H;��H;��H;��H;0�H;~�H;��H;d�H;�H;��H;��H;��H;��H;��H;`�H;�H;��H;��H;�H;k�H;�H;�I;�I;�I;I;XI;�I;�I;�I;�I;�I;�I;O!I;"I;{"I;h"I;'"I;      �I;�I;I;BI;I;sI;�I;�I;]I;�I;<I;�
I;�I;ZI;�I;> I;��H;Z�H;=�H;\�H;��H;��H;/�H;��H;��H;��H;��H;��H;�H;V�H;��H;z�H;�H;��H;��H;��H;o�H;��H;��H;��H;��H;|�H;��H;U�H;�H;��H;��H;��H;��H;��H;.�H;��H;��H;\�H;=�H;\�H;��H;; I;�I;WI;�I;�
I;9I;�I;_I;�I;�I;rI;I;BI;I;�I;      )I;I;�I;�I;�I;aI;�I;5I;HI;=	I;-I;I;�I;� I;c�H;Q�H;_�H;��H;��H;�H;n�H;��H;��H;��H;��H;��H;��H;�H;c�H;��H;]�H;��H;��H;t�H;C�H;&�H;�H;&�H;C�H;t�H;��H;��H;]�H;��H;d�H;�H;��H;��H;��H;��H;��H;��H;k�H;�H;��H;��H;\�H;O�H;b�H;� I;�I;I;*I;=	I;GI;5I;�I;bI;�I;�I;�I;I;      �I;�I;[I;�I;�
I;�	I;�I;II;�I;I;]I;� I;��H;��H;!�H;w�H;��H;"�H;��H;7�H;��H;��H;��H;��H;��H;��H;�H;o�H;��H;{�H;��H;��H;Z�H;2�H;��H;��H;��H;��H;��H;2�H;W�H;��H;��H;|�H;��H;o�H;�H;��H;��H;��H;��H;��H;��H;7�H;��H;$�H;��H;v�H;�H;��H;��H;� I;\I;I;�I;HI;�I;�	I;�
I;�I;ZI;�I;      �I;nI;I;�I;�I;�I;�I;�I;^I;��H;~�H;��H;��H;"�H;��H;,�H;��H;:�H;��H;��H;��H;��H;��H;��H;��H;T�H;��H;�H;��H;�H;��H;[�H;�H;��H;��H;��H;��H;��H;��H;��H;�H;^�H;��H;�H;��H;�H;��H;S�H;��H;��H;��H;��H;��H;��H;��H;;�H;��H;*�H;��H;$�H;��H;��H;{�H;��H;\I;�I;�I;�I;�I;�I;I;hI;      %I;I;�I;gI;�I;� I;7 I;9�H;9�H;�H;��H;��H;S�H;��H;��H;I�H;"�H;�H;��H;��H;��H;��H;	�H;L�H;y�H;��H;&�H;��H;/�H;��H;s�H;2�H;��H;��H;��H;��H;r�H;��H;��H;��H;��H;6�H;q�H;��H;2�H;��H;&�H;��H;z�H;J�H;	�H;��H;��H;��H;��H;	�H;�H;I�H;��H;��H;S�H;��H;��H;�H;<�H;9�H;7 I; I;�I;gI;�I;I;      � I;� I;B I;��H;y�H;��H;��H;�H;%�H;�H;��H;��H;��H;��H;b�H;C�H;9�H;�H;�H;�H;9�H;U�H;q�H;��H;�H;n�H;��H;n�H;��H;��H;@�H;��H;��H;��H;l�H;b�H;d�H;b�H;l�H;��H;��H; �H;@�H;��H;��H;n�H;��H;n�H;�H;��H;q�H;U�H;6�H;�H;�H;�H;6�H;C�H;a�H;��H;��H;��H;��H;�H;%�H;	�H;��H;��H;o�H;��H;B I;� I;      ��H;��H;��H;?�H;��H;$�H;��H;��H;��H;��H;��H;��H;��H;��H;��H;��H;��H;z�H;��H;��H;��H;�H;9�H;��H;��H;O�H;��H;@�H;��H;��H;$�H;��H;��H;��H;b�H;H�H;H�H;H�H;b�H;��H;��H;��H;$�H;��H;��H;@�H;��H;N�H;��H;��H;9�H;�H;��H;��H;��H;{�H;��H;��H;��H;��H;��H;��H;��H;��H;��H;��H;��H;(�H;��H;?�H;��H;��H;      ?�H;5�H;�H;��H;*�H;w�H;��H;0�H;?�H;o�H;��H;��H;��H;i�H;X�H;\�H;T�H;P�H;��H;��H;��H;��H;#�H;l�H;��H;@�H;��H;:�H;��H;q�H;�H;��H;��H;w�H;d�H;I�H;E�H;I�H;d�H;w�H;��H;��H;�H;s�H;��H;:�H;��H;A�H;��H;i�H;#�H;��H;��H;��H;��H;Q�H;R�H;\�H;X�H;j�H;��H;��H;��H;q�H;A�H;/�H;��H;|�H;�H;��H;�H;,�H;      ��H;��H;��H;?�H;��H;$�H;��H;��H;��H;��H;��H;��H;��H;��H;��H;��H;��H;z�H;��H;��H;��H;�H;8�H;��H;��H;O�H;��H;@�H;��H;��H;$�H;��H;��H;��H;b�H;H�H;H�H;H�H;b�H;��H;��H;��H;$�H;��H;��H;@�H;��H;N�H;��H;��H;9�H;�H;��H;��H;��H;{�H;��H;��H;��H;��H;��H;��H;��H;��H;��H;��H;��H;(�H;��H;?�H;��H;��H;      � I;� I;A I;��H;x�H;��H;��H;�H;%�H; �H;��H;��H;��H;��H;a�H;C�H;7�H;�H;�H;�H;:�H;U�H;q�H;��H;�H;n�H;��H;n�H;��H;��H;@�H;��H;��H;��H;l�H;b�H;d�H;b�H;l�H;��H;��H;�H;@�H;��H;��H;n�H;��H;n�H;�H;��H;q�H;U�H;6�H;�H;�H;�H;7�H;C�H;a�H;��H;��H;��H;��H;�H;%�H;	�H;��H;��H;o�H;��H;A I;� I;      &I;I;�I;gI;�I;� I;7 I;9�H;:�H;�H;��H;��H;S�H;��H;��H;I�H; �H;�H;��H;��H;��H;��H;	�H;L�H;z�H;��H;&�H;��H;.�H;��H;q�H;4�H;��H;��H;��H;��H;r�H;��H;��H;��H;��H;6�H;s�H;��H;2�H;��H;&�H;��H;y�H;J�H;	�H;��H;��H;��H;��H;	�H; �H;I�H;��H;��H;S�H;��H;��H;�H;<�H;:�H;7 I;I;�I;gI;�I;I;      �I;nI;I;�I;�I;�I;�I;�I;\I;��H;{�H;��H;��H;"�H;��H;*�H;��H;:�H;��H;��H;��H;��H;��H;��H;��H;T�H;��H;�H;��H;�H;��H;\�H;�H;��H;��H;��H;��H;��H;��H;��H;�H;_�H;��H;�H;��H;�H;��H;T�H;��H;��H;��H;��H;��H;��H;��H;:�H;��H;,�H;��H;"�H;��H;��H;~�H;��H;_I;�I;�I;�I;�I;�I;I;kI;      �I;�I;[I;�I;�
I;�	I;�I;KI;�I;I;\I;� I;��H;��H;�H;v�H;��H;"�H;��H;9�H;��H;��H;��H;��H;��H;��H;�H;o�H;��H;{�H;��H;��H;X�H;2�H;��H;��H;��H;��H;��H;2�H;W�H;��H;��H;|�H;��H;o�H;�H;��H;��H;��H;��H;��H;��H;7�H;��H;$�H;��H;w�H;�H;��H;��H;� I;]I;I;�I;II;�I;�	I;�
I;�I;[I;�I;      )I;I;�I;�I;�I;aI;�I;5I;GI;<	I;,I;I;�I;� I;b�H;P�H;\�H;��H;��H;�H;n�H;��H;��H;��H;��H;��H;��H;�H;a�H;��H;]�H;��H;��H;t�H;C�H;&�H;�H;&�H;C�H;t�H;��H;��H;]�H;��H;d�H;�H;��H;��H;��H;��H;��H;��H;k�H;�H;��H;��H;]�H;Q�H;c�H;� I;�I;I;,I;?	I;HI;6I;�I;bI;�I;�I;�I;I;      �I;�I;I;AI;I;nI;�I;�I;_I;�I;9I;�
I;�I;XI;�I;; I;��H;Z�H;=�H;]�H;��H;��H;/�H;��H;��H;��H;��H;��H;�H;V�H;��H;z�H;�H;��H;��H;��H;o�H;��H;��H;��H;�H;{�H;��H;U�H;
�H;��H;��H;��H;��H;��H;.�H;��H;��H;\�H;=�H;\�H;��H;? I;�I;XI;�I;�
I;<I;�I;`I;�I;�I;rI;I;AI;I;�I;      "I;,"I;k"I;y"I;"I;M!I;�I;�I;�I;�I;�I;�I;YI;I;�I;�I;�I;�H;k�H;�H;��H;��H;�H;`�H;��H;��H;��H;��H;��H;
�H;d�H;��H;�H;0�H;��H;��H;��H;��H;��H;0�H;�H;��H;d�H;�H;��H;��H;��H;��H;��H;_�H;�H;��H;��H;�H;k�H;�H;�I;�I;�I;I;YI;�I;�I;�I;�I;�I;�I;N!I;"I;u"I;m"I;+"I;      	�H;��H;�I;�	I;I;�I;�I;� I;�!I;� I;�I;�I;�I;)I;:I;r
I;�I;�I;l I;h�H;��H;l�H;G�H;P�H;i�H;��H;��H;��H;��H;��H;�H;o�H;	�H;��H;n�H;A�H;7�H;@�H;p�H;��H;
�H;q�H;�H;��H;��H;��H;��H;��H;f�H;P�H;F�H;l�H;��H;h�H;l I;�I;�I;u
I;<I;(I;�I;�I;�I;� I;�!I;� I;�I;�I;I;�	I;�I;��H;      �NH;�TH;�dH;�}H;��H;t�H;��H;��H;�I;FI;0 I;D!I;�I;fI;�I;PI;�I;�I;I;�I;@�H;B�H;��H;��H;T�H;��H;��H;��H;��H;��H;��H;�H;��H;*�H;��H;��H;��H;��H;��H;*�H;��H;�H;��H;��H;��H;��H;��H;��H;Q�H;��H;��H;A�H;<�H;�I;I;�I;�I;NI;�I;gI;�I;D!I;3 I;FI;�I;��H;��H;t�H;��H;�}H;�dH;�TH;      �IF;�YF;�F;�F;�'G;��G;��G;@CH;\�H;|�H;��H;I;I;!I;#I;.I;I;:I;�
I;CI;xI;��H;��H;��H;��H;��H;��H;��H;��H;��H;��H;��H;V�H;��H;r�H;V�H;G�H;V�H;u�H;��H;T�H;��H;��H;��H;��H;��H;��H;��H;��H;��H;��H;��H;tI;CI;�
I;;I;I;/I;%I;!I;I;I;��H;{�H;]�H;>CH;��G;��G;�'G; �F;�F;�YF;      EA;4lA;r�A;��B;kC;vaD;�\E;JF;�G;��G;�NH;a�H;�H;I;�I;� I;I;rI;I;�I;3I;I;W�H;��H;�H;��H;W�H;k�H;��H;��H;��H;��H;��H;��H;�H;��H;��H;��H;�H;��H;��H;��H;��H;��H;��H;k�H;V�H;��H;�H;��H;U�H;I;2I;�I;I;uI;I;� I;�I;I;�H;a�H;�NH;��G;�G; JF;�\E;vaD;kC;��B;r�A;2lA;      �J6;+�6;�7;�9;e;;/.=;mj?;x�A;J�C;{2E;�F;��G;�<H;��H;�H;�I;} I;OI;]I;tI;�I;�I;tI;j�H;��H;��H;��H;O�H;]�H;��H;��H;��H;��H;G�H;��H;��H;k�H;��H;��H;I�H;��H;��H;��H;��H;[�H;O�H;�H;��H;��H;h�H;rI;�I;�I;tI;[I;RI;| I;�I;�H;��H;�<H;��G;�F;x2E;K�C;{�A;mj?;1.=;t;;�9;�7;�6;      Wp ;!;"#;&;*;p.;�3;�7;��;;Bj?;mkB;?�D;�xF;�G;'dH;9�H;�
I;�I;�I;�I;VI;WI;�I;uI;S�H;��H;��H;H�H;�H;6�H;��H;��H;��H;	�H;v�H;;�H;&�H;;�H;v�H;�H;��H;��H;��H;2�H;�H;G�H;��H;��H;R�H;rI;�I;UI;PI;�I;�I;�I;�
I;9�H;)dH;�G;�xF;?�D;pkB;?j?;��;;�7;�3;p.;*;&;#;�!;      �t�:� �:}l�:M�;� 
;��;Nz;/P$;r�,;��3;6�9;2�>;A�B;K2E;5�F;�H;
�H;��H;AI;- I;]I;�I;UI;�I;I;��H;B�H;l�H;��H;��H;�H;��H;��H;��H;T�H;�H;��H;�H;U�H;��H;��H;��H;�H;��H;��H;l�H;>�H;��H;I;�I;QI;�I;ZI;. I;AI;��H;
�H;�H;6�F;K2E;A�B;4�>;4�9;��3;s�,;0P$;Mz;��;� 
;L�;}l�:� �:      �>:��G:(�b:���:V��:�4�:+�:�i;b�;b;5*;kr3;��:;�!@;��C;�IF;׿G;�H;C�H;�I;4 I;]I;UI;�I;0I;zI;=�H;��H;��H;��H;h�H;��H;��H;��H;2�H;��H;��H;��H;2�H;��H;��H;��H;h�H;��H;��H;��H;<�H;{I;0I;�I;SI;]I;2 I;�I;A�H;�H;տG;�IF;��C;�!@;��:;ir3;5*;b;c�;�i;+�:�4�:`��:���:,�b:��G:      毕�N���8tk�D� �����/694�!:�Ȋ:�4�:#�:��;;r�,;�6; �=;��B;��E;��G;}H;��H;�I;+ I;�I;tI;�I;DI;�I;e�H;�H;Z�H;�H;/�H;��H;��H;�H;��H;��H;��H;�H;��H;��H;0�H;�H;W�H;�H;e�H;�I;DI;�I;pI;�I;+ I;�I;��H;}H;��G;��E;��B; �=;�6;r�,;;��;�:�4�:�Ȋ:4�!:�/69x��D� �@tk�h���      "/�������x���X���/��� �����Xn칀:�9 �k:��:yo�:�B;&;l3;�<;O�A;�pE;ttG;}H;A�H;AI;�I;]I;I;�
I;I;n I;k�H;@�H;��H;��H;��H;��H;�H;��H;��H;��H;�H;��H;��H;��H;��H;=�H;h�H;n I;I;�
I;I;XI;�I;?I;>�H;}H;ttG;�pE;N�A;�<;l3;&;�B;yo�:��:$�k:�:�9Xn������� ���/���X���x����      ������q
����4�׻�+��®���;��lۺԖ �Q�9Ɋ:Y��:�;C!;��0;>;;ѓA;�pE;��G;�H;��H;�I;OI;pI;:I;�I;�I;�H;^�H;��H; �H;<�H;�H;�H;~�H;W�H;~�H;�H;�H;;�H;!�H;��H;]�H;�H;�I;�I;;I;pI;KI;�I;��H;ߎH;��G;�pE;ғA;>;;��0;F!;�;Y��:Ɋ:Q�9ؖ ��lۺ�;�®���+��2�׻����q
���      ����o8����>�k���O��3/�,B��׻����Q�@�P��0 ����>::5�:��;xb;��/;>;;O�A;��E;ԿG;	�H;�
I;} I;I;I;�I;�I;�I;��H;X�H;��H;��H;�H;/�H;��H;M�H;��H;/�H;�H;��H;��H;X�H;��H;�I;�I;�I;I;I;y I;�
I;	�H;ҿG;��E;O�A;@;;��/;xb;��;:5�:��>:0 ��P��S�@������׻,B��3/���O�>�k���p8��      >�� }�2�ݼ��˼d���,���}��G����<�һ����N��0/��:j׳:�;|b;£0;�<;��B;�IF;�H;:�H;�I;� I;/I;PI;r
I;�I;8 I;H�H;l�H;%�H;?�H;;�H;��H;U�H;��H;;�H;@�H;#�H;m�H;H�H;: I;�I;r
I;MI;2I;� I;�I;6�H;�H;�IF;��B;�<;ģ0;zb;�;j׳:�:0/�M������>�һ����G��}��,��d����˼2�ݼ}�      H�B�OR?��5���&��3��J��֮Ҽ#F����==� ?�.����/�Lnk�Ю�9b׳:��;B!;h3;�=;��C;1�F;'dH;�H;�I;%I;�I;:I;�I;�I;\�H;�H;��H;��H;\�H;��H;S�H;��H;[�H;��H;��H;�H;\�H;�I;�I;:I;�I;(I;�I;�H;"dH;2�F;��C;�=;h3;D!;��;b׳:Ю�9Lnk���/�.��?�>=���#F��֮Ҽ�J���3���&��5�PR?�      +��'W��뒐�%�����j�S`I���&����Fϼ�,���T[�i�cI��M;�<nk��:<5�:�;&;�6;�!@;H2E;�G;��H; I;!I;dI;%I;I;NI;� I;��H;�H;��H;z�H;��H;a�H;��H;z�H;��H;�H;��H;� I;PI;I;%I;cI;!I;I;��H;�G;H2E;�!@;�6;&;�;:5�:�:@nk�M;�cI��h��T[��,��Fϼ�����&�S`I���j�%���뒐�'W��      �J�����D��ͽ ���)�������L�'��'��
;���k����cI����/�0/���>:Y��:�B;r�,;��:;>�B;�xF;�<H;�H;I;�I;�I;XI;�I;�I;��H;��H;N�H;��H;��H;��H;��H;��H;N�H;��H;��H;�I;�I;UI;�I;�I;I;�H;�<H;�xF;?�B;��:;r�,;�B;_��:��>:0/���/�cI������k�
;��(��'����L����)�� ����ͽ�D����      T�:��*7���,�+���	�u�齅���#W����j�@�/��J���I���k�j�.��N��0 ��Ɋ:so�: ;hr3;.�>;<�D;{�G;Z�H;I;>!I;�I;�I;�
I;I;v I;��H;��H;��H;��H;y�H;��H;��H;��H;��H;v I;I;�
I;�I;�I;=!I;I;]�H;y�G;:�D;0�>;kr3; ;so�:
Ɋ:8 ��P��.��i��k��I���J��@�/���j�#W������t�齄�	�+���,��*7�      ^���p����4�l���M���,�Zl�T9ݽ�A���{� �5��J��
;���T[�?�����P���P�9��:��;1*;0�9;kkB;�F;�NH;��H;/ I;�I;�I;/I;!I;UI;w�H;��H;��H;��H;��H;��H;��H;��H;u�H;VI;"I;/I;�I;�I;- I;��H;�NH;݇F;ikB;0�9;2*;��;��:Q�9 P������?��T[�
;���J�� �5��{��A��T9ݽZl���,���M�4�l����p��      7m־S�Ѿ�>ľ����՗����{��I�+�����V���{�A�/�(���,��==�>�һR�@�ؖ �$�k:!�:b;��3;@j?;x2E;��G;|�H;CI;� I;�I;�I;4	I;I;��H;�H;��H;��H;m�H;��H;��H;�H;��H;I;4	I;�I;�I;� I;BI;|�H;��G;v2E;?j?;��3;b;�:$�k:Ԗ �S�@�>�һ==��,��(��A�/��{��V�����+��I���{�՗�������>ľS�Ѿ      E\�î�s5��z ��E۾ֳ�^��|�Z�N?#����A����j�'��Fϼ����������lۺh:�9�4�:_�;l�,;��;;D�C;�G;\�H;�I;�!I;�I;QI;:I;�I;TI;0�H;�H;��H;6�H;��H;�H;0�H;QI;�I;;I;QI;�I;�!I;�I;\�H;�G;C�C;��;;n�,;b�;�4�:X:�9�lۺ���������Fϼ'����j��A�����N?#�|�Z�^��ֳ��E۾�z �s5�î�      G�b��>]���M�Ŏ6�î�%���>ľ$q��|�Z�+�U9ݽ#W����L����#F���G��׻�;�`n��Ȋ:�i;&P$;�7;w�A;JF;ACH;��H;� I;zI;�I;+I;@I;�I;-�H;��H;��H;#�H;��H;��H;-�H;�I;@I;+I;�I;xI;� I;��H;@CH;JF;t�A;�7;(P$;�i;�Ȋ:`n��;��׻�G�#F�������L�#W��U9ݽ+�|�Z�$q���>ľ%��î�Ŏ6���M��>]�      p��򲗿���9�y�~�R���)�ov��>ľ^���I�Zl����������&�֮Ҽ�}�-B�®������4�!:+�:Dz;�3;ij?;�\E;��G;��H;}I;�I;�I;�I;�I;�I;0 I;��H;v�H;��H;v�H;��H;. I;�I;�I;�I;�I;�I;}I;��H;��G;�\E;fj?;�3;Dz;+�:0�!:����®��.B��}�֮Ҽ��&��������Zl��I�^���>ľov���)�~�R�9�y����򲗿      �˿�<ƿrL��B1����>]���)�%��ֳ���{���,�u��)��T`I��J���,���3/��+���� ��/69�4�:�;p.;..=;qaD;��G;r�H;�I;N!I;kI;`I;�	I;�I;� I;��H;&�H;v�H;'�H;��H;� I;�I;�	I;^I;hI;K!I;�I;q�H;��G;raD;(.=;p.;�;�4�:�/69�� ��+���3/��,���J��T`I�)��u�齦�,���{�ֳ�%����)��>]��B1��rL���<ƿ      ����>���X[忸˿�T���~�R�î��E۾՗����M���	� �����j��3�d����O�4�׻��/����`��:� 
;*;h;;�jC;�'G;��H;I;"I;I;�I;�
I;�I;�I;Y�H;��H;�H;��H;V�H;�I;�I;�
I;�I;�I;"I;I;��H;�'G;�jC;c;;*;� 
;f��:�����/�4�׻��O�d���3���j� �����	���M�՗���E۾î�~�R���T���˿X[�>���      O�7��v����˿B1��9�y�Ŏ6��z �����5�l�+��ͽ&�����&���˼?�k������X�@� ����:T�;&;�9;��B;�F;�}H;�	I;u"I;AI;�I;�I;�I;[I;��H;6�H;��H;6�H;��H;[I;�I;�I;�I;>I;r"I;�	I;�}H;�F;��B;�9; &;T�;���:H� ���X����@�k���˼��&�&����ͽ+�5�l������z �Ŏ6�9�y�B1���˿���v�7��      ��*��g&��#�v�X[�rL�������M�s5��>ľ����,��D�뒐��5�4�ݼ���q
��x�`tk� �b:_l�:#;՗7;��A;�F;�dH;�I;i"I;I;{I;QI;I;�I;3 I;��H;��H;��H;3 I;�I;I;QI;{I;I;f"I;�I;�dH;��F;��A;ϗ7;#;_l�:�b:htk��x��q
���4�ݼ�5�뒐��DὬ�,����>ľt5���M����rL��X[�v��#��g&�      ��8��4��g&�7��>����<ƿ򲗿�>]�î�S�Ѿ�p���*7����'W��PR?�}�p8�������p�����G:� �:�!;�6;&lA;�YF;�TH;{�H;)"I;�I;�I;�I;YI;I;s I;��H;"�H;��H;u I;I;WI;�I;�I;�I;'"I;{�H;�TH;�YF;&lA;�6;�!;� �:��G:r��������q8��}�PR?�'W�����*7��p��S�Ѿî��>]�򲗿�<ƿ>���7���g&��4�      ��!$������꿱�ſ�ޞ�(3s��2�@����� j���|HͽǸ����'�E<ͼq�n�e���1Q^�8-.�|��:�W;�S%;jo8;��A;hDF;�H;��H;��H;��H;V�H;N�H;V�H;��H; �H;��H;<�H;��H; �H;��H;U�H;O�H;V�H;��H;��H;��H;�H;gDF;��A;ho8;�S%;�W;���:<-.�1Q^�d���r�n�E<ͼ��'�Ǹ��|Hͽ�� j���@����2�(3s��ޞ���ſ������!$�      !$�������忉�����"cm�X�-�����Sh��Zde�$-�ڪɽ�v��*�$���ɼymj�8����X�d���ņ:x;K�%;9�8;uB;wRF;H;8�H;_�H;�H;y�H;R�H;H�H;��H;��H;��H;5�H;��H;��H;��H;G�H;T�H;y�H;�H;\�H;8�H;H;uRF;uB;6�8;P�%;x;�ņ:h���X�7���zmj���ɼ*�$��v��ڪɽ$-�Zde�Sh������X�-�"cm��������忞����      ��������� �ԿNw�����=�\�"����m��]0X�����;����w����������]� �黾F�`��ʒ:�;B�';ŏ9;)pB;�zF;�!H;��H;B�H;(�H;��H;X�H;N�H;��H;��H;��H; �H;��H;��H;��H;L�H;X�H;��H;&�H;?�H;��H;�!H;�zF;)pB;Ï9;D�';�;ʒ:h�깾F��黬�]����������w��;�����]0X�m�����"�=�\����Nw�� �Կ��𿞏�      ����� �Կp���ޞ�bF�j�C�/E�$�;�I���D���!"��j�c�~��֯���J��ѻ��)� }K�8��:$�
;�M*;z�:;�C;�F;�8H;`�H;��H;�H;��H;Q�H;L�H;��H;��H;��H;�H;��H;��H;��H;K�H;Q�H;��H;~�H;��H;`�H;�8H;�F;�C;w�:;�M*;$�
;:��: }K���)��ѻ��J��֯�~�j�c�!"�����D��I��$�;/E�j�C�bF��ޞ�p�� �Կ��      ��ſ���Nw���ޞ�����A�W�7�%�����jɰ��|x�i{+�ձ� ���J��  �϶��Y�1�&���+�#
9�:��;�-;��<;��C;�G;�TH;X�H;	�H;��H;��H;f�H;D�H;��H;��H;��H;�H;��H;��H;��H;B�H;g�H;��H;��H;�H;X�H;�TH;�G;��C;��<;�-;��;�:#
9+�$���Y�1�϶���  ��J� ��ձ�i{+��|x�jɰ�����7�%�A�W������ޞ�Nw�����      �ޞ�������bF�A�W�Y�-����BKɾ�G����O����ƽȸ��ф-���ۼㄼ44�ǐ��ζ��]:��:�;��1;�c>;x�D;�\G;MsH;��H;u�H;n�H;1�H;��H;:�H;}�H;��H;��H;��H;��H;��H;}�H;:�H;��H;1�H;k�H;q�H;��H;KsH;�\G;w�D;�c>;��1;�;��:�]:�ζ�ǐ�44�ㄼ��ۼф-�ȸ��ƽ�����O��G��BKɾ���Y�-�A�W�bF�������      (3s�!cm�<�\�j�C�7�%�����TҾm�� j��C(����aP����[�~������Y�4��WX��<���k:_��:� ;�5;NR@;nuE;�G;<�H;R�H;��H;�H;T�H;~�H;6�H;u�H;��H;j�H;��H;j�H;��H;u�H;7�H;�H;T�H;�H;��H;R�H;;�H;�G;kuE;LR@;�5;� ;a��:��k:�<�TX�4����Y����~���[�aP����콭C(� j�m���TҾ���7�%�j�C�<�\�!cm�      �2�X�-�"�.E�����BKɾm����s�:�5���y㻽�v��z0��;��+���*����!6��;S��M�:f�	;��(;$�9;�/B;�DF;^H;۫H;��H;��H;��H;��H;��H;#�H;E�H;R�H;N�H;m�H;N�H;S�H;E�H;"�H;��H;��H;��H;��H;��H;ثH;]H;|DF;�/B;&�9;��(;g�	;�M�:@;S�6�����*��+���;�z0��v��y㻽��:�5���s�m��BKɾ����.E�"�X�-�      @����������$�;jɰ��G�� j�:�5��	�Ҫɽ[����J�u���沼��]�����	x�,	���n:��:�v;��/;�-=;��C;O�F;*IH;��H;0�H;��H;.�H;��H;��H;��H;�H;!�H;)�H;9�H;)�H;!�H;�H;��H;��H;��H;-�H;��H;0�H;��H;*IH;M�F;��C;�-=;��/;�v;ݤ�:�n:*	���	x������]��沼u���J�[���Ҫɽ�	�:�5� j��G��jɰ�$�;��徹���      ��Sh��m���I���|x���O��C(���Ҫɽ����VDX�K��)<ͼ
ㄼ�X!��s���W�PtK�V��:�y;�#;I6;@R@;�PE;��G;��H;��H;=�H;��H;��H;��H;��H;��H;��H;��H;��H;��H;��H;��H;��H;��H;��H;��H;��H;��H;=�H;��H;��H;��G;�PE;>R@;I6;�#;�y;V��:@tK��W��s���X!�
ㄼ)<ͼK��VDX�����Ҫɽ���C(���O��|x��I��m��Sh��       j�Yde�\0X��D�i{+�������y㻽\���VDX������ۼ̾����;�B>ۻX���y�H?":��:��;�-;��;;�B;�zF;�H;��H;��H;2�H;��H;�H;��H;��H;��H;��H;��H;��H;��H;��H;��H;��H;��H;��H;��H;�H;��H;2�H;��H;��H;�H;�zF;��B;��;;�-;��;��:T?":��y�X�B>ۻ��;�̾����ۼ���VDX�[���y㻽��콄��i{+��D�\0X�Yde�      ��$-������ձ�ƽaP���v���J�J����ۼ��c�J�����~+��\rѺ*
9N�:��;� $;�5;�?;��D;l\G;fH; �H;��H;��H;��H;.�H;�H;i�H;��H;r�H;k�H;x�H;Q�H;x�H;m�H;r�H;��H;k�H;�H;/�H;��H;��H;��H;��H;fH;k\G;��D;�?;�5;� $;��;N�: *
9^rѺ~+������c�J�����ۼJ���J��v��aP��ƽձ轅����$-�      |Hͽڪɽ�;�� "�� ��ȸ����[�z0�u��*<ͼ̾��d�J�����j��f*��,��:lb�:^�;��/;�L<;C;9mF;��G;�H;�H; �H; �H;V�H;f�H;�H;<�H;H�H;5�H;/�H;�H;�H;�H;/�H;3�H;G�H;=�H;�H;f�H;T�H; �H;�H;�H;�H;��G;6mF;C;�L<;��/;^�;rb�:*��:��f*��j�����d�J�̾��)<ͼu��z0���[�ȸ�� �� "���;��ڪɽ      Ǹ���v����w�i�c��J�ф-�~��;缈沼
ㄼ��;������j���5����d?Q:���:pi;�M*;��8;��@;�PE;�uG;LiH;��H;��H;%�H;7�H;��H;��H;��H;�H;��H;��H;��H;��H;��H;��H;��H;��H;��H;�H;��H;��H;��H;9�H;"�H;��H;��H;IiH;�uG;�PE;��@;��8;�M*;ri;}��:d?Q:��깑5��j��������;�
ㄼ�沼�;�~�ф-��J�i�c���w��v��      ��'�*�$����~��  ���ۼ����+����]��X!�B>ۻ+��g*����8�>:��: �;B�%;��5;��>;�(D;�F;�!H;D�H;f�H;�H;��H;��H;�H;��H;��H;��H;��H;��H;��H;i�H;��H;i�H;��H;��H;��H;��H;��H;��H; �H;��H;��H;�H;d�H;@�H;�!H;�F;�(D;��>;��5;E�%;�;��:8�>:���g*�+��B>ۻ�X!���]��+�������ۼ�  �~����*�$�      D<ͼ��ɼ�����֯�϶��ㄼ��Y��*�����s��X�\rѺ�\?Q:��:��
;]�#;q�3;�c=;$C;7DF;�G;$�H;��H;%�H;O�H;�H;p�H;=�H;�H;��H;{�H;S�H;m�H;'�H;�H;$�H;�H;'�H;m�H;Q�H;}�H;��H;�H;9�H;p�H;�H;P�H;$�H;��H; �H;�G;3DF;$C;�c=;s�3;[�#;��
;��:h?Q:�\rѺX��s������*���Y�ㄼ϶���֯�������ɼ      q�n�vmj���]���J�Z�1�34�0������	x��W���y� *
9*��:}��: �;Y�#;d�2;�<;~pB;:�E;čG;�eH;�H;K�H;��H;�H;��H;��H;W�H;e�H;T�H;+�H;�H;��H;��H;��H;��H;��H;��H;��H;�H;-�H;T�H;c�H;T�H;��H;��H;�H;��H;G�H;�H;�eH;��G;;�E;|pB;�<;f�2;Y�#; �;}��:*��:*
9��y��W��	x����0��24�Y�1���J���]�xmj�      f���7������ѻ&���ǐ�WX�"6�*	��ptK�T?":N�:nb�:ni;C�%;q�3;�<;U0B;��E;�\G;�HH;Z�H;��H;v�H;�H;R�H;X�H;��H;4�H;6�H; �H;��H;��H;~�H;p�H;o�H;L�H;o�H;p�H;}�H;��H;��H; �H;5�H;1�H;��H;V�H;S�H;�H;q�H;��H;Z�H;�HH;�\G;��E;W0B;�<;p�3;C�%;pi;nb�:N�:X?":@tK�$	��$6�WX�ǐ�#����ѻ��<���      &Q^��X��F���)�+��ζ���<� <S��n:T��:���:��;^�;�M*;��5;�c=;|pB;��E;�JG;h8H;��H;��H;*�H;E�H;��H;��H;��H;�H;�H;��H;��H;��H;u�H;"�H;�H;�H;��H;�H;�H; �H;s�H;��H;��H;��H;�H;�H;��H;��H;��H;A�H;'�H;��H;�H;k8H;�JG;��E;|pB;�c=;��5;�M*;^�;��;���:T��:�n: <S���<��ζ�
+���)��F��X�      ,-.�$��H���|K��"
9�]:��k:�M�:ۤ�:�y;��;� $;��/;��8;��>;$C;9�E;�\G;f8H;ۥH;�H;:�H;��H;Q�H;��H;p�H;��H;��H;��H;��H;Z�H;1�H;�H;��H;��H;��H;��H;��H;��H;��H;�H;3�H;Z�H;��H;��H;��H;��H;p�H;��H;K�H;��H;;�H;�H;ݥH;f8H;�\G;:�E;$C;��>;��8;��/;� $;��;�y;ۤ�:�M�:��k:�]:�#
9�|K�H��H��      ���:Ɔ:ʒ:*��:�:!��:a��:d�	;�v;�#;�-;�5;�L<;��@;�(D;4DF;čG;�HH;��H;�H;��H;g�H;��H;|�H;>�H;��H;��H;��H;��H;C�H;&�H;��H;��H;��H;R�H;E�H;E�H;E�H;R�H;��H;��H;��H;&�H;A�H;~�H;��H;��H;��H;>�H;x�H;��H;g�H;��H; �H;��H;�HH;ÍG;4DF;�(D;��@;�L<;�5;�-;�#;�v;f�	;a��:'��:�:.��:
ʒ:�ņ:      �W;�x;�;�
;��;�;� ;��(;��/;I6;��;;	�?;C;�PE;#�F;�G;�eH;\�H;��H;=�H;g�H;��H;N�H;�H;��H;��H;��H;��H;�H;��H;��H;j�H;A�H;/�H;��H;��H;��H;��H;��H;/�H;>�H;j�H;��H;��H;�H;��H;��H;��H;��H;�H;L�H;��H;e�H;>�H;��H;]�H;�eH;�G;#�F;�PE;C;	�?;��;;I6;��/;��(;� ;�;̅;�
;�;�x;      �S%;O�%;C�';�M*;�-;��1;�5;$�9;�-=;@R@;�B;��D;9mF;�uG;�!H;#�H;
�H;��H;,�H;��H;��H;O�H;#�H;��H;��H;��H;]�H;�H;��H;��H;I�H;�H;��H;��H;��H;��H;{�H;��H;��H;��H;��H;�H;I�H;��H;��H;�H;X�H;��H;��H;��H;%�H;P�H;��H;��H;,�H;��H;
�H;!�H;�!H;�uG;9mF;��D;�B;>R@;�-=;$�9;�5;��1;�-;�M*;F�';B�%;      �o8;I�8;̏9;|�:;��<;�c>;XR@;�/B;��C;�PE;�zF;o\G;��G;OiH;F�H;��H;J�H;w�H;E�H;O�H;x�H;�H;��H;��H;��H;o�H;�H;��H;��H;9�H;��H;��H;��H;V�H;Q�H;D�H;!�H;D�H;R�H;U�H;��H;��H;��H;6�H;��H;��H;�H;o�H;��H;��H;��H;�H;u�H;O�H;E�H;x�H;J�H;��H;F�H;OiH;��G;n\G;�zF;�PE;��C;�/B;VR@;�c>;��<;|�:;Ϗ9;;�8;      ��A;�B;pB;�C;��C;z�D;nuE;DF;Q�F;��G;�H;fH;�H;��H;j�H;*�H;��H;�H;��H;��H;A�H;��H;��H;��H;O�H;��H;��H;��H;/�H;��H;��H;m�H;:�H;�H;��H;��H;��H;��H;��H;�H;9�H;n�H;��H;��H;/�H;��H;��H;��H;P�H;��H;��H;��H;A�H;��H;��H;�H;��H;(�H;j�H;��H;�H;fH;�H;��G;O�F;DF;nuE;z�D;��C;�C;pB;�B;      sDF;�RF;�zF;�F;�G;�\G;�G;XH;,IH;��H;��H;�H;�H;��H;�H;O�H;�H;P�H;��H;o�H;��H;��H;��H;n�H;��H;��H;��H;(�H;��H;��H;H�H;	�H;��H;��H;��H;��H;��H;��H;��H;��H;��H;�H;J�H;��H;��H;)�H;��H;��H;��H;l�H;��H;��H;��H;p�H;��H;P�H;�H;M�H;�H;��H;�H;�H;��H;��H;,IH;XH;�G;�\G;�G;�F;�zF;xRF;      �H;H;�!H;�8H;�TH;RsH;C�H;ޫH;��H;��H;��H;��H;�H;&�H;��H;�H;��H;V�H;��H;��H;��H;��H;Z�H;�H;��H;��H;�H;��H;x�H;H�H;��H;��H;��H;w�H;^�H;9�H;M�H;9�H;\�H;v�H;��H;��H;�H;G�H;x�H;��H;�H;��H;��H;�H;X�H;��H;��H;��H;��H;W�H;��H;�H;��H;&�H;�H;��H;��H;��H;��H;ܫH;E�H;OsH;�TH;�8H;�!H;H;      ��H;;�H;��H;]�H;[�H;��H;Y�H;��H;8�H;E�H;9�H;��H;"�H;=�H;��H;p�H;��H;��H; �H;��H;��H;��H;�H;��H;��H;)�H;��H;��H;7�H;��H;��H;z�H;T�H;!�H;�H;�H;�H;�H;�H;!�H;Q�H;z�H;��H;��H;6�H;��H;��H;)�H;��H;��H;�H;��H;��H;��H; �H;��H;��H;p�H;��H;;�H;"�H;��H;7�H;C�H;8�H;��H;[�H;��H;e�H;]�H;��H;H�H;      �H;d�H;>�H;��H;	�H;w�H;��H;��H;��H;�H;��H;��H;W�H;��H;�H;?�H;X�H;1�H;�H;��H;��H;�H;��H;��H;(�H;��H;t�H;7�H;��H;��H;l�H;5�H; �H;��H;��H;��H;��H;��H;��H;��H;��H;6�H;l�H;��H;��H;7�H;u�H;��H;*�H;��H;��H;�H;��H;��H;�H;2�H;W�H;=�H;�H;��H;W�H;��H;��H;��H;��H;��H;��H;u�H;�H;��H;A�H;[�H;      �H;�H;2�H;��H;	�H;u�H;�H;��H;:�H;��H;�H;<�H;o�H;��H;��H;��H;h�H;2�H;��H;��H;B�H;��H;��H;9�H;��H;��H;D�H;��H;��H;c�H;2�H;��H;��H;��H;��H;��H;w�H;��H;��H;��H;��H;��H;2�H;b�H;��H;��H;A�H;��H;��H;9�H;��H;��H;A�H;��H;��H;4�H;f�H;��H;��H;��H;o�H;<�H;�H;��H;;�H;��H;�H;u�H;�H;��H;.�H;�H;      [�H;��H;��H;��H;�H;5�H;b�H;��H;��H;��H;�H;�H;�H;�H;��H;��H;Z�H;�H;��H;`�H;*�H;��H;H�H;��H;��H;J�H;��H;��H;j�H;5�H;��H;��H;��H;y�H;V�H;`�H;^�H;`�H;V�H;y�H;��H;��H;��H;4�H;l�H;��H;��H;H�H;��H;��H;G�H;��H;'�H;`�H;��H;�H;Z�H;��H;��H;�H;�H;�H;�H;��H;��H;��H;b�H;6�H;�H;��H;��H;��H;      [�H;d�H;_�H;\�H;p�H;��H;��H;��H;��H;��H;��H;t�H;A�H;�H;��H;��H;5�H;��H;��H;:�H;��H;n�H;�H;��H;j�H;	�H;��H;{�H;4�H;��H;��H;��H;z�H;F�H;1�H;0�H;3�H;0�H;1�H;F�H;w�H;��H;��H;��H;5�H;{�H;��H;�H;k�H;��H;�H;n�H;��H;:�H;��H;��H;4�H;��H;��H;�H;C�H;t�H;��H;��H;��H;��H;��H;��H;n�H;\�H;_�H;`�H;      ]�H;^�H;Y�H;Z�H;U�H;=�H;=�H;/�H;�H;��H;��H;��H;N�H;��H;��H;X�H;�H;��H;w�H;�H;��H;@�H;��H;��H;5�H;��H;��H;U�H;�H;��H;��H;|�H;4�H;)�H;)�H;�H;��H;�H;)�H;)�H;1�H;~�H;��H;��H;�H;W�H;��H;��H;6�H;��H;��H;@�H;��H;�H;w�H;��H;�H;X�H;��H;��H;M�H;��H;��H;��H;�H;/�H;=�H;@�H;N�H;Z�H;Y�H;W�H;      ��H;��H;��H;��H;��H;|�H;�H;R�H;"�H;�H;��H;{�H;9�H;��H;��H;t�H;��H;~�H;%�H;��H;��H;/�H;��H;[�H;�H;��H;s�H; �H;��H;��H;w�H;H�H;%�H;�H;�H;��H;��H;��H;�H;�H;#�H;J�H;w�H;��H;��H; �H;s�H;��H;�H;Y�H;��H;/�H;��H;��H;%�H;��H;��H;t�H;��H;��H;9�H;{�H;��H;�H;#�H;R�H;�H;�H;��H;��H;��H;��H;      �H;�H;��H;��H;��H;��H;��H;c�H;-�H;��H;��H;{�H;9�H;��H;��H;1�H;��H;n�H;�H;��H;Y�H;��H;��H;T�H;��H;��H;X�H;�H;��H;��H;T�H;5�H;'�H;�H;��H;��H;��H;��H;��H;�H;&�H;8�H;T�H;��H;��H;�H;W�H;��H;��H;R�H;��H;��H;V�H;��H;�H;o�H;��H;1�H;��H;��H;9�H;{�H;��H;��H;-�H;a�H;��H;��H;��H;��H;��H;�H;      ��H;��H;��H;��H;��H;��H;v�H;^�H;9�H;��H;��H;��H;%�H;��H;o�H;�H;��H;k�H;�H;��H;I�H;��H;��H;H�H;��H;��H;6�H;�H;��H;��H;`�H;4�H;�H;��H;��H;��H;��H;��H;��H;��H;�H;8�H;`�H;��H;��H;�H;5�H;��H;��H;F�H;��H;��H;H�H;��H;�H;l�H;��H;�H;p�H;��H;%�H;��H;��H;��H;9�H;]�H;v�H;��H;��H;��H;��H;��H;      A�H;F�H;7�H;�H;�H;��H;��H;y�H;B�H;��H;��H;\�H;�H;��H;��H;-�H;��H;E�H;��H;��H;E�H;��H;u�H;"�H;��H;��H;I�H;	�H;��H;z�H;a�H;:�H;��H;��H;��H;��H;��H;��H;��H;��H;��H;;�H;a�H;z�H;��H;	�H;G�H;��H;��H; �H;w�H;��H;E�H;��H;��H;F�H;��H;-�H;��H;��H;�H;]�H;��H;��H;E�H;x�H;��H;��H;�H;�H;5�H;>�H;      ��H;��H;��H;��H;��H;��H;v�H;^�H;9�H;��H;��H;��H;%�H;��H;p�H;�H;��H;k�H;�H;��H;K�H;��H;��H;G�H;��H;��H;6�H;�H;��H;��H;`�H;5�H;�H;��H;��H;��H;��H;��H;��H;��H;�H;7�H;`�H;��H;��H;�H;5�H;��H;��H;F�H;��H;��H;H�H;��H;�H;l�H;��H;�H;o�H;��H;%�H;��H;��H;��H;9�H;]�H;v�H;��H;��H;��H;��H;��H;      �H;�H;��H;��H;��H;��H;��H;c�H;-�H;��H;��H;{�H;9�H;��H;��H;1�H;��H;n�H;�H;��H;Z�H;��H;��H;T�H;��H;��H;X�H;�H;��H;��H;T�H;5�H;'�H;�H;��H;��H;��H;��H;��H;�H;&�H;:�H;T�H;��H;��H;�H;W�H;��H;��H;Q�H;��H;��H;V�H;��H;�H;o�H;��H;1�H;��H;��H;9�H;{�H;��H;��H;-�H;a�H;��H;��H;��H;��H;��H;�H;      ��H;��H;��H;��H;��H;{�H;�H;R�H;"�H;�H;��H;{�H;9�H;��H;��H;t�H;��H;~�H;%�H;��H;��H;/�H;��H;[�H;�H;��H;s�H; �H;��H;��H;w�H;H�H;%�H;�H;�H;��H;��H;��H;�H;�H;#�H;J�H;w�H;��H;��H; �H;t�H;��H;�H;Y�H;��H;/�H;��H;��H;%�H;��H;��H;t�H;��H;��H;9�H;{�H;��H;�H;#�H;R�H;�H;��H;��H;��H;��H;��H;      `�H;]�H;Z�H;]�H;S�H;=�H;>�H;-�H;�H;��H;��H;��H;M�H;��H;��H;X�H;�H;��H;w�H;�H;��H;@�H;��H;��H;6�H;��H;��H;W�H;�H;��H;��H;|�H;3�H;'�H;)�H;�H;��H;�H;)�H;'�H;1�H;��H;��H;��H;�H;U�H;��H;��H;5�H;��H;��H;@�H;��H;�H;w�H;��H;�H;X�H;��H;��H;M�H;��H;��H;��H;�H;,�H;>�H;@�H;L�H;]�H;V�H;\�H;      [�H;d�H;`�H;[�H;p�H;��H;��H;��H;��H;��H;��H;t�H;A�H;�H;��H;��H;4�H;��H;��H;;�H;��H;n�H;�H;��H;k�H;	�H;��H;{�H;2�H;��H;��H;��H;y�H;F�H;1�H;0�H;3�H;0�H;1�H;F�H;w�H;��H;��H;��H;5�H;{�H;��H;�H;j�H;��H;�H;n�H;��H;:�H;��H;��H;4�H;��H;��H;�H;A�H;t�H;��H;��H;��H;��H;��H;��H;n�H;[�H;_�H;`�H;      [�H;��H;��H;��H;�H;4�H;b�H;��H;��H;��H;�H;�H;�H;�H;��H;��H;X�H;�H;��H;`�H;,�H;��H;H�H;��H;��H;J�H;��H;��H;j�H;5�H;��H;��H;��H;y�H;V�H;`�H;^�H;`�H;V�H;y�H;��H;��H;��H;4�H;l�H;��H;��H;H�H;��H;��H;E�H;��H;'�H;`�H;��H;�H;Z�H;��H;��H;�H;�H;�H;�H;��H;��H;��H;b�H;6�H;�H;��H;��H;��H;      �H;�H;1�H;��H;�H;p�H;�H;��H;;�H;��H;�H;<�H;o�H;��H;��H;��H;h�H;2�H;��H;��H;E�H;��H;��H;9�H;��H;��H;D�H;��H;��H;c�H;2�H;��H;��H;��H;��H;��H;w�H;��H;��H;��H;��H;��H;2�H;b�H;��H;��H;A�H;��H;��H;9�H;��H;��H;A�H;��H;��H;4�H;f�H;��H;��H;��H;o�H;<�H;�H;��H;<�H;��H;�H;t�H;�H;��H;1�H;�H;      
�H;`�H;D�H;��H;�H;q�H;��H;��H;��H;��H;��H;��H;W�H;��H;�H;=�H;X�H;1�H;�H;��H;��H;�H;��H;��H;*�H;��H;t�H;7�H;��H;��H;l�H;4�H;��H;��H;��H;��H;��H;��H;��H;��H;��H;6�H;l�H;��H;��H;7�H;u�H;��H;(�H;��H;��H;�H;��H;��H;�H;2�H;X�H;@�H;�H;��H;W�H;��H;��H;�H;��H;��H;��H;u�H;�H;��H;F�H;`�H;      ��H;<�H;��H;]�H;[�H;��H;[�H;��H;7�H;C�H;9�H;��H;"�H;;�H;��H;p�H;��H;��H; �H;��H;��H;��H;�H;��H;��H;)�H;��H;��H;7�H;��H;��H;z�H;S�H; �H;�H;�H;�H;�H;�H;!�H;S�H;{�H;��H;��H;7�H;��H;��H;)�H;��H;��H;�H;��H;��H;��H; �H;��H;��H;r�H;��H;:�H;"�H;��H;7�H;E�H;;�H;��H;Y�H;��H;g�H;]�H;��H;E�H;      �H;H;�!H;�8H;�TH;NsH;C�H;ޫH;��H;��H;��H;��H;�H;&�H;��H;�H;��H;V�H;��H;��H;��H;��H;Z�H;�H;��H;��H;�H;��H;x�H;H�H;�H;��H;��H;v�H;\�H;9�H;M�H;8�H;^�H;v�H;��H;��H;��H;G�H;w�H;��H;�H;��H;��H;�H;X�H;��H;��H;��H;��H;W�H;��H;�H;��H;&�H;�H;��H;��H;��H;��H;ޫH;B�H;MsH;�TH;�8H;�!H;H;      yDF;�RF;�zF;�F;�G;�\G;�G;[H;*IH;��H;��H;�H;�H;��H;�H;O�H;�H;O�H;��H;p�H;��H;��H;��H;n�H;��H;��H;��H;)�H;��H;��H;J�H;	�H;��H;��H;��H;��H;��H;��H;��H;��H;��H;�H;H�H;��H;��H;(�H;��H;��H;��H;l�H;��H;��H;��H;o�H;��H;R�H;�H;O�H;�H;��H;�H;�H;��H;��H;*IH;ZH;�G;�\G;�G;�F;�zF;tRF;      ��A;�B;pB;�C;��C;z�D;nuE;DF;O�F;��G;�H;fH;�H;��H;j�H;*�H;��H;�H;��H;��H;C�H;��H;��H;��H;P�H;��H;��H;��H;/�H;��H;��H;m�H;9�H;�H;��H;��H;��H;��H;��H;�H;9�H;p�H;��H;��H;,�H;��H;��H;��H;O�H;��H;��H;��H;?�H;��H;��H;�H;��H;*�H;j�H;��H;�H;fH;�H;��G;Q�F;�DF;nuE;z�D;��C;�C;pB;�B;      �o8;F�8;ԏ9;y�:;��<; d>;RR@;�/B;��C;�PE;�zF;n\G;��G;OiH;F�H;��H;J�H;v�H;E�H;O�H;y�H;�H;��H;��H;��H;n�H;�H;��H;��H;9�H;��H;��H;��H;T�H;O�H;F�H;!�H;D�H;R�H;V�H;��H;��H;��H;6�H;��H;��H;�H;o�H;��H;��H;��H;�H;u�H;O�H;E�H;x�H;I�H;��H;F�H;OiH;��G;o\G;�zF;�PE;��C;�/B;RR@;d>;��<;w�:;׏9;9�8;      �S%;^�%;R�';�M*;�-;��1;�5;$�9;�-=;>R@;�B;��D;8mF;�uG;�!H;#�H;
�H;��H;,�H;��H;��H;P�H;&�H;��H;��H;��H;]�H;�H;��H;��H;I�H;�H;��H;��H;��H;��H;{�H;��H;��H;��H;��H;�H;I�H;��H;��H;�H;Z�H;��H;��H;��H;"�H;O�H;��H;��H;,�H;��H;�H;#�H;�!H;�uG;8mF;��D;�B;=R@;�-=;&�9;�5;��1;�-;�M*;J�';L�%;      �W;�x;�;�
;��;�;� ;��(;��/;I6;��;;	�?;C;�PE;"�F;�G;�eH;\�H;��H;=�H;g�H;��H;N�H;�H;��H;��H;��H;��H;�H;��H;��H;j�H;@�H;/�H;��H;��H;��H;��H;��H;/�H;@�H;j�H;��H;��H;�H;��H;��H;��H;��H;�H;K�H;��H;e�H;>�H;��H;]�H;�eH;�G;$�F;�PE;C;�?;��;;I6;��/;��(;� ;�;Ѕ;�
;�;�x;      ���:Ɔ:ʒ:.��:�:��:g��:i�	;�v;�#;�-;�5;�L<;��@;�(D;4DF;čG;�HH;��H; �H;��H;g�H;��H;|�H;>�H;��H;��H;��H;��H;C�H;&�H;��H;��H;��H;R�H;E�H;E�H;E�H;R�H;��H;��H;��H;&�H;A�H;~�H;��H;��H;��H;>�H;x�H;��H;g�H;��H;�H;��H;�HH;ÍG;4DF;�(D;��@;�L<;�5;�-;�#;�v;g�	;g��:!��:
�:,��:ʒ:�ņ:      4-.� ��(�� }K�P#
9�]:��k:�M�:ݤ�:�y;��;� $;��/;��8;��>;$C;9�E;�\G;f8H;ۥH;�H;;�H;��H;Q�H;��H;p�H;��H;��H;��H;��H;Z�H;1�H;�H;��H;��H;��H;��H;��H;��H;��H;�H;3�H;Z�H;��H;��H;��H;��H;p�H;��H;K�H;��H;:�H;�H;ݥH;f8H;�\G;:�E;$C;��>;��8;��/;� $;��;�y;��:�M�:��k:�]:�#
9 }K�0��T��      &Q^��X��F���)�+��ζ���<��;S��n:T��:���:��;^�;�M*;��5;�c=;~pB;��E;�JG;i8H;��H;��H;,�H;E�H;��H;��H;��H;�H;�H;��H;��H;��H;u�H; �H;�H;�H;��H;�H;�H;"�H;s�H;��H;��H;��H;�H;�H;��H;��H;��H;?�H;&�H;��H;�H;k8H;�JG;��E;|pB;�c=;��5;�M*;^�;��;���:T��:�n:�;S���<��ζ�	+���)��F��X�      d���8������ѻ&���ǐ�UX�"6�&	��@tK�T?":N�:nb�:ni;C�%;p�3;�<;U0B;��E;�\G;�HH;Z�H;��H;v�H;�H;P�H;X�H;��H;4�H;6�H; �H;��H;��H;}�H;p�H;o�H;L�H;o�H;p�H;~�H;��H;��H; �H;5�H;1�H;��H;V�H;S�H;�H;p�H;��H;Z�H;�HH;�\G;��E;W0B;�<;q�3;C�%;ni;nb�:N�:T?":ptK�$	��"6�UX�ǐ�"����ѻ��<���      q�n�vmj���]���J�Y�1�34�/������	x��W���y� *
9*��:}��: �;Y�#;f�2;�<;|pB;;�E;ÍG;�eH;
�H;K�H;��H;�H;��H;��H;U�H;e�H;T�H;-�H;�H;��H;��H;��H;��H;��H;��H;��H;�H;-�H;T�H;c�H;T�H;��H;��H;�H;��H;G�H;�H;�eH;ÍG;=�E;~pB;�<;d�2;Y�#; �;}��:*��: *
9��y��W��	x����0��24�X�1���J���]�ymj�      D<ͼ��ɼ�����֯�϶��ㄼ��Y��*�����s��X�\rѺ�d?Q:��:��
;]�#;q�3;�c=;$C;4DF;�G;#�H;��H;$�H;O�H;�H;p�H;=�H;~�H;��H;{�H;S�H;m�H;'�H;�H;$�H;�H;'�H;m�H;Q�H;}�H;��H;�H;9�H;p�H;�H;P�H;%�H;��H; �H;�G;4DF;$C;�c=;s�3;[�#;��
;��:\?Q:�\rѺX��s������*���Y�ㄼ϶���֯�������ɼ      ��'�*�$����~��  ���ۼ����+����]��X!�B>ۻ+��g*����8�>:��: �;B�%;��5;��>;�(D;�F;�!H;D�H;d�H;�H;��H;��H;�H;��H;��H;��H;��H;��H;��H;i�H;��H;i�H;��H;��H;��H;��H;��H;��H; �H;��H;��H;�H;f�H;@�H;�!H;�F;�(D;��>;��5;E�%;�;��:8�>:���g*�+��B>ۻ�X!���]��+�������ۼ�  �~����*�$�      Ǹ���v����w�i�c��J�ф-�~��;缈沼
ㄼ��;������j���5����d?Q:���:pi;�M*;��8;��@;�PE;�uG;LiH;��H;��H;%�H;9�H;��H;��H;��H;�H;��H;��H;��H;��H;��H;��H;��H;��H;��H;�H;��H;��H;��H;7�H;#�H;��H;��H;IiH;�uG;�PE;��@;��8;�M*;ri;}��:d?Q:��깑5��j��������;�
ㄼ�沼�;�~�ф-��J�i�c���w��v��      |Hͽڪɽ�;�� "�� ��ȸ����[�z0�u��)<ͼ̾��d�J�����j��f*��*��:nb�:^�;��/;�L<;C;;mF;��G;�H;�H; �H; �H;T�H;f�H;�H;<�H;G�H;3�H;/�H;�H;�H;�H;/�H;5�H;G�H;<�H;�H;f�H;S�H; �H;�H;�H;�H;��G;5mF;C;�L<;��/;^�;rb�:*��:�d*��j�����d�J�̾��)<ͼu��z0���[�ȸ�� �� "���;��ڪɽ      ��$-������ձ�ƽaP���v���J�J����ۼ��c�J�����~+��^rѺ*
9N�:��;� $;�5;�?;��D;n\G;fH;��H;��H;��H;��H;/�H;�H;i�H;��H;t�H;m�H;z�H;Q�H;z�H;k�H;r�H;��H;j�H;�H;/�H;��H;��H;��H;��H;fH;i\G;��D;�?;�5;� $;��;N�: *
9^rѺ~+������c�J�����ۼJ���J��v��aP��ƽձ轅����$-�       j�Yde�\0X��D�i{+�������y㻽\���VDX������ۼ̾����;�B>ۻX���y�P?":��:��;�-;��;;�B;�zF;�H;��H;��H;2�H;��H;�H;��H;��H;��H;��H;��H;��H;��H;��H;��H;��H;��H;��H;��H;�H;��H;2�H;��H;��H;�H;�zF;��B;��;;�-;��;��:T?":��y�X�A>ۻ��;�̾����ۼ���VDX�\���y㻽��콄��i{+��D�]0X�Yde�      ��Sh��m���I���|x���O��C(���Ҫɽ����VDX�K��)<ͼ
ㄼ�X!��s���W�PtK�V��:�y;�#;I6;@R@;�PE;��G;��H;��H;=�H;��H;��H;��H;��H;��H;��H;��H;��H;��H;��H;��H;��H;��H;��H;��H;��H;��H;=�H;��H;��H;��G;�PE;>R@;I6;�#;�y;V��:@tK��W��s���X!�
ㄼ)<ͼK��VDX�����Ҫɽ���C(���O��|x��I��m��Sh��      @����������$�;jɰ��G�� j�:�5��	�Ҫɽ[����J�u���沼��]�����	x�,	���n:��:�v;��/;�-=;��C;M�F;*IH;��H;0�H;��H;-�H;��H;��H;��H;�H;!�H;)�H;9�H;)�H;!�H;�H;��H;��H;��H;-�H;��H;0�H;��H;*IH;O�F;��C;�-=;��/;�v;ݤ�:�n:*	���	x������]��沼u���J�\���Ҫɽ�	�:�5� j��G��jɰ�$�;��徹���      �2�X�-�"�.E�����BKɾm����s�:�5���y㻽�v��z0��;��+���*����!6�@;S��M�:d�	;��(;&�9;�/B;|DF;]H;٫H;��H;��H;��H;��H;��H;#�H;G�H;U�H;N�H;m�H;P�H;R�H;G�H;"�H;��H;��H;��H;��H;��H;٫H;[H;�DF;�/B;$�9;��(;g�	;�M�:�;S�6�����*��+���;�z0��v��y㻽��:�5���s�m��BKɾ����.E�"�X�-�      (3s�!cm�<�\�j�C�7�%�����TҾm�� j��C(����aP����[�~������Y�2��UX��<���k:[��:� ;�5;OR@;kuE;�G;<�H;R�H;��H;�H;T�H;~�H;9�H;v�H;��H;j�H;��H;j�H;��H;u�H;4�H;~�H;T�H;�H;��H;R�H;;�H;�G;nuE;LR@;	�5;� ;a��:��k:�<�TX�4����Y����~���[�aP����콭C(� j�m���TҾ���7�%�j�C�<�\�!cm�      �ޞ�������bF�A�W�Y�-����BKɾ�G����O����ƽȸ��ф-���ۼㄼ34�ǐ��ζ��]:��:�;��1;�c>;w�D;�\G;MsH;��H;u�H;n�H;1�H;��H;;�H;}�H;��H;��H;��H;��H;��H;}�H;9�H;��H;1�H;k�H;q�H;��H;KsH;�\G;x�D;�c>;��1;�;��:�]:�ζ�ǐ�44�ㄼ��ۼф-�ȸ��ƽ�����O��G��BKɾ���Y�-�A�W�bF�������      ��ſ���Nw���ޞ�����A�W�7�%�����jɰ��|x�i{+�ձ� ���J��  �϶��Y�1�%���+�#
9�:��;�-;��<;��C;�G;�TH;X�H;	�H;��H;��H;f�H;D�H;��H;��H;��H;�H;��H;��H;��H;B�H;g�H;��H;��H;�H;X�H;�TH;�G;��C;��<;�-;��;�:�"
9+�$���Y�1�϶���  ��J� ��ձ�i{+��|x�jɰ�����7�%�A�W������ޞ�Nw�����      ����� �Կp���ޞ�bF�j�C�/E�$�;�I���D���!"��j�c�~��֯���J��ѻ��)��|K�4��:$�
;�M*;z�:;�C;�F;�8H;`�H;��H;��H;��H;Q�H;L�H;��H;��H;��H;�H;��H;��H;��H;K�H;O�H;��H;~�H;��H;`�H;�8H;�F;�C;v�:;�M*;$�
;:��: }K���)��ѻ��J��֯�~�j�c�!"�����D��I��$�;/E�j�C�bF��ޞ�p�� �Կ��      ��������� �ԿNw�����<�\�"����m��]0X�����;����w����������]��黾F�h�� ʒ:�;B�';Ə9;)pB;�zF;�!H;��H;B�H;(�H;��H;X�H;N�H;��H;��H;��H; �H;��H;��H;��H;L�H;X�H;��H;&�H;?�H;��H;�!H;�zF;)pB;9;D�';�;ʒ:h�깾F��黬�]����������w��;�����]0X�m�����"�<�\����Nw�� �Կ��𿞏�      !$�������忊�����"cm�X�-�����Sh��Zde�$-�ڪɽ�v��*�$���ɼymj�8����X�d���ņ:x;K�%;9�8;uB;wRF;H;8�H;_�H;�H;y�H;R�H;H�H;��H;��H;��H;5�H;��H;��H;��H;G�H;T�H;y�H;�H;\�H;8�H;H;uRF;uB;6�8;P�%;x;�ņ:h���X�7���zmj���ɼ*�$��v��ڪɽ$-�Zde�Sh������X�-�"cm��������忞����      gܿ5�ֿ�aǿ?^��1���\o���7����iþ�(���-=��` �A���_�3]�1p����I�R�ѻx�)���R���:E�
;�*;%�:;ܣB;HIF;6�G;�lH;;�H;��H;q�H;��H;��H;��H;��H;<�H;��H;<�H;��H;��H;��H;��H;q�H;��H;8�H;�lH;7�G;HIF;ܣB;"�:;�*;E�
;��:��R�x�)�P�ѻ��I�1p��3]��_�A���` ��-=��(���iþ����7�\o�1���?^���aǿ5�ֿ      5�ֿFpѿ�¿������bXi�ҕ3��
�XD��Hl��C�9��.���R��&\� �gx��1�E��ͻ�$�`��፨:S�;��*;>�:;�B;)UF;��G;[nH;֡H;�H;��H;��H;��H;��H;��H;Q�H;��H;Q�H;��H;��H;��H;��H;��H;�H;ԡH;[nH;��G;(UF;�B;9�:;��*;S�;㍨:����$��ͻ2�E�gx�� �&\��R���.��C�9�Hl��XD���
�ҕ3�bXi��������¿Fpѿ      �aǿ�¿����������"Y��f'�����:o���.}��k/����(ڟ�&<Q�0#�ע��(;�,���*�� 77�	�:�;�,;��;;�C;HwF;*�G;�rH;b�H;ǸH;G�H;+�H;'�H;��H;��H;}�H;�H;}�H;��H;��H;&�H;-�H;G�H;ŸH;_�H;�rH;*�G;GwF;�C;��;;�,;�;	�: 87�*��,����(;�ע�0#�&<Q�(ڟ�����k/��.}�:o�������f'��"Y�����������¿      ?^������m���\o���@�+�'�޾����<ce�2��¯ڽ����g@������R���O*�FG������`F^9>��:;�d.;�<;ǐC;=�F;��G;�yH;ͥH;?�H;T�H;��H;��H;�H;#�H;��H;G�H;��H;#�H;�H;��H;��H;T�H;=�H;˥H;�yH;��G;=�F;ƐC;�<;�d.;;@��:PF^9����FG���O*��R������g@�����¯ڽ2��<ce�����'�޾+���@�\o�m�������      1����������\o��!J�M�#��\��XD������}PH�����b��"C��� +���ټ*����꿐������:?��:a�;�Y1;>;�0D;��F;|H;v�H;�H;3�H;��H;��H;;�H;��H;��H;��H;��H;��H;~�H;��H;9�H;��H;��H;0�H;�H;v�H;~H;��F;�0D;>;�Y1;a�;A��:�:����꿐���)����ټ� +�"C���b�����}PH�����XD���\��M�#��!J�\o��������      \o�bXi��"Y���@�M�#��
��о�A���i���(����yr���_��5��ɺ�t�`��<��^�d��\���X:�P�: a; �4;ҧ?;��D;�8G;�0H;ˋH;��H;��H;9�H;��H;��H;,�H;��H;@�H;��H;@�H;��H;,�H;��H;��H;9�H;��H;��H;ˋH;�0H;�8G;��D;̧?;��4; a;�P�:��X:�\�\�d��<��t�`��ɺ��5��_�yr�������(��i��A���о�
�M�#���@��"Y�bXi�      ��7�ҕ3��f'�+��\���о�����.}��-=�~
���Ľ^��.:����������7�GĻ��$�pN����:�{;�D&;',8;1JA;+�E;��G;�LH;�H;��H;[�H;�H;9�H;��H;��H;Q�H;��H;I�H;��H;Q�H;��H;��H;;�H;�H;Z�H;��H;�H;�LH;��G;'�E;/JA;$,8;�D&;�{;��:pN����$�GĻ�7���������.:�^����Ľ~
��-=��.}������о�\��+��f'�ҕ3�      ���
�����&�޾XD���A���.}�+�D�jt���ڽ�!��\����_�ļ�
v�=��¿���Iɺ�S�9��:1(;�-;��;;��B;�IF;��G;CfH;ϝH;#�H;V�H;��H;��H;��H;��H;��H;#�H;��H;#�H;��H;��H;��H;��H;��H;V�H; �H;ΝH;AfH;��G;�IF;��B;��;;�-;2(;��:�S�9�Iɺ¿��=���
v�_�ļ���\��!����ڽjt�+�D��.}��A��XD��&�޾�����
�      �iþXD��:o�����������i��-=�jt����R��mys�} +����{񗼔(;�(�ѻ�s@���!�p4j:Q�:�;�D3;g�>;8FD;��F;�	H;c|H;ťH;��H;`�H;'�H;'�H;��H;P�H;f�H;��H;�H;��H;f�H;O�H;��H;*�H;'�H;`�H;��H;ƥH;`|H;�	H;��F;5FD;f�>;�D3;�;Q�:p4j:��!��s@�(�ѻ�(;�{����} +�mys��R����kt��-=��i���������:o��XD��      �(��Hl���.}�<ce�}PH���(�~
���ڽ�R���{�F�6�� �/p��b�`�̨��,��IҺ�M^9ɇ�:�;�~(;U�8;JA;+|E;DjG;�=H;p�H;
�H;Y�H;��H;]�H;��H;��H;�H;��H;%�H;~�H;%�H;��H;�H;��H;��H;]�H;��H;U�H;
�H;p�H;�=H;AjG;(|E;JA;U�8;�~(;�;ɇ�:�M^9IҺ�,��̨�b�`�/p��� �F�6��{��R����ڽ~
���(�}PH�<ce��.}�Hl��      �-=�C�9��k/�2��������Ľ�!��mys�F�6�&#��ɺ��vz����<^��X�$��}�r:>��:
�;�Y1;$I=;\xC;QwF;S�G;6fH;w�H;��H;��H;��H;��H;�H;�H;��H;��H;��H;��H;��H;��H;��H;�H;�H;��H;��H;��H;��H;v�H;5fH;Q�G;LwF;YxC;$I=;�Y1;�;>��:��r: ~�Y�$�<^������vz��ɺ�&#�F�6�mys��!����Ľ����2���k/�C�9�      �` ��.�����¯ڽ�b��yr��^��\�} +�� ��ɺ�B��O*�Bͻ�5R��ƅ�4�:[��:��;�);u8;��@;�*E;�8G;v$H;{�H;r�H;)�H;]�H;��H;��H;��H;4�H;��H;'�H;�H;W�H;�H;'�H;��H;4�H;��H;��H;��H;\�H;)�H;o�H;x�H;t$H;�8G;�*E;��@;u8;�);��;a��:4�:�ƅ��5R�Aͻ�O*�A��ɺ�� �} +�\�^��yr���b��¯ڽ��.��      A���R��(ڟ�����"C���_�/:�������/p���vz��O*��4ֻk������09r�:$1;w� ;�D3;m�=;ԐC;lF;��G;�\H;ЗH;��H;7�H;v�H;��H;��H;�H;1�H;A�H;��H;��H;��H;��H;��H;A�H;1�H;�H;��H;��H;u�H;7�H;}�H;ΗH;�\H;��G;lF;ԐC;m�=;�D3;w� ;&1;p�:��09���k��4ֻ�O*��vz�.p����輧��.:��_�"C������(ڟ��R��      �_�%\�%<Q�g@�� +��5�����^�ļz�a�`����Aͻk��Hɺ o6�r�:Q�:F�;e.;w�:;I�A;X|E;�NG;u'H;5�H; �H;��H;��H;c�H;��H;��H;j�H;/�H;��H;F�H;��H;7�H;��H;F�H;��H;/�H;m�H;��H;��H;`�H;��H;��H; �H;4�H;t'H;�NG;X|E;I�A;w�:;e.;I�;Q�:r�: n6��Hɺk�@ͻ���`�`�z�_�ļ�����5�� +�g@�%<Q�%\�      3]� �/#�������ټ�ɺ������
v��(;�ͨ�=^���5R���� q6����:��:�;E�*;,8;�!@;��D;��F;+�G;	fH;��H;ưH;׿H;��H;�H;��H;Z�H;��H;�H;��H;��H;`�H;��H;`�H;��H;��H;�H;��H;Z�H;��H;�H;��H;ֿH;ưH;��H;fH;&�G;��F;��D;�!@;,8;H�*;�;��:���: q6�����5R�=^��̨��(;��
v������ɺ���ټ����/#� �      0p��fx��ע��R��)��t�`� �7�>��&�ѻ�,��W�$��ƅ���09p�:#��:�;�~(;�Z6;��>;��C;!IF;�G;EH;�H;�H;�H;H�H;c�H;N�H;2�H;�H;��H;��H;I�H;$�H;��H;��H;��H;$�H;G�H;��H;��H;�H;2�H;H�H;c�H;F�H;�H;�H;{�H;EH;�G;IF;��C;��>;�Z6;�~(;�;#��:r�:��09�ƅ�W�$��,��&�ѻ>�� �7�s�`�)���R��ע�gx��      ��I�.�E��(;��O*����<��GĻ¿���s@�IҺ�}�4�:l�:Q�:�;�~(;3�5;�>;fC;f�E;�cG;p$H;/|H;q�H;W�H;��H;��H;t�H;�H;X�H;��H;��H;��H;��H;{�H;�H;-�H;�H;{�H;��H;��H;��H;��H;W�H;�H;t�H;��H;��H;V�H;l�H;*|H;q$H;�cG;h�E;fC;�>;5�5;�~(;�;Q�:l�:4�: ~�IҺ�s@�¿��GĻ�<�����O*��(;�1�E�      S�ѻ�ͻ*���EG��뿐�h�d���$��Iɺ��!��M^9��r:[��:$1;F�;G�*;�Z6;�>;a�B;��E;9G;�	H;6nH;P�H;�H;߽H;��H;��H;�H;��H;=�H;��H;��H;9�H;6�H;��H;@�H;c�H;>�H;��H;6�H;8�H;��H;��H;;�H;��H;�H;��H;��H;߽H;z�H;L�H;6nH;�	H;9G;��E;a�B;�>;�Z6;G�*;G�;$1;[��:��r:�M^9��!��Iɺ��$�d�d�鿐�DG��)����ͻ      m�)��$�!����������\�PN���S�9t4j:Ň�:B��:��;w� ;e.;,8;��>;cC;��E;�)G;��G;JdH;��H;ϫH;��H;��H;r�H;�H;�H;��H;��H;��H;��H;��H;��H;:�H;o�H;��H;o�H;:�H;��H;��H;��H;��H;��H;��H;�H;�H;t�H;��H;��H;˫H;��H;FdH;��G;�)G;��E;cC;��>;,8;e.;w� ;��;>��:ɇ�:|4j:�S�9@N�� �\�򬷺���!���$�      ��R�`�� 57�PF^9�:�X:��:��:Q�:�;
�;�);�D3;s�:;�!@;��C;f�E;9G;��G;�`H;��H;R�H;T�H;��H;|�H;q�H;��H;��H;��H;�H;��H;F�H;'�H;��H;h�H;��H;��H;��H;h�H;��H;%�H;G�H;��H;�H;��H;��H;��H;q�H;}�H;��H;Q�H;R�H;��H;�`H;��G;9G;f�E;��C;�!@;s�:;�D3;�);
�;�;Q�:��:��:��X:8�:PF^9 57� ��      ��:��:�:0��:-��:�P�:�{;0(;�;�~(;�Y1;u8;m�=;K�A;��D;IF;�cG;�	H;JdH;��H;��H;�H;k�H;/�H;�H;|�H;��H;��H;b�H;#�H;��H;��H;��H;%�H;��H;��H;��H;��H;��H;#�H;��H;��H;��H;!�H;_�H;��H;��H;|�H;	�H;,�H;m�H;�H;~�H;��H;JdH;�	H;�cG;IF;��D;K�A;m�=;u8;�Y1;�~(;�;0(;�{;�P�:1��:2��:�:፨:      K�
;o�;�;;a�;a;�D&;�-;�D3;V�8;*I=;��@;אC;[|E;��F;�G;q$H;8nH;��H;T�H;�H;��H;t�H;Z�H;��H;��H;!�H;��H;��H;F�H;^�H;3�H;��H;\�H;��H;��H;��H;��H;��H;\�H;��H;3�H;^�H;B�H;��H;��H;�H;��H;��H;W�H;t�H;��H;�H;U�H;��H;8nH;q$H;�G;��F;[|E;אC;��@;*I=;X�8;�D3;�-;�D&;a;v�;;�;j�;      �*;��*;�,;�d.;�Y1; �4;*,8;��;;i�>;JA;_xC;�*E;lF;�NG;+�G;EH;.|H;P�H;ϫH;W�H;m�H;w�H;��H;7�H;5�H;��H;J�H;(�H;��H;�H;��H;��H;!�H;x�H;��H;��H;��H;��H;��H;x�H;!�H;��H;��H;�H;��H;(�H;H�H;��H;6�H;5�H;��H;x�H;j�H;Z�H;ϫH;P�H;,|H;EH;+�G;�NG;lF;�*E;\xC;JA;i�>;��;;+,8;�4;�Y1;�d.;�,;��*;      9�:;I�:;��;;�<;>;Ч?;:JA;��B;9FD;)|E;RwF;�8G;��G;x'H;	fH;}�H;p�H;��H;��H;��H;,�H;Z�H;6�H;!�H;W�H;��H;��H;q�H;��H;��H;U�H;��H;Z�H;��H;��H;��H;�H;��H;��H;��H;Y�H;��H;U�H;��H;��H;r�H;��H;��H;X�H;�H;5�H;[�H;*�H;��H;��H;��H;n�H;}�H;	fH;x'H;��G;�8G;QwF;)|E;9FD;��B;8JA;Ч?;#>;�<;��;;<�:;      �B;(�B;�C;ʐC;�0D;��D;)�E;�IF;��F;DjG;S�G;z$H;�\H;9�H;��H;�H;]�H;�H;��H;��H;�H;��H;:�H;\�H;��H;��H;9�H;��H;h�H;5�H;��H;�H;n�H;��H;��H;��H;��H;��H;��H;��H;m�H;�H;��H;5�H;f�H;��H;9�H;��H;��H;[�H;9�H;��H;�H;��H;��H;�H;Z�H;�H;��H;8�H;�\H;z$H;S�G;AjG;��F;�IF;)�E;��D;�0D;͐C;�C;)�B;      UIF;7UF;=wF;:�F;��F;�8G;��G;��G;�	H;�=H;6fH;|�H;ΗH; �H;İH;�H;��H;��H;q�H;q�H;y�H;��H;��H;��H;��H;6�H;e�H;J�H;��H;��H;�H;`�H;u�H;��H;��H;��H;��H;��H;��H;��H;r�H;a�H;�H;��H;��H;J�H;d�H;9�H;��H;��H;��H;��H;u�H;q�H;q�H;��H;��H;�H;İH; �H;ΗH;|�H;6fH;�=H;�	H;��G;��G;�8G;��F;;�F;@wF;*UF;      C�G;��G;*�G;��G;�H;�0H;�LH;DfH;f|H;r�H;w�H;t�H;}�H;��H;׿H;J�H;��H;��H;�H;��H;��H;!�H;I�H;��H;3�H;h�H;<�H;��H;��H;��H;!�H;n�H;��H;��H;��H;��H;��H;��H;��H;��H;��H;n�H;!�H;��H;��H;��H;;�H;h�H;9�H;��H;H�H;!�H;��H;��H;�H;��H;��H;G�H;׿H;��H;}�H;t�H;w�H;p�H;g|H;CfH;�LH;�0H;�H;��G;+�G;��G;      �lH;^nH;�rH;�yH;w�H;΋H;�H;ٝH;̥H;�H;��H;0�H;8�H;��H;��H;d�H;t�H;�H;�H;��H;��H;��H;(�H;t�H;z�H;J�H;��H;q�H;��H;*�H;G�H;x�H;��H;��H;��H;��H;��H;��H;��H;��H;��H;x�H;H�H;&�H;��H;r�H;��H;L�H;}�H;t�H;(�H;��H;��H;��H;�H;�H;r�H;d�H;��H;��H;7�H;/�H;��H;�H;ͥH;ٝH;�H;͋H;��H;�yH;�rH;hnH;      P�H;ܡH;^�H;ҥH;�H;��H;��H;(�H;��H;\�H;��H;c�H;x�H;c�H;�H;N�H;�H;��H;��H;��H;b�H;��H;��H;��H;a�H;��H;��H;��H;	�H;N�H;k�H;��H;��H;��H;��H;��H;��H;��H;��H;��H;��H;��H;k�H;L�H;
�H;��H;��H;��H;c�H;��H;��H;��H;_�H;��H;��H;��H;�H;N�H;�H;c�H;x�H;`�H;��H;Y�H;��H;'�H;��H;��H;�H;ҥH;`�H;ҡH;      ��H;�H;ѸH;A�H;C�H;��H;e�H;^�H;k�H;��H;��H;��H;��H;��H;��H;6�H;[�H;9�H;��H;�H;"�H;C�H;�H;��H;+�H;��H;��H;&�H;L�H;a�H;��H;�H;��H;��H;��H;��H;��H;��H;��H;��H;��H;��H;��H;`�H;K�H;&�H;��H;��H;,�H;��H;�H;C�H;"�H;�H;��H;9�H;Z�H;4�H;��H;��H;��H;��H;��H;��H;m�H;a�H;c�H;��H;A�H;A�H;͸H;�H;      x�H;��H;U�H;`�H;��H;:�H;�H;�H;1�H;d�H;��H;��H;��H;��H;_�H;�H;��H;��H;��H;��H;��H;^�H;��H;Y�H;��H;�H;�H;H�H;j�H;��H;��H;��H;{�H;}�H;��H;��H;m�H;��H;��H;}�H;x�H;��H;��H;��H;k�H;H�H;�H;�H;��H;X�H;��H;^�H;��H;��H;��H;��H;��H;�H;^�H;��H;��H;��H;��H;d�H;2�H;�H;�H;=�H;��H;b�H;V�H;��H;      ��H;��H;5�H;��H;��H;��H;?�H;��H;0�H;��H;�H;��H;�H;r�H;��H;��H;��H;��H;��H;P�H;��H;7�H;��H;��H;�H;^�H;k�H;x�H;��H;��H;��H;��H;|�H;v�H;��H;n�H;d�H;n�H;��H;v�H;y�H;��H;��H;��H;��H;x�H;k�H;]�H;�H;��H;��H;7�H;��H;P�H;��H;��H;��H;��H;��H;t�H;�H;��H;�H;��H;1�H;��H;?�H;��H;��H;��H;6�H;��H;      ��H;��H;3�H;��H;I�H;��H;��H;��H;��H;��H;�H;?�H;6�H;6�H;
�H;��H;��H;5�H;��H;+�H;��H;��H;!�H;^�H;g�H;t�H;��H;��H;��H;��H;{�H;�H;��H;�H;]�H;]�H;��H;]�H;]�H;�H;}�H;��H;{�H;��H;��H;��H;��H;r�H;h�H;^�H;�H;��H;��H;,�H;��H;8�H;��H;��H;	�H;6�H;5�H;>�H;�H;��H;��H;��H;��H;��H;B�H;��H;3�H;��H;      ��H;��H;��H;�H;��H;)�H;��H;��H;W�H;�H;��H;��H;E�H;�H;��H;Q�H;��H;6�H;��H;��H;(�H;]�H;v�H;��H;��H;��H;��H;��H;��H;��H;|�H;x�H;{�H;h�H;Y�H;^�H;c�H;^�H;Y�H;h�H;y�H;{�H;|�H;��H;��H;��H;��H;��H;��H;��H;v�H;]�H;(�H;��H;��H;7�H;��H;Q�H;��H;�H;E�H;��H;��H;�H;Z�H;��H;��H;.�H;��H;�H;��H;��H;      ��H;��H;��H;.�H;��H;��H;^�H;��H;q�H;��H;��H;5�H;��H;N�H;��H;.�H;��H;��H;:�H;o�H;��H;��H;��H;��H;��H;��H;��H;��H;��H;��H;��H;��H;\�H;Y�H;d�H;Y�H;=�H;Y�H;d�H;Z�H;Y�H;��H;��H;��H;��H;��H;��H;��H;��H;��H;��H;��H;��H;o�H;:�H;��H;��H;.�H;��H;N�H;��H;5�H;��H; �H;q�H;��H;^�H;��H;��H;0�H;��H;��H;      9�H;_�H;��H;��H;��H;=�H;��H;2�H;��H;)�H;��H;$�H;��H;��H;g�H;��H;�H;9�H;q�H;��H;��H;��H;��H;��H;��H;��H;��H;��H;��H;��H;��H;r�H;\�H;c�H;Z�H;V�H;E�H;V�H;Z�H;`�H;Z�H;u�H;��H;��H;��H;��H;��H;��H;��H;��H;��H;��H;��H;��H;q�H;:�H;�H;��H;f�H;��H;��H;$�H;��H;,�H;��H;0�H;��H;A�H;��H;��H;��H;W�H;      ��H;�H;�H;M�H;��H;��H;R�H;��H;#�H;��H;��H;c�H;��H;@�H;��H;��H;3�H;Z�H;��H;��H;��H;��H;��H;�H;��H;��H;��H;��H;��H;��H;o�H;k�H;��H;e�H;=�H;G�H;@�H;G�H;=�H;e�H;��H;m�H;o�H;��H;��H;��H;��H;��H;��H;�H;��H;��H;��H;��H;��H;\�H;2�H;��H;��H;@�H;��H;c�H;��H;��H;%�H;��H;R�H;��H;��H;M�H;�H;��H;      9�H;_�H;��H;��H;��H;=�H;��H;2�H;��H;)�H;��H;$�H;��H;��H;f�H;��H;�H;9�H;q�H;��H;��H;��H;��H;��H;��H;��H;��H;��H;��H;��H;��H;r�H;\�H;c�H;Z�H;V�H;E�H;V�H;Z�H;`�H;Z�H;u�H;��H;��H;��H;��H;��H;��H;��H;��H;��H;��H;��H;��H;q�H;:�H;�H;��H;g�H;��H;��H;$�H;��H;*�H;��H;0�H;��H;A�H;��H;��H;��H;U�H;      ��H;��H;��H;0�H;��H;��H;\�H;��H;q�H;��H;��H;5�H;��H;N�H;��H;.�H;��H;��H;:�H;o�H;��H;��H;��H;��H;��H;��H;��H;��H;��H;��H;��H;��H;\�H;Z�H;d�H;Y�H;=�H;Y�H;d�H;Y�H;Y�H;��H;��H;��H;��H;��H;��H;��H;��H;��H;��H;��H;��H;o�H;:�H;��H;��H;.�H;��H;N�H;��H;5�H;��H; �H;q�H;��H;^�H;��H;��H;0�H;��H;��H;      ��H;��H;��H;�H;��H;)�H;��H;��H;W�H;�H;��H;��H;E�H;�H;��H;Q�H;��H;6�H;��H;��H;*�H;]�H;v�H;��H;��H;��H;��H;��H;��H;��H;|�H;x�H;{�H;h�H;Y�H;^�H;c�H;^�H;Y�H;h�H;y�H;{�H;|�H;��H;��H;��H;��H;��H;��H;��H;v�H;]�H;(�H;��H;��H;7�H;��H;Q�H;��H;�H;E�H;��H;��H;�H;X�H;��H;��H;.�H;��H;�H;��H;��H;      ��H;��H;4�H;��H;I�H;��H;��H;��H;��H;��H;�H;>�H;5�H;6�H;	�H;��H;��H;5�H;��H;+�H;��H;��H;!�H;^�H;h�H;t�H;��H;��H;��H;��H;{�H;�H;�H;}�H;]�H;]�H;��H;\�H;]�H;}�H;}�H;��H;{�H;��H;��H;��H;��H;r�H;g�H;]�H;�H;��H;��H;,�H;��H;6�H;��H;��H;
�H;6�H;5�H;?�H;�H;��H;��H;��H;��H;��H;@�H;��H;0�H;��H;      ��H;��H;6�H;��H;��H;��H;C�H;��H;0�H;��H;�H;��H;�H;r�H;��H;��H;��H;��H;��H;P�H;��H;7�H;��H;��H;�H;^�H;k�H;x�H;��H;��H;��H;��H;y�H;v�H;��H;n�H;d�H;n�H;��H;v�H;y�H;��H;��H;��H;��H;x�H;k�H;]�H;�H;��H;��H;7�H;��H;P�H;��H;��H;��H;��H;��H;r�H;�H;��H;�H;��H;1�H;��H;B�H;��H;��H;��H;6�H;��H;      x�H;��H;U�H;b�H;��H;:�H;�H;�H;2�H;c�H;��H;��H;��H;��H;^�H;�H;��H;��H;��H;��H;��H;^�H;��H;[�H;��H;�H;�H;H�H;h�H;��H;��H;��H;y�H;}�H;��H;��H;m�H;��H;��H;}�H;x�H;��H;��H;��H;k�H;H�H;�H;�H;��H;X�H;��H;^�H;��H;��H;��H;��H;��H;�H;_�H;��H;��H;��H;��H;e�H;2�H;	�H;�H;=�H;��H;`�H;U�H;��H;      ��H;�H;иH;@�H;A�H;��H;f�H;a�H;k�H;��H;��H;��H;��H;��H;��H;4�H;[�H;7�H;��H;�H;%�H;C�H;�H;��H;,�H;��H;��H;&�H;K�H;a�H;��H;�H;��H;��H;��H;��H;��H;��H;��H;��H;��H;��H;��H;`�H;L�H;&�H;��H;��H;+�H;��H;�H;C�H;"�H;�H;��H;:�H;Z�H;7�H;��H;��H;��H;��H;��H;��H;n�H;b�H;f�H;��H;?�H;A�H;иH;�H;      I�H;ءH;c�H;ХH;�H;��H;��H;(�H;��H;Y�H;��H;a�H;x�H;c�H;�H;N�H;�H;��H;��H;��H;e�H;��H;��H;��H;c�H;�H;��H;��H;	�H;N�H;k�H;��H;��H;��H;��H;��H;��H;��H;��H;��H;��H;��H;k�H;L�H;	�H;��H;��H;��H;a�H;��H;��H;��H;a�H;��H;��H;��H;�H;O�H;�H;c�H;x�H;c�H;��H;[�H;��H;(�H;��H;��H;�H;̥H;g�H;աH;      �lH;^nH;�rH;�yH;y�H;͋H;�H;ٝH;̥H;�H;��H;/�H;7�H;��H;��H;d�H;t�H;
�H;�H;��H;��H;��H;(�H;t�H;}�H;J�H;��H;r�H;��H;*�H;H�H;x�H;��H;��H;��H;��H;��H;��H;��H;��H;��H;y�H;G�H;(�H;��H;q�H;��H;J�H;z�H;t�H;'�H;��H;��H;��H;�H;�H;r�H;e�H;��H;��H;8�H;/�H;��H;�H;ͥH;۝H;�H;ˋH;��H;�yH;�rH;hnH;      =�G;��G;+�G;��G;�H;�0H;�LH;DfH;f|H;q�H;w�H;t�H;}�H;��H;׿H;H�H;��H;��H;�H;��H;��H;!�H;I�H;��H;9�H;h�H;<�H;��H;��H;��H;!�H;n�H;��H;��H;��H;��H;��H;��H;��H;��H;��H;o�H;!�H;��H;��H;��H;;�H;h�H;3�H;��H;H�H;!�H;��H;��H;�H;��H;��H;H�H;׿H;��H;}�H;t�H;z�H;q�H;g|H;DfH;�LH;�0H;�H;��G;(�G;��G;      ZIF;4UF;HwF;=�F;��F;�8G;��G;��G;�	H;�=H;6fH;y�H;ΗH; �H;ðH;�H;��H;��H;q�H;q�H;{�H;��H;��H;��H;��H;7�H;g�H;J�H;��H;��H;�H;`�H;t�H;��H;��H;��H;��H;��H;��H;��H;r�H;a�H;�H;��H;��H;J�H;d�H;7�H;��H;��H;��H;��H;v�H;q�H;q�H;��H;��H;�H;İH; �H;͗H;|�H;6fH;�=H;�	H;��G;��G;�8G;��F;;�F;HwF;&UF;      �B;(�B;�C;͐C;�0D;��D;)�E;�IF;��F;BjG;U�G;z$H;�\H;8�H;��H;�H;[�H;�H;��H;��H;�H;��H;:�H;\�H;��H;��H;:�H;��H;i�H;6�H;��H;�H;m�H;��H;��H;��H;��H;��H;��H;��H;m�H;�H;��H;3�H;e�H;��H;7�H;��H;��H;\�H;9�H;��H;�H;��H;��H;�H;Z�H;�H;��H;8�H;�\H;z$H;S�G;BjG;��F;�IF;)�E;��D;�0D;ʐC;�C;(�B;      ;�:;H�:;��;;�<;>;ԧ?;6JA;��B;;FD;,|E;RwF;�8G;��G;x'H;	fH;}�H;p�H;�H;��H;��H;-�H;[�H;6�H;!�H;X�H;��H;��H;r�H;��H;��H;U�H;��H;Z�H;��H;��H;��H;�H;��H;��H;��H;Y�H;��H;U�H;��H;��H;q�H;��H;��H;W�H; �H;5�H;Z�H;*�H;��H;��H;��H;n�H;}�H;	fH;w'H;��G;�8G;QwF;(|E;;FD;��B;4JA;֧?;'>;�<;��;;9�:;      �*;��*;�,;�d.;�Y1;�4;/,8;��;;i�>;JA;\xC;�*E;lF;�NG;+�G;EH;.|H;M�H;ϫH;X�H;p�H;x�H;��H;7�H;6�H;��H;J�H;(�H;��H;�H;��H;��H;!�H;x�H;��H;��H;��H;��H;��H;x�H;�H;��H;��H;�H;��H;(�H;H�H;��H;5�H;5�H;��H;w�H;i�H;X�H;ϫH;R�H;.|H;EH;-�G;�NG;lF;�*E;]xC;	JA;i�>;��;;/,8;�4;�Y1;�d.;�,;��*;      K�
;o�;�;;d�;
a;�D&;�-;�D3;X�8;*I=;��@;אC;[|E;��F;�G;p$H;6nH;��H;T�H;�H;��H;u�H;[�H;��H;��H;!�H;��H;��H;F�H;^�H;3�H;��H;\�H;��H;��H;��H;��H;��H;\�H;��H;3�H;^�H;B�H;��H;��H;�H;��H;��H;W�H;q�H;��H;�H;U�H;��H;9nH;p$H;�G;��F;[|E;אC;��@;*I=;V�8;�D3;�-;�D&;a;w�;;�;j�;      ��:���:�:2��:1��:�P�:�{;2(;�;�~(;�Y1;u8;l�=;K�A;��D;IF;�cG;�	H;JdH;��H;��H;�H;n�H;0�H;	�H;|�H;��H;��H;a�H;#�H;��H;��H;��H;"�H;��H;��H;��H;��H;��H;%�H;��H;��H;��H;!�H;_�H;��H;��H;|�H;�H;*�H;j�H;�H;~�H;��H;JdH;�	H;�cG;IF;��D;K�A;n�=;u8;�Y1;�~(;�;2(;�{;�P�:9��:0��:�:ߍ�:      ��R�`�� 17�0F^9$�:�X:��:��:Q�:�;�;�);�D3;s�:;�!@;��C;f�E;9G;��G;�`H;��H;R�H;T�H;��H;}�H;q�H;��H;��H;��H;�H;��H;F�H;'�H;��H;h�H;��H;��H;��H;h�H;��H;%�H;G�H;��H;�H;��H;��H;��H;q�H;|�H;��H;Q�H;R�H;��H;�`H;��G;9G;f�E;��C;�!@;s�:;�D3;�);�;�;Q�:��:��:��X:@�:0F^9 17���      m�)��$� ����������\�@N���S�9t4j:ɇ�:B��:��;w� ;e.;,8;��>;cC;��E;�)G;��G;HdH;��H;ϫH;��H;��H;r�H;�H;�H;��H;��H;��H;��H;��H;��H;:�H;o�H;��H;o�H;:�H;��H;��H;��H;��H;��H;��H;�H;�H;r�H;��H;��H;˫H;��H;GdH;��G;�)G;��E;aC;��>;,8;e.;w� ;��;B��:Ň�:|4j:�S�9PN�� �\�𬷺���!���$�      R�ѻ�ͻ*���EG��쿐�i�d���$��Iɺ��!��M^9��r:[��:&1;F�;G�*;�Z6;�>;`�B;��E;9G;�	H;6nH;P�H;�H;߽H;��H;��H;�H;��H;=�H;��H;��H;9�H;6�H;��H;@�H;c�H;@�H;��H;6�H;8�H;��H;��H;;�H;��H;�H;��H;��H;߽H;{�H;M�H;6nH;�	H;9G;��E;a�B;�>;�Z6;G�*;F�;$1;[��:��r:�M^9��!��Iɺ��$�e�d�运�FG��*����ͻ      ��I�/�E��(;��O*����<��GĻ¿���s@�IҺ�}�4�:l�:Q�:�;�~(;5�5;�>;dC;g�E;�cG;q$H;/|H;p�H;V�H;��H;��H;t�H;�H;X�H;��H;��H;��H;��H;{�H;�H;-�H;�H;{�H;��H;��H;��H;��H;W�H;�H;t�H;��H;��H;W�H;m�H;*|H;p$H;�cG;h�E;fC;�>;5�5;�~(;�;Q�:l�:4�:�}�IҺ�s@�����GĻ�<�����O*��(;�1�E�      0p��fx��ע��R��)��t�`� �7�=��&�ѻ�,��W�$��ƅ���09p�:#��:�;�~(;�Z6;��>;��C;IF;�G;EH;�H;�H;�H;H�H;c�H;M�H;2�H;�H;��H;��H;G�H;$�H;��H;��H;��H;$�H;I�H;��H;��H;�H;2�H;J�H;c�H;F�H;�H;�H;{�H;EH;�G;IF;��C;��>;�Z6;�~(;�;#��:p�:��09�ƅ�W�$��,��&�ѻ=�� �7�s�`�)���R��ע�gx��      3]� �/#�������ټ�ɺ������
v��(;�̨�=^���5R���� q6����:��:�;D�*;,8;�!@;��D;��F;-�G;fH;��H;ðH;׿H;��H;�H;��H;Z�H;��H;�H;��H;��H;`�H;��H;`�H;��H;��H;�H;��H;Z�H;��H;�H;��H;ֿH;ǰH;��H;fH;&�G;��F;��D;�!@;,8;H�*;�;��:���: q6�����5R�<^��ͨ��(;��
v������ɺ���ټ����/#� �      �_�%\�%<Q�g@�� +��5�����_�ļz�a�`����Bͻk��Hɺ n6�r�:Q�:G�;e.;w�:;H�A;X|E;�NG;w'H;4�H;��H;��H;��H;a�H;��H;��H;j�H;0�H;��H;F�H;��H;7�H;��H;F�H;��H;.�H;k�H;��H;��H;a�H;��H;��H;�H;5�H;r'H;�NG;X|E;K�A;w�:;e.;I�;Q�:r�: o6��Hɺk�Aͻ���a�`�z�_�ļ�����5�� +�g@�%<Q�%\�      A���R��(ڟ�����"C���_�.:�������.p���vz��O*��4ֻk������09r�:$1;w� ;�D3;l�=;ԐC;lF;��G;�\H;ΗH;��H;7�H;v�H;��H;��H;�H;1�H;A�H;��H;��H;��H;��H;��H;A�H;/�H;�H;��H;��H;t�H;7�H;}�H;їH;�\H;��G;lF;ԐC;m�=;�D3;w� ;&1;p�:��09���k��4ֻ�O*��vz�/p����輧��/:��_�"C������(ڟ��R��      �` ��.�����¯ڽ�b��yr��^��\�} +�� ��ɺ�A��O*�Bͻ�5R��ƅ�4�:_��:��;�);u8;��@;�*E;�8G;t$H;y�H;r�H;)�H;]�H;��H;��H;��H;5�H;��H;'�H;�H;W�H;�H;'�H;��H;3�H;��H;��H;��H;\�H;)�H;p�H;y�H;v$H;�8G;�*E;��@;u8;�);��;a��:0�:�ƅ��5R�Bͻ�O*�A��ɺ�� �} +�\�^��yr���b��¯ڽ��.��      �-=�C�9��k/�2��������Ľ�!��mys�F�6�&#��ɺ��vz����<^��Y�$��}�r:>��:
�;�Y1;$I=;\xC;QwF;Q�G;6fH;w�H;��H;��H;��H;��H;�H;�H;��H;��H;��H;��H;��H;��H;��H;�H;�H;��H;��H;��H;��H;v�H;6fH;S�G;LwF;YxC;$I=;�Y1;�;>��:��r: ~�Z�$�<^������vz��ɺ�&#�F�6�mys��!����Ľ����2���k/�C�9�      �(��Hl���.}�<ce�}PH���(�~
���ڽ�R���{�F�6�� �/p��b�`�̨��,��IҺ�M^9ɇ�:�;�~(;U�8;JA;+|E;AjG;�=H;q�H;
�H;X�H;��H;]�H;��H;��H;�H;��H;%�H;~�H;%�H;��H;�H;��H;��H;]�H;��H;U�H;
�H;n�H;�=H;DjG;(|E;JA;U�8;�~(;�;ɇ�:�M^9IҺ�,��̨�b�`�/p��� �F�6��{��R����ڽ~
���(�}PH�<ce��.}�Hl��      �iþXD��:o�����������i��-=�jt����R��mys�} +����{񗼔(;�(�ѻ�s@���!�p4j:Q�:�;�D3;g�>;8FD;��F;�	H;c|H;ƥH;��H;`�H;'�H;)�H;��H;O�H;f�H;��H;�H;��H;f�H;P�H;��H;'�H;'�H;^�H;��H;ťH;`|H;�	H;��F;7FD;f�>;�D3;�;Q�:p4j:��!��s@�(�ѻ�(;�{����} +�mys��R����jt��-=��i���������:o��XD��      ���
�����&�޾XD���A���.}�+�D�jt���ڽ�!��\����_�ļ�
v�=��¿���Iɺ�S�9��:0(;�-;��;;��B;�IF;��G;CfH;ΝH;#�H;V�H;��H;��H;��H;��H;��H;#�H;��H;%�H;��H;��H;��H;��H;��H;V�H; �H;ϝH;AfH;��G;�IF;��B;��;;�-;2(;��:�S�9�Iɺÿ��=���
v�_�ļ���\��!����ڽjt�+�D��.}��A��XD��&�޾�����
�      ��7�ҕ3��f'�+��\���о�����.}��-=�~
���Ľ^��.:����������7�GĻ��$�pN����:�{;�D&;',8;3JA;'�E;��G;�LH;�H;��H;[�H;�H;9�H;��H;��H;Q�H;��H;I�H;��H;Q�H;��H;��H;9�H;�H;Z�H;��H;�H;�LH;��G;+�E;/JA;%,8;�D&;�{;��:pN����$�GĻ�7���������.:�^����Ľ~
��-=��.}������о�\��+��f'�ҕ3�      \o�bXi��"Y���@�M�#��
��о�A���i���(����yr���_��5��ɺ�t�`��<��]�d��\���X:�P�: a;��4;Ч?;��D;�8G;�0H;ˋH;��H;��H;9�H;��H;��H;,�H;��H;@�H;��H;A�H;��H;,�H;��H;��H;9�H;��H;��H;ˋH;�0H;�8G;��D;ͧ?; �4; a;�P�:��X:�\�\�d��<��t�`��ɺ��5��_�yr�������(��i��A���о�
�M�#���@��"Y�bXi�      1����������\o��!J�M�#��\��XD������}PH�����b��"C��� +���ټ*����꿐������:9��:a�;�Y1;>;�0D;��F;|H;v�H;�H;3�H;��H;��H;;�H;��H;��H;��H;��H;��H;~�H;��H;9�H;��H;��H;0�H;�H;v�H;~H;��F;�0D;>;�Y1;a�;A��:�:����꿐���*����ټ� +�"C���b�����}PH�����XD���\��M�#��!J�\o��������      ?^������m���\o���@�+�'�޾����<ce�2��¯ڽ����g@������R���O*�FG������`F^9<��:;�d.;�<;ƐC;=�F;��G;�yH;̥H;@�H;T�H;��H;��H;�H;#�H;��H;G�H;��H;#�H;�H;��H;��H;T�H;=�H;˥H;�yH;��G;=�F;ǐC;	�<;�d.;;@��:PF^9����FG���O*��R������g@�����¯ڽ2��<ce�����'�޾+���@�\o�m�������      �aǿ�¿����������"Y��f'�����:o���.}��k/����(ڟ�&<Q�/#�ע��(;�,���*�� 87��:�;�,;��;;�C;HwF;*�G;�rH;b�H;ǸH;G�H;+�H;'�H;��H;��H;}�H;�H;}�H;��H;��H;&�H;-�H;G�H;ŸH;_�H;�rH;*�G;GwF;�C;��;;�,;�;	�: 87�*��,����(;�ע�0#�&<Q�(ڟ�����k/��.}�:o�������f'��"Y�����������¿      5�ֿFpѿ�¿������bXi�ҕ3��
�XD��Hl��C�9��.���R��&\� �gx��1�E��ͻ�$�p��፨:S�;��*;>�:;�B;)UF;��G;[nH;֡H;�H;��H;��H;��H;��H;��H;Q�H;��H;Q�H;��H;��H;��H;��H;��H;�H;ԡH;[nH;��G;(UF;�B;;�:;��*;S�;㍨:����$��ͻ2�E�gx�� �&\��R���.��C�9�Hl��XD���
�ҕ3�bXi��������¿Fpѿ      �?��~h��?v��� ��:�X��O/�1y�D�;㰖��+X����ѽ����dn;�a�������B(�ܚ��D���e9 �:;�Y.;[�<;�WC;/[F;�G;30H;zjH;]�H;|�H;��H;X�H;��H;��H;��H;��H;��H;��H;��H;V�H;��H;|�H;[�H;wjH;30H;�G;.[F;�WC;Y�<;�Y.;;"�:��e9D��ښ���B(�����a��dn;������ѽ���+X�㰖�D�;1y��O/�:�X�� ��?v��~h��      ~h��1���c�����y�YvS�rM+��v�9ɾ�����T�"]�\ν����|\8�����x��%�P���`�뺠�9u-�:}�;��.;%�<;oC;�dF;��G;�1H;(kH;ΌH;ڤH;�H;��H;�H;��H; �H;��H; �H;��H;�H;��H;�H;ڤH;ʌH;%kH;�1H;��G;�dF;oC;!�<;��.;}�;y-�:��9`��P���%��x�����|\8�����\ν#]��T�����9ɾ�v�rM+�YvS���y�c���1���      ?v��c���X ��c�h�9E�Z��m���㼾���nH�Ո�}�ý�Ȅ��s/��o��#�����&J��к�
�9`g�:�l;^0;+]=;�C;'�F;��G;M6H;dmH;O�H;إH;��H;/�H;u�H;�H;8�H;�H;8�H;�H;u�H;-�H;��H;إH;J�H;amH;O6H;��G;%�F;�C;']=;a0;�l;`g�:�
�9к$J������#���o��s/��Ȅ�}�ýՈ��nH���㼾m���Z��9E�c�h�X ��c���      � ����y�c�h��N��O/����E�߾B���*|��6�s}�䳽nSt�@�!�urμGF{��_��X�������:6��:[;�2;�O>;�D;s�F;��G;J=H;�pH;��H;�H;�H;�H;�H;��H;��H;��H;��H;��H;�H;�H;�H;}�H;��H;�pH;J=H;��G;p�F;�D;�O>;�2;[;<��:�:�����X���_�GF{�urμ@�!�nSt�䳽s}��6��*|�B��E�߾����O/��N�c�h���y�      :�X�YvS�9E��O/��S�KW����������OS\��� ���=����Y�~��ԃ����]�����"�b�`�Y���Y:��:~`;n�4;��?;j�D;�F;(�G;7FH;�uH;�H;éH;��H;F�H;��H;V�H;L�H;,�H;L�H;T�H;��H;D�H;��H;éH;�H;�uH;7FH;)�G;�F;h�D;��?;p�4;~`;��:��Y:h�Y�!�b�������]�ԃ��~���Y�=����彔� �OS\���������KW���S��O/�9E�YvS�      �O/�rM+�Z�����JW��9ɾD���Mw�� :�l��{�ý M��`n;�d���wv���E<��˻��-�����y�:�^;�%;��7;��@;E5E;�"G;)�G;lPH;<{H;�H;��H;��H;��H;+�H;D�H;�H;��H;�H;D�H;)�H;��H;��H;��H;�H;8{H;lPH;'�G;�"G;C5E;��@;��7;�%;�^;�y�:�����-��˻�E<�wv��c���`n;� M��{�ýl��� :��Mw�D��9ɾJW�����Z��rM+�      1y��v�m���E�߾����D��A����nH���Gὠu����d�3O�nrμL"�����	�����`s89�;�:p�;�+;�|:;�7B;�E;?bG;�H; [H;��H;S�H;ϯH;,�H;y�H;{�H;<�H;�H;��H;�H;<�H;y�H;y�H;.�H;ϯH;Q�H;��H; [H;�H;>bG;�E;�7B;�|:;�+;q�;�;�:`s89���	�����L"��nrμ3O���d��u��G����nH�A���D������E�߾m����v�      C�;9ɾ㼾B�������Mw��nH�����Z�䳽͕��u\8�t#������^N�N����b��Hx��5:3��:B�; �0;O]=;_�C;�[F;�G;*H;fH;��H;M�H;t�H;��H;M�H;�H;b�H;�H;��H; �H;b�H;�H;K�H;��H;r�H;M�H;��H;fH;*H;�G;�[F;[�C;O]=; �0;D�;1��:�5:�Hx���b�M��^N�����t#��u\8�͕��䳽�Z񽳯��nH��Mw�����B��㼾9ɾ      㰖��������*|�OS\�� :����Z�o$�������K�x���Oļ����������2&� ��r/�:�^;��#;�G6;m�?;�D;~�F;��G;+@H;�pH;�H;��H;E�H;��H;^�H;��H;��H;	�H;��H;	�H;��H;��H;^�H;��H;E�H;��H;�H;�pH;)@H;��G;z�F;�D;k�?;�G6;��#;�^;r/�:���2&������������Oļx���K�����o$���Z���� :�PS\��*|�������      �+X��T��nH��6��� �l��G�䳽�����mR����ټ�����E<��?ݻ/d\�����8!:�d�:��;B�,;��:;�7B;��E;�LG;iH;�SH;�{H;��H;�H;G�H;r�H;��H;B�H;��H;%�H;��H;%�H;��H;A�H;��H;u�H;G�H;�H;��H;�{H;�SH;hH;�LG;��E;�7B;��:;D�,;��;�d�:<!:����0d\��?ݻ�E<�����ټ����mR�����䳽G�l���� ��6��nH��T�      ��"]�Ո�r}���{�ý�u��͕���K�����o�mv���&R�!��T^��d�� <>�"��:|B;f";��4;��>;qD;��F;)�G;*H;�dH;��H;E�H;��H;^�H;a�H;��H;��H;T�H;A�H; �H;@�H;T�H;��H;��H;c�H;]�H;��H;B�H;��H;�dH;*H;&�G;��F;oD;��>;��4;d";zB;&��: @>�f��T^��!���&R�lv���o�����K�͕���u��{�ý��r}�Ո�"]�      �ѽ\ν|�ý䳽=��� M����d�u\8�x��ټlv����Y��_����3��p[� �Y:���:jm;�r-;,�:;��A;boE;�"G;��G;�GH;�sH;�H;��H;�H;]�H;L�H;��H;��H;��H;Z�H;�H;Z�H;��H;��H;��H;M�H;\�H;�H;��H;�H;�sH;�GH;�G;�"G;]oE;��A;,�:;�r-;jm;���:��Y:t[�2������_���Y�lv��ټx��u\8���d� M��=���䳽|�ý\ν      ���������Ȅ�nSt��Y�`n;�3O�t#���Oļ�����&R��_������N3���Y�84:<�:�;@&;�G6;�X?;�D;[xF;�G;e!H;�^H;��H;!�H;�H;s�H;7�H;/�H;�H;C�H;�H;��H;C�H;��H;�H;B�H;�H;2�H;9�H;s�H;�H;!�H;��H;�^H;a!H;�G;WxF;�D;�X?;�G6;@&;�;8�:84:��Y��N3������_��&R������Oļu#��3O�`n;��Y�nSt��Ȅ�����      cn;�|\8��s/�?�!�}��c���nrμ��������E<� ������N3�Hx�X�9 �: _;l ;N2;��<;�B;ղE;`5G;3�G;cFH;�qH;юH;z�H;�H;~�H;��H;��H;0�H;��H;N�H;��H;=�H;��H;N�H;��H;0�H;��H;��H;~�H;�H;z�H;юH;�qH;`FH;1�G;[5G;ղE;�B;��<;N2;m ; _; �:`�9Hx��N3���� ���E<��������nrμb���}��?�!��s/�|\8�      `������o�trμՃ��wv��L"��^N�����?ݻT^��5����Y�H�9�:��:��;m�.;�|:;?A;��D;U�F;߶G;*H;LaH;G�H;��H;�H;m�H;N�H;k�H;��H;+�H;L�H;��H;��H;�H;��H;��H;L�H;+�H;��H;j�H;K�H;h�H;�H;��H;H�H;IaH;*H;ڶG;U�F;��D;?A;�|:;n�.;��;��:�:H�9��Y�5��T^���?ݻ���^N�L"��vv��ԃ��trμ�o����      �����x���#��EF{���]��E<����O�뻦���/d\�d��p[�84:�:��:�[;��,;�8;D!@;�0D;�[F;L{G;#H;sPH;FvH;�H;p�H;.�H;_�H;��H;��H;
�H;�H;��H;��H;��H;��H;��H;��H;��H;�H;�H;��H;��H;Z�H;.�H;o�H;�H;FvH;mPH;H;L{G;�[F;�0D;D!@;	�8;��,;�[;��: �:84:t[�d��-d\�����P�뻥���E<���]�EF{��#���x��      �B(�%�����_������˻�����b�1&����� 8>� �Y:8�: _;�;��,;0`8;��?;�C;�F;GG;v�G; @H;VkH;0�H;6�H;#�H;��H;��H;��H;��H;L�H;��H;�H;��H;��H;��H;��H;��H;�H;��H;M�H;��H;��H;��H;��H;�H;7�H;0�H;SkH;@H;v�G;GG;�F;�C;��?;2`8;��,;��; _;8�: �Y: @>�����/&���b�����˻�����_����%�      ܚ��P���"J���X��$�b���-�����Hx� ��8!:&��:���:�;l ;m�.;�8;��?;�C;��E;c#G;�G;
2H;bH;w�H;��H;��H;ݷH;�H;��H;J�H;h�H;j�H;�H;I�H;��H;k�H;��H;k�H;��H;H�H;�H;j�H;h�H;H�H;��H;�H;ڷH;��H;��H;u�H;bH;
2H;�G;d#G;��E; �C;�?;�8;m�.;o ;�;���:*��:<!:����Hx������-��b��X��"J��T���      0��b��к����|�Y�����s89�5:r/�:�d�:|B;jm;@&;P2;�|:;A!@;�C;��E;�G;�G;�(H;)[H;�zH;m�H;�H;ӳH;��H;��H;��H;��H;��H;+�H;��H;_�H;~�H;/�H;��H;/�H;~�H;_�H;�H;-�H;��H;��H;��H;��H;��H;ӳH;�H;j�H;�zH;)[H;�(H;	�G;�G;��E;�C;A!@;�|:;P2;@&;lm;|B;�d�:x/�:|5:�s89h��d�Y����� к`��      �e9 �9�
�9�:��Y:�y�:�;�:'��:�^;��;d";�r-;�G6;��<;?A;�0D;�F;`#G;�G;%H;�WH;�vH;��H;q�H;y�H;��H;A�H;��H;��H;l�H;�H;��H;��H;\�H;A�H;��H;,�H;��H;@�H;\�H;��H;��H;�H;i�H;��H;��H;?�H;��H;w�H;o�H;��H;�vH;�WH;%H;�G;b#G;�F;�0D;?A;��<;�G6;�r-;d";��;�^;'��:�;�:�y�: �Y:�:�
�9��9      4�:�-�:hg�:(��:��:�^;r�;B�;��#;D�,;��4;)�:;�X?;�B;��D;�[F;GG;�G;�(H;�WH;�uH;��H;E�H;.�H;V�H;-�H;��H;!�H;�H;��H;��H;�H;��H;#�H; �H;��H;��H;��H; �H;#�H;��H;�H;��H;��H;�H;!�H;��H;-�H;U�H;)�H;E�H;��H;�uH;�WH;�(H;�G;GG;�[F;��D;�B;�X?;)�:;��4;D�,;��#;A�;t�;�^;��:2��:hg�:y-�:      ;��;
m;�Z;~`;�%;�+;�0;�G6;��:;��>;��A;�D;ղE;W�F;J{G;v�G;
2H;*[H;�vH;��H;��H;��H; �H;��H;��H;��H;��H;��H;�H;r�H;m�H;��H;��H;��H;��H;�H;��H;��H;��H;��H;m�H;r�H;�H;��H;��H;��H;��H;��H;��H;��H;��H;��H;�vH;+[H;2H;u�G;I{G;X�F;ֲE;�D;��A;��>;��:;�G6;�0;�+;�%;�`;�Z;
m;��;      �Y.;��.;^0;�2;h�4;��7;�|:;O]=;n�?;�7B;sD;boE;ZxF;a5G;߶G;!H;@H;bH;�zH;��H;G�H;��H;~�H;�H;��H;��H;��H;+�H;T�H;��H;��H;��H;��H;}�H;$�H;W�H;�H;U�H;$�H;}�H;��H;��H;��H;��H;S�H;-�H;��H;��H;��H;��H;}�H;��H;B�H;��H;�zH;bH;@H;H;޶G;`5G;ZxF;coE;qD;�7B;n�?;O]=;�|:;��7;r�4;�2;_0;��.;      n�<;/�<;0]=;�O>;��?;��@;�7B;\�C;�D;��E;��F;�"G;�G;5�G;*H;qPH;VkH;|�H;m�H;q�H;)�H;��H;�H;j�H;h�H;o�H;��H;��H;X�H;s�H;2�H;G�H;C�H;�H;z�H;��H;��H;��H;{�H;�H;A�H;H�H;2�H;p�H;V�H;��H;��H;p�H;k�H;j�H;�H;��H;'�H;q�H;m�H;|�H;TkH;qPH;*H;3�G;�G;�"G;��F;��E;�D;\�C;�7B;��@;�?;�O>;3]=;$�<;      �WC;oC;�C;�D;k�D;H5E;�E;�[F;}�F;�LG;)�G;��G;e!H;gFH;OaH;JvH;7�H;��H;�H;~�H;Y�H;��H;��H;o�H;-�H;A�H;{�H;��H;"�H;��H;�H;��H;��H;o�H;��H;�H;�H;�H;��H;m�H;��H;��H;�H;��H;�H;��H;x�H;A�H;0�H;o�H;��H;��H;X�H;��H;�H;��H;4�H;HvH;MaH;dFH;b!H;��G;'�G;�LG;~�F;�[F;�E;I5E;m�D;�D;��C;oC;      9[F;�dF;�F;o�F;�F;�"G;?bG;�G;��G;kH;*H;�GH;�^H;�qH;F�H;�H;6�H;��H;гH;��H;*�H;��H;��H;n�H;:�H;c�H;��H;��H;��H;��H;��H;��H;^�H;��H;�H;M�H;M�H;M�H;�H;��H;[�H;��H;��H;��H;��H;��H;��H;d�H;<�H;n�H;��H;��H;&�H;��H;гH;��H;5�H;�H;F�H;�qH;�^H;�GH;*H;iH;��G;�G;?bG;�"G;�F;p�F;�F;�dF;      �G;��G;��G;��G;,�G;+�G;�H;
*H;+@H;�SH;�dH;�sH;��H;ҎH;��H;q�H;%�H;ڷH;��H;D�H;��H;��H;��H;��H;r�H;��H;��H;z�H;��H;��H;��H;4�H;��H;�H;=�H;p�H;��H;p�H;<�H;�H;��H;4�H;��H;��H;��H;z�H;��H;��H;v�H;��H;��H;��H;��H;D�H;��H;۷H;#�H;p�H;��H;ҎH;��H;�sH;�dH;�SH;.@H;	*H;�H;*�G;1�G;��G;��G; �G;      )0H;�1H;T6H;G=H;7FH;mPH;&[H;fH;�pH;�{H;��H;!�H;#�H;~�H;�H;/�H;��H;�H;��H;��H;!�H;��H;-�H;��H;��H;��H;x�H;��H;��H;��H;9�H;��H;��H;J�H;|�H;��H;��H;��H;|�H;H�H;��H;��H;9�H;��H;��H;��H;x�H;��H;��H;��H;-�H;��H;�H;��H;��H;�H;��H;/�H;�H;|�H;!�H; �H;��H;�{H;�pH;fH;&[H;mPH;CFH;E=H;V6H;�1H;      �jH;*kH;amH;�pH;�uH;9{H;��H;��H;�H;��H;G�H;ŦH;�H;�H;m�H;_�H;��H;��H;��H;��H;�H;��H;Q�H;[�H;�H;��H;��H;��H;��H;'�H;��H;��H;/�H;m�H;��H;��H;��H;��H;��H;m�H;,�H;��H;��H;&�H;��H;��H;��H;��H;�H;\�H;P�H;��H;�H;��H;��H;��H;��H;_�H;k�H;�H;�H;æH;E�H;��H;�H;��H;��H;<{H;�uH;�pH;bmH; kH;      h�H;ԌH;X�H;��H;��H;�H;[�H;U�H;��H;�H;��H;(�H;y�H;��H;Q�H;��H;��H;F�H;��H;o�H;��H;�H;��H;r�H;��H;��H;��H;��H;&�H;��H;��H;6�H;k�H;��H;��H;��H;��H;��H;��H;��H;i�H;7�H;��H;��H;$�H;��H;��H;��H;��H;s�H;��H;�H;��H;o�H;��H;G�H;��H;��H;O�H;��H;y�H;&�H;��H;�H;��H;W�H;[�H;�H;��H;��H;U�H;ьH;      ��H;�H;�H;��H;ԩH;��H;گH;}�H;O�H;O�H;e�H;h�H;>�H;��H;n�H;��H;��H;h�H;��H;�H;��H;t�H;��H;5�H;�H;��H;��H;9�H;��H;��H;/�H;b�H;��H;��H;��H;��H;��H;��H;��H;��H;��H;c�H;/�H;��H;��H;;�H;��H;��H;�H;5�H;��H;t�H;��H;�H;��H;h�H;��H;��H;n�H;��H;>�H;g�H;d�H;O�H;O�H;}�H;گH;��H;ѩH;��H;�H;�H;      еH;�H;ʶH;�H;ƹH;��H;0�H;��H;��H;u�H;i�H;T�H;3�H;��H;��H;�H;S�H;k�H;1�H;��H;�H;q�H;��H;I�H;��H;��H;/�H;��H;��H;6�H;]�H;{�H;��H;��H;��H;��H;��H;��H;��H;��H;��H;|�H;_�H;7�H;��H;��H;1�H;��H;��H;I�H;��H;q�H;�H;��H;1�H;m�H;S�H;�H;��H;��H;3�H;V�H;i�H;u�H;��H;��H;0�H;��H;ĹH;�H;˶H;�H;      `�H;��H;:�H;�H;S�H;��H;~�H;X�H;g�H;��H;��H;��H;�H;6�H;/�H;�H;��H;�H;��H;��H;��H;��H;��H;H�H;��H;\�H;��H;��H;0�H;p�H;��H;��H;��H;��H;��H;��H;��H;��H;��H;��H;��H;��H;��H;q�H;2�H;��H;��H;[�H;��H;F�H;��H;��H;��H;��H;��H;�H;��H;�H;.�H;6�H;�H;��H;��H;��H;h�H;V�H;~�H;��H;L�H;�H;:�H;��H;      ��H;�H;t�H;�H;�H;(�H;��H;�H;��H;E�H;�H;��H;F�H;��H;Q�H;��H;�H;H�H;c�H;c�H;)�H;��H;y�H;�H;e�H;��H;�H;F�H;j�H;��H;��H;��H;��H;��H;��H;��H;��H;��H;��H;��H;��H;��H;��H;��H;m�H;F�H;�H;��H;f�H;�H;y�H;��H;(�H;c�H;c�H;I�H;�H;��H;P�H;��H;F�H;��H;�H;E�H;��H;�H;��H;,�H; �H;�H;t�H;�H;      ��H;��H;�H;��H;t�H;A�H;I�H;q�H;��H; �H;[�H;��H;�H;T�H;��H;��H;��H;��H;�H;H�H;�H;��H; �H;}�H;��H;�H;9�H;{�H;��H;��H;��H;��H;��H;��H;��H;��H;��H;��H;��H;��H;��H;��H;��H;��H;��H;{�H;6�H;�H;��H;{�H; �H;��H;�H;H�H;�H;��H;��H;��H;��H;T�H;�H;��H;Z�H;�H;��H;p�H;I�H;E�H;i�H;��H;�H;��H;      ��H;�H;C�H;��H;^�H;�H;�H;�H;�H;'�H;I�H;e�H;��H;��H;��H;��H;��H;f�H;0�H;��H;��H;��H;T�H;��H;	�H;H�H;m�H;��H;��H;��H;��H;��H;��H;��H;��H;��H;��H;��H;��H;��H;��H;��H;��H;��H;��H;��H;k�H;G�H;�H;��H;T�H;��H;��H;��H;0�H;g�H;��H;��H;��H;��H;��H;e�H;H�H;+�H;�H;�H;�H;�H;S�H;��H;C�H;�H;      ��H;��H;(�H;��H;A�H;��H;��H;��H;��H;��H;�H;*�H;G�H;E�H;�H;��H;��H;��H;��H;1�H;��H;�H;{�H;��H;�H;H�H;��H;��H;��H;��H;��H;��H;��H;��H;��H;��H;��H;��H;��H;��H;��H;��H;��H;��H;��H;��H;��H;J�H;�H;��H;{�H;�H;��H;1�H;��H;��H;��H;��H;�H;E�H;G�H;*�H;�H;��H;��H;��H;��H;��H;5�H;��H;'�H;��H;      ��H;�H;C�H;��H;_�H;�H;�H;�H;�H;(�H;I�H;e�H;��H;��H;��H;��H;��H;f�H;0�H;��H;��H;��H;T�H;��H;�H;H�H;m�H;��H;��H;��H;��H;��H;��H;��H;��H;��H;��H;��H;��H;��H;��H;��H;��H;��H;��H;��H;k�H;H�H;	�H;��H;T�H;��H;��H;��H;0�H;g�H;��H;��H;��H;��H;��H;e�H;I�H;(�H;�H;�H;�H;�H;S�H;��H;A�H;�H;      ��H;��H;�H;��H;t�H;A�H;I�H;s�H;��H;�H;Z�H;��H;�H;T�H;��H;��H;��H;��H;�H;H�H;�H;��H; �H;}�H;��H;�H;7�H;{�H;��H;��H;��H;��H;��H;��H;��H;��H;��H;��H;��H;��H;��H;��H;��H;��H;��H;{�H;6�H;�H;��H;z�H; �H;��H;�H;H�H;�H;��H;��H;��H;��H;T�H;�H;��H;Z�H;�H;��H;p�H;I�H;E�H;j�H;��H;�H;��H;      ��H;�H;t�H;�H;�H;(�H;��H;�H;��H;E�H;�H;��H;F�H;��H;P�H;��H;�H;H�H;c�H;c�H;,�H;��H;y�H;�H;f�H;��H;�H;F�H;j�H;��H;��H;��H;��H;��H;��H;��H;��H;��H;��H;��H;��H;��H;��H;��H;m�H;F�H;�H;��H;e�H;�H;y�H;��H;(�H;c�H;c�H;I�H;�H;��H;P�H;��H;F�H;��H;�H;E�H;��H;�H;��H;,�H;��H;�H;r�H;�H;      b�H;��H;:�H;�H;Q�H;��H;~�H;V�H;h�H;��H;��H;��H;�H;6�H;.�H;�H;��H;�H;��H;��H;��H;��H;��H;F�H;��H;\�H;��H;��H;0�H;p�H;��H;��H;��H;��H;��H;��H;��H;��H;��H;��H;��H;��H;��H;q�H;2�H;��H;��H;[�H;��H;E�H;��H;��H;��H;��H;��H;�H;��H;�H;/�H;6�H;�H;��H;��H;��H;g�H;T�H;~�H;��H;J�H;�H;7�H;��H;      еH;�H;̶H;�H;ǹH;��H;5�H;��H;��H;t�H;h�H;T�H;3�H;��H;��H;�H;S�H;k�H;1�H;��H;�H;q�H;��H;I�H;��H;��H;1�H;��H;��H;6�H;_�H;{�H;��H;��H;��H;��H;��H;��H;��H;��H;��H;|�H;]�H;7�H;��H;��H;/�H;��H;��H;I�H;��H;q�H;�H;��H;1�H;m�H;S�H;�H;��H;��H;3�H;V�H;h�H;u�H;��H;��H;5�H;��H;ĹH;�H;˶H;�H;      ��H;�H;�H;��H;ԩH;��H;گH;}�H;O�H;N�H;e�H;g�H;>�H;��H;n�H;��H;��H;g�H;��H;�H;��H;t�H;��H;6�H;�H;��H;��H;;�H;��H;��H;/�H;b�H;��H;��H;��H;��H;��H;��H;��H;��H;��H;c�H;/�H;��H;��H;9�H;��H;��H;�H;5�H;��H;t�H;��H;�H;��H;h�H;��H;��H;n�H;��H;>�H;h�H;d�H;P�H;O�H;}�H;گH;��H;ѩH;��H;�H;�H;      a�H;ԌH;X�H;��H;��H;�H;^�H;W�H;��H;�H;��H;&�H;y�H;��H;O�H;��H;��H;F�H;��H;p�H;��H;�H;��H;s�H;��H;��H;��H;��H;$�H;��H;��H;6�H;j�H;��H;��H;��H;��H;��H;��H;��H;j�H;7�H;��H;��H;&�H;��H;��H;��H;��H;r�H;��H;�H;��H;o�H;��H;G�H;��H;��H;Q�H;��H;y�H;(�H;��H;�H;��H;X�H;]�H;�H;��H;��H;V�H;ӌH;      �jH;&kH;hmH;�pH;�uH;6{H;��H;��H;�H;��H;G�H;ĦH;�H;�H;k�H;_�H;��H;��H;��H;��H;�H;��H;S�H;\�H;�H;��H;��H;��H;��H;'�H;��H;��H;.�H;m�H;��H;��H;��H;��H;��H;m�H;.�H;��H;��H;&�H;��H;��H;��H;��H;�H;[�H;P�H;��H;�H;��H;��H;��H;��H;a�H;k�H;�H;�H;ŦH;G�H;��H;�H;��H;��H;8{H;�uH;�pH;imH;&kH;      )0H;�1H;T6H;E=H;9FH;mPH;&[H;fH;�pH;�{H;��H; �H;!�H;}�H;�H;/�H;��H;�H;��H;��H;$�H;��H;.�H;��H;��H;��H;x�H;��H;��H;��H;9�H;��H;��H;G�H;{�H;��H;��H;��H;|�H;J�H;��H;��H;9�H;��H;��H;��H;x�H;��H;��H;��H;+�H;��H;�H;��H;��H;�H;��H;1�H;�H;|�H;#�H;!�H;��H;�{H;�pH;fH;&[H;jPH;DFH;G=H;V6H;�1H;      �G; �G;��G;��G;*�G;'�G;�H;	*H;+@H;�SH;�dH;�sH;��H;ҎH;��H;q�H;%�H;ٷH;��H;D�H;��H;��H;��H;��H;v�H;��H;��H;z�H;��H;��H;��H;4�H;��H;�H;<�H;p�H;��H;n�H;=�H;�H;��H;5�H;��H;��H;��H;z�H;��H;��H;r�H;��H;��H;��H;��H;D�H;��H;۷H;#�H;p�H;��H;ҎH;��H;�sH;�dH;�SH;-@H;
*H;�H;'�G;,�G;��G;��G;��G;      ?[F;�dF;%�F;s�F;�F;�"G;?bG;�G;��G;kH;*H;�GH;�^H;�qH;D�H;�H;6�H;��H;гH;��H;,�H;��H;��H;o�H;<�H;c�H;��H;��H;��H;��H;��H;��H;\�H;��H;	�H;M�H;M�H;M�H;�H;��H;[�H;��H;��H;��H;��H;��H;��H;d�H;:�H;l�H;��H;��H;&�H;��H;гH;��H;5�H;�H;F�H;�qH;�^H;�GH;*H;iH;��G;�G;@bG;�"G;�F;p�F;%�F;�dF;      �WC;oC;�C;�D;m�D;H5E;�E;�[F;}�F;�LG;)�G;��G;b!H;dFH;MaH;JvH;5�H;��H;�H;��H;[�H;��H;��H;q�H;0�H;?�H;{�H;��H;"�H;��H;�H;��H;��H;m�H;��H;�H;�H;�H;��H;m�H;��H;��H;�H;��H;�H;��H;x�H;A�H;-�H;o�H;��H;��H;X�H;��H;�H;��H;4�H;JvH;OaH;fFH;e!H;��G;)�G;�LG;}�F;�[F;�E;H5E;k�D;�D;��C;oC;      q�<;-�<;9]=;�O>;��?;��@;�7B;_�C;�D;��E;��F;�"G;�G;3�G;*H;qPH;VkH;y�H;m�H;q�H;+�H;��H;�H;l�H;k�H;o�H;��H;��H;Y�H;s�H;2�H;G�H;B�H;�H;x�H;��H;��H;��H;{�H;�H;B�H;H�H;2�H;p�H;U�H;��H;��H;o�H;h�H;j�H;��H;��H;'�H;q�H;m�H;}�H;TkH;qPH;*H;5�G;�G;�"G;��F;��E;�D;_�C;�7B;��@;	�?;�O>;9]=;"�<;      �Y.;��.;p0;�2;h�4;��7;�|:;O]=;n�?;�7B;qD;coE;XxF;`5G;޶G; H;@H;bH;�zH;��H;H�H;��H;~�H;�H;��H;��H; �H;-�H;T�H;��H;��H;��H;��H;}�H;$�H;W�H;�H;U�H;$�H;}�H;��H;��H;��H;��H;Q�H;+�H;��H;��H;��H;��H;}�H;��H;B�H;��H;�zH;bH; @H;!H;�G;a5G;XxF;coE;qD;�7B;n�?;O]=;�|:;��7;n�4;�2;e0;��.;      ;��;
m;�Z;�`;�%;�+;�0;�G6;��:;��>;��A;�D;ֲE;W�F;J{G;u�G;2H;+[H;�vH;��H;��H;��H; �H;��H;��H;��H;��H;��H;�H;r�H;m�H;��H;��H;��H;��H;�H;��H;��H;��H;��H;m�H;r�H;�H;��H;��H;��H;��H;��H;��H;��H;��H;��H;�vH;*[H;2H;u�G;J{G;X�F;ղE;�D;��A;��>;��:;�G6;�0;�+;�%;�`;�Z;
m;��;      (�:�-�:pg�:2��:��:�^;w�;D�;��#;D�,;��4;)�:;�X?;�B;��D;�[F;GG;�G;�(H;�WH;�uH;��H;G�H;.�H;U�H;,�H;��H;!�H;�H;��H;��H;�H;��H;"�H; �H;��H;��H;��H; �H;#�H;��H;�H;��H;��H;�H;!�H;��H;-�H;V�H;)�H;D�H;��H;�uH;�WH;�(H;�G;GG;�[F;��D;�B;�X?;)�:;��4;B�,;��#;D�;t�;�^;��:,��:pg�:s-�:      �e90�9�
�9�:��Y:�y�:�;�:+��:�^;��;d";�r-;�G6;��<;?A;�0D;�F;`#G;�G;%H;�WH;�vH;��H;s�H;w�H;��H;A�H;��H;��H;l�H;�H;��H;��H;\�H;@�H;��H;,�H;��H;A�H;\�H;��H;��H;�H;i�H;��H;��H;?�H;��H;y�H;m�H;��H;�vH;�WH;%H;�G;b#G;�F;�0D;?A;��<;�G6;�r-;b";��;�^;-��:�;�:�y�:�Y:�:�
�9��9      0��b�� к����t�Y�����s89�5:r/�:�d�:|B;jm;@&;P2;�|:;A!@;�C;��E;�G;�G;�(H;)[H;�zH;n�H;�H;ҳH;��H;��H;��H;��H;��H;+�H;��H;_�H;~�H;/�H;��H;/�H;~�H;_�H;�H;-�H;��H;��H;��H;��H;��H;ԳH;�H;i�H;�zH;)[H;�(H;	�G;�G;��E;�C;A!@;�|:;N2;@&;jm;|B;�d�:x/�:�5:�s89p��`�Y����� к`��      ܚ��P���"J���X��$�b���-�����Hx����<!:&��:���:�;l ;m�.;�8;��?;�C;��E;c#G;�G;
2H;bH;w�H;��H;��H;ݷH;�H;��H;J�H;h�H;h�H;�H;H�H;��H;k�H;��H;k�H;��H;I�H;�H;k�H;h�H;H�H;��H;�H;ڷH;��H;��H;u�H;bH;
2H;�G;d#G;��E; �C;�?;�8;m�.;l ;�;���:&��:8!:����Hx������-��b��X��"J��T���      �B(�%�����_������˻�����b�1&����� 8>� �Y:8�: _;��;��,;2`8;��?;�C;�F;GG;v�G; @H;WkH;0�H;6�H;#�H;��H;��H;��H;��H;M�H;��H;�H;��H;��H;��H;��H;��H;�H;��H;M�H;��H;��H;��H;��H;�H;6�H;0�H;RkH;@H;v�G;GG;�F;�C;��?;0`8;��,;�; _;8�: �Y: 8>�����0&���b�����˻�����_����%�      �����x���#��EF{���]��E<����O�뻦���-d\�d��p[�84:�:��:�[;��,;�8;D!@;�0D;�[F;L{G; H;qPH;FvH;�H;q�H;.�H;^�H;��H;��H;
�H;�H;��H;��H;��H;��H;��H;��H;��H;�H;�H;��H;��H;Z�H;.�H;m�H;�H;FvH;oPH;H;L{G;�[F;�0D;D!@;	�8;��,;�[;��:�:84:p[�d��/d\�����N�뻥���E<���]�EF{��#���x��      `������o�trμԃ��wv��L"��^N�����?ݻT^��5����Y�H�9�:��:��;l�.;�|:;?A;��D;U�F;߶G;*H;IaH;G�H;��H;�H;m�H;M�H;j�H;��H;-�H;L�H;��H;��H;�H;��H;��H;M�H;+�H;��H;k�H;M�H;j�H;�H;��H;G�H;LaH;*H;ڶG;U�F;��D;?A;�|:;n�.;��;��:�:@�9��Y�5��T^���?ݻ���^N�L"��vv��ԃ��trμ�o����      cn;�|\8��s/�?�!�}��c���nrμ��������E<� ������N3�Hx�`�9 �: _;l ;N2;��<;�B;ղE;`5G;3�G;`FH;�qH;ҎH;z�H;�H;~�H;��H;��H;2�H;��H;N�H;��H;=�H;��H;N�H;��H;/�H;��H;��H;~�H;�H;z�H;ώH;�qH;cFH;1�G;[5G;ղE;�B;��<;N2;o ; _; �:X�9Hx��N3���� ���E<��������nrμb���}��?�!��s/�|\8�      ���������Ȅ�nSt��Y�`n;�3O�t#���Oļ�����&R��_������N3���Y�44:<�:�;@&;�G6;�X?;�D;[xF;�G;a!H;�^H;��H;!�H;�H;s�H;9�H;0�H;�H;B�H;�H;��H;C�H;��H;�H;C�H;�H;/�H;7�H;s�H;��H;!�H;��H;�^H;e!H;�G;WxF;�D;�X?;�G6;@&;�;8�:84:��Y��N3������_��&R������Oļt#��3O�`n;��Y�nSt��Ȅ�����      �ѽ\ν|�ý䳽=��� M����d�u\8�x��ټlv����Y��_����1��t[� �Y:���:jm;�r-;)�:;��A;`oE;�"G;�G;�GH;�sH;�H;��H;�H;\�H;J�H;��H;��H;��H;[�H;�H;[�H;��H;��H;��H;M�H;]�H;�H;��H;�H;�sH;�GH;��G;�"G;]oE;��A;,�:;�r-;jm;���:��Y:x[�2������_���Y�lv��ټx��u\8���d� M��=���䳽|�ý\ν      ��"]�Ո�r}���{�ý�u��͕���K�����o�mv���&R�!��T^��f�� <>�$��:zB;f";��4;��>;qD;��F;&�G;*H;�dH;��H;E�H;��H;]�H;a�H;��H;��H;T�H;@�H; �H;A�H;T�H;��H;��H;c�H;^�H;��H;B�H;��H;�dH;*H;)�G;��F;oD;��>;��4;e";|B;&��: D>�h��T^��!���&R�mv���o�����K�͕���u��{�ý��r}�Ո�"]�      �+X��T��nH��6��� �l��G�䳽�����mR����ټ�����E<��?ݻ0d\�����0!:�d�:��;B�,;��:;�7B;��E;�LG;iH;�SH;�{H;��H;�H;G�H;t�H;��H;A�H;��H;%�H;��H;%�H;��H;B�H;��H;r�H;G�H;�H;��H;�{H;�SH;iH;�LG;��E;�7B;��:;B�,;��;�d�:<!:����0d\��?ݻ�E<�����ټ����mR�����䳽G�l���� ��6��nH��T�      㰖��������*|�OS\�� :����Z�o$�������K�x���Oļ����������0&� ��r/�:�^;��#;�G6;m�?;�D;z�F;��G;*@H;�pH;�H;��H;E�H;��H;`�H;��H;��H;	�H;��H;	�H;��H;��H;]�H;��H;E�H;��H;�H;�pH;)@H;��G;~�F;�D;k�?;�G6;��#;�^;r/�:���3&������������Oļx���K�����o$���Z���� :�PS\��*|�������      C�;9ɾ㼾B�������Mw��nH�����Z�䳽͕��u\8�t#������^N�N����b��Hx��5:3��:A�; �0;O]=;^�C;�[F;�G;*H;fH;��H;M�H;r�H;��H;M�H;�H;c�H; �H;��H;�H;b�H;�H;K�H;��H;t�H;M�H;��H;fH;*H;�G;�[F;[�C;O]=; �0;D�;1��:�5:�Hx���b�N��^N�����t#��u\8�͕��䳽�Z񽳯��nH��Mw�����B��㼾9ɾ      1y��v�m���E�߾����D��A����nH���Gὠu����d�3O�nrμL"����� 	�����`s89�;�:n�;�+;�|:;�7B;�E;>bG;�H; [H;��H;S�H;ϯH;+�H;z�H;{�H;<�H;�H;��H;�H;<�H;{�H;w�H;,�H;ϯH;Q�H;��H; [H;�H;>bG;�E;�7B;�|:;�+;q�;�;�:`s89���	�����L"��nrμ3O���d��u��G����nH�A���D������E�߾m����v�      �O/�rM+�Z�����JW��9ɾD���Mw�� :�l��{�ý M��`n;�d���wv���E<��˻��-�����y�:�^;�%;��7;��@;C5E;�"G;)�G;lPH;:{H;�H;��H;��H;��H;)�H;D�H;�H;��H;�H;D�H;+�H;��H;��H;��H;�H;8{H;lPH;'�G;�"G;E5E;��@;��7;�%;�^;�y�:�����-��˻�E<�wv��d���`n;� M��{�ýl��� :��Mw�D��9ɾJW�����Z��rM+�      :�X�YvS�9E��O/��S�KW����������OS\��� ���=����Y�~��ԃ����]�����"�b�h�Y���Y:��:~`;n�4;��?;h�D;�F;(�G;7FH;�uH;�H;éH;��H;F�H;��H;U�H;L�H;,�H;L�H;U�H;��H;D�H;��H;éH;�H;�uH;7FH;)�G;�F;j�D;��?;p�4;~`;��:��Y:`�Y�!�b�������]�ԃ��~���Y�=����彔� �OS\���������KW���S��O/�9E�YvS�      � ����y�c�h��N��O/����E�߾B���*|��6�s}�䳽nSt�@�!�urμGF{��_��X�������:4��:[;�2;�O>;�D;q�F;��G;J=H;�pH;��H;}�H;�H;�H;�H;��H;��H;��H;��H;��H;�H;�H;�H;�H;��H;�pH;J=H;��G;q�F;�D;�O>;�2;[;<��:�:�����X���_�GF{�urμ@�!�nSt�䳽s}��6��*|�B��E�߾����O/��N�c�h���y�      ?v��c���X ��c�h�9E�Z��m���㼾���nH�Ո�}�ý�Ȅ��s/��o��#�����%J��к�
�9\g�:�l;^0;+]=;�C;'�F;��G;O6H;dmH;N�H;إH;��H;/�H;u�H;�H;7�H;�H;8�H;�H;u�H;-�H;��H;إH;K�H;amH;M6H;��G;%�F;�C;']=;a0;�l;`g�:�
�9к%J������#���o��s/��Ȅ�}�ýՈ��nH���㼾m���Z��9E�c�h�X ��c���      ~h��1���c�����y�YvS�rM+��v�9ɾ�����T�"]�\ν����|\8�����x��%�P���`�뺠�9u-�:}�;��.;%�<;oC;�dF;��G;�1H;(kH;ΌH;ڤH;�H;��H;�H;��H;��H;��H; �H;��H;�H;��H;�H;ڤH;̌H;%kH;�1H;��G;�dF;oC;"�<;��.;}�;y-�:��9b��P���%��x�����|\8�����\ν#]��T�����9ɾ�v�rM+�YvS���y�c���1���      IEb�c]��N���7����v� ���˾��,�j��!,�t���O��Jm�/��=,˼Ūx�]���1��������:s�:�;P�1;@,>;��C;�wF;�G;� H;?H;�hH;b�H;��H;L�H;,�H;��H;<�H;��H;>�H;��H;,�H;J�H;��H;b�H;�hH;?H;� H;�G;�wF;��C;=,>;T�1;�;w�:��:�����1��^��Ūx�=,˼/��Jm�O��t����!,�,�j�����˾v� ������7��N�c]�      c]�g�W��TI�v3� E�������Ǿy����f�:)�*��w;���Fi��k���Ǽ�[t�O�	�.Ȅ�X��d�:
��:��;dJ2;\Z>;S	D;�F;P�G;&H;�?H;�iH;��H;�H;��H;I�H;��H;h�H;��H;h�H;��H;I�H;��H;�H;��H;�iH;�?H;&H;P�G;�F;T	D;YZ>;jJ2;��;��:\�:X��-Ȅ�P�	��[t���Ǽ�k��Fi�w;��*��:)��f�y�����Ǿ���� E�v3��TI�g�W�      �N��TI���;�1�'�l��쾂���z󐾶Z��K ��s�D����&^���"����g����ըu�� ��X3<:��:;qg3;��>;�BD;F;��G;�H;YBH;�kH;d�H;�H;<�H;�H;~�H;��H;V�H;��H;}�H;�H;;�H;�H;d�H;�kH;UBH;�H;��G;��F;�BD;��>;tg3;;!��:P3<:� ��Ԩu������g��"����&^�D����s潨K ��Z�z󐾂�����l�1�'���;��TI�      ��7�v3�1�'����v� ��{Ծ"���J���|�F�����ӽ���c�L�Nv��뮼VT����PV�t�=��)i:~��:�z ;�$5;��?;�D;ٺF;�G;�H;�FH;�nH;��H;��H;�H;�H;F�H;e�H;�H;e�H;F�H;�H;~�H;��H;��H;�nH;�FH;�H;�G;ٺF;�D;��?;�$5;�z ;���:�)i:x�=��PV���VT��뮼Mv�c�L�����ӽ���|�F�J���"����{Ծv� ����1�'�v3�      ��� E�l�v� �Y�ݾm���X͓��f��>/�����'���섽T�6��t�w��b�:�'Tʻ~.��ڷ��t�:�;��$;�Y7;d�@;
E;)�F;F�G;�H;JLH;�rH;��H;ڤH;1�H;,�H;@�H;X�H;��H;V�H;?�H;,�H;0�H;ۤH;��H;�rH;HLH;�H;G�G;)�F;
E;a�@;�Y7;��$;�;�t�:�ڷ�}.�(Tʻb�:�w���t�T�6��섽�'������>/��f�X͓�m���Y�ݾv� �l� E�      u� ��������{Ծm���x���^�x��SC��^���޽C���}�e�+��H�Ѽ)G������R������ߤ8��:�Y;^�);��9;
�A;ȄE;�G;+�G;u!H;NSH;�wH;��H;��H;N�H;��H;��H;��H;��H;��H;��H;��H;N�H;��H;��H;�wH;ISH;u!H;*�G;�G;ȄE;�A;��9;^�);�Y;��:�ߤ8����R�����)G��H�Ѽ+��}�e�C�����޽�^��SC�^�x�x���m����{Ծ�쾤���      ��˾��Ǿ����"���X͓�^�x���J��K �r���!������?����뮼0�[�#���3|��W����:��:�';{/;rg<;�C;zF;�NG;��G;<-H;|[H;�}H;ӗH;֪H;ɸH;��H;	�H;��H;�H;��H;	�H;��H;ɸH;تH;ӗH;�}H;y[H;<-H;��G;�NG;wF;�C;rg<;|/;�';��:��:�W��3|�#���0�[��뮼���?����!��r����K ���J�^�x�X͓�"���������Ǿ      ��y���z�J����f��SC��K �rn���Ž����Z��k�$}ռ0X��ey-�/���i.�H���P�:�+�:��;+4;D�>;D;�wF;@�G;��G;�9H;edH;��H;��H;n�H;|�H;��H;��H;_�H;|�H;_�H;��H;��H;{�H;p�H;��H;��H;bdH;�9H;��G;@�G;�wF;D;E�>;,4;��;�+�:�P�:8��i.�.���ey-�0X��$}ռ�k��Z�����Žsn���K ��SC��f�J���z�y���      ,�j��f��Z�|�F��>/��^�r����ŽI ���Fi��Q+��t�sT��t�W�����1��Ⱥ�X�9�P�:�Y;��(;�8;	A;�E;�F;x�G;�H;�FH;�mH;��H;ΡH;M�H;z�H;��H;��H;�H; �H;�H;��H;��H;z�H;N�H;͡H;��H;�mH;�FH;�H;x�G;�F;�E;	A;�8;��(;�Y;�P�:�X�9Ⱥ�1�����t�W�sT���t�Q+��Fi�I ���Žr����^��>/�|�F��Z��f�      �!,�;)��K ���������޽!������Fi��0����鷼��x�����.��N�(����8+i:���:N�;��0;Z�<;�C;��E;=G;
�G;%H;pTH;�wH;��H;#�H;[�H;��H;L�H;��H;��H;��H;��H;��H;L�H;��H;\�H;#�H;��H;�wH;pTH;%H;�G;=G;��E;�C;\�<;��0;N�;���:@+i:���O�(��.�������x�鷼����0��Fi����!����޽�������K �;)�      t���)��s��ӽ�'��C�������Z��Q+�����"�� G��Ļ0���׻˕b�*W��pY�9::`;�*';�Y7;$@;8�D;�F;%�G;��G;E8H;bH;�H;f�H;��H;��H;��H;��H;��H;\�H;H�H;\�H;��H;��H;��H;��H;��H;f�H;	�H;bH;D8H;��G;"�G;�F;5�D;$@;�Y7;�*';:`;���:hY�9(W��˕b���׻Ļ0� G���"������Q+��Z����C����'���ӽ�s�)��      O��w;��D�������섽}�e��?��k��t�鷼 G���e7���� Ȅ�d0���t�Fu�:",�:�;�1;d�<;s�B;7�E;G;�G;oH;�JH;koH;�H;��H;"�H;��H;��H;,�H;��H;�H;��H;�H;��H;+�H;��H;��H;"�H;��H;�H;koH;JH;mH; �G;G;5�E;s�B;d�<;�1;�;*,�:Du�: �t�f0� Ȅ���껈e7� G��鷼�t��k��?�}�e��섽���D���w;��      Jm��Fi��&^�c�L�T�6�+����$}ռsT����x�Ļ0���������@ط�,o`:��:+�;8�*;L�8;�@;I�D;x�F;~G;��G;�1H;�[H;}|H;ΕH;�H;��H;��H;��H;��H;��H;��H;��H;��H;��H;��H;��H;��H;��H;�H;˕H;}|H;�[H;�1H;��G;�}G;t�F;I�D;!�@;J�8;9�*;/�;��:0o`:8ط���������Ļ0���x�rT��$}ռ��+��T�6�c�L��&^��Fi�      /���k��Mv��t�H�Ѽ�뮼0X��s�W������׻�Ǆ������45<:}��:�Y;�t%;%5;�Z>;aC;��E;E*G;v�G;$H;HH;}lH;�H;�H;үH;߼H;��H;��H;�H;��H;}�H;=�H;}�H;��H;�H;��H;��H;�H;ЯH;�H;�H;zlH;HH;#H;q�G;@*G;��E;aC;�Z>;%5;�t%;�Y;}��:<5<:������Ǆ���׻���r�W�0X���뮼G�Ѽ�t�Mv���k�      <,˼��Ǽ�"���뮼w��(G��0�[�fy-�����.��˕b�h0�Hط�45<:M�:�\;��!;�J2;�g<;_0B;=CE;<�F;^�G;�G;�4H;�\H;|H;��H;��H;i�H;��H;O�H;��H;^�H;`�H;�H;��H;�H;a�H;_�H;��H;R�H;��H;f�H;��H;��H;|H;�\H;�4H; �G;W�G;<�F;<CE;a0B;�g<;�J2;��!;�\;M�:45<:Hط�h0�˕b��.�����fy-�0�[�(G��w���뮼�"����Ǽ      Īx��[t���g�UT�b�:���� ���0����1��N�(�,W����t�,o`:{��:�\;{ ;��0;m;;=A;(�D;�wF;�cG;d�G;�!H;�MH;�oH;��H;��H;ԯH;��H;u�H;��H;j�H;}�H;�H;��H;4�H;��H;�H;|�H;h�H;��H;t�H;��H;ϯH;��H;��H;�oH;�MH;�!H;`�G;�cG;�wF;(�D;=A;o;;��0;{ ;�\;}��:,o`:��t�,W��M�(��1��0��� ������b�:�UT���g��[t�      ]��L�	������)Tʻ�R��3|�h.�Ⱥ���xY�9Du�:��:�Y;��!;��0;��:;��@;CD;�2F;�8G;��G;�H;y@H;5dH;ԀH;��H;U�H;Y�H;\�H;��H; �H;��H;}�H;��H;�H;��H;�H;��H;}�H;��H;�H;��H;[�H;U�H;T�H;��H;րH;5dH;u@H;�H;��G;�8G;�2F;CD;ŵ@;��:;��0;��!;�Y;��:Fu�:hY�9���Ⱥj.�3|��R��'Tʻ�����O�	�      �1��-Ȅ�Шu��PV��.�����W��P��X�98+i:���:",�:+�;�t%;�J2;k;;��@;~D;F;9G;��G;�H;�5H;�ZH;ExH;P�H;:�H;'�H;%�H;h�H;~�H;*�H;?�H;9�H;M�H;i�H;��H;i�H;M�H;7�H;>�H;,�H;|�H;h�H;!�H;(�H;9�H;P�H;CxH;�ZH;�5H;�H;��G;9G;F;D;��@;k;;�J2;�t%;+�;",�:���:@+i:�X�9`��W�����y.��PV�Шu�2Ȅ�      楥�X��� ��p�=� ۷��ߤ8��:�P�:�P�:���::`;�;7�*;%5;�g<;=A;CD;F;�G;��G;v�G;�-H;*SH;iqH;��H;НH;��H;%�H;J�H;�H;�H;��H;d�H;��H;��H;��H;��H;��H;��H;��H;b�H;��H;�H; �H;H�H;'�H;��H;ҝH;�H;eqH;&SH;�-H;s�G;��G;�G; F;CD;=A;�g<;%5;7�*;�;:`;���:�P�:�P�:��:`�8�ڷ�l�=�� ��X��      ��:��:d3<:�)i:�t�:��:��:�+�:�Y;N�;�*';�1;H�8;�Z>;_0B;"�D;�2F;6G;��G;+�G;�)H;�NH;�lH;[�H;w�H;��H;��H;?�H;��H;�H;I�H;;�H;B�H;k�H;��H;��H;��H;��H;��H;k�H;B�H;<�H;J�H;�H;��H;?�H;��H;��H;w�H;W�H;�lH;�NH;�)H;-�G;��G;6G;�2F;"�D;_0B;�Z>;H�8;�1;�*';N�;�Y;�+�:��:��:�t�:�)i:d3<:��:      ��:(��:1��:r��:�;�Y;�';��;��(;��0;�Y7;b�<;�@;aC;<CE;�wF;�8G;��G;w�G;�)H;�LH;jH;F�H;m�H;��H;�H;̾H;t�H;7�H;��H;&�H;g�H;��H;��H;��H;��H;��H;��H;��H;��H;��H;h�H;&�H;��H;5�H;u�H;̾H;�H;��H;j�H;D�H;jH;�LH;�)H;w�G;��G;�8G;�wF;;CE;aC;�@;b�<;�Y7;��0;��(;��;�';�Y;�;v��:-��:��:      �;��;;�z ;��$;h�);�/;54;�8;]�<;"$@;t�B;J�D;��E;=�F;�cG;��G;�H;�-H;�NH;jH;Z�H;ƔH;��H;�H;ѼH;��H;��H;]�H;�H;��H;B�H;^�H;��H;��H;~�H;��H;~�H;��H;��H;\�H;B�H;��H;��H;Y�H;��H;��H;ԼH;�H;��H;ÔH;Z�H;jH;�NH;�-H;�H;��G;�cG;>�F;��E;J�D;v�B; $@;^�<;�8;24;�/;i�);��$;�z ;;��;      X�1;hJ2;rg3;�$5;�Y7;��9;vg<;G�>;A;�C;8�D;9�E;w�F;E*G;]�G;c�G;�H;�5H;*SH;�lH;F�H;ǔH;<�H;�H;��H;}�H;u�H;G�H;�H;��H;��H;��H;��H;��H;��H;>�H;��H;>�H;��H;��H;��H;��H;��H;��H;�H;G�H;q�H;~�H;��H;�H;;�H;ǔH;C�H;�lH;*SH;�5H;�H;b�G;\�G;E*G;w�F;9�E;8�D;�C;A;E�>;xg<;��9;�Y7;�$5;ug3;YJ2;      R,>;fZ>;�>;��?;d�@;�A;�C;	D;�E;��E;	�F;G;�}G;t�G;�G;�!H;w@H;�ZH;hqH;[�H;i�H;��H;�H;0�H;��H;��H;`�H;*�H;�H;�H;~�H;M�H;��H;��H;x�H;��H;�H;��H;y�H;��H;��H;O�H;|�H;�H;�H;*�H;]�H;��H;��H;-�H;�H;��H;g�H;\�H;hqH;�ZH;u@H;�!H;�G;t�G;�}G;G;�F;��E;�E;	D;�C;�A;k�@;��?;�>;ZZ>;      ��C;Z	D;rBD;�D;
E;˄E;wF;�wF;�F;=G;"�G;�G;��G;'H;�4H;�MH;;dH;FxH;��H;~�H;��H;�H;��H;��H;_�H;�H;��H;��H;��H;��H;��H;��H;��H;q�H;�H;s�H;}�H;s�H;�H;o�H;��H;��H;��H;��H;��H;��H;��H;�H;_�H;��H;��H;�H;��H;��H;��H;IxH;8dH;�MH;�4H;'H;��G;�G;"�G;=G;�F;�wF;wF;̈́E;
E;�D;rBD;[	D;      �wF;�F;��F;׺F;)�F;�G;�NG;;�G;x�G;
�G;��G;pH;�1H;HH;�\H;�oH;ӀH;O�H;͝H;��H;�H;ѼH;z�H;��H;
�H;��H;Q�H;L�H;��H;��H;I�H;��H;g�H;*�H;��H;��H;��H;��H;��H;*�H;d�H;��H;I�H;��H;��H;L�H;O�H;��H;�H;��H;z�H;ѼH;ݳH;��H;͝H;O�H;ӀH;�oH;�\H;HH;�1H;pH;��G;�G;y�G;;�G;�NG;�G;0�F;ٺF;��F;�F;      �G;Q�G;��G;�G;G�G;/�G;��G;��G;�H;%H;G8H;�JH;�[H;|lH;|H;��H;��H;7�H;��H;��H;ϾH;��H;t�H;b�H;��H;T�H;6�H;��H;|�H;*�H;i�H;D�H;�H;��H;�H;9�H;G�H;9�H;�H;��H;�H;B�H;i�H;(�H;{�H;��H;3�H;S�H;��H;a�H;r�H;��H;̾H;��H;��H;9�H;��H;��H;|H;|lH;�[H;�JH;G8H; %H;�H;��G;��G;-�G;N�G;�G;��G;S�G;      � H;'H;�H;�H;�H;u!H;@-H;�9H; GH;vTH;bH;qoH;~|H;�H;��H;��H;T�H;$�H;$�H;B�H;t�H;��H;I�H;-�H;��H;N�H;��H;��H;�H;:�H;:�H;�H;��H;�H;M�H;��H;��H;��H;M�H;�H;��H;�H;:�H;7�H;	�H;��H;��H;N�H;��H;-�H;G�H;��H;r�H;B�H;$�H;$�H;S�H;��H;��H;�H;}|H;qoH;bH;uTH;GH;�9H;@-H;s!H;�H;�H;�H;1H;      ?H;�?H;UBH;�FH;HLH;KSH;�[H;hdH;�mH;�wH;�H;�H;ΕH;�H;��H;ԯH;Z�H;!�H;I�H;��H;7�H;[�H;�H;�H;��H;��H;y�H;�H;V�H;(�H;��H;��H;�H;l�H;��H;��H;��H;��H;��H;l�H;�H;��H;��H;&�H;V�H;�H;y�H;��H;��H;�H;�H;\�H;5�H;��H;I�H;"�H;Y�H;ԯH;��H;�H;ΕH;�H;	�H;�wH;�mH;gdH;�[H;LSH;OLH;�FH;UBH;�?H;      iH;�iH;�kH;�nH;�rH;�wH;�}H;��H;��H;��H;n�H;ʡH;�H;ٯH;k�H;��H;_�H;d�H;��H; �H;��H;��H;��H;�H;��H;��H;'�H;9�H;&�H;�H;��H;�H;Z�H;��H;��H;��H;��H;��H;��H;��H;U�H;�H;��H;�H;%�H;7�H;$�H;��H;��H;�H;��H; �H;��H; �H;��H;e�H;]�H;��H;k�H;ׯH;�H;ɡH;n�H;��H;��H;��H;�}H;�wH;�rH;�nH;�kH;�iH;      g�H;�H;q�H;��H;ЏH;��H;ݗH;ÜH;סH;*�H;��H;.�H;��H;�H;��H;|�H;��H;~�H;�H;P�H;*�H;��H;��H;�H;��H;L�H;f�H;;�H;��H;��H;�H;h�H;��H;��H;�H; �H; �H; �H;�H;��H;��H;i�H;�H;��H;��H;;�H;f�H;I�H;��H;��H;��H;��H;'�H;N�H;�H;|�H;��H;{�H;��H;�H;��H;,�H;��H;*�H;סH;H;ݗH;��H;͏H;��H;r�H;	�H;      ��H;��H;��H;��H;ߤH;��H;٪H;w�H;Q�H;\�H;��H;��H;��H;��H;V�H;��H;�H;,�H;��H;B�H;k�H;F�H;��H;P�H;��H;��H;B�H;�H;��H;�H;c�H;��H;��H;�H;�H;<�H;X�H;<�H;�H;�H;��H;��H;e�H;�H;��H;�H;A�H;��H;��H;Q�H;��H;D�H;j�H;B�H;��H;-�H;�H;��H;U�H;��H;��H;��H;��H;\�H;R�H;u�H;ڪH;��H;ޤH;��H;��H;��H;      S�H;��H;F�H;��H;;�H;N�H;͸H;��H;��H;��H;��H;��H;��H;��H;��H;n�H;��H;;�H;f�H;H�H;��H;]�H;��H;��H;��H;h�H;�H;��H;�H;_�H;��H;��H;�H;0�H;U�H;J�H;=�H;J�H;U�H;/�H;�H;��H;��H;_�H;�H;��H;�H;e�H;��H;��H;��H;\�H;��H;I�H;f�H;<�H;��H;n�H;��H;��H;��H;��H;��H;��H;��H;��H;͸H;R�H;4�H;��H;G�H;��H;      <�H;X�H;�H;��H;7�H;��H;��H;��H;��H;N�H;��H;2�H;��H;�H;c�H;��H;��H;9�H;��H;r�H;��H;��H;��H;��H;g�H;)�H;��H;�H;i�H;��H;��H;�H;(�H;=�H;g�H;u�H;T�H;u�H;g�H;=�H;'�H;	�H;��H;��H;m�H;�H;��H;&�H;j�H;��H;��H;��H;��H;r�H;��H;:�H;��H;��H;c�H;�H;��H;2�H;��H;N�H;��H;��H;��H;��H;-�H;��H;�H;P�H;      ��H;�H;��H;N�H;\�H;��H;�H;��H;��H;��H;��H;��H;��H;��H;g�H;�H;��H;J�H;��H;��H;��H;��H;��H;{�H;�H;��H;��H;L�H;��H;��H;�H;�H;R�H;j�H;M�H;j�H;��H;j�H;M�H;j�H;O�H; �H;�H;��H;��H;L�H;��H;��H;�H;y�H;��H;��H;��H;��H;��H;L�H;��H;�H;e�H;��H;��H;��H;��H;��H;��H;��H;�H;��H;Q�H;P�H;��H;�H;      8�H;r�H;��H;i�H;j�H;��H;��H;m�H;�H;��H;d�H;&�H;��H;��H;!�H;��H;�H;d�H;��H;��H;��H;~�H;=�H;��H;l�H;��H;6�H;��H;��H;��H;�H;?�H;G�H;x�H;j�H;b�H;q�H;b�H;j�H;t�H;F�H;A�H;�H;��H;��H;��H;5�H;��H;n�H;��H;=�H;~�H;��H;��H;��H;f�H;�H;��H;!�H;��H;��H;&�H;c�H;��H;�H;j�H;��H;��H;]�H;i�H;��H;h�H;      ��H;��H;g�H;�H;��H;��H;�H;��H;	�H;��H;O�H;��H;��H;F�H;��H;:�H;��H;��H;��H;��H;��H;��H;��H;�H;u�H;��H;D�H;��H;��H;�H; �H;]�H;<�H;X�H;��H;r�H;_�H;r�H;��H;X�H;9�H;_�H; �H;�H;��H;��H;C�H;��H;u�H;
�H;��H;��H;��H;��H;��H;��H;��H;:�H;��H;F�H;��H;��H;O�H;��H;�H;��H;�H;��H;��H;�H;g�H;��H;      8�H;r�H;��H;j�H;k�H;��H;��H;m�H;�H;��H;d�H;&�H;��H;��H;!�H;��H;�H;d�H;��H;��H;��H;~�H;=�H;��H;n�H;��H;6�H;��H;��H;��H;�H;?�H;G�H;x�H;j�H;b�H;q�H;b�H;j�H;u�H;F�H;A�H;�H;��H;��H;��H;5�H;��H;l�H;��H;=�H;~�H;��H;��H;��H;f�H;�H;��H;!�H;��H;��H;&�H;d�H;��H;�H;j�H;��H;��H;_�H;i�H;��H;h�H;      ��H;�H;��H;P�H;\�H;��H;�H;��H;��H;��H;��H;��H;��H;��H;e�H;�H;��H;J�H;��H;��H;��H;��H;��H;{�H;�H;��H;��H;L�H;��H;��H;�H;�H;R�H;j�H;M�H;j�H;��H;j�H;M�H;j�H;O�H;!�H;�H;��H;��H;L�H;��H;��H;�H;x�H;��H;��H;��H;��H;��H;L�H;��H;�H;e�H;��H;��H;��H;��H;��H;��H;��H;�H;��H;Q�H;N�H;��H;�H;      >�H;X�H;�H;��H;7�H;��H;��H;��H;��H;N�H;��H;2�H;��H;�H;c�H;��H;��H;9�H;��H;q�H;��H;��H;��H;��H;j�H;'�H;��H;�H;j�H;��H;��H;�H;(�H;=�H;g�H;u�H;T�H;t�H;g�H;=�H;'�H;	�H;��H;��H;l�H;�H;��H;)�H;g�H;��H;��H;��H;��H;r�H;��H;:�H;��H;��H;c�H;�H;��H;2�H;��H;N�H;��H;��H;��H;��H;,�H;��H;�H;P�H;      V�H;��H;G�H;��H;:�H;O�H;͸H;��H;��H;��H;��H;��H;��H;��H;��H;n�H;��H;;�H;f�H;H�H;��H;\�H;��H;��H;��H;g�H;�H;��H;�H;_�H;��H;��H;�H;.�H;U�H;J�H;=�H;J�H;U�H;/�H;�H;��H;��H;a�H;�H;��H;�H;g�H;��H;��H;��H;]�H;��H;I�H;f�H;;�H;��H;n�H;��H;��H;��H;��H;��H;��H;��H;��H;͸H;T�H;1�H;��H;D�H;��H;      ��H; �H;��H;��H;�H;��H;ߪH;x�H;R�H;\�H;��H;��H;��H;��H;U�H;��H;�H;,�H;��H;C�H;n�H;D�H;��H;Q�H;��H;��H;A�H;�H;��H;�H;e�H;��H;��H;�H;�H;<�H;X�H;<�H;�H;�H;��H;��H;c�H;�H;��H;�H;A�H;��H;��H;P�H;��H;F�H;j�H;B�H;��H;-�H;�H;��H;U�H;��H;��H;��H;��H;]�H;T�H;u�H;ݪH;��H;ޤH;��H;��H;��H;      g�H;�H;q�H;��H;ЏH;��H;ݗH;ÜH;סH;)�H;��H;,�H;��H;�H;��H;|�H;��H;{�H;�H;N�H;,�H;��H;��H;��H;��H;J�H;f�H;;�H;��H;��H;�H;h�H;��H;��H;�H; �H; �H;�H;�H;��H;��H;i�H;�H;��H;��H;;�H;f�H;J�H;��H;�H;��H;��H;'�H;P�H;�H;~�H;��H;|�H;��H;�H;��H;.�H;��H;,�H;סH;ÜH;ݗH;��H;͏H;��H;q�H;	�H;       iH;�iH;�kH;�nH;�rH;�wH;�}H;��H;��H;��H;n�H;ʡH;�H;ٯH;k�H;��H;_�H;d�H;��H; �H;��H; �H;��H;�H;��H;��H;&�H;7�H;&�H;�H;��H;�H;W�H;��H;��H;��H;��H;��H;��H;��H;W�H;�H;��H;�H;&�H;9�H;$�H;��H;��H;�H;��H;��H;��H; �H;��H;e�H;]�H;��H;k�H;ׯH;�H;ʡH;n�H;��H;��H;��H;�}H;�wH;�rH;�nH;�kH;�iH;      ?H;�?H;\BH;�FH;OLH;HSH;�[H;idH;�mH;�wH;�H;�H;ΕH;�H;��H;ԯH;Z�H;!�H;I�H;��H;:�H;\�H;�H;�H;��H;��H;y�H;�H;V�H;(�H;��H;��H;�H;l�H;��H;��H;��H;��H;��H;l�H;�H;��H;��H;&�H;V�H;�H;{�H;��H;��H;�H;�H;[�H;5�H;��H;I�H;"�H;Y�H;֯H;��H;�H;ΕH;�H;�H;�wH;�mH;hdH;�[H;KSH;JLH;�FH;]BH;�?H;      � H;'H;�H;�H;�H;s!H;@-H;�9H; GH;uTH;bH;qoH;}|H;�H;��H;��H;T�H;"�H;$�H;B�H;x�H;��H;I�H;-�H;��H;N�H;��H;��H;�H;:�H;:�H;�H;��H;�H;L�H;��H;��H;��H;M�H;�H;��H;�H;:�H;7�H;�H;��H;��H;O�H;��H;-�H;G�H;��H;q�H;B�H;$�H;$�H;S�H;��H;��H;�H;~|H;qoH;bH;vTH;GH;�9H;@-H;r!H;�H;�H;�H;2H;      �G;S�G;��G; �G;G�G;+�G;��G;��G;�H;%H;G8H;�JH;�[H;|lH;|H;��H;��H;7�H;��H;��H;ҾH;��H;t�H;a�H;��H;S�H;6�H;��H;|�H;*�H;i�H;B�H;�H;��H;�H;9�H;G�H;8�H;�H;��H;�H;E�H;i�H;(�H;{�H;��H;4�H;T�H;��H;a�H;r�H;��H;̾H;��H;��H;9�H;��H;��H;|H;|lH;�[H;�JH;H8H;%H;�H;��G;��G;*�G;I�G; �G;��G;J�G;      �wF;�F;��F;ܺF;,�F;�G;�NG;>�G;v�G;�G;��G;oH;�1H;HH;�\H;�oH;ӀH;M�H;͝H;��H;�H;ѼH;|�H;��H;�H;��H;Q�H;L�H;��H;��H;I�H;��H;e�H;*�H;��H;��H;��H;��H;��H;*�H;d�H;��H;I�H;��H;��H;L�H;P�H;��H;
�H;��H;z�H;ѼH;۳H;��H;͝H;O�H;рH;�oH;�\H;HH;�1H;pH;��G;�G;x�G;<�G;�NG;�G;0�F;ٺF;��F;�F;      ��C;Z	D;qBD;�D;
E;˄E;wF;�wF;�F;=G;$�G;�G;��G;'H;�4H;�MH;:dH;FxH;��H;�H;��H;�H;��H;��H;_�H;�H;��H;��H;��H;��H;��H;��H;��H;o�H;�H;u�H;}�H;s�H;�H;o�H;��H;��H;��H;��H;��H;��H;��H;�H;_�H;��H;��H;�H;��H;�H;��H;IxH;8dH;�MH;�4H;&H;��G;�G;"�G;=G;�F;�wF;wF;˄E;
E;�D;rBD;Z	D;      U,>;dZ>;�>;��?;`�@;
�A;�C;D;�E;��E;	�F;G;�}G;t�G;�G;�!H;w@H;�ZH;hqH;\�H;k�H;��H;�H;0�H;��H;��H;`�H;*�H;�H;�H;|�H;M�H;��H;��H;v�H;��H;�H;��H;y�H;��H;��H;O�H;~�H;�H;�H;*�H;^�H;��H;��H;0�H;�H;��H;f�H;[�H;hqH;�ZH;u@H;�!H;�G;t�G;�}G;G;�F;��E;�E;D;�C;�A;o�@;��?;�>;YZ>;      Q�1;uJ2;�g3;�$5;�Y7;�9;|g<;G�>;A;�C;8�D;:�E;v�F;E*G;]�G;c�G;�H;�5H;*SH;�lH;H�H;ǔH;>�H;�H;��H;}�H;u�H;G�H;�H;��H;��H;��H;��H;��H;��H;>�H;��H;>�H;��H;��H;��H;��H;��H;��H;�H;G�H;r�H;~�H;��H;�H;:�H;ǔH;A�H;�lH;*SH;�5H;�H;c�G;^�G;E*G;v�F;9�E;8�D;�C;A;E�>;zg<;�9;�Y7;�$5;yg3;eJ2;      �;��;;�z ;��$;h�);�/;54;�8;^�<;"$@;v�B;J�D;��E;=�F;�cG;��G;�H;�-H;�NH;jH;Z�H;ƔH;¤H;�H;ӼH;��H;��H;\�H;�H;��H;B�H;]�H;��H;��H;~�H;��H;~�H;��H;��H;]�H;C�H;��H;��H;Y�H;��H;��H;ӼH;�H;��H;H;Z�H;jH;�NH;�-H;�H;��G;�cG;>�F;��E;J�D;v�B; $@;]�<;�8;34;�/;h�);��$;�z ;;��;      {�:��:;��:v��:�;�Y;�';��;��(;��0;�Y7;b�<;�@;aC;<CE;�wF;�8G;��G;w�G;�)H;�LH;jH;F�H;m�H;��H;�H;ξH;u�H;7�H;��H;&�H;g�H;��H;��H;��H;��H;��H;��H;��H;��H;��H;j�H;&�H;��H;3�H;t�H;˾H;�H;��H;i�H;D�H;jH;�LH;�)H;w�G;��G;�8G;�wF;<CE;aC;�@;b�<;�Y7;��0;��(;��;�';�Y;�;v��:5��:��:      ��:��:x3<:�)i:�t�:��:��:�+�:�Y;N�;�*';�1;H�8;�Z>;_0B;"�D;�2F;5G;��G;+�G;�)H;�NH;�lH;[�H;w�H;��H;��H;?�H;��H;�H;J�H;;�H;B�H;k�H;��H;��H;��H;��H;��H;k�H;A�H;<�H;I�H;�H;��H;?�H;��H;��H;w�H;X�H;�lH;�NH;�)H;-�G;��G;7G;�2F;"�D;_0B;�Z>;H�8;�1;�*';N�;�Y;�+�:��:��:�t�:�)i:d3<:��:      楥�X��� ��l�=��ڷ��ߤ8��:�P�:�P�:���::`;�;7�*;%5;�g<;=A;CD;F;�G;��G;v�G;�-H;*SH;hqH;�H;ѝH;��H;'�H;J�H;�H;�H;��H;c�H;��H;��H;��H;��H;��H;��H;��H;c�H;��H;�H;��H;H�H;%�H;��H;ѝH;��H;eqH;&SH;�-H;u�G;��G;�G; F;CD;=A;�g<;%5;7�*;�;:`;���:�P�:�P�:��:��8�ڷ�p�=�� ��X��      �1��-Ȅ�Шu��PV��.�����W��P��X�9@+i:���:",�:+�;�t%;�J2;k;;��@;~D;F;9G;��G;�H;�5H;�ZH;CxH;O�H;;�H;(�H;$�H;j�H;|�H;*�H;?�H;7�H;M�H;i�H;��H;i�H;M�H;9�H;>�H;,�H;~�H;g�H;!�H;'�H;7�H;Q�H;ExH;�ZH;�5H;�H;��G;:G;F;D;��@;k;;�J2;�t%;+�;",�:���:8+i:�X�9X��W�����z.��PV�Шu�2Ȅ�      ]��M�	������(Tʻ�R��3|�h.�Ⱥ���xY�9Fu�:��:�Y;��!;��0;��:;��@;CD;�2F;�8G;��G;�H;y@H;5dH;ӀH;��H;T�H;W�H;\�H;��H;�H;��H;}�H;��H;�H;��H;�H;��H;~�H;��H;�H;��H;[�H;V�H;U�H;��H;րH;5dH;u@H;�H;��G;�8G;�2F;CD;ĵ@;��:;��0;��!;�Y;��:Du�:pY�9���Ⱥi.�3|��R��'Tʻ�����O�	�      Īx��[t���g�UT�b�:���� ���0����1��M�(�,W����t�,o`:{��:�\;{ ;��0;m;;=A;(�D;�wF;�cG;c�G;�!H;�MH;�oH;��H;��H;ӯH;��H;t�H;��H;j�H;|�H;�H;��H;4�H;��H;�H;}�H;h�H;��H;u�H;��H;ЯH;��H;��H;�oH;�MH;�!H;`�G;�cG;�wF;(�D;=A;o;;��0;{ ;�\;{��:,o`: �t�,W��O�(��1��0��� ������b�:�UT���g��[t�      <,˼��Ǽ�"���뮼w��)G��0�[�fy-�����.��̕b�h0�Hط�45<:M�:�\;��!;�J2;�g<;`0B;<CE;<�F;]�G;�G;�4H;�\H;|H;��H;��H;g�H;��H;N�H;��H;_�H;a�H;�H;��H;�H;`�H;_�H;��H;R�H;��H;g�H;��H;��H;|H;�\H;�4H; �G;Y�G;<�F;<CE;`0B;�g<;�J2;��!;�\;M�:05<:Hط�h0�˕b��.�����fy-�0�[�(G��w���뮼�"����Ǽ      /���k��Mv��t�H�Ѽ�뮼0X��s�W������׻ Ȅ������<5<:}��:�Y;�t%;%5;�Z>;aC;��E;E*G;t�G;#H;HH;|lH;�H;�H;үH;�H;��H;��H;�H;��H;}�H;=�H;}�H;��H;�H;��H;��H;߼H;үH;�H;�H;|lH;HH;$H;q�G;@*G;��E;aC;�Z>;%5;�t%;�Y;}��:85<:������Ǆ���׻���s�W�0X���뮼G�Ѽ�t�Mv���k�      Jm��Fi��&^�c�L�T�6�+����$}ռsT����x�Ļ0���������8ط�,o`:��:-�;9�*;J�8;�@;I�D;x�F;~G;��G;�1H;�[H;}|H;͕H;�H;��H;��H;��H;��H;��H;��H;��H;��H;��H;��H;��H;��H;��H;�H;˕H;}|H;�[H;�1H;��G;�}G;t�F;I�D;�@;J�8;8�*;-�;��:,o`:@ط���������Ļ0���x�sT��$}ռ��+��T�6�c�L��&^��Fi�      O��w;��D�������섽}�e��?��k��t�鷼 G���e7���� Ȅ�d0� �t�Fu�:$,�:�;�1;b�<;s�B;7�E;G; �G;mH;�JH;koH;�H;��H;"�H;��H;��H;,�H;��H;�H;��H;�H;��H;,�H;��H;��H;"�H;��H;�H;koH;�JH;mH;�G;G;5�E;s�B;d�<;�1;�;(,�:Du�: �t�d0� Ȅ���껈e7� G��鷼�t��k��?�}�e��섽���D���w;��      t���)��s��ӽ�'��C�������Z��Q+�����"�� G��Ļ0���׻˕b�(W��hY�9���::`;�*';�Y7;$@;8�D;�F;"�G;��G;E8H;bH;�H;f�H;��H;�H;��H;��H;��H;\�H;H�H;\�H;��H;��H;��H;��H;��H;f�H;	�H;bH;E8H;��G;%�G;�F;5�D;$@;�Y7;�*';:`;���:hY�9,W��˕b���׻Ļ0� G���"������Q+��Z����C����'���ӽ�s�)��      �!,�:)��K ���������޽!������Fi��0����鷼��x�����.��O�(����8+i:���:N�;��0;\�<;�C;��E;=G;�G;%H;pTH;�wH;��H;#�H;Y�H;��H;L�H;��H;��H;��H;��H;��H;L�H;��H;[�H;#�H;��H;�wH;pTH;%H;�G;=G;��E;�C;Z�<;��0;L�;���:@+i:���O�(��.�������x�鷼����0��Fi����!����޽�������K �;)�      ,�j��f��Z�|�F��>/��^�q����ŽI ���Fi��Q+��t�sT��t�W�����1��Ⱥ�X�9�P�:�Y;��(;�8;A;�E;�F;v�G;�H;�FH;�mH;��H;͡H;K�H;{�H;��H;��H;�H; �H;�H;��H;��H;x�H;M�H;ΡH;��H;�mH;�FH;�H;v�G;�F;�E;	A;�8;��(;�Y;�P�:�X�9Ⱥ�1�����t�W�sT���t�Q+��Fi�I ���Žr����^��>/�|�F��Z��f�      ��y���z�J����f��SC��K �rn���Ž����Z��k�$}ռ0X��ey-�/���h.�@���P�:�+�:��;,4;E�>;D;�wF;@�G;��G;�9H;edH;��H;��H;n�H;|�H;��H;��H;_�H;|�H;`�H;��H;��H;{�H;n�H;��H;��H;bdH;�9H;��G;?�G;�wF;D;E�>;+4;��;�+�:�P�:8��k.�/���ey-�0X��$}ռ�k��Z�����Žrn���K ��SC��f�J���z�y���      ��˾��Ǿ����"���X͓�^�x���J��K �r���!������?����뮼0�[�#���3|��W����:��:�';|/;tg<;�C;wF;�NG;��G;<-H;|[H;�}H;ӗH;֪H;ʸH;��H;	�H;��H;�H;��H;	�H;��H;ǸH;֪H;ӗH;�}H;{[H;<-H;��G;�NG;zF;�C;rg<;{/;�';��:��:�W��3|�$���0�[��뮼���?����!��r����K ���J�^�x�X͓�"���������Ǿ      u� ��������{Ծm���x���^�x��SC��^���޽C���}�e�+��H�Ѽ)G������R������ߤ8��:�Y;^�);��9;�A;ȄE;�G;+�G;u!H;NSH;�wH;��H;��H;O�H;��H;��H;��H;��H;��H;��H;��H;M�H;��H;��H;�wH;ISH;u!H;*�G;�G;ȄE;�A;��9;^�);�Y;��:�ߤ8����R�����)G��H�Ѽ+��}�e�C�����޽�^��SC�^�x�x���m����{Ծ�쾤���      ��� E�l�v� �Y�ݾm���X͓��f��>/�����'���섽T�6��t�w��b�:�'Tʻ~.��ڷ��t�:�;��$;�Y7;f�@;
E;+�F;F�G;�H;JLH;�rH;��H;ڤH;1�H;,�H;@�H;V�H;��H;X�H;?�H;,�H;0�H;ۤH;��H;�rH;ILH;�H;G�G;(�F;
E;a�@;�Y7;��$;�;�t�:�ڷ�}.�(Tʻb�:�w���t�T�6��섽�'������>/��f�X͓�m���Y�ݾv� �l� E�      ��7�v3�1�'����v� ��{Ծ"���J���|�F�����ӽ���c�L�Mv��뮼VT����PV�x�=��)i:z��:�z ;�$5;��?;�D;ٺF;�G;�H;�FH;�nH;��H;��H;�H;�H;F�H;e�H;�H;e�H;F�H;�H;~�H;��H;��H;�nH;�FH;�H;�G;ٺF;�D;��?;�$5;�z ;���:�)i:t�=��PV���VT��뮼Mv�c�L�����ӽ���|�F�J���"����{Ծv� ����1�'�v3�      �N��TI���;�1�'�l��쾂���z󐾶Z��K ��s�D����&^���"����g����Ԩu�� ��P3<:��:;qg3;��>;�BD;F;��G;�H;XBH;�kH;d�H;�H;<�H;�H;~�H;��H;V�H;��H;~�H;�H;;�H;�H;d�H;�kH;VBH;�H;��G;��F;�BD;��>;ug3;;!��:P3<:� ��Ԩu������g��"����&^�D����s潨K ��Z�z󐾂�����l�1�'���;��TI�      c]�g�W��TI�v3� E�������Ǿy����f�:)�*��w;���Fi��k���Ǽ�[t�O�	�.Ȅ�X��d�:��:��;dJ2;]Z>;T	D;�F;P�G;&H;�?H;�iH;��H;�H;��H;I�H;��H;h�H;��H;h�H;��H;I�H;��H;�H;��H;�iH;�?H;&H;N�G;�F;S	D;XZ>;jJ2;��;
��:\�:X��-Ȅ�P�	��[t���Ǽ�k��Fi�w;��*��:)��f�y�����Ǿ���� E�v3��TI�g�W�      4�$��� ����%��C��*�þ�*��5Dx���=�����Pν
���)'K��c�%��v�V����E^���S�x[:���:e;e�4;O`?;�mD;��F;avG;G�G;�H;�OH;�sH;�H;��H;��H;+�H;��H;X�H;��H;+�H;��H;��H;��H;�sH;�OH;�H;G�G;avG;��F;�mD;K`?;g�4;e;���:x[:��S�E^����w�V�%���c�)'K�
����Pν�����=�5Dx��*��*�þC��%������� �      �� ����T��P��2������0��8�s�ڀ:�j9�!�ʽ5Z���G��8�.���5S����0X�d�D��Bd:�B�: ;,�4;ӈ?;D;Y�F;$yG;��G;� H;QPH;PtH;G�H;��H;��H;i�H;��H;j�H;��H;j�H;��H;��H;I�H;PtH;OPH;� H;��G;$yG;X�F;D;ψ?;1�4; ;�B�:�Bd:d�D�0X���껴5S�.���8��G�5Z��!�ʽj9�ڀ:�8�s��0�����2��P��T�����      ���T��;�
������Yؾ"���॒���f���0�][�R8��Ӑ����>�����PȤ��6H�e�ܻrF������}:���:t";e�5;�?;��D;�F;�G;��G;v#H;�RH;�uH;��H;��H;��H;�H;%�H;��H;%�H; �H;��H;��H;��H;�uH;�RH;t#H;��G; �G;�F;��D;��?;h�5;t";���:��}:���rF�f�ܻ�6H�PȤ�������>�Ӑ��R8��][���0���f�॒�"����Yؾ����:�
�T��      %��P������AI�*�þ�R��=���wS��Q"��s������}��0��켍�����6�J�ƻ<}*�Ȇ���:�x;l%;m7;�@;��D;�F;��G;��G;8(H;VH;�xH;��H;z�H;ֲH;�H;��H;��H;��H;�H;زH;x�H;��H;�xH;VH;5(H;��G;��G;�F;��D;�@;m7;l%;�x;�:Ȇ��:}*�J�ƻ��6��������0���}�����s��Q"�wS�=����R��*�þAIᾧ���P��      C��2�很Yؾ+�þĪ�~쏾�k�ڀ:����ؽ�����c�ay���Ҽ���H� �j�-�� +(7��:��
;�(;�_9;ƘA;�\E;��F;ٝG;��G;�.H;�ZH;"|H;*�H;}�H;��H;I�H;�H;��H;�H;G�H;��H;|�H;+�H;"|H;�ZH;�.H;��G;۝G;��F;�\E;��A;�_9;�(;��
;��: +(7,��j�H� ������Ҽay��c������ؽ��ڀ:��k�~쏾Ī�+�þ�Yؾ3��      *�þ���"����R��~쏾9�s��H�����������Ґ����D��c�����E�f�W,�����P����9��:�;<j-;��;;��B;�E;�G;��G;��G;�6H;�`H;��H;��H;�H;��H;ݾH;��H;�H;��H;ݾH;��H;�H;��H;��H;�`H;�6H;��G;��G;�G;�E;��B;��;;<j-;�;��:��9�P�����W,�E�f������c���D�Ґ�������������H�9�s�~쏾�R��"������      �*���0��॒�=����k��H��#%�][��Pνt��f�f�7/%���伊���{�=��?ػ�FL���D���R::�:B�;O2;��=;ԚC;�0F;�GG;��G;VH;@H;�gH;��H;i�H;�H;̸H;��H;'�H;��H;'�H;��H;̸H;�H;k�H;��H;�gH;@H;VH;��G;�GG;�0F;њC;��=;O2;C�;6�:��R:��D��FL��?ػ{�=��������7/%�f�f�t���Pν][��#%��H��k�=���॒��0��      5Dx�8�s���f�wS�ڀ:����][��7ս�榽��}���;��8�Z�����r����>G����`̬�G��:0�;�}$;��6;2�?;�D;��F;�pG;��G;H;_JH;joH;u�H;��H;3�H;q�H;��H;��H;`�H;��H;��H;q�H;1�H;��H;u�H;joH;]JH;H;��G;�pG;��F;�D;2�?;�6;�}$;.�;G��: ̬���=G�������r�Z����8���;���}��榽�7ս][����ڀ:�wS���f�8�s�      ��=�ڀ:���0��Q"��������Pν�榽C���G�5����Ҽ	 ��OE:�B�ܻ�D^������i:j��:�;N|,;ϡ:;��A;ciE;��F;T�G;��G;�(H;oUH;�wH;��H;_�H;ɳH;,�H;�H;��H;M�H;��H;�H;+�H;ȳH;a�H;��H;�wH;mUH;�(H;��G;U�G;��F;`iE;��A;ϡ:;Q|,;�;j��:�i:�����D^�B�ܻOE:�	 ����Ҽ6���G�C���榽�Pν�������Q"���0�ڀ:�      ���j9�^[��s��ؽ���t����}��G������4c��]�V�J,��*����� ����:B��:x ;~�3;�0>;��C;
F;9G;i�G;�H;%8H;�`H;5�H;&�H;3�H;�H;#�H;��H;�H;M�H;�H;��H;#�H;|�H;6�H;&�H;5�H;�`H;&8H;�H;j�G;9G;F;��C;�0>;}�3;v ;B��:��: ������*��I,�]�V�4c��������G���}�t�������ؽ�s�^[�j9�      �Pν �ʽR8���������Ґ��f�f���;�6�����HȤ�:�f�-��Rߵ�Wo5���D�~�-:e��:�>;�+;�_9;�A;��D;K�F;�vG;�G;MH;�GH;�lH;�H;̞H;-�H;c�H;.�H;��H;<�H;`�H;<�H;��H;-�H;a�H;0�H;̞H;�H;�lH;�GH;MH;�G;�vG;E�F;��D;�A;�_9;�+;�>;i��:v�-:��D�Wo5�Qߵ�-��:�f�GȤ����6����;�f�f�Ґ���������R8�� �ʽ      
���5Z��Ґ����}��c���D�7/%��8���Ҽ4c��:�f�����ƻ�/X�R���討9-�:M�;�";��3;^>;kYC;��E;G;!�G;��G;�,H;:WH;JxH;��H;j�H;"�H;H�H;&�H;l�H;{�H;k�H;{�H;n�H;&�H;H�H;%�H;l�H;��H;JxH;;WH;�,H;��G;�G;G;��E;mYC;^>;��3;�";P�;+�:�9R����/X��ƻ���:�f�4c����Ҽ�8�7/%���D��c���}�Ґ��5Z��      ('K��G���>��0�by��c����Z���	 ��]�V�-���ƻ�od�|�º �(7�4�:���:��;Q.;�:;5zA;X�D;��F;}nG;r�G;'H;�@H;[fH;��H;c�H;�H;�H;!�H;'�H;��H;��H;u�H;��H;��H;%�H;"�H;�H;�H;c�H;��H;\fH;�@H;*H;q�G;ynG;��F;Z�D;5zA;��:;Q.;��;���:�4�: �(7x�º�od��ƻ,��\�V�	 ��Z�����伙c�by��0���>��G�      �c��8���������Ҽ����������r�OE:�I,�Pߵ��/X�z�º�Ŭ���}:)�:;_�);Fm7;>�?;��C;2F;�)G;B�G;��G;<*H;�SH;�tH;��H;��H;+�H;�H;��H;�H;L�H;��H;��H;��H;L�H;�H;��H;�H;,�H;��H;��H;�tH;�SH;=*H;�G;A�G;�)G;2F;��C;<�?;Gm7;b�);;)�:��}:�Ŭ�x�º/X�Pߵ�H,�NE:���r�����������Ҽ�켽����8�      $��.��PȤ��������E�f�{�=����C�ܻ�*��Xo5�T��� �(7��}:�n�:A�;�>&;��4;�=;��B;�E;?�F;āG;&�G;hH;�AH;�eH;u�H;�H;��H;�H;��H;\�H;��H;��H;��H;��H;��H;��H;��H;[�H;��H;�H;��H;�H;w�H;�eH;�AH;fH;"�G;��G;@�F;�E;��B;�=;��4;�>&;A�;�n�:��}: �(7R���Wo5��*��B�ܻ���{�=�D�f��������PȤ�.��      u�V��5S��6H���6�H� �X,��?ػ?G���D^������D�討9�4�:'�:B�; %;��3;8�<;|B;�E;+�F;�XG;7�G;| H;�0H;�WH;�vH;)�H;��H;��H;˽H;�H;��H;��H;��H;��H;v�H;��H;��H;��H;��H;�H;˽H;��H;��H;*�H;�vH;�WH;�0H;w H;4�G;�XG;*�F;�E;~B;;�<;��3; %;B�;)�:�4�:討9��D�����D^�@G���?ػW,�H� ���6��6H��5S�      ��ﻭ��e�ܻK�ƻk󩻹���FL����������~�-:+�:���:;�>&;��3;v9<;3�A;�D;tZF;N5G;-�G;�G;�!H;jJH;kkH;܅H;��H;��H;׸H;%�H;��H;��H;�H;��H;��H;/�H;��H;��H;�H;��H;��H;%�H;ԸH;��H;��H;مH;mkH;jJH;�!H;�G;/�G;N5G;uZF;�D;6�A;v9<;��3;�>&;;���:+�:v�-:����������FL����j�K�ƻe�ܻ���      E^�0X�rF�8}*�0���P����D��̬��i:��:i��:M�;��;\�);��4;6�<;2�A;E�D;�9F; G;��G;x�G;rH;P?H;�aH;N}H;��H;��H;ԳH;�H;��H;��H;��H;W�H;��H;^�H;��H;^�H;��H;V�H;��H;��H;��H;�H;ҳH;��H;��H;P}H;�aH;N?H;pH;y�G;��G;G;�9F;H�D;2�A;6�<;��4;_�);��;N�;i��:��:�i:�̬���D��P��*��6}*�rF�0X�      d�S�l�D����Ȇ�� ((7��9��R:C��:l��:B��:�>;�";
Q.;Gm7;�=;{B;�D;�9F;LG;O�G;��G;�H;�6H;�YH;vH;[�H;*�H;:�H;=�H;��H;^�H;��H;U�H;s�H;��H;��H;2�H;��H;��H;s�H;T�H;��H;]�H;��H;:�H;9�H;&�H;\�H;vH;�YH;�6H;�H;��G;R�G;NG;�9F;�D;{B;�=;Fm7;
Q.;�";�>;B��:p��:C��:��R:��9 .(7Ȇ�����h�D�      x[:4Cd:��}:�:��:
��:4�:-�;�;x ;�+;��3;��:;7�?;��B;�E;pZF;�G;M�G;��G;vH;�1H;TH;�pH;�H;��H;"�H;��H;��H;��H;:�H;�H;��H;]�H;1�H;Q�H;��H;Q�H;1�H;\�H;��H;�H;:�H;��H;��H;��H;�H;��H;�H;�pH;
TH;�1H;tH;��G;N�G;�G;qZF;�E;��B;7�?;��:;��3;�+;x ;�;-�;6�:��:��:�:��}:Cd:      ���:�B�:��:yx;��
;�;E�;�}$;M|,;~�3;�_9;[>;3zA;��C;�E;+�F;N5G;��G;��G;xH;�/H;+QH;=mH;��H;חH;ϧH;��H;7�H;��H;T�H;��H;��H;��H; �H;��H;��H;��H;��H;��H;�H;��H;��H;��H;Q�H;��H;7�H;��H;ϧH;חH;��H;;mH;+QH;�/H;zH;��G;��G;M5G;+�F;�E;��C;2zA;[>;�_9;}�3;P|,;�}$;F�;�;��
;|x;���:�B�:      )e;2 ;�";d%;�(;Cj-;Y2;�6;ҡ:;�0>;�A;kYC;V�D;4F;B�F;�XG;-�G;{�G;�H;�1H;*QH;lH;��H;��H;s�H;j�H;�H;��H;��H;K�H;��H;�H;��H;��H;��H;��H;��H;��H;��H;��H;��H;�H;��H;G�H;��H;��H;�H;k�H;s�H;��H;��H;lH;(QH;�1H;�H;{�G;-�G;�XG;C�F;2F;X�D;kYC;�A;�0>;ա:;�6;W2;Fj-;�(;e%;�";, ;      m�4;-�4;e�5;m7;�_9;��;;��=;2�?;��A;��C;��D;��E;��F;�)G;āG;7�G;�G;uH;�6H;TH;=mH;��H;�H;E�H;��H;��H;d�H;o�H;�H;��H;T�H;)�H;q�H;��H; �H;��H;��H;��H; �H;��H;n�H;)�H;T�H;��H;�H;o�H;a�H;��H;��H;C�H;�H;��H;9mH;TH;�6H;vH;�G;4�G;āG;�)G;��F;��E;��D;��C;��A;1�?;��=;��;;�_9;m7;h�5;�4;      a`?;ۈ?;
�?;�@;ƘA;��B;ۚC;�D;aiE;F;H�F;G;ynG;A�G;%�G;z H;�!H;S?H;�YH;�pH;��H;��H;E�H;��H;˺H;g�H;��H;C�H;��H;��H;��H;��H;��H;�H;��H;t�H;��H;r�H;��H;�H;��H;��H;��H;��H;��H;C�H;��H;g�H;̺H;~�H;B�H;��H;��H;�pH;�YH;S?H;�!H;z H;%�G;A�G;ynG;G;H�F;F;aiE;�D;ښC;��B;͘A;�@;�?;ш?;      �mD;D;t�D;��D;�\E;�E;�0F;��F;��F;9G;�vG;!�G;q�G;��G;hH;�0H;pJH;�aH;"vH;�H;ۗH;w�H;��H;ӺH;)�H;�H;��H;O�H;&�H;7�H;��H;|�H;��H;�H;��H;#�H;g�H;"�H;��H;�H;��H;}�H;��H;6�H;#�H;O�H;��H;�H;*�H;ѺH;��H;w�H;ڗH; �H;"vH;�aH;nJH;�0H;hH;��G;p�G;!�G;�vG;9G;��F;��F;�0F;�E;�\E;��D;r�D;D;      ��F;d�F;ծF; �F;��F;�G;�GG;�pG;S�G;i�G;�G;��G;'H;:*H;�AH;�WH;jkH;L}H;X�H;��H;̧H;i�H;��H;e�H;��H;t�H;��H;��H;��H;Q�H;N�H;��H;��H;��H;u�H;��H;�H;��H;v�H;��H;��H;��H;N�H;P�H;��H;��H;��H;u�H;�H;d�H;��H;i�H;ȧH;��H;X�H;M}H;hkH;�WH;�AH;:*H;'H;��G;�G;g�G;T�G;�pG;�GG;�G;��F;�F;ծF;Y�F;      lvG;&yG;�G;��G;۝G;��G;��G;��G;��G;�H;LH;�,H;�@H;�SH;�eH;�vH;ޅH;��H;)�H;#�H;��H;�H;d�H;��H;��H; �H;��H;��H;�H;�H;��H;��H;��H;��H;�H;b�H;b�H;b�H;�H;��H;��H;��H;��H;�H;�H;��H;��H;��H;��H;��H;b�H;�H;��H;%�H;*�H;��H;ޅH;�vH;�eH;�SH;�@H;�,H;LH;�H;��G;��G;��G;��G;�G;��G;�G;$yG;      <�G;��G;��G;��G;��G;��G;ZH;$H;�(H;)8H;�GH;@WH;\fH;�tH;w�H;)�H;��H;��H;7�H;��H;7�H;��H;q�H;F�H;J�H;��H;��H;��H; �H;��H;��H;��H;��H;�H;��H;��H;��H;��H;��H;�H;��H;��H;��H;��H;��H;��H;��H;��H;L�H;H�H;o�H;��H;4�H;��H;7�H;��H;�H;*�H;w�H;�tH;[fH;@WH;�GH;)8H;�(H;$H;ZH;��G;��G;��G;��G;��G;      �H;� H;t#H;;(H;�.H;�6H; @H;`JH;pUH;�`H;�lH;OxH;��H;��H;�H;��H;��H;ҳH;=�H;��H;��H;��H;�H;��H;�H;��H;�H; �H;r�H;��H;��H;��H;-�H;��H;��H;�H;/�H;�H;��H;��H;*�H;��H;��H;��H;p�H; �H;�H;��H; �H;��H;�H;��H;��H;��H;=�H;ҳH;��H;��H;�H;��H;��H;MxH;�lH;�`H;sUH;`JH; @H;�6H;�.H;;(H;t#H;� H;      �OH;WPH;�RH;VH;�ZH;�`H;�gH;qoH;�wH;>�H;��H;͑H;i�H;��H;��H;��H;׸H;�H;��H;��H;T�H;H�H;��H;��H;-�H;N�H;�H;��H;��H;��H;��H;*�H;��H;	�H;<�H;_�H;t�H;_�H;<�H;	�H;��H;*�H;��H;��H;��H;��H;�H;L�H;/�H;��H;��H;H�H;R�H;��H;��H;�H;ָH;��H;��H;��H;i�H;͑H;��H;>�H;�wH;roH;�gH;�`H;�ZH;VH;�RH;TPH;      �sH;atH;�uH;�xH;1|H;��H;ąH;�H;��H;*�H;ҞH;v�H;�H;0�H;�H;ҽH;)�H;��H;^�H;?�H;��H;��H;T�H;��H;��H;O�H;��H;��H;��H;��H;�H;��H;�H;P�H;��H;��H;��H;��H;��H;P�H;�H;��H;�H;��H;��H;��H;��H;N�H;��H;��H;P�H;��H;��H;?�H;`�H;��H;(�H;ѽH;�H;/�H;�H;t�H;ҞH;,�H;��H;}�H;ƅH;��H;.|H;�xH;�uH;atH;       �H;S�H;��H;��H;1�H;��H;n�H;��H;c�H;5�H;4�H;*�H;�H;�H;��H;
�H;�H;��H;��H;�H;��H;"�H;)�H;��H;x�H;��H;��H;��H;��H;,�H;��H;�H;L�H;��H;��H;��H;��H;��H;��H;��H;I�H;�H;��H;-�H;��H;��H;��H;��H;{�H;��H;'�H;"�H;��H;�H;��H;��H;�H;
�H;��H;�H;�H;,�H;4�H;5�H;e�H;��H;n�H;��H;.�H;��H;��H;O�H;      ��H;�H; �H;��H;��H;�H;�H;<�H;ϳH;�H;d�H;P�H;%�H;��H;]�H;��H;��H;��H;U�H;��H;��H;��H;q�H;��H;��H;��H;��H;��H;1�H;��H;	�H;P�H;��H;��H;��H;��H;�H;��H;��H;��H;��H;Q�H;�H;��H;3�H;��H;��H;��H;��H;��H;p�H;��H;��H;��H;U�H;��H;��H;��H;\�H;��H;%�H;O�H;d�H;��H;ϳH;:�H;�H;�H;}�H;��H;�H;�H;      ǰH;�H;��H;ܲH;��H;��H;ӸH;{�H;2�H;&�H;4�H;,�H;(�H;�H;��H;��H;�H;U�H;t�H;d�H;&�H;��H;��H;�H;�H;��H;}�H;�H;��H;	�H;M�H;��H;��H;��H;��H;�H;�H;�H;��H;��H;��H;��H;L�H;	�H;��H;�H;}�H;��H;�H;�H;��H;��H;$�H;d�H;t�H;V�H;�H;��H;��H;�H;(�H;,�H;3�H;&�H;3�H;y�H;ӸH;��H;��H;ݲH;��H;�H;      +�H;�H;�H;��H;c�H;ھH;��H;��H;�H;��H;��H;w�H;��H;Q�H;��H;��H;��H;��H;��H;8�H;��H;��H;��H;��H;��H;t�H;�H;��H;��H;?�H;��H;��H;��H;��H;�H;�H;�H;�H;�H;��H;��H;��H;��H;?�H;��H;��H;�H;t�H;��H;��H;��H;��H;��H;8�H;��H;��H;��H;��H;��H;Q�H;��H;w�H;��H;��H;�H;��H;��H;߾H;X�H;��H;�H;w�H;      ��H;��H;.�H;��H;(�H;��H;1�H;�H; �H;�H;C�H;��H;��H;��H;��H;��H;��H;W�H;��H;Y�H;��H;��H;��H;u�H;�H;��H;a�H;��H;�H;a�H;��H;��H;��H;�H;�H;0�H;(�H;0�H;�H;�H;��H;��H;��H;b�H;�H;��H;`�H;��H;�H;u�H;��H;��H;��H;Y�H;��H;Y�H;��H;��H;��H;��H;��H;��H;C�H;�H;��H;��H;1�H;��H;�H;��H;0�H;��H;      \�H;s�H;��H;��H;��H;�H;��H;g�H;U�H;M�H;g�H;u�H;z�H;��H;��H;|�H;5�H;��H;2�H;��H;��H;��H;��H;��H;a�H;�H;a�H;��H;1�H;{�H;��H;��H;�H;�H;�H;)�H;3�H;)�H;�H;�H;�H;��H;��H;{�H;4�H;��H;`�H;�H;a�H;��H;��H;��H;��H;��H;2�H;��H;3�H;|�H;��H;��H;z�H;u�H;g�H;P�H;V�H;d�H;��H;�H;��H;��H;��H;i�H;      ��H;��H;.�H;��H;(�H;��H;1�H;�H;��H;�H;C�H;��H;��H;��H;��H;��H;��H;W�H;��H;Y�H;��H;��H;��H;w�H;�H;��H;a�H;��H;�H;a�H;��H;��H;��H;�H;�H;0�H;(�H;0�H;�H;�H;��H;��H;��H;b�H;�H;��H;`�H;��H;�H;u�H;��H;��H;��H;Y�H;��H;Y�H;��H;��H;��H;��H;��H;��H;D�H;�H; �H;��H;2�H;��H;�H;��H;-�H;��H;      )�H;�H;�H;��H;c�H;ھH;��H;��H;�H;��H;��H;w�H;��H;Q�H;��H;��H;��H;��H;��H;8�H;��H;��H;��H;��H;��H;t�H;�H;��H;��H;?�H;��H;��H;��H;��H;�H;�H;�H;�H;�H;��H;��H;��H;��H;@�H;��H;��H;�H;u�H;��H;��H;��H;��H;��H;8�H;��H;��H;��H;��H;��H;Q�H;��H;w�H;��H;��H;�H;��H;��H;߾H;X�H;��H;�H;u�H;      ɰH;�H;��H;ݲH;��H;��H;ӸH;{�H;2�H;&�H;4�H;,�H;(�H;�H;��H;��H;�H;U�H;t�H;c�H;(�H;��H;��H;�H;�H;��H;}�H;�H;��H;�H;L�H;��H;��H;��H;��H;�H;�H;�H;��H;��H;��H;��H;M�H;	�H;��H;�H;}�H;��H;�H;�H;��H;��H;$�H;d�H;t�H;W�H;�H;��H;��H;�H;(�H;,�H;4�H;&�H;3�H;y�H;ӸH;��H;��H;ܲH;��H;�H;      ��H;�H;�H;��H;��H;	�H;�H;;�H;ϳH;�H;d�H;O�H;#�H;��H;\�H;��H;��H;��H;U�H;��H;��H;��H;q�H;��H;��H;��H;��H;��H;1�H;��H;�H;P�H;��H;��H;��H;��H;�H;��H;��H;��H;��H;S�H;	�H;��H;3�H;��H;��H;��H;��H;��H;p�H;��H;��H;��H;U�H;��H;��H;��H;]�H;��H;#�H;P�H;d�H;��H;ϳH;8�H;�H;�H;|�H;��H;��H;	�H;       �H;S�H;��H;��H;1�H;��H;p�H;��H;c�H;6�H;4�H;*�H;�H;�H;��H;
�H;�H;��H;��H;�H;��H;"�H;*�H;��H;{�H;��H;��H;��H;��H;,�H;��H;�H;J�H;��H;��H;��H;��H;��H;��H;��H;I�H;�H;��H;-�H;��H;��H;��H;��H;x�H;��H;'�H;"�H;��H;�H;��H;��H;�H;�H;��H;�H;�H;,�H;4�H;6�H;e�H;��H;p�H;��H;-�H;��H;��H;O�H;      �sH;atH;�uH;�xH;1|H;��H;ƅH;�H;��H;*�H;ҞH;t�H;�H;0�H;�H;ҽH;(�H;��H;`�H;?�H;��H;��H;T�H;��H;��H;O�H;��H;��H;��H;��H;�H;��H;�H;P�H;��H;��H;��H;��H;��H;P�H;�H;��H;�H;��H;��H;��H;��H;N�H;��H;��H;Q�H;��H;��H;?�H;^�H;��H;(�H;ҽH;�H;0�H;�H;v�H;ўH;,�H;��H;�H;ąH;��H;.|H;�xH;�uH;`tH;      �OH;VPH;�RH;VH;�ZH;�`H;�gH;toH;�wH;<�H;��H;͑H;i�H;��H;��H;��H;׸H;�H;��H;��H;V�H;H�H;��H;��H;/�H;M�H;�H;��H;��H;��H;��H;*�H;��H;�H;<�H;_�H;t�H;_�H;<�H;	�H;��H;,�H;��H;��H;��H;��H;�H;M�H;-�H;��H;��H;H�H;R�H;��H;��H;�H;ָH;��H;��H;��H;i�H;͑H;��H;<�H;�wH;toH;�gH;�`H;�ZH;VH;�RH;VPH;      �H;� H;{#H;:(H;�.H;�6H;%@H;bJH;pUH;�`H;�lH;OxH;��H;��H;�H;��H;��H;гH;=�H;��H;��H;��H;�H;��H; �H;��H;�H; �H;p�H;��H;��H;��H;,�H;��H;��H;�H;/�H;�H;��H;��H;,�H;��H;��H;��H;p�H; �H;�H;��H;�H;��H;�H;��H;��H;��H;=�H;ӳH;��H;��H;�H;��H;��H;OxH;�lH;�`H;qUH;`JH;#@H;�6H;�.H;7(H;{#H;� H;      <�G;��G;��G;��G;��G;��G;ZH;%H;�(H;)8H;�GH;@WH;[fH;�tH;w�H;*�H;��H;��H;7�H;��H;:�H;��H;q�H;F�H;L�H;��H;��H;��H; �H;��H;��H;��H;��H;�H;��H;��H;��H;��H;��H;�H;��H;��H;��H;��H;��H;��H;��H;��H;J�H;H�H;o�H;��H;6�H;��H;7�H;��H;�H;*�H;w�H;�tH;\fH;@WH;�GH;)8H;�(H;$H;ZH;��G;��G;��G;��G;��G;      gvG;'yG; �G;��G;ڝG;��G;��G;��G;��G;�H;LH;�,H;�@H;�SH;�eH;�vH;ޅH;��H;*�H;%�H;��H;�H;d�H;��H;��H; �H;��H;��H;�H;�H;��H;��H;��H;��H;�H;b�H;b�H;a�H;�H;��H;��H;��H;��H;�H;�H;��H;��H; �H;��H;��H;b�H;�H;��H;#�H;)�H;��H;܅H;�vH;�eH;�SH;�@H;�,H;MH;�H;��G;��G;��G;��G;ݝG;��G;�G;yG;      ��F;`�F;߮F;�F;��F;�G;�GG;�pG;S�G;i�G;�G;��G;'H;:*H;�AH;�WH;jkH;L}H;X�H;��H;ͧH;i�H;��H;d�H;�H;t�H;��H;��H;��H;Q�H;N�H;��H;��H;��H;t�H;��H;�H;��H;v�H;��H;��H;��H;N�H;N�H;��H;��H;��H;u�H;��H;d�H;��H;i�H;ȧH;��H;X�H;M}H;hkH;�WH;�AH;:*H;'H;��G;�G;g�G;S�G;�pG;�GG;�G;��F; �F;߮F;V�F;      �mD;D;r�D;��D;�\E;�E;�0F;��F;��F;9G;�vG;!�G;p�G;��G;hH;�0H;nJH;�aH;"vH; �H;ݗH;w�H;��H;ҺH;*�H;�H;��H;O�H;&�H;7�H;��H;|�H;��H;�H;��H;#�H;g�H;"�H;��H;�H;��H;�H;��H;6�H;#�H;O�H;��H;�H;)�H;ҺH;��H;w�H;ڗH; �H;"vH;�aH;mJH;�0H;hH;��G;q�G;!�G;�vG;9G;��F;��F;�0F;�E;�\E;��D;r�D;D;      g`?;ڈ?;�?;�@;��A;��B;ךC;�D;ciE;F;I�F;G;znG;A�G;%�G;z H;�!H;P?H;�YH;�pH;��H;��H;E�H;��H;̺H;e�H;��H;C�H;��H;��H;��H;��H;��H;	�H;��H;t�H;��H;r�H;��H;�H;��H;��H;��H;��H;��H;C�H;��H;g�H;˺H;��H;B�H;��H;��H;�pH;�YH;U?H;�!H;z H;%�G;A�G;ynG;G;G�F;F;ciE;�D;ךC;��B;јA;�@;�?;ψ?;      f�4;9�4;w�5;m7;�_9;��;;��=;2�?;��A;��C;��D;��E;��F;�)G;āG;5�G;�G;rH;�6H;TH;?mH;��H;�H;E�H;��H;��H;d�H;o�H;�H;��H;T�H;)�H;q�H;��H; �H;��H;��H;��H; �H;��H;p�H;)�H;T�H;��H;�H;o�H;b�H;��H;��H;C�H;�H;��H;9mH;TH;�6H;vH;�G;7�G;ƁG;�)G;��F;��E;��D;��C;��A;1�?;��=;��;;�_9;m7;l�5;*�4;      )e;2 ;�";e%;�(;Dj-;W2;�6;ҡ:;�0>;�A;kYC;X�D;4F;B�F;�XG;,�G;y�G;�H;�1H;+QH;lH;��H;��H;s�H;j�H;�H;��H;��H;K�H;��H;�H;��H;��H;��H;��H;��H;��H;��H;��H;��H;�H;��H;G�H;��H;��H;�H;k�H;s�H;��H;��H;lH;*QH;�1H;�H;|�G;,�G;�XG;C�F;2F;V�D;mYC;�A;�0>;ա:;�6;Y2;Cj-;�(;d%;�";, ;      ���:�B�:��:|x;��
;�;I�;�}$;M|,;}�3;�_9;[>;3zA;��C;�E;+�F;N5G;��G;��G;xH;�/H;+QH;<mH;��H;חH;ͧH;��H;7�H;��H;T�H;��H;��H;��H;�H;��H;��H;��H;��H;��H; �H;��H;��H;��H;Q�H;��H;7�H;��H;ϧH;חH;��H;<mH;+QH;�/H;zH;��G;��G;M5G;+�F;�E;��C;3zA;[>;�_9;{�3;N|,;�}$;I�;�;��
;zx;��:�B�:      x[:<Cd:��}:�:��:
��::�:.�;�;y ;�+;��3;��:;7�?;��B;�E;qZF;�G;N�G;��G;xH;�1H;TH;�pH;�H;��H;"�H;��H;��H;��H;:�H;�H;��H;\�H;1�H;R�H;��H;R�H;1�H;]�H;��H;�H;:�H;��H;��H;��H;�H;��H;�H;�pH;
TH;�1H;tH;��G;M�G;�G;pZF;�E;��B;7�?;��:;��3;�+;x ;�;.�;8�:��:��:�:��}:Cd:      d�S�h�D����Ȇ�� ((7��9��R:E��:l��:B��:�>;�";
Q.;Fm7;�=;{B;�D;�9F;NG;Q�G;��G;�H;�6H;�YH;vH;Z�H;)�H;9�H;=�H;��H;]�H;��H;U�H;s�H;��H;��H;2�H;��H;��H;s�H;T�H;��H;^�H;��H;:�H;:�H;'�H;\�H;vH;�YH;�6H;�H;��G;Q�G;LG;�9F;�D;{B;�=;Fm7;
Q.;�";�>;B��:p��:C��:��R:��9 .(7Ȇ�����h�D�      E^�0X�rF�7}*�1���P����D��̬��i:��:i��:N�;��;]�);��4;6�<;3�A;G�D;�9F; G;��G;y�G;sH;R?H;�aH;M}H;��H;��H;ӳH;�H;��H;��H;��H;V�H;��H;^�H;��H;^�H;��H;W�H;��H;��H;��H;�H;ҳH;��H;��H;P}H;�aH;L?H;oH;x�G;��G;G;�9F;G�D;0�A;6�<;��4;\�);��;M�;i��:��:�i:�̬���D��P��*��8}*�	rF�0X�      ��ﻮ��f�ܻK�ƻj󩻺���FL����������~�-:+�:���:;�>&;��3;x9<;3�A;�D;uZF;N5G;/�G;�G;�!H;jJH;kkH;ޅH;��H;��H;׸H;%�H;��H;��H;�H;��H;��H;/�H;��H;��H;�H;��H;��H;%�H;ָH;��H;��H;؅H;mkH;jJH;�!H;�G;-�G;M5G;uZF;�D;5�A;v9<;��3;�>&;;���:+�:~�-:���������FL����j�K�ƻf�ܻ���      u�V��5S��6H���6�H� �X,��?ػ?G���D^������D�討9�4�:'�:B�; %;��3;:�<;~B;�E;+�F;�XG;7�G;| H;�0H;�WH;�vH;*�H;��H;��H;˽H;�H;��H;��H;��H;��H;v�H;��H;��H;��H;��H;�H;˽H;��H;��H;)�H;�vH;�WH;�0H;w H;2�G;�XG;*�F;�E;|B;:�<;��3; %;D�;%�:�4�:討9��D�����D^�?G���?ػV,�H� ���6��6H��5S�      $��.��PȤ��������E�f�{�=����D�ܻ�*��Xo5�R��� �(7��}:�n�:A�;�>&;��4;�=;��B;�E;@�F;ƁG;(�G;fH;�AH;�eH;w�H;�H;��H;�H;��H;]�H;��H;��H;��H;��H;��H;��H;��H;\�H;��H;�H;��H;�H;u�H;�eH;�AH;hH;"�G;��G;?�F;�E;��B;�=;��4;�>&;A�;�n�:��}: �(7T���Xo5��*��C�ܻ���{�=�D�f��������PȤ�.��      �c��8���������Ҽ����������r�OE:�H,�Pߵ��/X�x�º�Ŭ���}:)�:;`�);Gm7;;�?;��C;2F;�)G;C�G;�G;<*H;�SH;�tH;��H;��H;,�H;�H;��H;�H;L�H;��H;��H;��H;L�H;�H;��H;�H;+�H;��H;��H;�tH;�SH;<*H;��G;?�G;�)G;2F;��C;;�?;Fm7;b�);;)�:��}: Ƭ�z�º�/X�Pߵ�I,�NE:���r�����������Ҽ�켽����8�      ('K��G���>��0�ay��c����Z���	 ��]�V�,���ƻ�od�x�º �(7�4�:���:��;Q.;��:;3zA;Z�D;��F;~nG;q�G;(H;�@H;\fH;��H;c�H;�H;�H;"�H;%�H;��H;��H;u�H;��H;��H;'�H;�H;�H;�H;c�H;��H;[fH;�@H;*H;r�G;vnG;��F;X�D;5zA;��:;Q.;��;���:�4�: �(7|�º�od��ƻ-��]�V�	 ��Z�����伙c�by��0���>��G�      
���5Z��Ґ����}��c���D�7/%��8���Ҽ4c��:�f�����ƻ�/X�P����9-�:N�;�";��3;[>;mYC;��E;G;�G;��G;�,H;;WH;LxH;��H;l�H;"�H;I�H;(�H;n�H;|�H;k�H;|�H;l�H;&�H;G�H;#�H;j�H;��H;IxH;:WH;�,H;��G;!�G;G;��E;kYC;_>;��3;�";P�;+�:ب�9P����/X��ƻ���:�f�4c����Ҽ�8�7/%���D��c���}�Ґ��5Z��      �Pν �ʽR8���������Ґ��f�f���;�6�����GȤ�:�f�-��Rߵ�Wo5���D�z�-:g��:�>;�+;�_9;�A;��D;K�F;�vG;�G;OH;�GH;�lH;�H;̞H;-�H;c�H;-�H;��H;<�H;`�H;<�H;��H;.�H;a�H;/�H;̞H;�H;�lH;�GH;LH;�G;�vG;E�F;��D;�A;�_9;�+;�>;i��:v�-:��D�Wo5�Rߵ�-��:�f�HȤ����6����;�f�f�Ґ���������R8�� �ʽ      ���j9�^[��s��ؽ���t����}��G������4c��]�V�J,��*���������:B��:x ;{�3;�0>;��C;F;9G;j�G;�H;&8H;�`H;5�H;&�H;3�H;�H;#�H;��H;�H;M�H;�H;��H;#�H;}�H;5�H;&�H;5�H;�`H;%8H;�H;i�G;9G;F;��C;�0>;~�3;v ;B��:��: ������*��J,�]�V�5c��������G���}�t�������ؽ�s�^[�j9�      ��=�ڀ:���0��Q"��������Pν�榽C���G�5����Ҽ	 ��OE:�B�ܻ�D^������i:j��:�;N|,;ϡ:;��A;diE;��F;U�G;��G;�(H;pUH;�wH;��H;_�H;˳H;+�H;�H;��H;M�H;��H;�H;,�H;ȳH;_�H;��H;�wH;lUH;�(H;��G;T�G;��F;^iE;��A;ϡ:;P|,;�;j��:�i:�����D^�B�ܻOE:�	 ����Ҽ6���G�C���榽�Pν�������Q"���0�ڀ:�      5Dx�8�s���f�wS�ڀ:����][��7ս�榽��}���;��8�Z�����r����>G����@̬�G��:0�;�}$;�6;2�?;�D;��F;�pG;��G;H;`JH;joH;u�H;��H;3�H;r�H;��H;��H;`�H;��H;��H;r�H;1�H;��H;u�H;joH;\JH;H;��G;�pG;��F;�D;2�?;��6;�}$;.�;G��:@̬���>G�������r�Z����8���;���}��榽�7ս][����ڀ:�wS���f�8�s�      �*���0��॒�=����k��H��#%�][��Pνt��f�f�7/%���伊���{�=��?ػ�FL���D���R::�:@�;O2;��=;՚C;�0F;�GG;��G;VH;@H;�gH;��H;i�H;�H;͸H;��H;'�H;��H;'�H;��H;̸H;�H;i�H;��H;�gH;@H;VH;��G;�GG;�0F;њC;��=;O2;C�;6�:��R:��D��FL��?ػ{�=��������7/%�f�f�t���Pν][��#%��H��k�=���॒��0��      *�þ���"����R��~쏾9�s��H�����������Ґ����D��c�����E�f�W,�����P����9��:�;<j-;��;;��B;�E;�G;��G;��G;�6H;�`H;��H;��H;	�H;��H;ݾH;��H;�H;��H;ݾH;��H;�H;��H;��H;�`H;�6H;��G;��G;�G;�E;��B;��;;<j-;�;��:��9�P�����W,�E�f������c���D�Ґ�������������H�9�s�~쏾�R��"������      C��2�很Yؾ+�þĪ�~쏾�k�ڀ:����ؽ�����c�ay���Ҽ���H� �j�-�� +(7��:��
;�(;�_9;ƘA;�\E;��F;ڝG;��G;�.H;�ZH;"|H;*�H;}�H;��H;I�H;�H;��H;�H;G�H;��H;|�H;+�H;"|H;�ZH;�.H;��G;ڝG;��F;�\E;ØA;�_9;�(;��
;��: +(7,��k�H� ������Ҽay��c������ؽ��ڀ:��k�~쏾Ī�+�þ�Yؾ3��      %��P������AI�*�þ�R��=���wS��Q"��s������}��0��켍�����6�J�ƻ:}*�Ȇ���:x;l%;
m7;�@;��D;�F;��G;��G;8(H;VH;�xH;��H;z�H;زH;�H;��H;��H;��H;�H;ֲH;x�H;��H;�xH;VH;5(H;��G;��G;�F;��D;�@;m7;l%;�x;�:Ȇ��:}*�K�ƻ��6��������0���}�����s��Q"�wS�=����R��*�þAIᾧ���P��      ���T��:�
������Yؾ"���॒���f���0�][�R8��Ґ����>�����PȤ��6H�f�ܻrF������}:��:t";e�5;�?;��D;�F; �G;��G;v#H;�RH;�uH;��H;��H;��H;�H;%�H;��H;%�H;�H;��H;��H;��H;�uH;�RH;t#H;��G;�G;�F;��D;��?;h�5;t";���:��}:���rF�f�ܻ�6H�PȤ�������>�Ӑ��R8��][���0���f�॒�"����Yؾ����:�
�T��      �� ����T��P��2������0��8�s�ڀ:�j9�!�ʽ5Z���G��8�.���5S����0X�d�D��Bd:�B�: ;,�4;ӈ?;D;Y�F;$yG;��G;� H;QPH;PtH;G�H;��H;��H;i�H;��H;j�H;��H;j�H;��H;��H;I�H;PtH;OPH;� H;��G;#yG;X�F;D;Ј?;1�4; ;�B�:�Bd:d�D�0X���껴5S�.���8��G�5Z��!�ʽj9�ڀ:�8�s��0�����2��P��T�����      IF�Zh����YVھ:�������~���S��#��o��<S��s₽7�6�w���ny��\FB��Eֻ�A?���	��Y�:���:w�";�46;g@;��D;ةF;�nG;�G;BH;;@H;gH;��H;d�H;ĩH;�H;�H;��H;�H;�H;ĩH;c�H;��H;gH;:@H;?H;�G;�nG;ةF;��D;c@;�46;w�";���:�Y�:��	��A?��Eֻ]FB�ny��w���7�6�s₽<S���o���#��S��~������:��YVھ��Zh��      Zh���b���쾪*־�v��+���*��*�O�X� �s��r���؀�L�3���Eݜ�B�>�W�ѻ�9�����`o�:=% ;�M#;y�6;XA@;�D;үF;,qG;z�G;VH;AH;�gH;�H;ĚH;�H;P�H;,�H;�H;,�H;P�H;�H;ÚH;�H;�gH;AH;TH;z�G;,qG;үF;�D;RA@;�6;�M#;>% ;^o�:�����9�X�ѻB�>�Eݜ���L�3��؀��r��s�X� �*�O�*��+����v���*־���b��      ���쾷�޾25ʾP;���:��,�v��E�b'����v����u���+��W��A����4���Ļ$9)�0j���W�:b�;%;l7;1�@;�D;�F;xG;��G;xH;gCH;aiH;Q�H;țH;ڪH;��H;ʺH;��H;ʺH;�H;ڪH;ƛH;Q�H;aiH;cCH;vH;��G;xG;�F;�D;-�@;l7;%;a�;�W�:0j��"9)���Ļ��4��A���W缈�+���u�v�����b'��E�,�v��:��P;��25ʾ��޾��      YVھ�*־25ʾu��������M���9b��5�����ս����Xc�
��Җռ�I��[�$�oT���Z��[��N�:�;}�';R�8;,RA;�9E;��F;܂G;�G;�H;0GH;HlH;��H;p�H;�H;�H;ɻH;��H;ɻH;��H;�H;o�H;��H;HlH;/GH;�H;�G;܂G;��F;�9E;'RA;W�8;}�';�;L�:�[���Z�oT��[�$��I��Җռ
���Xc������ս���5��9b��M������u���25ʾ�*־      :���v��O;������UP��I�r�}�H�X� ���9@��Փ����K�e�־���s�x���񕻥ܺ�5u9Q&�:)�;D�+;��:;�"B;��E;�F;�G;�G;qH;`LH;3pH;|�H;��H;٭H;r�H;�H;��H;�H;q�H;ۭH;��H;}�H;1pH;[LH;pH;�G;�G;�F;��E;�"B;��:;D�+;*�;O&�:�5u9�ܺ��w����s�־�e���K�Փ��9@����X� �}�H�I�r�UP������O;���v��      ����+����:���M��I�r�*�O�#,�[�
��gٽtĥ���u�|1�q���/Ϥ���P�[�.o�lp��r:���:Q;U�/;l�<;C;J�E;�!G;U�G;4�G;�%H;�RH;uH;4�H;{�H;�H;=�H;��H;;�H;��H;?�H;�H;{�H;7�H;uH;�RH;�%H;4�G;S�G;�!G;J�E;C;m�<;U�/;Q;���:n:jp���.o�[򻲎P�/Ϥ�q���|1���u�tĥ��gٽ[�
�#,�*�O�I�r��M���:��+���      �~��*��,�v��9b�}�H�#,�PZ����;S��{^����N������μ�I���%+����؝.�p����j~:���:<m;��3;L�>;W�C;rPF;�FG;t�G; �G;�/H;.ZH;�zH;��H;��H;��H;Z�H;`�H;�H;^�H;\�H;��H;��H;��H;�zH;,ZH;�/H; �G;r�G;�FG;oPF;Q�C;M�>;��3;=m;���:�j~:X���؝.�����%+��I����μ�����N�{^��;S�����PZ�#,�}�H��9b�,�v�*��      �S�*�O��E��5�X� �[�
���罨9��+l���Xc���(��������[�����ݎ�6ܺ�;9F��:T�	;Xd';� 8;p�@;��D;�F;UjG;��G;�H;�:H;nbH;�H;C�H;h�H;}�H;��H;p�H;�H;p�H;��H;}�H;f�H;E�H;�H;mbH;�:H;�H;��G;VjG;�F;��D;p�@;� 8;Yd';R�	;H��:�;99ܺ�ݎ������[��������(��Xc�+l���9�����[�
�X� ��5��E�*�O�      �#�X� �b'������gٽ;S��+l��T�j�H�3��i��վ����(���ĻdA?�p�B�.�@:�[�:/Q;�.;�;;�tB;=�E;��F;e�G;'�G;H;�FH;UkH;��H;\�H;F�H;��H;H�H;��H;/�H;��H;H�H;��H;F�H;^�H;��H;SkH;�FH;H;%�G;f�G;��F;;�E;�tB;�;;�.;.Q;�[�:6�@:p�B�bA?���Ļ(�����վ��i�H�3�T�j�+l��;S���gٽ����b'�X� �      �o��s��罯�ս9@��tĥ�{^���Xc�H�3���	�Ќ˼�]��XFB�[򻱜��eӺ���8��:�;�M#;�=5;:?;��C;�@F;=:G;(�G;O�G;h'H;�RH;�tH;�H;��H;b�H;�H;��H;	�H;}�H;	�H;��H;�H;a�H;��H;�H;�tH;�RH;h'H;M�G;)�G;<:G;�@F;�C;:?;�=5;�M#;�;��:���8eӺ����[�XFB��]��Ќ˼��	�H�3��Xc�{^��tĥ�9@����ս���s�      <S���r��v�����Փ����u���N���(��i�ό˼�A����P�ks��<|� ����\:P�:��;�n-;�:;�A;�,E;��F;coG;+�G;�H;8H;{_H;=~H;(�H;<�H;��H;K�H;��H;v�H;��H;t�H;��H;I�H;��H;?�H;(�H;<~H;x_H;8H;�H;-�G;aoG;��F;�,E;�A;�:;�n-;��;V�:�\: ���;|��ks���P��A��ό˼�i���(���N���u�Փ�����v���r��      s₽�؀���u��Xc���K�}1�������վ��]����P����DT����9���o�4�9�&�:p�	;x%;u�5;��>;ѻC;�F;�!G;ךG;�G;xH;�HH;lH;ׇH;��H;ͭH;�H;��H;��H;��H;�H;��H;��H;��H;�H;ЭH;��H;ׇH;lH;�HH;vH;	�G;ԚG;�!G;�F;ѻC;��>;r�5;x%;s�	;�&�:4�9��o���9�DT�������P��]���վ�����|1���K��Xc���u��؀�      7�6�K�3���+�
��e�p�����μ������XFB�ks�DT��(�D��{��P;u9�q�:���:�Y;
u0;�;;B;:E;�F;1hG;�G;A�G;�0H;�XH;hxH;Z�H;��H;=�H;3�H;�H;O�H;f�H;t�H;f�H;N�H;�H;3�H;>�H;��H;Z�H;exH;�XH;�0H;D�G;�G;.hG;�F; :E;B;�;;
u0;�Y;���:�q�:`;u9�{��(�D�DT��js�WFB�~��������μp���f�
����+�L�3�      v�����W�іռ־�/Ϥ��I����[�(�[����9��{��0<9pX�:�X�:XQ;W,;��8;�A@;5BD;�@F;�,G;��G;��G;�H;	EH;ZhH;o�H;��H;��H;��H;]�H;[�H;�H;��H;��H;��H;�H;X�H;]�H;��H;��H;��H;l�H;XhH;EH;�H;��G;��G;�,G;�@F;5BD;�A@;��8;Z,;WQ;�X�:tX�:P<9�{����9�� [�(���[��I��.Ϥ�־�іռ�W���      ny��Eݜ��A���I����s���P��%+������Ļ����<|���o�@;u9nX�:,�:n;�);�6;��>;�PC;��E;%�F;�xG;b�G;�H;�1H;QXH;=wH;�H;P�H;?�H;��H;T�H;}�H;��H;#�H;��H;#�H;��H;}�H;T�H;��H;?�H;O�H;�H;;wH;PXH;�1H;�H;_�G;�xG;&�F;��E;�PC;��>;��6;�);m;,�:pX�:@;u9��o�;|�������Ļ����%+���P���s��I���A��Fݜ�      [FB�B�>���4�[�$�x��[�����ݎ�bA?�eӺ��� 4�9�q�:}X�:n;��';�=5;��=;-�B;LGE;x�F;�UG;W�G;�G;�H;�HH;NjH;4�H;��H;��H;o�H;��H;�H;|�H;I�H;Z�H;�H;Z�H;I�H;{�H;�H;��H;o�H;��H;��H;4�H;JjH;�HH;�H;�G;T�G;�UG;u�F;MGE;-�B;��=;�=5;��';p;�X�:�q�: 4�9���dӺbA?��ݎ����[�x��Z�$���4�C�>�      �EֻQ�ѻ��ĻpT���񕻺.o�ҝ.�6ܺp�B� ��8�\:�&�:���:UQ;�);�=5;
;=;H#B;��D;vF; 7G;��G;��G;�H;�:H;N^H;�zH;6�H;��H;�H;F�H;�H;��H;X�H;��H;g�H;��H;e�H;��H;X�H;��H;�H;F�H;��H;��H;5�H;�zH;O^H;�:H;�H;��G;��G;7G;vF;��D;L#B;;=;�=5;�);WQ;���:�&�:�\:@��8h�B�9ܺҝ.��.o���pT����ĻW�ѻ      �A?��9� 9)��Z��ܺ�p��h����;9.�@:��:T�:q�	;�Y;V,;�6;��=;F#B;��D;�XF;"G;��G;S�G;�H;//H;�SH;�qH;�H;�H;��H;��H;��H;�H;��H;	�H;��H;W�H;��H;U�H;��H;	�H;��H;�H;��H;��H;��H;�H;�H;�qH;�SH;,/H;�H;S�G;��G;"G;�XF;��D;F#B;��=;�6;W,;�Y;q�	;V�:��::�@:�;9h���|p���ܺ�Z� 9)��9�      ��	������i���[��`5u9v:�j~:F��:�[�:�;��;z%;	u0;��8;��>;*�B;��D;�XF;gG;��G;��G;��G;.&H;AKH;�iH;!�H;ƗH;u�H;��H;E�H;��H;��H;��H;n�H;��H;�H;��H;�H;��H;m�H;��H;��H;��H;B�H;��H;u�H;ėH;"�H;�iH;>KH;+&H;��G;��G;��G;hG;�XF;��D;+�B;��>;��8;	u0;z%;��;�;�[�:B��:k~:�:�5u9`[���i������      �Y�:�o�:�W�:P�:M&�:���:���:Q�	;-Q;�M#;�n-;p�5;�;;�A@;�PC;FGE;vF;�!G;��G;�G;N�G;� H;IEH;�cH;x}H;��H;��H;ޱH;�H;��H;��H;f�H;��H;��H;��H;��H;*�H;��H;��H;��H;��H;g�H;��H;��H;��H;ܱH;�H;��H;z}H;�cH;DEH;� H;M�G;�G;��G;"G;vF;FGE;�PC;�A@;�;;p�5;�n-;�M#;.Q;Q�	;���:���:c&�:P�:�W�:po�:      ���:K% ;j�;��;$�;Q;@m;Vd';�.;�=5;�:;��>;�B;2BD;��E;w�F;7G;��G;��G;P�G;�H;$BH;E`H;�yH;��H;`�H;��H;�H;��H;�H;��H;j�H;��H;|�H;.�H;�H;��H;�H;.�H;|�H;��H;l�H;��H;�H;��H;�H;��H;a�H;��H;�yH;E`H;$BH;�H;Q�G;��G;��G;7G;u�F;��E;2BD;�B;��>; �:;�=5;�.;Vd';@m;Q;'�;��;f�;;% ;      �";�M#;(%;t�';D�+;^�/;��3;� 8;�;;=?;�A;ѻC; :E;�@F;&�F;�UG;��G;U�G;��G;� H;"BH;�^H;�wH;X�H;ÝH;�H;̷H;j�H;<�H;d�H;]�H;&�H;��H;�H;��H;��H;��H;��H;��H;�H;��H;&�H;]�H;`�H;9�H;l�H;ɷH;�H;ĝH;V�H;�wH;�^H;!BH;� H;��G;V�G;�G;�UG;'�F;�@F; :E;ѻC;�A;=?;�;;� 8;��3;^�/;\�+;t�';&%;�M#;      �46;|�6;l7;K�8;��:;l�<;P�>;p�@;�tB;~�C;�,E;�F;�F;�,G;�xG;V�G;��G;�H;.&H;JEH;E`H;�wH;m�H;s�H;��H;'�H;׿H;��H;�H;:�H;h�H;|�H;��H;��H;��H;��H;��H;��H;��H;��H;��H;{�H;h�H;7�H;�H;��H;ֿH;)�H;��H;p�H;m�H;�wH;B`H;LEH;.&H;�H;��G;T�G;�xG;�,G;�F;�F;�,E;~�C;�tB;o�@;P�>;o�<;��:;K�8;l7;n�6;      y@;bA@;8�@;'RA;�"B;C;[�C;��D;;�E;�@F;��F;�!G;+hG;��G;_�G;�G;�H;//H;@KH;�cH;�yH;W�H;p�H;�H;C�H;��H;��H;�H;N�H;��H;��H;��H;z�H;��H;�H;��H;��H;��H;�H;��H;x�H;��H;��H;��H;M�H;�H;��H;��H;F�H;��H;p�H;W�H;�yH;�cH;@KH;0/H;�H;�G;_�G;��G;+hG;�!G;��F;�@F;=�E;��D;Y�C;C;�"B;(RA;8�@;XA@;      ��D;!�D;�D;�9E;��E;M�E;nPF;�F;��F;::G;_oG;ךG;�G;��G;�H;�H;�:H;�SH;�iH;}H;��H;ǝH;��H;L�H;x�H;!�H;k�H;��H;��H;l�H; �H;F�H;��H;(�H;��H;]�H;��H;_�H;��H;'�H;��H;G�H; �H;j�H;��H;��H;l�H;!�H;x�H;I�H;��H;ɝH;��H;�}H;�iH;�SH;�:H;�H;�H;��G;�G;ؚG;`oG;9:G;��F;�F;oPF;M�E;��E;�9E;�D;!�D;      �F;ܯF;�F;��F;�F;�!G;�FG;RjG;c�G;(�G;)�G;	�G;@�G;�H;�1H;�HH;M^H;�qH;�H;��H;]�H;�H;$�H;��H;�H;L�H;[�H;��H;��H;��H;��H;��H;-�H;�H;��H;�H;I�H;�H;��H;�H;*�H;��H;��H;��H;��H;��H;\�H;L�H;�H;��H;$�H;�H;X�H;��H;�H;�qH;K^H;�HH;�1H;�H;A�G;�G;*�G;&�G;e�G;RjG;�FG;�!G;�F;��F;�F;үF;      �nG;,qG;xG;߂G;�G;W�G;x�G;��G;&�G;L�G;�H;{H;�0H;EH;PXH;NjH;�zH;�H;ƗH;��H;��H;̷H;ֿH;��H;e�H;_�H;}�H;��H;��H;��H;��H;�H; �H;��H;r�H;��H;��H;��H;q�H;��H;�H;�H;��H;��H;��H;��H;{�H;^�H;g�H;��H;ԿH;̷H;��H;��H;ƗH;�H;�zH;MjH;PXH;EH;�0H;{H;�H;L�G;)�G;��G;x�G;V�G;��G;݂G;xG;+qG;      �G;{�G;��G;�G;�G;3�G;$�G;�H;H;n'H;8H;�HH;�XH;[hH;=wH;4�H;5�H;�H;r�H;�H;�H;j�H;��H;�H;��H;��H;��H;y�H;��H;��H;��H;�H;��H;��H;�H;B�H;S�H;A�H;�H;��H;��H;�H;��H;��H;��H;x�H;��H;��H;��H;�H;��H;j�H;�H;�H;s�H;�H;3�H;4�H;>wH;ZhH;�XH;�HH;8H;n'H;H;�H;$�G;3�G;%�G;�G;��G;��G;      WH;RH;wH;�H;pH;�%H;�/H;�:H;�FH;�RH;x_H;lH;gxH;n�H;�H;��H;��H;��H;��H;�H;��H;;�H;�H;R�H;��H; �H;��H;��H;`�H;��H;�H;��H;��H; �H;��H;��H;��H;��H;��H; �H;��H;��H;�H;��H;`�H;��H;��H;��H;��H;R�H;�H;;�H;��H;�H;��H;��H;��H;��H;�H;n�H;hxH;
lH;v_H;�RH;�FH;�:H;�/H;�%H;vH;�H;vH;HH;      E@H;AH;nCH;4GH;oLH;�RH;2ZH;rbH;ZkH;�tH;D~H;�H;_�H;��H;S�H;��H;�H;��H;A�H;��H;�H;a�H;6�H;��H;b�H;��H;��H;��H;��H;�H;��H;��H;8�H;��H;��H;�H;�H;�H;��H;��H;4�H;��H;��H;�H;��H;��H;��H;��H;c�H;��H;4�H;a�H;�H;��H;B�H;��H;�H;��H;S�H;��H;_�H;�H;F~H;�tH;]kH;tbH;2ZH;�RH;kLH;4GH;hCH;AH;      gH;�gH;liH;QlH;>pH;uH;�zH;��H;ćH;�H;+�H;��H;��H;��H;A�H;v�H;J�H;��H;��H;��H;��H;]�H;h�H;��H;�H;��H;��H;��H;�H;��H;��H;C�H;��H;��H;�H;J�H;f�H;J�H;�H;��H;��H;E�H;��H;��H;�H;��H;��H;��H;�H;��H;e�H;]�H;��H;��H;��H;��H;J�H;u�H;A�H;��H;��H;��H;,�H;�H;ŇH;�H;�zH;uH;;pH;SlH;liH;�gH;      ��H;��H;[�H;��H;��H;7�H;��H;J�H;_�H;��H;A�H;ԭH;@�H;��H;��H;��H;�H;�H;��H;n�H;s�H;*�H;~�H;��H;A�H;��H;�H;�H;��H;��H;A�H;��H;��H;<�H;e�H;��H;��H;��H;e�H;<�H;��H;��H;A�H;��H;��H;�H;�H;��H;D�H;��H;{�H;*�H;p�H;p�H;��H;�H;�H;��H;��H;��H;@�H;ԭH;B�H;��H;a�H;H�H;��H;:�H;�H;��H;\�H;��H;      i�H;ΚH;ЛH;t�H;��H;{�H;��H;p�H;J�H;a�H;��H;�H;5�H;`�H;V�H;�H;��H;��H;��H;��H;��H;��H;��H;�H;��H;/�H;$�H;��H;��H;?�H;��H;��H;?�H;w�H;��H;��H;��H;��H;��H;w�H;<�H;��H;��H;A�H;��H;��H; �H;-�H;��H;�H;��H;��H;��H;��H;��H;��H;��H;�H;T�H;`�H;3�H;�H;��H;b�H;J�H;o�H;��H;~�H;��H;t�H;ЛH;ǚH;      ԩH;$�H;ӪH;"�H;�H;�H;��H;��H;��H;�H;O�H;��H;�H;^�H;��H;��H;]�H;�H;o�H;��H;��H;�H;��H;��H; �H;�H;��H;��H;�H;��H;��H;<�H;p�H;��H;��H;��H;��H;��H;��H;��H;o�H;?�H;��H;��H; �H;��H;��H;�H;!�H;��H;��H;�H;��H;��H;o�H;	�H;\�H;��H;��H;^�H;�H;��H;N�H;�H;��H;��H;��H;�H;٭H;"�H;ժH;�H;      �H;d�H;��H;�H;��H;<�H;c�H;ǽH;O�H;��H;��H;��H;S�H;�H;��H;P�H;��H;��H;��H;��H;6�H;��H;��H;�H;��H;��H;n�H;�H;��H;��H;�H;h�H;��H;��H;��H;��H;��H;��H;��H;��H;��H;j�H;�H;��H;��H;�H;m�H;��H;��H;	�H;��H;��H;5�H;��H;��H;��H;��H;P�H;��H;�H;R�H;��H;��H;��H;O�H;ĽH;c�H;@�H;��H;�H; �H;[�H;      ��H;3�H;ѺH;˻H;�H;��H;i�H;z�H;��H;�H;{�H;��H;i�H;��H;&�H;_�H;m�H;P�H;�H;��H;%�H;��H;��H;��H;X�H;�H;��H;A�H;��H;�H;I�H;��H;��H;��H;��H;��H;��H;��H;��H;��H;��H;��H;I�H;�H;��H;A�H;��H;�H;Y�H;��H;��H;��H;$�H;��H;�H;Q�H;k�H;_�H;&�H;��H;i�H;��H;z�H;
�H;��H;w�H;h�H;��H;�H;˻H;ӺH;+�H;      ��H;�H;��H;��H;ʾH;<�H;�H;�H;9�H;|�H;��H;#�H;u�H;��H;��H;�H;��H;��H;��H;/�H;��H;��H;��H;��H;��H;D�H;��H;W�H;��H;�H;h�H;��H;��H;��H;��H;��H;��H;��H;��H;��H;��H;��H;h�H; �H;��H;W�H;��H;E�H;��H;��H;��H;��H;��H;/�H;��H;��H;��H;�H;��H;��H;u�H;#�H;��H;~�H;9�H;�H;�H;A�H;��H;��H;��H;�H;      ��H;5�H;ѺH;˻H;�H;��H;i�H;z�H;��H;�H;{�H;��H;i�H;��H;&�H;_�H;m�H;P�H;�H;��H;'�H;��H;��H;��H;Y�H;�H;��H;A�H;��H;�H;I�H;��H;��H;��H;��H;��H;��H;��H;��H;��H;��H;��H;I�H;�H;��H;A�H;��H;�H;X�H;��H;��H;��H;$�H;��H;�H;Q�H;k�H;_�H;&�H;��H;i�H;��H;{�H;	�H;��H;w�H;i�H;��H;�H;˻H;ϺH;(�H;      �H;d�H;��H;�H;��H;<�H;c�H;ǽH;O�H;��H;��H;��H;S�H;�H;��H;P�H;��H;��H;��H;��H;9�H;��H;��H;�H;��H;��H;n�H;�H;��H;��H;�H;h�H;��H;��H;��H;��H;��H;��H;��H;��H;��H;l�H;�H;��H;��H;�H;m�H;��H;��H;�H;��H;��H;4�H;��H;��H;��H;��H;P�H;��H;�H;S�H;��H;��H;��H;O�H;ĽH;c�H;@�H;��H;�H;��H;[�H;      թH;$�H;ժH;"�H;�H;�H;��H;��H;��H;�H;O�H;��H;�H;^�H;��H;��H;]�H;�H;o�H;��H;��H;�H;��H;��H;!�H;�H;��H;��H;�H;��H;��H;<�H;p�H;��H;��H;��H;��H;��H;��H;��H;o�H;?�H;��H;��H; �H;��H;��H;�H; �H;��H;��H;�H;��H;��H;o�H;	�H;\�H;��H;��H;^�H;�H;��H;O�H;�H;��H;��H;��H;�H;حH;"�H;ժH;�H;      k�H;ΚH;ЛH;v�H;��H;{�H;��H;o�H;J�H;a�H;��H;�H;3�H;`�H;T�H;�H;��H;��H;��H;��H;��H;��H;��H;�H;��H;.�H;"�H;��H;��H;?�H;��H;��H;=�H;v�H;��H;��H;��H;��H;��H;v�H;<�H;��H;��H;A�H;��H;��H;!�H;.�H;��H;~�H;��H;��H;��H;��H;��H;��H;��H;�H;U�H;`�H;3�H;�H;��H;b�H;J�H;l�H;��H;�H;��H;v�H;ϛH;ʚH;      ��H;��H;\�H;��H;��H;7�H;��H;J�H;_�H;��H;A�H;ԭH;@�H;��H;��H;��H;�H;�H;��H;q�H;v�H;*�H;~�H;��H;D�H;��H;�H;�H;��H;��H;A�H;��H;��H;<�H;e�H;��H;��H;��H;e�H;<�H;��H;��H;A�H;��H;��H;�H;�H;��H;A�H;��H;|�H;*�H;q�H;n�H;��H;�H;�H;��H;��H;��H;@�H;ԭH;A�H;��H;a�H;H�H;��H;9�H;}�H;��H;]�H;��H;      gH;�gH;liH;SlH;>pH;uH;�zH;��H;ŇH;�H;,�H;��H;��H;��H;A�H;v�H;J�H;��H;��H;��H;��H;]�H;h�H;��H;�H;��H;��H;��H;�H;��H;��H;C�H;��H;��H;�H;J�H;f�H;J�H;�H;��H;��H;E�H;��H;��H;�H;��H;��H;��H;�H;��H;e�H;]�H;��H;��H;��H;��H;H�H;v�H;A�H;��H;��H;��H;)�H;�H;ŇH;�H;�zH;uH;;pH;QlH;liH;�gH;      ?@H;	AH;mCH;4GH;kLH;�RH;5ZH;ubH;\kH;�tH;D~H;�H;^�H;��H;S�H;��H;�H;��H;A�H;��H;�H;a�H;6�H;��H;c�H;��H;��H;��H;��H;�H;��H;��H;7�H;��H;��H;�H;�H;�H;��H;��H;7�H;��H;��H;�H;��H;��H;��H;��H;b�H;��H;4�H;a�H;�H;��H;A�H;��H;�H;��H;S�H;��H;_�H;�H;D~H;�tH;^kH;ubH;5ZH;�RH;iLH;6GH;kCH;AH;      PH;NH;}H;�H;tH;�%H;�/H;�:H;�FH;�RH;x_H;lH;gxH;n�H;�H;��H;��H;��H;��H;�H;��H;;�H;�H;Q�H;��H; �H;��H;��H;`�H;��H;�H;��H;��H; �H;��H;��H;��H;��H;��H; �H;��H;��H;�H;��H;`�H;��H;��H;��H;��H;R�H;�H;;�H;��H;�H;��H;��H;��H;��H;�H;n�H;gxH;lH;x_H;�RH;�FH;�:H;�/H;�%H;qH;�H;}H;OH;      �G;{�G;��G;�G;�G;3�G;$�G;�H;H;n'H;
8H;�HH;�XH;[hH;>wH;4�H;5�H;�H;s�H;�H;"�H;j�H;��H;�H;��H;��H;��H;x�H;��H;��H;��H;�H;��H;��H;�H;B�H;S�H;B�H;�H;��H;��H;�H;��H;��H;��H;y�H;��H;��H;��H;�H;��H;j�H;�H;�H;r�H;�H;3�H;5�H;=wH;XhH;�XH;�HH;8H;n'H;H;�H;$�G;0�G;%�G;�G;��G;��G;      �nG;.qG;xG;؂G;�G;S�G;v�G;��G;&�G;M�G;�H;{H;�0H;EH;PXH;NjH;�zH;�H;ƗH;��H;��H;̷H;ֿH;��H;g�H;_�H;~�H;��H;��H;��H;��H;�H; �H;��H;q�H;��H;��H;��H;r�H;��H;�H;�H;��H;��H;��H;��H;{�H;_�H;e�H;��H;ԿH;̷H;��H;��H;ƗH;�H;�zH;MjH;PXH;EH;�0H;{H;�H;M�G;&�G;��G;v�G;R�G;�G;؂G;xG;$qG;      �F;دF;�F;��F;�F;�!G;�FG;UjG;b�G;(�G;*�G;�G;A�G;�H;�1H;�HH;M^H;�qH;�H;��H;^�H;�H;$�H;��H;�H;L�H;^�H;��H;��H;��H;��H;��H;+�H;�H;��H;�H;I�H;�H;��H;�H;*�H;��H;��H;��H;��H;��H;[�H;L�H;�H;��H;$�H;�H;X�H;��H;�H;�qH;K^H;�HH;�1H;�H;@�G;	�G;*�G;&�G;c�G;RjG;�FG;�!G;�F;��F;�F;ίF;      ��D;!�D;�D;�9E;��E;M�E;oPF;�F;��F;::G;aoG;ؚG;�G;��G;�H;�H;�:H;�SH;�iH;�}H;ÎH;ɝH;��H;L�H;x�H; �H;n�H;��H;��H;l�H; �H;F�H;��H;'�H;��H;_�H;��H;]�H;��H;'�H;��H;H�H; �H;j�H;��H;��H;k�H;!�H;x�H;J�H;��H;ǝH;��H;�}H;�iH;�SH;�:H;�H;�H;��G;�G;ךG;_oG;9:G;��F;�F;nPF;M�E;��E;�9E;�D;!�D;      @;_A@;>�@;%RA;�"B;C;X�C;��D;=�E;�@F;��F;�!G;-hG;��G;_�G;�G;�H;-/H;@KH;�cH;�yH;W�H;r�H;�H;F�H;��H;��H;�H;O�H;��H;��H;��H;z�H;��H;�H;��H;��H;��H;�H;��H;x�H;��H;��H;��H;K�H;�H;��H;��H;C�H;��H;o�H;W�H;�yH;�cH;@KH;0/H;�H;�G;_�G;��G;+hG;�!G;��F;�@F;=�E;��D;X�C;C;�"B;%RA;;�@;UA@;      �46;��6;/l7;K�8;��:;q�<;T�>;p�@;�tB;~�C;�,E;�F;�F;�,G;�xG;V�G;��G;�H;.&H;JEH;H`H;�wH;n�H;s�H;��H;(�H;ٿH;��H;�H;:�H;h�H;{�H;��H;��H;��H;��H;��H;��H;��H;��H;��H;|�H;h�H;7�H;�H;��H;ԿH;(�H;��H;r�H;m�H;�wH;B`H;LEH;.&H;�H;��G;V�G;�xG;�,G;�F;�F;�,E;{�C;�tB;o�@;V�>;q�<;��:;J�8;#l7;y�6;      �";�M#;*%;t�';F�+;^�/;��3;� 8;�;;=?;�A;ѻC; :E;�@F;&�F;�UG;�G;S�G;��G;� H;$BH;�^H;�wH;Z�H;ĝH;�H;̷H;l�H;=�H;d�H;]�H;&�H;��H;�H;��H;��H;��H;��H;��H;�H;��H;&�H;]�H;`�H;8�H;j�H;ɷH;�H;ÝH;V�H;�wH;�^H;"BH;� H;��G;V�G;�G;�UG;'�F;�@F; :E;һC;�A;=?;�;;� 8;��3;^�/;\�+;t�';'%;�M#;      ���:F% ;n�;��;$�;Q;Dm;Yd';�.;�=5;�:;��>;�B;2BD;��E;u�F;7G;��G;��G;P�G;�H;$BH;F`H;�yH;��H;a�H;��H;�H;��H;�H;��H;j�H;��H;{�H;.�H;�H;��H;�H;.�H;|�H;��H;m�H;��H;�H;��H;�H;��H;`�H;��H;�yH;C`H;$BH;�H;P�G;��G;��G;7G;u�F;��E;2BD;�B;��>; �:;�=5;�.;Xd';Cm;Q;+�;��;l�;:% ;      �Y�:�o�:�W�:L�:U&�:���:���:R�	;.Q;�M#;�n-;p�5;�;;�A@;�PC;FGE;vF; "G;��G;�G;P�G;� H;IEH;�cH;z}H;��H;�H;ܱH;�H;��H;��H;f�H;��H;��H;��H;��H;*�H;��H;��H;��H;��H;g�H;��H;��H;��H;ޱH;�H;��H;x}H;�cH;FEH;� H;L�G;�G;��G; "G;vF;FGE;�PC;�A@;�;;o�5;�n-;�M#;.Q;R�	;���:���:c&�:L�:�W�:po�:      ��	������i��`[��p5u9v:k~:F��:�[�:�;��;z%;	u0;��8;��>;+�B;��D;�XF;hG;��G;��G;��G;/&H;AKH;�iH;�H;ƗH;u�H;��H;E�H;��H;��H;��H;m�H;��H;�H;��H;�H;��H;n�H;��H;��H;��H;B�H;��H;u�H;ŗH;"�H;�iH;>KH;)&H;��G;��G;��G;gG;�XF;��D;*�B;��>;��8;	u0;z%;��;�;�[�:F��:�j~:�:�5u9�[���i������      �A?��9� 9)��Z��ܺ�p��h����;9.�@:��:V�:q�	;�Y;U,;�6;��=;H#B;��D;�XF;"G;��G;S�G;�H;0/H;�SH;�qH;�H;�H;��H;��H;��H;�H;��H;	�H;��H;U�H;��H;U�H;��H;	�H;��H;�H;��H;��H;��H;�H;�H;�qH;�SH;*/H;�H;S�G;��G;"G;�XF;��D;E#B;��=;�6;U,;�Y;q�	;T�:��::�@:�;9h���|p���ܺ�Z�!9)��9�      �EֻR�ѻ��ĻpT���񕻻.o�ҝ.�6ܺp�B�@��8�\:�&�:���:WQ;�);�=5;;=;I#B;��D;vF; 7G;��G;��G;�H;�:H;N^H;�zH;5�H;��H;�H;F�H;�H;��H;X�H;��H;g�H;��H;g�H;��H;Y�H;��H;�H;F�H; �H;��H;6�H;�zH;O^H;�:H;�H;��G;��G;7G;vF;��D;J#B;
;=;�=5;�);UQ;���:�&�:�\:���8l�B�9ܺҝ.��.o���pT����ĻW�ѻ      \FB�B�>���4�Z�$�x��[�����ݎ�bA?�bӺ���4�9�q�:}X�:p;��';�=5;��=;-�B;MGE;w�F;�UG;W�G;�G;�H;�HH;MjH;4�H;��H;��H;o�H;��H;�H;{�H;I�H;Z�H;�H;Z�H;I�H;|�H;�H;��H;o�H;��H;��H;4�H;KjH;�HH;�H;�G;T�G;�UG;u�F;LGE;-�B;��=;�=5;��';p;{X�:�q�: 4�9���fӺbA?��ݎ����[�x��[�$���4�D�>�      ny��Eݜ��A���I����s���P��%+������Ļ����<|���o�@;u9pX�:,�:m;�);�6;��>;�PC;��E;&�F;�xG;d�G;�H;�1H;QXH;;wH;�H;P�H;?�H;��H;U�H;}�H;��H;#�H;��H;#�H;��H;~�H;T�H;��H;?�H;O�H;�H;=wH;PXH;�1H;�H;^�G;�xG;%�F;��E;�PC;��>;��6;�);n;,�:nX�:@;u9��o�<|�������Ļ����%+���P���s��I���A��Fݜ�      v�����W�іռ־�/Ϥ��I����[�(� [����9��{��@<9tX�:�X�:XQ;Y,;��8;�A@;3BD;�@F;�,G;��G;��G;�H;	EH;XhH;n�H;��H;��H;��H;_�H;Z�H;�H;��H;��H;��H;�H;Z�H;\�H;��H;��H;��H;n�H;ZhH;EH;�H;��G;��G;�,G;�@F;6BD;�A@;��8;Z,;WQ;�X�:pX�: <9�{����9�� [�(���[��I��.Ϥ�־�іռ�W���      7�6�K�3���+�
��e�p�����μ���~���XFB�js�DT��(�D��{��`;u9�q�:���:�Y;
u0;�;;B; :E;�F;2hG;�G;C�G;�0H;�XH;gxH;Z�H;��H;=�H;3�H;�H;N�H;f�H;t�H;f�H;O�H;�H;2�H;>�H;��H;Z�H;exH;�XH;�0H;D�G;�G;+hG;�F;:E;B;�;;
u0;�Y;���:�q�:P;u9�{��(�D�DT��ks�XFB�~��������μp���e�
����+�L�3�      s₽�؀���u��Xc���K�|1�������վ��]����P����DT����9���o�4�9�&�:q�	;x%;s�5;��>;ѻC;�F;�!G;ԚG;�G;xH;�HH;lH;ׇH;��H;ͭH;�H;��H;��H;��H;�H;��H;��H;��H;�H;έH;��H;ׇH;lH;�HH;xH;�G;ךG;�!G;�F;ѻC;��>;s�5;x%;s�	;�&�: 4�9��o���9�DT�������P��]���վ�����|1���K��Xc���u��؀�      <S���r��v�����Փ����u���N���(��i�ό˼�A����P�ks��;|� ����\:T�:��;�n-;�:;�A;�,E;��F;aoG;-�G;�H;8H;{_H;=~H;(�H;;�H;��H;I�H;��H;v�H;��H;v�H;��H;K�H;��H;?�H;(�H;<~H;x_H;8H;�H;+�G;coG;��F;�,E;�A;�:;�n-;��;V�:�\:���;|��ks���P��A��ό˼�i���(���N���u�Փ�����v���r��      �o��s��罯�ս9@��tĥ�{^���Xc�H�3���	�Ќ˼�]��XFB�[򻰜��eӺ ��8��:�;�M#;�=5;:?;��C;�@F;<:G;)�G;O�G;h'H;�RH;�tH;�H;��H;b�H;�H;��H;	�H;}�H;	�H;��H;�H;a�H;��H;�H;�tH;�RH;h'H;M�G;(�G;=:G;�@F;�C;:?;�=5;�M#;�;��:���8fӺ����[�XFB��]��Ќ˼��	�H�3��Xc�{^��tĥ�9@����ս���s�      �#�X� �b'������gٽ;S��+l��T�j�H�3��i��վ����(���ĻbA?�h�B�2�@:�[�:/Q;�.;�;;�tB;>�E;��F;f�G;'�G;H;�FH;SkH;��H;\�H;G�H;��H;H�H;��H;/�H;��H;F�H;��H;D�H;\�H;��H;SkH;�FH;H;%�G;e�G;��F;:�E;�tB;�;;�.;.Q;�[�:6�@:x�B�dA?���Ļ(�����վ��i�H�3�T�j�+l��;S���gٽ����b'�X� �      �S�*�O��E��5�X� �[�
���罨9��+l���Xc���(��������[�����ݎ�5ܺ�;9H��:T�	;Vd';� 8;p�@;��D;�F;VjG;��G;�H;�:H;nbH;�H;C�H;i�H;~�H;��H;p�H;�H;q�H;��H;~�H;f�H;C�H;�H;nbH;�:H;�H;��G;SjG;�F;��D;p�@;� 8;Yd';R�	;F��:�;9;ܺ�ݎ������[��������(��Xc�+l���9�����[�
�X� ��5��E�*�O�      �~��*��,�v��9b�}�H�#,�PZ����;S��{^����N������μ�I���%+����֝.�`����j~:���::m;��3;M�>;W�C;qPF;�FG;t�G; �G;�/H;.ZH;�zH;��H;��H;��H;\�H;^�H;�H;`�H;Z�H;��H;��H;��H;�zH;,ZH;�/H; �G;r�G;�FG;rPF;R�C;L�>;��3;=m;���:�j~:X���؝.�����%+��I����μ�����N�{^��;S�����PZ�#,�}�H��9b�,�v�*��      ����+����:���M��I�r�*�O�#,�[�
��gٽtĥ���u�|1�q���/Ϥ���P�[�.o�lp��n:���:Q;U�/;l�<;C;J�E;�!G;U�G;4�G;�%H;�RH;uH;4�H;|�H;�H;?�H;��H;;�H;��H;=�H;�H;z�H;7�H;uH;�RH;�%H;4�G;S�G;�!G;J�E;C;l�<;U�/;Q;���:r:jp���.o�[򻲎P�/Ϥ�q���|1���u�tĥ��gٽ[�
�#,�*�O�I�r��M���:��+���      :���v��O;������UP��I�r�}�H�X� ���9@��Փ����K�e�־���s�x���񕻥ܺ�5u9O&�:'�;D�+;��:;�"B;��E;�F;�G;�G;sH;`LH;1pH;|�H;��H;ۭH;r�H;�H;��H;�H;q�H;٭H;��H;}�H;3pH;]LH;pH;�G;�G;�F;��E;�"B;��:;D�+;*�;O&�:�5u9�ܺ��x����s�־�e���K�Փ��9@����X� �}�H�I�r�UP������O;���v��      YVھ�*־25ʾu��������M���9b��5�����ս����Xc�
��Җռ�I��[�$�oT���Z��[��P�:�;}�';R�8;,RA;�9E;��F;܂G;�G;�H;2GH;HlH;��H;p�H;�H;��H;ɻH;��H;ɻH;��H;�H;o�H;��H;HlH;/GH;�H;�G;܂G;��F;�9E;'RA;W�8;}�';�;L�:�[���Z�pT��[�$��I��Җռ
���Xc������ս���5��9b��M������u���25ʾ�*־      ���쾶�޾25ʾP;���:��,�v��E�b'����v����u���+��W��A����4���Ļ#9)�0j���W�:`�;%;l7;1�@;�D;�F;xG;��G;xH;eCH;aiH;Q�H;țH;ڪH;��H;ʺH;��H;ʺH;��H;ڪH;ƛH;Q�H;aiH;cCH;vH;��G;xG;�F;�D;-�@;l7;%;b�;�W�:0j��"9)���Ļ��4��A���W缈�+���u�v�����b'��E�,�v��:��P;��25ʾ��޾��      Zh���b���쾪*־�v��+���*��*�O�X� �s��r���؀�L�3���Eݜ�B�>�W�ѻ�9�����`o�:=% ;�M#;y�6;YA@;�D;үF;,qG;z�G;VH;AH;�gH;�H;ĚH;�H;P�H;,�H;�H;,�H;Q�H;�H;ÚH;�H;�gH;AH;TH;z�G;+qG;үF;�D;TA@;�6;�M#;>% ;^o�:�����9�X�ѻB�>�Eݜ���L�3��؀��r��s�X� �*�O�*��+����v���*־���b��      ���
^�X_ݾ��ɾl*���{x�)G�R,�����b��d@{���/�����䙼�J;�P�ͻ��4��V�L��:8;��#;S�6;[@;^�D;ܱF;�lG;��G;H;�:H;�bH;!�H;c�H;j�H;�H;*�H;�H;*�H;�H;j�H;a�H;$�H;�bH;�:H;|H;��G;�lG;ܱF;^�D;[@;V�6;��#;9;H��:�V���4�R�ͻ�J;��䙼����/�d@{��b�����R,�)G�{x��l*����ɾX_ݾ
^�      
^�7���:پ~�žj�����9t�s�C������誫�]`w�L-����/`����7�9Sɻ�K/��xƹ���:�/;�f$;�7;�~@;y�D;��F;�nG;%�G;hH;�;H;�cH;��H;��H;��H;G�H;a�H;Y�H;a�H;H�H;��H;��H;��H;�cH;�;H;eH;%�G;�nG;��F;y�D;�~@;�7;�f$;�/;�:�xƹ�K/�:Sɻ��7�/`�����L-�]`w�誫������s�C�9t���j���~�ž�:پ7��      X_ݾ�:پ�V;+���Ƥ�Na����g��$:��Z�tݽ�ƣ��l�j.%��߼l���9.�ʹ��SV��0p�5A�:x;_(&;j�7;I�@;-E;.�F;�uG;S�G;�H;>H;�eH;	�H;��H;��H;�H;�H;�H;�H;�H;��H;��H;
�H;�eH;>H;�H;S�G;�uG;.�F;-E;C�@;m�7;^(&;x;1A�:�0p�RV�δ���9.�l���߼j.%��l��ƣ�tݽ�Z��$:���g�Na���Ƥ�+���V;�:پ      ��ɾ~�ž+��sת��#�����T��J+�=��2̽�s���yZ����Tμky����^Ϩ�P,� .�6W��: �
;r�(;�N9;�A;�NE;u�F;�G;�G;�H;�AH;lhH;+�H;w�H;�H;�H;ܹH;��H;ܹH;�H;�H;u�H;+�H;khH;�AH;�H;�G;�G;u�F;�NE;�A;�N9;p�(;�
;S��: .�6O,�^Ϩ���ky��Sμ����yZ��s���2̽=��J+���T�#����sת�+��~�ž      l*��j����Ƥ���/��B�c��G=����zｔж��ɇ�V�C���)"��y;k��&��-��o�˺�Y�9���:9;i,;�	;;QB;��E;G;��G;�G;�H;9GH;�lH;A�H;ќH;ϫH;w�H;;�H;�H;;�H;v�H;ͫH;МH;B�H;�lH;6GH;�H;�G;��G;G;��E;QB;�	;;i,;9;���:�Y�9n�˺�-���&�y;k�)"����V�C��ɇ��ж��z����G=�B�c��/����Ƥ�j���      ����Na��#���B�c�t�C�}#� ��VvϽ�����l�ig*����
���I���軼\c�퀺u,:6��:��;�_0;��<;�1C;�E;�#G;t�G;A�G;O H;�MH;qqH;�H;��H;�H;h�H;ּH;��H;ּH;j�H;�H;��H;�H;qqH;�MH;J H;A�G;s�G;�#G;�E;�1C;��<;�_0; �;4��:�t,:퀺�\c�����I��
�����ig*��l�����VvϽ ��}#�s�C�B�c�#���Na����      {x�9t���g���T��G=�}#�6�sݽ�b������GG�����Ǽly��O�$�h����$��uƹr��:'�:š ;h4;��>;jD;�[F;�FG;��G;9�G;@*H;�UH;2wH;:�H;!�H;��H;��H;��H;e�H;��H;��H;��H;!�H;<�H;3wH;�UH;=*H;9�G;��G;�FG;�[F;fD;��>;h4;ǡ ;'�:r��:�uƹ�$�h���O�$�ly���Ǽ���GG������b��sݽ6�}#��G=���T���g�9t�      )G�s�C��$:��J+��� ��sݽ`���0I���yZ���"����׫��jT��� �M����˺m9dٶ:��;`(;.�8;��@;��D;�F;�hG;��G;�H;p5H;(^H;�}H;'�H;��H;��H;�H;��H;r�H;��H;�H;��H;�H;*�H;�}H;(^H;l5H;�H;��G;�hG;�F;��D;��@;.�8;`(;��;dٶ: m9��˺M���� �iT�׫�������"��yZ�0I��a���sݽ �����J+��$:�s�C�      R,����Z�=��z�VvϽ�b��0I��k]a�K-�l� �&"���{�I�!�������4�lP(�6oQ:�L�:$�;��/;�'<;�B;�E;�F;ɇG;��G;lH;{AH;HgH;��H;q�H;�H;ҶH;��H;3�H;��H;3�H;��H;ҶH;�H;r�H;��H;GgH;xAH;jH;��G;ɇG;�F;�E;�B;�'<;�/;"�;�L�::oQ:lP(���4�����I�!�~�{�&"��l� �K-�k]a�1I���b��VvϽ�z�=��Z���      ������tݽ�2̽�ж����������yZ�K-�ٷ�4aļ\O���J;����}�|���º�O@9ガ:X�;�f$;��5;�N?;pD;�LF;1;G;ۤG;'�G;�!H;NH;�pH;ƋH;�H;d�H;)�H;~�H;��H;��H;��H;~�H;)�H;c�H;�H;ƋH;�pH;NH;�!H;%�G;ܤG;0;G;�LF;nD;�N?;��5;�f$;X�;炬:pO@9��º|�|�����J;�\O��4aļٷ�K-��yZ����������ж��2̽tݽ���      �b��誫��ƣ��s���ɇ��l�GG���"�l� �3aļf���I��C��ۙ�@��tƹ��k:���:+�;k>.;;
;;��A;BE;��F;GmG;��G;��G;�2H;&[H;�zH;�H;ɥH;ͳH;��H;k�H;8�H;N�H;8�H;k�H;��H;̳H;ͥH;�H;�zH;"[H;�2H;��G;��G;DmG;��F;
BE;��A;:
;;i>.;+�;���:��k:�tƹ?��ۙ��C��I�f��3aļl� ���"�GG��l��ɇ��s���ƣ�誫�      d@{�]`w��l��yZ�V�C�ig*�������'"��\O���I�A|�;Ϩ�lK/�X$T�jQ:���:��;�(&;$6;�%?;��C;�#F;+$G;X�G;��G;�H;dCH; hH;��H;��H;��H;"�H;-�H;]�H;��H;��H;��H;^�H;+�H; �H;��H;��H;��H;hH;dCH;�H;��G;U�G;*$G;�#F;��C;�%?;$6;�(&;��;���:nQ:X$T�jK/�;Ϩ�A|��I�\O��'"����鼲��ig*�V�C��yZ��l�^`w�      ��/�K-�j.%����������Ǽث��~�{��J;��C�<Ϩ�FO:������[�9���:�;��;_.1;.(<;�5B;OE;E�F;dfG;�G;n�G;/+H;TH;uH;X�H;��H;Z�H;��H;��H;$�H;8�H;]�H;8�H;"�H;��H;��H;[�H;��H;Y�H;uH;TH;,+H;p�G;�G;afG;B�F;OE;�5B;-(<;_.1;��;�;���:�[�9����FO:�;Ϩ��C��J;�~�{�ث���Ǽ��������j.%�K-�      ������߼Sμ("���
��ky��iT�I�!���軿ۙ�jK/������m9B�:���:N�;[�,;�N9;q@;�^D;�LF;�.G;�G;��G;H;�?H;TdH;T�H;��H;D�H;նH;��H;�H;�H;��H;��H;��H;�H;�H;��H;ضH;F�H;��H;S�H;VdH;�?H;H;��G;�G;�.G;�LF;�^D;q@;�N9;^�,;L�;���:B�:�m9����iK/��ۙ����H�!�iT�ky���
��)"��Sμ�߼���      �䙼0`��l��ky��z;k��I�P�$��� �����|�|�@�\$T��[�9B�:���::�;9�);E7;�>;�tC;E�E;�F;vG;R�G;��G;>,H;�SH;�sH;H;��H;J�H;�H;��H;r�H;��H;/�H;�H;/�H;��H;t�H;��H;�H;L�H;��H;��H;�sH;�SH;?,H;��G;N�G;vG;�F;E�E;�tC;�>;H7;7�);:�;���:B�:�[�9X$T�@�z�|������� �P�$��I�z;k�ky��l��0`��      �J;���7��9.����&����f���M����4���º�tƹjQ:���:���::�;��(;��5;��=;��B;�[E;r�F;UG;ߩG;��G;�H;�CH;NfH;�H;��H;.�H;ȶH; �H;��H;��H;5�H;v�H;^�H;v�H;5�H;��H;��H;�H;ʶH;/�H;��H;�H;MfH;�CH;�H;��G;کG;UG;o�F;�[E;��B;��=;��5;��(;:�;���:���:jQ:�tƹ��º��4�M��f�����軬&����9.���7�      P�ͻ3Sɻʹ��`Ϩ��-���\c��$���˺pP(��O@9��k:���:�;L�;:�);��5;n�=;GQB;�E;"�F;X8G;t�G;��G;�	H;�5H;�YH;�wH;�H;�H;�H;μH;��H;��H;^�H;��H;��H;`�H;��H;��H;_�H;��H;��H;μH;�H;�H;�H;|wH;�YH;�5H;�	H;}�G;t�G;W8G;#�F;�E;KQB;o�=;��5;:�);L�;�;���:��k:�O@9hP(���˺�$��\c��-��`Ϩ�ʹ��9Sɻ      ��4��K/�QV�L,�x�˺퀺�uƹ�m92oQ:催:���:��;��;X�,;C7;��=;DQB;��D;�cF;R$G; �G;�G;�G;�)H;�NH;nH;�H;�H;d�H;P�H;N�H;�H;��H;�H;�H;��H;Q�H;��H;�H;�H;��H;�H;N�H;O�H;c�H;�H;�H;nH;�NH;�)H;�G;�G;��G;T$G;�cF;��D;EQB;��=;E7;[�,;��;��;���:炬:>oQ:�m9�uƹ퀺j�˺L,�RV��K/�      �VṨxƹ 0p� 0�6pY�9u,:|��:`ٶ:�L�:X�;,�;�(&;_.1;�N9;�>;��B;�E;�cF;G;d�G;��G;�G;� H;(FH;�eH;�H;��H;�H;��H;žH;L�H;�H;��H;��H;*�H;��H;��H;��H;+�H;��H;��H;�H;K�H;þH;�H;�H;��H;�H;�eH;$FH;� H;�G;�G;e�G;G;�cF;�E;��B;�>;�N9;_.1;�(&;,�;X�;�L�:`ٶ:|��:"u,:�Y�9 0�6 0p��xƹ      N��:��:5A�:W��:���:0��:'�:��; �;�f$;h>.;$6;)(<;h@;�tC;�[E;�F;N$G;`�G;�G;S�G;�H;@H;�_H;0zH;��H;^�H;��H;r�H;��H;��H;��H;��H;��H;�H;:�H;��H;:�H;�H;��H;��H;��H;��H;��H;m�H;��H;[�H;��H;0zH;�_H;@H;�H;P�G;�G;`�G;P$G;�F;�[E;�tC;h@;)(<;$6;i>.;�f$;"�;��;'�:6��:���:W��:3A�:��:      B;�/;x;��
;9;�;ȡ ;`(;�/;��5;7
;;�%?;�5B;�^D;B�E;q�F;W8G; �G;��G;V�G;	H;�<H;�[H;(vH;ŋH;��H;y�H;}�H;��H;��H;��H;��H;J�H;��H;��H;��H;�H;��H;��H;��H;I�H;��H;��H;��H;��H;|�H;w�H;��H;ŋH;$vH;�[H;�<H;H;V�G;��G;�G;U8G;q�F;B�E;�^D;�5B;�%?;6
;;��5;�/;`(;ˡ ;�;9;��
;x;�/;      ��#;�f$;n(&;i�(;i,;�_0;r4;5�8;�'<;�N?;��A;��C;OE;�LF;�F;UG;t�G;�G;�G;�H;�<H;�ZH;tH;8�H;ߚH;ʩH;�H;�H;��H;V�H;|�H;q�H;��H;��H;+�H;�H;S�H;�H;+�H;��H;��H;o�H;}�H;R�H;��H;�H;�H;˩H;��H;4�H;tH;�ZH;�<H;�H;�G;!�G;s�G;UG; �F;�LF;OE;��C;��A;�N?;�'<;5�8;r4;�_0;i,;i�(;l(&;�f$;      [�6;�7;m�7;�N9;�	;;��<;��>;��@;�B;mD;BE;�#F;B�F;�.G;vG;ݩG;~�G;�G;� H;@H;�[H;tH;u�H;��H;0�H;i�H;@�H;d�H;;�H;c�H;��H;��H;��H;k�H;y�H;0�H;p�H;0�H;x�H;k�H;��H;��H;��H;`�H;8�H;c�H;=�H;i�H;0�H;��H;s�H;tH;�[H;@H;� H;�G;}�G;ܩG;vG;�.G;C�F;�#F;BE;mD;�B;��@;��>;��<;�	;;�N9;m�7;�7;      .[@;�~@;P�@;
�A;QB;�1C;nD;��D;�E;�LF;��F;*$G;_fG;�G;O�G;��G;�	H;�)H;'FH;�_H;$vH;5�H;��H;��H;y�H;[�H;i�H;�H;��H;��H;L�H;�H;�H;��H;��H;9�H;��H;9�H;��H;��H;�H;�H;J�H;��H;��H;�H;i�H;[�H;y�H;��H;��H;5�H;!vH;�_H;'FH;�)H;�	H;��G;O�G;�G;_fG;+$G;��F;�LF;�E;��D;mD;�1C;QB;�A;N�@;�~@;      m�D;|�D;E;�NE;��E;�E;�[F;�F;�F;-;G;AmG;W�G;�G;��G;��G;�H;�5H;�NH;�eH;7zH;ȋH;�H;5�H;��H;�H;��H;j�H;��H;8�H;��H;��H;��H;��H;��H;��H;0�H;N�H;/�H;��H;��H;��H;��H;��H;��H;5�H;��H;g�H;��H;�H;�H;3�H;�H;ƋH;9zH;�eH;�NH;�5H;�H;��G;��G;�G;X�G;AmG;,;G;�F;�F;�[F;�E;��E;�NE;E;|�D;      �F;��F; �F;t�F;G;�#G;�FG;~hG;ƇG;٤G;��G;��G;k�G; H;:,H;�CH;�YH;nH;�H;��H;��H;ɩH;g�H;Z�H;��H;3�H;v�H;��H;T�H;^�H;��H;E�H;��H;��H;��H; �H;��H; �H;��H;��H;��H;G�H;��H;]�H;S�H;��H;v�H;3�H;��H;X�H;e�H;ǩH;��H;��H;�H;nH;�YH;�CH;;,H; H;l�G;��G;��G;ؤG;ȇG;}hG;�FG;�#G;G;t�F;�F;��F;      �lG;�nG;uG;�G;��G;w�G;��G;��G;��G;"�G;��G;�H;,+H;�?H;�SH;NfH;wH;�H;��H;_�H;z�H;�H;?�H;m�H;a�H;y�H;��H;�H;�H;j�H;]�H;��H;��H;��H;@�H;��H;��H;��H;>�H;��H;��H;��H;]�H;i�H;�H;�H;��H;w�H;d�H;l�H;?�H;�H;w�H;a�H;��H;�H;wH;NfH;�SH;�?H;,+H;�H;��G;"�G;��G;��G;��G;v�G;�G;�G;uG;�nG;      ��G;$�G;Y�G;�G;�G;@�G;;�G;�H;lH;�!H;�2H;gCH;TH;WdH;�sH;�H;�H;��H;�H;��H;|�H;�H;c�H;�H;��H;��H;�H;��H;N�H;�H;��H;��H;��H;y�H;��H;�H;X�H;�H;��H;{�H;��H;��H;��H;�H;N�H;��H;�H;��H;��H;�H;c�H;�H;z�H;��H;�H;��H;�H;�H;�sH;TdH;TH;gCH;�2H;�!H;mH;�H;;�G;@�G;�G;�G;W�G;/�G;      �H;dH;�H;�H;�H;M H;A*H;o5H;zAH;NH;#[H;"hH;uH;Q�H;��H;��H;�H;a�H;��H;r�H;��H;��H;8�H;��H;/�H;T�H; �H;N�H;�H;��H;��H;��H;t�H;��H;S�H;��H;��H;��H;T�H;��H;q�H;��H;��H;��H;�H;N�H;�H;T�H;1�H;��H;6�H;��H;��H;r�H;��H;c�H;�H;��H;��H;Q�H;uH; hH;"[H;NH;}AH;o5H;A*H;M H;�H;�H;�H;ZH;      �:H;�;H;>H;�AH;GGH;�MH;�UH;,^H;OgH;�pH;�zH;��H;]�H;��H;��H;1�H;�H;J�H;þH;��H;��H;R�H;_�H;��H;��H;Z�H;h�H;�H;��H;��H;��H;j�H; �H;s�H;��H;��H;��H;��H;��H;s�H;��H;j�H;��H;��H;��H;�H;f�H;Y�H;��H;��H;]�H;R�H;��H;��H;þH;L�H;�H;1�H;��H;��H;]�H;��H;�zH;�pH;RgH;/^H;�UH;�MH;BGH;�AH;	>H;�;H;      �bH;�cH;�eH;shH;�lH;pqH;7wH;�}H;��H;ˋH;�H;��H;��H;J�H;M�H;϶H;ԼH;M�H;L�H;��H;��H;|�H;��H;M�H;��H;��H;Z�H;��H;��H;��H;�H;��H;g�H;��H;�H;.�H;P�H;.�H;�H;��H;d�H;��H;}�H;��H;��H;��H;Z�H;��H;��H;M�H;��H;|�H;��H;��H;L�H;M�H;ӼH;ζH;M�H;I�H;��H;��H;�H;̋H;��H;�}H;7wH;qqH;�lH;uhH;�eH;�cH;      2�H;��H;�H;.�H;C�H;�H;;�H;.�H;u�H;�H;ХH;��H;^�H;ܶH;
�H;�H;��H;�H;�H;��H;��H;r�H;��H;�H;��H;D�H;��H;��H;��H;k�H;��H;}�H;��H;+�H;Q�H;~�H;m�H;}�H;Q�H;+�H;��H;}�H;��H;m�H;��H;��H;��H;B�H;��H;�H;��H;r�H;��H;��H;�H;�H;��H;�H;
�H;ܶH;^�H;��H;ХH;�H;w�H;-�H;;�H;�H;B�H;-�H;�H;��H;      e�H;��H;��H;z�H;؜H;��H;!�H;��H;�H;c�H;ϳH;)�H;��H;��H;��H;��H;��H;��H;��H;��H;P�H;��H;��H;�H;��H;��H;��H;��H;x�H;�H;h�H;��H;9�H;S�H;��H;��H;p�H;��H;��H;S�H;6�H;��H;h�H;�H;y�H;��H;��H;��H;��H;�H;��H;��H;O�H;��H;��H;��H;��H;��H;��H;��H;��H;'�H;ϳH;d�H;	�H;��H;!�H;��H;ќH;z�H;��H;��H;      u�H;��H;��H;�H;׫H;�H;°H;��H;ֶH;,�H;��H;1�H;��H;�H;v�H;��H;e�H;�H;��H;��H;��H;��H;j�H;��H;��H;��H;��H;x�H;��H;s�H;��H;+�H;L�H;��H;��H;��H;��H;��H;��H;��H;J�H;-�H;��H;u�H;��H;x�H;��H;��H;��H;��H;j�H;��H;��H;��H;��H;�H;c�H;��H;v�H;�H;��H;1�H;��H;,�H;ֶH;��H;°H;�H;ͫH;�H;��H;��H;      �H;[�H;�H;�H;��H;g�H;��H;�H;ľH;�H;p�H;e�H;'�H;�H;��H;=�H;��H;��H;-�H;�H;��H;,�H;v�H;��H;��H;��H;:�H;��H;S�H;��H;�H;T�H;��H;��H;��H;��H;��H;��H;��H;��H;��H;W�H;�H;��H;T�H;��H;9�H;��H;��H;��H;v�H;,�H;��H;�H;-�H;��H;��H;=�H;��H;�H;'�H;e�H;o�H;��H;ľH;�H;��H;k�H;��H;�H;��H;R�H;      &�H;g�H;��H;޹H;K�H;ѼH;þH;��H;=�H;��H;>�H;��H;<�H;��H;3�H;}�H;��H;��H;��H;B�H;��H;�H;0�H;=�H;(�H;��H;��H;�H;��H;��H;-�H;�H;��H;��H;��H;��H;��H;��H;��H;��H;��H;��H;-�H;��H;��H;�H;��H;��H;)�H;<�H;0�H;�H;��H;B�H;��H;��H;��H;}�H;2�H;��H;<�H;��H;>�H;��H;=�H;��H;þH;ּH;>�H;߹H;��H;^�H;      �H;_�H;��H;��H;�H;��H;i�H;w�H;��H;��H;T�H;��H;`�H;��H;�H;e�H;e�H;G�H;��H;��H;�H;U�H;n�H;��H;G�H;��H;��H;[�H;��H;��H;Q�H;s�H;o�H;��H;��H;��H;��H;��H;��H;��H;l�H;t�H;Q�H;��H;��H;[�H;��H;��H;G�H;��H;n�H;U�H;�H;��H;��H;I�H;d�H;e�H;�H;��H;`�H;��H;T�H;��H;��H;t�H;i�H;��H;�H;��H;��H;V�H;      &�H;h�H;��H;߹H;K�H;ѼH;þH;��H;=�H;��H;>�H;��H;<�H;��H;2�H;}�H;��H;��H;��H;B�H;��H;�H;0�H;=�H;)�H;��H;��H;�H;��H;��H;-�H;�H;��H;��H;��H;��H;��H;��H;��H;��H;��H;��H;-�H;��H;��H;�H;��H;��H;(�H;<�H;0�H;�H;��H;B�H;��H;��H;��H;}�H;2�H;��H;<�H;��H;?�H;��H;>�H;��H;þH;ּH;>�H;߹H;��H;]�H;      �H;[�H;�H;�H;��H;g�H;��H;�H;ľH;�H;n�H;e�H;'�H;�H;��H;=�H;��H;��H;-�H;�H;��H;,�H;v�H;��H;��H;��H;:�H;��H;S�H;��H;�H;T�H;��H;��H;��H;��H;��H;��H;��H;��H;��H;X�H;�H;��H;T�H;��H;9�H;��H;��H;��H;v�H;,�H;��H;�H;-�H;��H;��H;=�H;��H;�H;'�H;e�H;o�H;��H;ľH;�H;��H;j�H;��H;�H;�H;R�H;      v�H;��H;��H;�H;׫H;�H;°H;��H;ֶH;,�H;��H;1�H;��H;�H;v�H;��H;e�H;�H;��H;��H;��H;��H;j�H;��H;��H;��H;��H;x�H;��H;s�H;��H;*�H;L�H;��H;��H;��H;��H;��H;��H;��H;J�H;.�H;��H;u�H;��H;x�H;��H;��H;��H;��H;j�H;��H;��H;��H;��H;�H;c�H;��H;v�H;�H;��H;1�H;��H;,�H;ضH;��H;°H;�H;̫H;�H;��H;��H;      h�H;��H;��H;{�H;לH;��H;!�H;��H;	�H;c�H;ϳH;'�H;��H;��H;��H;��H;��H;��H;��H;��H;Q�H;��H;��H;�H;��H;��H;��H;��H;x�H;�H;h�H;��H;8�H;Q�H;��H;��H;p�H;��H;��H;Q�H;6�H;��H;h�H;�H;y�H;��H;��H;��H;��H;�H;��H;��H;O�H;��H;��H;��H;��H;��H;��H;��H;��H;)�H;ϳH;d�H;�H;��H;!�H;��H;ΜH;{�H;��H;��H;      2�H;��H;�H;+�H;C�H;�H;>�H;/�H;u�H;�H;ХH;��H;^�H;ܶH;
�H;�H;��H;�H;�H;��H;��H;r�H;��H;�H;��H;D�H;��H;��H;��H;k�H;��H;}�H;��H;+�H;Q�H;~�H;m�H;}�H;Q�H;+�H;��H;~�H;��H;m�H;��H;��H;��H;B�H;��H;�H;��H;r�H;��H;��H;�H;�H;��H;�H;
�H;ܶH;\�H;��H;ХH;�H;w�H;+�H;>�H;�H;A�H;+�H;�H;��H;      �bH;�cH;�eH;uhH;�lH;pqH;7wH;�}H;��H;ˋH;�H;��H;��H;J�H;M�H;϶H;ӼH;K�H;L�H;��H;��H;|�H;��H;N�H;��H;��H;Z�H;��H;��H;��H;}�H;��H;e�H;��H;�H;.�H;P�H;.�H;�H;��H;d�H;��H;�H;��H;��H;��H;Z�H;��H;��H;M�H;��H;|�H;��H;��H;L�H;M�H;ӼH;϶H;M�H;J�H;��H;��H;�H;̋H;��H;�}H;7wH;sqH;�lH;shH;�eH;�cH;      �:H;�;H;>H;�AH;AGH;�MH;�UH;/^H;PgH;�pH;�zH;��H;]�H;��H;��H;1�H;�H;J�H;þH;��H;��H;R�H;_�H;��H;��H;Z�H;h�H;�H;��H;��H;��H;h�H;��H;r�H;��H;��H;��H;��H;��H;s�H;��H;k�H;��H;��H;��H;�H;f�H;Y�H;��H;��H;]�H;R�H;��H;��H;þH;L�H;�H;2�H;��H;��H;]�H;��H;�zH;�pH;RgH;/^H;�UH;�MH;@GH;�AH;>H;�;H;      �H;aH;�H;�H;�H;H H;D*H;q5H;{AH;NH;#[H;"hH;uH;Q�H;H;��H;�H;a�H;��H;t�H;��H;��H;8�H;��H;1�H;V�H; �H;N�H;�H;��H;��H;��H;r�H;��H;S�H;��H;��H;��H;S�H;��H;r�H;��H;��H;��H;�H;N�H;�H;S�H;/�H;��H;6�H;��H;��H;r�H;��H;c�H;�H;��H;��H;Q�H;uH;"hH;#[H;NH;}AH;o5H;D*H;L H;�H;�H;�H;aH;      ��G;$�G;Y�G;�G;�G;@�G;;�G;�H;lH;�!H;�2H;gCH;TH;WdH;�sH;�H;�H;��H;�H;��H;��H;�H;d�H;�H;��H;��H;�H;��H;P�H;�H;��H;��H;��H;y�H;��H;�H;X�H;�H;��H;y�H;��H;��H;��H;�H;M�H;��H;�H;��H;��H;�H;b�H;�H;y�H;��H;�H;��H;�H;�H;�sH;TdH;TH;gCH;�2H;�!H;mH;�H;;�G;=�G;�G;�G;Y�G;1�G;      �lG;�nG;�uG;�G;��G;s�G;��G;��G;��G;$�G;��G;�H;,+H;�?H;�SH;OfH;�wH;�H;��H;b�H;}�H;�H;@�H;m�H;d�H;y�H;��H;�H;�H;j�H;]�H;��H;��H;��H;>�H;��H;��H;��H;@�H;��H;��H;��H;]�H;i�H; �H;�H;��H;y�H;a�H;l�H;=�H;�H;w�H;_�H;��H;�H;}wH;NfH;�SH;�?H;,+H;�H;��G;$�G;��G;��G;��G;q�G;��G;�G;uG;�nG;      �F;��F;*�F;u�F;G;�#G;�FG;hG;ŇG;٤G;��G;��G;l�G; H;;,H;�CH;�YH;nH;�H;��H;��H;ǩH;g�H;Z�H;��H;4�H;v�H;��H;T�H;^�H;��H;E�H;��H;��H;��H; �H;��H; �H;��H;��H;��H;G�H;��H;\�H;S�H;��H;u�H;3�H;��H;Z�H;g�H;ɩH;��H;��H;�H;nH;�YH;�CH;:,H; H;k�G;��G;��G;ؤG;ƇG;}hG;�FG;�#G;G;u�F;*�F;��F;      m�D;}�D;E;�NE;��E;�E;�[F;�F;�F;-;G;CmG;X�G;�G;��G;��G;�H;�5H;�NH;�eH;9zH;ˋH;�H;5�H;��H;�H;��H;h�H;��H;8�H;��H;��H;��H;��H;��H;��H;/�H;N�H;0�H;��H;��H;��H;��H;��H;��H;5�H;��H;g�H;��H;�H;��H;3�H;�H;ȋH;9zH;�eH;�NH;�5H;�H;��G;��G;�G;W�G;AmG;,;G;�F;�F;�[F;�E;��E;�NE;E;|�D;      6[@;�~@;R�@;�A;	QB;�1C;lD;��D;�E;�LF;��F;+$G;`fG;�G;O�G;��G;�	H;�)H;'FH;�_H;%vH;5�H;��H;��H;y�H;[�H;j�H;�H;��H;��H;J�H;�H;�H;��H;��H;9�H;��H;9�H;��H;��H;�H;�H;L�H;��H;��H;�H;i�H;[�H;y�H;��H;��H;5�H;!vH;�_H;'FH;�)H;�	H;��G;O�G;�G;_fG;*$G;��F;�LF;�E;��D;lD;�1C;QB;�A;Q�@;�~@;      V�6;�7;|�7;�N9;�	;;��<;��>;��@;�B;mD;BE;�#F;B�F;�.G;vG;ݩG;~�G;�G;� H;@H;�[H;tH;u�H;��H;0�H;h�H;@�H;c�H;9�H;c�H;��H;��H;��H;k�H;x�H;0�H;p�H;0�H;y�H;k�H;��H;��H;��H;`�H;8�H;d�H;?�H;i�H;0�H;��H;s�H;tH;�[H;@H;� H;�G;~�G;ݩG;vG;�.G;@�F;�#F;
BE;jD;�B;��@;��>;��<;�	;;�N9;q�7;�7;      ��#;�f$;n(&;i�(;i,;�_0;r4;6�8;�'<;�N?;��A;��C;OE;�LF;�F;UG;s�G;�G;�G;�H;�<H;�ZH;tH;8�H;��H;ʩH;�H;�H;��H;V�H;}�H;q�H;��H;��H;+�H;�H;S�H;�H;+�H;��H;��H;q�H;|�H;R�H;��H;�H;�H;˩H;ߚH;5�H;tH;�ZH;�<H;�H;�G;�G;s�G;UG; �F;�LF;OE;��C;��A;�N?;�'<;5�8;r4;�_0;i,;i�(;m(&;�f$;      :;�/;"x;��
;9;��;Ρ ; `(;�/;��5;8
;;�%?;�5B;�^D;B�E;q�F;W8G; �G;��G;U�G;	H;�<H;�[H;(vH;ŋH;��H;y�H;|�H;��H;��H;��H;��H;J�H;��H;��H;��H;�H;��H;��H;��H;J�H;��H;��H;��H;��H;}�H;w�H;��H;ŋH;%vH;�[H;�<H;H;V�G;��G;�G;U8G;q�F;B�E;�^D;�5B;�%?;7
;;��5;�/;`(;̡ ;�;9;��
; x;�/;      L��:��:?A�:S��:���:0��:'�:��;"�;�f$;i>.;$6;)(<;h@;�tC;�[E;�F;N$G;`�G;�G;U�G;�H;@H;�_H;0zH;��H;^�H;��H;r�H;��H;��H;��H;��H;��H;�H;;�H;��H;;�H;�H;��H;��H;��H;��H;��H;m�H;��H;\�H;��H;0zH;�_H;@H;�H;R�G;�G;`�G;P$G;�F;�[E;�tC;h@;'(<;$6;g>.;�f$;"�;��;'�:6��:���:S��:5A�:��:      �VṨxƹ 0p� 0�6pY�9u,:|��:bٶ:�L�:X�;,�;�(&;_.1;�N9;�>;��B;�E;�cF;G;d�G;��G;�G;� H;(FH;�eH;�H;��H;�H;��H;žH;K�H;�H;��H;��H;*�H;��H;��H;��H;*�H;��H;��H;�H;L�H;þH;�H;�H;��H; �H;�eH;%FH;� H;�G;�G;e�G;G;�cF;�E;��B;�>;�N9;_.1;�(&;,�;X�;�L�:^ٶ:|��:"u,:�Y�9 0�6 0p��xƹ      ��4��K/�PV�L,�y�˺ 퀺�uƹ�m92oQ:炬:���:��;��;X�,;E7;��=;EQB;��D;�cF;R$G; �G;�G;�G;�)H;�NH;nH;�H;�H;e�H;P�H;N�H;�H;��H;�H;�H;��H;Q�H;��H;�H;�H;��H;�H;N�H;O�H;c�H;�H;�H;nH;�NH;�)H;�G;�G;��G;T$G;�cF;��D;BQB;��=;C7;X�,;��;��;���:催:>oQ:�m9�uƹ퀺m�˺N,�RV��K/�      P�ͻ4Sɻʹ��`Ϩ��-���\c��$���˺pP(��O@9��k:���:�;L�;:�);��5;q�=;GQB;�E;"�F;X8G;t�G;��G;�	H;�5H;�YH;�wH;�H;�H;�H;μH;��H;��H;_�H;��H;��H;`�H;��H;��H;_�H;��H;��H;μH;�H;�H;�H;}wH;�YH;�5H;�	H;}�G;t�G;W8G;#�F;�E;HQB;n�=;��5;:�);L�;�;���:��k:pO@9hP(���˺�$��\c��-��`Ϩ�δ��9Sɻ      �J;���7��9.����&����f���M����4���º�tƹjQ:���:���::�;��(;��5;��=;��B;�[E;q�F;UG;ܩG;��G;�H;�CH;OfH;�H;��H;/�H;ʶH; �H;��H;��H;5�H;v�H;^�H;v�H;5�H;��H;��H;�H;ȶH;.�H;��H;�H;KfH;�CH;�H;��G;ܩG;UG;q�F;�[E;��B;��=;��5;��(;:�;���:���:jQ:�tƹ��º��4�M��f�����軬&����9.���7�      �䙼0`��l��ky��z;k��I�P�$��� �����z�|�@�X$T��[�9B�:���::�;9�);E7;�>;�tC;E�E;�F;vG;R�G;��G;>,H;�SH;�sH;ŌH;��H;L�H;�H;��H;t�H;��H;/�H;�H;/�H;��H;t�H;��H;�H;J�H;��H;��H;�sH;�SH;?,H;��G;N�G;vG;�F;E�E;�tC;�>;H7;7�);:�;���:B�:�[�9`$T�@�|�|������� �P�$��I�z;k�ky��l��1`��      ������߼Sμ("���
��ky��iT�I�!���軾ۙ�jK/������m9B�:���:N�;]�,;�N9;o@;�^D;�LF;�.G;�G;��G;H;�?H;VdH;T�H;��H;F�H;նH;��H;�H;�H;��H;��H;��H;�H;�H;��H;ֶH;D�H;��H;S�H;TdH;�?H;H;��G;�G;�.G;�LF;�^D;o@;�N9;^�,;L�;���:B�:�m9����jK/��ۙ����H�!�jT�ky���
��)"��Sμ�߼���      ��/�K-�j.%����������Ǽث��~�{��J;��C�;Ϩ�FO:������[�9���:�;��;_.1;-(<;�5B;OE;F�F;ffG;�G;n�G;/+H;TH;uH;Y�H;��H;Z�H;��H;��H;"�H;8�H;]�H;8�H;"�H;��H;��H;Z�H;��H;X�H;uH;TH;,+H;r�G;�G;_fG;@�F;OE;�5B;-(<;_.1;��;�;���:�[�9����FO:�<Ϩ��C��J;�~�{�ث���Ǽ��������j.%�K-�      d@{�^`w��l��yZ�V�C�ig*�������'"��\O���I�A|�;Ϩ�kK/�X$T�nQ:���:��;�(&;$6;�%?;��C;�#F;-$G;U�G;��G;�H;dCH;hH;��H;��H;��H;#�H;-�H;^�H;��H;��H;��H;]�H;-�H; �H;��H;��H;��H;hH;dCH;�H;��G;X�G;'$G;�#F;��C;�%?;$6;�(&;��;���:fQ:X$T�lK/�;Ϩ�A|��I�\O��'"����鼲��ig*�V�C��yZ��l�^`w�      �b��誫��ƣ��s���ɇ��l�HG���"�l� �3aļf���I��C��ۙ�?��tƹ��k:���:+�;k>.;8
;;��A;BE;��F;DmG;��G;��G;�2H;%[H;�zH;�H;ʥH;ͳH;��H;k�H;8�H;N�H;8�H;k�H;��H;̳H;˥H;�H;�zH;#[H;�2H;��G;��G;GmG;��F;
BE;��A;:
;;i>.;+�;���:��k:�tƹ@��ۙ��C��I�f��3aļl� ���"�HG��l��ɇ��s���ƣ�誫�      ������tݽ�2̽�ж����������yZ�K-�ٷ�4aļ\O���J;����|�|���º�O@9催:X�;�f$;��5;�N?;pD;�LF;0;G;ۤG;'�G;�!H;NH;�pH;ƋH;�H;d�H;)�H;~�H;��H;��H;��H;~�H;)�H;c�H;�H;ƋH;�pH;NH;�!H;%�G;ܤG;1;G;�LF;nD;�N?;��5;�f$;X�;炬:pO@9��º|�|�����J;�\O��4aļٷ�K-��yZ����������ж��2̽tݽ���      R,����Z�=��z�WvϽ�b��0I��k]a�K-�l� �&"��~�{�I�!�������4�hP(�6oQ:�L�:$�;�/;�'<;�B;!�E;�F;ɇG;��G;jH;{AH;GgH;��H;q�H;�H;ҶH;��H;3�H;��H;3�H;��H;ҶH;�H;q�H;��H;GgH;xAH;lH;��G;ɇG;�F;�E;�B;�'<;�/;"�;�L�:6oQ:pP(���4�����I�!��{�&"��l� �K-�k]a�0I���b��VvϽ�z�=��Z���      )G�s�C��$:��J+��� ��sݽ`���0I���yZ���"����׫��jT��� �M����˺m9dٶ:��;`(;.�8;��@;��D;�F;�hG;��G;�H;p5H;(^H;�}H;'�H;��H;��H;�H;��H;r�H;��H;�H;��H;�H;(�H;�}H;(^H;m5H;�H;��G;hG;�F;��D;��@;.�8;`(;��;dٶ:m9��˺M���� �jT�׫�������"��yZ�0I��a���sݽ �����J+��$:�s�C�      {x�9t���g���T��G=�}#�6�sݽ�b������GG�����Ǽly��O�$�h����$��uƹr��:'�:ġ ;h4;��>;lD;�[F;�FG;��G;9�G;@*H;�UH;3wH;;�H;"�H;��H;��H;��H;e�H;��H;��H;��H;�H;:�H;2wH;�UH;?*H;9�G;��G;�FG;�[F;fD;��>;h4;ȡ ;'�:r��:�uƹ�$�h���O�$�ly���Ǽ���GG������b��sݽ6�}#��G=���T���g�9t�      ����Na��#���B�c�s�C�}#� ��VvϽ�����l�ig*����
���I���軼\c�퀺�t,:4��:��;�_0;��<;�1C;�E;�#G;t�G;A�G;O H;�MH;qqH;�H;��H;�H;j�H;ּH;��H;ؼH;h�H;�H;��H;�H;qqH;�MH;J H;A�G;s�G;�#G;�E;�1C;��<;�_0; �;4��:u,:퀺�\c�����I��
�����ig*��l�����VvϽ ��}#�s�C�B�c�#���Na����      l*��j����Ƥ���/��B�c��G=����zｔж��ɇ�V�C���)"��y;k��&��-��o�˺�Y�9���:9;i,;�	;;QB;��E;G;��G;�G;�H;9GH;�lH;A�H;ќH;ͫH;w�H;;�H;�H;;�H;v�H;ϫH;МH;B�H;�lH;6GH;�H;�G;��G;G;��E;QB;�	;;i,;9;���:�Y�9n�˺�-���&�y;k�)"����V�C��ɇ��ж��z����G=�B�c��/����Ƥ�j���      ��ɾ~�ž+��sת��#�����T��J+�=��2̽�s���yZ����Tμky����^Ϩ�O,� .�6U��: �
;p�(;�N9;�A;�NE;u�F;�G;�G;�H;�AH;khH;+�H;w�H;�H;�H;ܹH;��H;ܹH;�H;�H;u�H;*�H;lhH;�AH;�H;�G;�G;u�F;�NE;�A;�N9;r�(;�
;U��: .�6O,�_Ϩ���ky��Sμ����yZ��s���2̽=��J+���T�#����sת�+��~�ž      X_ݾ�:پ�V;+���Ƥ�Na����g��$:��Z�tݽ�ƣ��l�j.%��߼l���9.�ʹ��SV��0p�1A�:x;^(&;h�7;I�@;-E;-�F;�uG;S�G;�H;>H;�eH;
�H;��H;��H;�H;�H;�H;�H;�H;��H;��H;	�H;�eH;>H;�H;S�G;�uG;-�F;-E;D�@;m�7;_(&;x;3A�:�0p�RV�δ���9.�l���߼j.%��l��ƣ�tݽ�Z��$:���g�Na���Ƥ�+���V;�:پ      
^�7���:پ~�žj�����9t�s�C������誫�]`w�L-����0`����7�9Sɻ�K/��xƹ���:�/;�f$;�7;�~@;y�D;��F;�nG;%�G;hH;�;H;�cH;��H;��H;��H;G�H;a�H;Y�H;a�H;H�H;��H;��H;��H;�cH;�;H;eH;%�G;�nG;��F;y�D;�~@;�7;�f$;�/;�:�xƹ�K/�:Sɻ��7�0`�����K-�]`w�誫������s�C�9t���j���~�ž�:پ7��      HF�Zh����XVھ:�������~���S��#��o��<S��r₽6�6�v���my��[FB��Eֻ�A?���	��Y�:���:z�";�46;j@;��D;کF;�nG;"�G;BH;>@H;!gH;��H;f�H;ƩH;�H;�H;��H;�H;�H;ƩH;d�H;��H;!gH;<@H;?H;"�G;�nG;۩F;��D;g@;�46;z�";���:�Y�:��	��A?��Eֻ[FB�my��v���6�6�r₽<S���o���#��S��~������:��XVھ��Zh��      Zh���b���쾪*־�v��+���*��*�O�X� �s��r���؀�K�3���Dݜ�@�>�R�ѻ�9�p���ho�:A% ;�M#;}�6;[A@;!�D;ԯF;,qG;~�G;VH;	AH;�gH;�H;ŚH;�H;Q�H;.�H;�H;.�H;S�H;�H;ĚH;��H;�gH;AH;TH;~�G;,qG;ԯF;!�D;VA@;��6;�M#;A% ;fo�:x���ޡ9�S�ѻ@�>�Dݜ���K�3��؀��r��s�X� �*�O�*��+����v���*־���b��      ���쾶�޾25ʾO;���:��,�v��E�b'����t����u���+��W��A����4���Ļ9)�j���W�:g�;%;!l7;5�@; �D;�F;xG;��G;zH;jCH;ciH;R�H;țH;ڪH;��H;˺H;��H;˺H;��H;ڪH;ƛH;R�H;ciH;gCH;wH;��G;xG;�F; �D;0�@;#l7;%;f�;�W�:j��9)���Ļ��4��A���W缇�+���u�t�����b'��E�,�v��:��O;��25ʾ��޾��      XVھ�*־25ʾu��������M���9b��5�����ս����Xc�	��Жռ�I��X�$�kT���Z��Z��V�:�;��';X�8;.RA;�9E;��F;݂G;"�G;�H;4GH;JlH;��H;p�H;�H;�H;˻H;��H;˻H;�H;�H;o�H;��H;LlH;2GH;�H;!�G;݂G;��F;�9E;(RA;[�8;��';�;R�: [���Z�lT��Y�$��I��Жռ	���Xc������ս���5��9b��M������u���25ʾ�*־      :���v��O;������UP��I�r�~�H�X� ���8@��ԓ����K�e� ־���s�u���񕻘ܺ�5u9Y&�:-�;H�+;��:;�"B;��E;�F;�G;�G;sH;dLH;3pH;|�H;��H;ܭH;u�H;�H;��H;�H;r�H;ۭH;��H;�H;3pH;aLH;qH;�G;��G;�F;��E;�"B;��:;H�+;.�;W&�:�5u9�ܺ��u����s� ־�e���K�ԓ��8@����X� �~�H�I�r�UP������O;���v��      ����+����:���M��I�r�*�O�#,�Z�
��gٽtĥ���u�|1�o���.Ϥ���P�[�.o�bp���:���:Q;Y�/;p�<;C;M�E;�!G;V�G;7�G;�%H;�RH;uH;7�H;|�H;�H;@�H;��H;>�H;��H;@�H;�H;|�H;9�H;uH;�RH;�%H;7�G;U�G;�!G;L�E;C;p�<;X�/;Q;���:�:^p���.o�[򻯎P�.Ϥ�o���|1���u�tĥ��gٽZ�
�#,�*�O�I�r��M���:��+���      �~��*��,�v��9b�~�H�#,�OZ����:S��z^����N������μ�I���%+����ҝ.�@���k~:���:@m;��3;R�>;X�C;uPF;�FG;v�G;#�G;�/H;/ZH;�zH;��H;��H;��H;]�H;b�H;�H;b�H;]�H;��H;��H;��H;�zH;.ZH;�/H;#�G;u�G;�FG;rPF;T�C;P�>;��3;Am;���:k~:(���ҝ.�����%+��I����μ�����N�z^��:S�����OZ�#,�~�H��9b�,�v�*��      �S�*�O��E��5�X� �Z�
���罨9��+l���Xc���(��������[�����ݎ�)ܺ <9P��:X�	;\d';� 8;s�@;��D;�F;YjG;��G;�H;�:H;nbH;�H;C�H;i�H;��H;��H;q�H;�H;q�H;��H;�H;h�H;F�H;�H;nbH;�:H;�H;��G;YjG;�F;��D;s�@;� 8;]d';W�	;P��:@<9)ܺ�ݎ������[��������(��Xc�+l���9�����Z�
�X� ��5��E�*�O�      �#�X� �b'������gٽ:S��+l��T�j�G�3��i��վ�}���(���Ļ]A?�\�B�B�@:�[�:4Q;!�.;�;;�tB;>�E;��F;g�G;)�G;H;�FH;VkH;��H;^�H;G�H;��H;H�H;��H;2�H;��H;I�H;��H;G�H;_�H;��H;SkH;�FH;H;&�G;g�G;��F;=�E;�tB;�;;"�.;4Q;�[�:J�@:X�B�]A?���Ļ
(�}����վ��i�G�3�S�j�+l��:S���gٽ����b'�X� �      �o��s��置�ս9@��tĥ�{^���Xc�G�3���	�Ό˼�]��VFB��Z򻭜��XӺ���8��:��;�M#;�=5;=?;��C;�@F;@:G;+�G;Q�G;k'H;�RH;�tH;�H;��H;b�H;�H;��H;
�H;}�H;
�H;��H;�H;a�H;��H;�H;�tH;�RH;m'H;O�G;,�G;=:G;�@F;��C;=?;�=5;�M#;��;��:���8XӺ�����Z�VFB��]��Ό˼��	�G�3��Xc�{^��tĥ�9@����ս���s�      <S���r��t�����ԓ����u���N���(��i�Ό˼�A����P�is��5|������\:Z�:��;�n-;	�:;�A;�,E;��F;foG;.�G;�H;8H;|_H;=~H;)�H;>�H;��H;L�H;��H;v�H;��H;v�H;��H;K�H;��H;A�H;)�H;=~H;y_H;8H;�H;0�G;doG;��F;�,E;�A;�:;�n-;��;`�:�\:����5|��hs���P��A��Ό˼�i���(���N���u�ԓ�����t���r��      r₽�؀���u��Xc���K�|1�������վ��]����P����AT����9���o�44�9�&�:t�	;}%;w�5;��>;һC;�F;�!G;ښG;�G;yH;�HH;
lH;هH;��H;ͭH;�H;��H;��H;��H;�H;��H;��H;��H;�H;ЭH;��H;هH;lH;�HH;yH;�G;ךG;�!G;�F;ԻC;��>;v�5;}%;x�	;�&�:<4�9��o���9�@T�������P��]���վ�����|1���K��Xc���u��؀�      6�6�J�3���+�	��e�o�����μ���}���VFB�hs�AT��$�D��{���;u9�q�:���:�Y;u0;�;;B;":E;�F;4hG;�G;D�G;�0H;�XH;hxH;[�H;��H;>�H;5�H;�H;O�H;g�H;t�H;g�H;O�H;�H;5�H;@�H;��H;[�H;gxH;�XH;�0H;G�G;�G;0hG;�F;$:E;B;�;;u0;�Y;���:�q�:�;u9�{��$�D�AT��hs�VFB�}��������μo���e�	����+�K�3�      u�����W�Жռ ־�.Ϥ��I����[�
(��Z����9��{���<9tX�:�X�:[Q;Z,;��8;�A@;6BD;�@F;�,G;��G;��G;�H;EH;[hH;o�H;��H;��H;��H;_�H;\�H;�H;��H;��H;��H;�H;Z�H;_�H;��H;��H;��H;n�H;ZhH;EH;�H;��G;��G;�,G;�@F;6BD;�A@;��8;],;[Q;�X�:xX�:�<9�{����9���Z�	(���[��I��.Ϥ� ־�Жռ�W���      my��Dݜ��A���I����s���P��%+������Ļ����6|���o��;u9tX�:,�:q;�);�6;��>;�PC;��E;)�F;�xG;e�G;�H;�1H;SXH;>wH;�H;S�H;@�H;��H;V�H;~�H;��H;%�H;��H;%�H;��H;��H;U�H;��H;@�H;P�H;�H;>wH;QXH;�1H;�H;b�G;�xG;)�F;��E;�PC;��>;�6;�);q;,�:tX�:�;u9��o�5|�������Ļ����%+���P���s��I���A��Eݜ�      ZFB�@�>���4�Y�$�u��[�����ݎ�]A?�XӺ����,4�9�q�:�X�:s;��';�=5;��=;.�B;QGE;{�F;�UG;[�G;�G;�H;�HH;OjH;5�H;��H;��H;p�H;��H;�H;}�H;K�H;[�H;�H;[�H;K�H;|�H;�H;��H;p�H;��H;��H;5�H;MjH;IH;�H;�G;W�G;�UG;x�F;NGE;.�B;��=;�=5;��';s;�X�:�q�:<4�9����ZӺ[A?��ݎ����[�v��X�$���4�B�>�      �EֻM�ѻ��ĻmT���񕻴.o�̝.�(ܺ\�B����8\:�&�:���:ZQ;);�=5;;=;J#B;��D;vF;!7G;��G;��G;�H;�:H;O^H;�zH;7�H;��H;�H;G�H;�H;��H;Y�H;��H;h�H;��H;h�H;��H;[�H;��H;	�H;G�H; �H;��H;7�H;�zH;Q^H;�:H;�H;��G;��G; 7G;vF;��D;M#B;;=;�=5;);ZQ;���:�&�:�\:���8T�B�)̝ܺ.��.o���mT����ĻR�ѻ      �A?��9�9)��Z��ܺzp��H��� <9B�@:��:\�:t�	;�Y;V,;�6;��=;I#B;�D;�XF;"G;��G;V�G;�H;0/H;�SH;�qH;�H;��H;��H;��H;��H;�H;��H;�H;��H;X�H;��H;W�H;��H;�H;��H;!�H;��H;��H;��H;��H;�H;�qH;�SH;-/H;�H;V�G;��G;"G;�XF;�D;H#B;��=;�6;Z,;�Y;t�	;^�:��:J�@:�;9@���rp���ܺ�Z�9)��9�      ��	������i���Z���5u9�:k~:J��:�[�:��;��;}%;u0;��8;��>;.�B;��D;�XF;hG;��G;��G;��G;/&H;DKH;�iH;"�H;ȗH;v�H;��H;F�H;��H;��H;��H;o�H;��H;�H;��H;�H;��H;o�H;��H;��H;��H;C�H;��H;v�H;ŗH;#�H;�iH;AKH;,&H;��G;��G;��G;hG;�XF;��D;.�B;��>;��8;u0;~%;��;��;�[�:J��:k~:�:06u9�Z���i��x���      �Y�:�o�:�W�:T�:U&�:���:���:T�	;/Q;�M#;�n-;s�5;�;;�A@;�PC;IGE;vF;"G;��G;
�G;P�G;� H;IEH;�cH;z}H;��H;��H;߱H;�H;��H;��H;i�H;��H;��H;��H;��H;+�H;��H;��H;��H;��H;j�H;��H;��H;��H;ޱH;�H;��H;z}H;�cH;GEH;� H;N�G;�G;��G;"G;vF;JGE;�PC;�A@;�;;s�5;�n-;�M#;1Q;U�	;���:���:k&�:V�:�W�:vo�:      ���:N% ;m�; �;)�;Q;Am;[d';�.;�=5;�:;��>;B;5BD;��E;x�F; 7G;��G;��G;Q�G;�H;%BH;H`H;�yH;��H;a�H;��H;!�H;��H;�H;��H;o�H;��H;|�H;/�H;�H;��H;�H;/�H;|�H;��H;p�H;��H;�H;��H; �H;��H;a�H;��H;�yH;E`H;'BH;�H;T�G;��G;��G;7G;x�F;��E;5BD;B;��>;�:;�=5;!�.;Yd';Cm;Q;+�;�;l�;>% ;      ��";�M#;-%;x�';H�+;`�/;��3;� 8;�;;>?; �A;һC;":E;�@F;)�F;�UG;��G;V�G;��G;� H;$BH;�^H;�wH;Z�H;ĝH;�H;ͷH;l�H;=�H;e�H;^�H;'�H;��H;�H;��H;��H;��H;��H;��H;�H;��H;'�H;^�H;a�H;9�H;l�H;˷H;�H;ƝH;V�H;�wH;�^H;$BH;� H;��G;Y�G;��G;�UG;*�F;�@F;":E;ԻC;�A;??;�;;� 8;��3;b�/;`�+;x�';*%;�M#;      �46;��6;"l7;N�8;��:;q�<;S�>;r�@;�tB;��C;�,E;�F;�F;�,G;�xG;W�G;��G;�H;.&H;LEH;F`H;�wH;n�H;s�H;��H;(�H;ٿH;��H;�H;;�H;j�H;~�H;��H;��H;��H;��H;��H;��H;��H;��H;��H;~�H;j�H;9�H;�H;��H;ֿH;)�H;��H;r�H;m�H;�wH;B`H;MEH;/&H;�H;��G;V�G;�xG;�,G;�F;�F;�,E;�C;�tB;s�@;S�>;s�<;��:;N�8;#l7;u�6;      |@;gA@;<�@;)RA;�"B;C;\�C;��D;=�E;�@F;��F;�!G;.hG;��G;a�G;�G;�H;0/H;AKH;�cH;�yH;X�H;r�H;�H;D�H;��H;��H;�H;O�H;��H;��H;��H;{�H;��H;�H;��H;��H;��H;	�H;��H;x�H;��H;��H;��H;M�H;�H;��H;��H;F�H;��H;p�H;W�H;�yH;�cH;AKH;2/H;�H;�G;a�G;��G;.hG;�!G;��F;�@F;>�E;��D;[�C;C;�"B;(RA;;�@;\A@;      ��D;#�D;�D;�9E;��E;P�E;qPF;�F;��F;<:G;aoG;ؚG;�G;��G;�H;�H;�:H;�SH;�iH;�}H;ÎH;ɝH;��H;M�H;x�H;!�H;k�H;��H;��H;m�H;"�H;G�H;��H;*�H;��H;_�H;��H;_�H;��H;'�H;��H;G�H;"�H;l�H;��H;��H;k�H;!�H;z�H;J�H;��H;ɝH;��H;�}H;�iH;�SH;�:H;�H;�H;��G;�G;ښG;aoG;::G;��F;�F;qPF;O�E;��E;�9E;�D;#�D;      �F;߯F;�F;��F;�F;�!G;�FG;UjG;b�G;(�G;*�G;�G;A�G;�H;�1H;�HH;N^H;�qH;�H;��H;^�H;�H;%�H;��H;�H;M�H;\�H;��H; �H;��H;��H;��H;/�H;�H;��H;�H;K�H;�H;��H;�H;-�H;��H;��H;��H;��H;��H;\�H;M�H;�H;��H;%�H;�H;Z�H;��H;�H;�qH;M^H;�HH;�1H;�H;A�G;�G;+�G;(�G;e�G;SjG;�FG;�!G;�F;��F;�F;ׯF;      �nG;.qG;xG;߂G;��G;Y�G;y�G;��G;%�G;L�G;�H;{H;�0H;	EH;QXH;OjH;�zH;�H;ȗH;��H;��H;ͷH;׿H;��H;g�H;_�H;~�H;��H;��H;��H;��H;�H;"�H;��H;t�H;��H;��H;��H;r�H;��H; �H;�H;��H;��H;��H;��H;}�H;^�H;h�H;��H;ֿH;ͷH;��H;��H;ȗH;�H;�zH;NjH;QXH;	EH;�0H;{H;�H;L�G;'�G;��G;y�G;V�G;��G;߂G;xG;,qG;      �G;~�G;��G;�G;�G;4�G;&�G;�H;H;k'H;8H;�HH;�XH;]hH;=wH;5�H;6�H;�H;s�H;�H; �H;l�H;��H;�H;��H;��H;��H;{�H;��H;��H;��H;�H;��H;��H;�H;B�H;V�H;B�H;�H;��H;��H;�H;��H;��H;��H;{�H;��H;��H;��H;�H;��H;j�H;�H;�H;s�H;�H;5�H;5�H;@wH;[hH;�XH;�HH;8H;k'H;H;�H;$�G;5�G;)�G;�G;��G;��G;      XH;TH;xH;�H;pH;�%H;�/H;�:H;�FH;�RH;y_H;lH;gxH;n�H;�H;��H;��H;��H;��H;�H;��H;<�H;�H;T�H;��H;�H;��H;��H;a�H;��H;�H;��H;��H; �H;��H;��H;��H;��H;��H; �H;��H;��H;�H;��H;a�H;��H;��H; �H;��H;T�H;�H;<�H;��H;�H;��H;��H;��H;��H;�H;o�H;hxH;
lH;y_H;�RH;�FH;�:H;�/H;�%H;wH;�H;wH;HH;      H@H;AH;nCH;6GH;pLH;�RH;2ZH;tbH;\kH;�tH;D~H;�H;_�H;��H;S�H;��H;�H;�H;B�H;��H;�H;a�H;6�H;��H;b�H;��H;��H;��H;��H;�H;��H;��H;7�H;��H;��H;�H;�H;�H;��H;��H;4�H;��H;��H;�H;��H;��H;��H;��H;e�H;��H;4�H;c�H;�H;��H;B�H;��H;�H;��H;S�H;��H;_�H;�H;F~H;�tH;^kH;ubH;2ZH;�RH;nLH;6GH;jCH;AH;      gH;�gH;miH;PlH;<pH;uH;�zH;��H;ŇH;�H;,�H;��H;��H;��H;A�H;v�H;K�H;��H;��H;��H;��H;]�H;j�H;��H;�H;��H;��H;��H;�H;��H;��H;C�H;��H;��H;�H;J�H;f�H;J�H;�H;��H;��H;E�H;��H;��H;�H;��H;��H;��H;�H;��H;e�H;[�H;��H;��H;��H;��H;J�H;u�H;A�H;��H;��H;��H;.�H;�H;ƇH;��H;�zH;uH;:pH;QlH;miH;�gH;      ��H;��H;\�H;��H;��H;7�H;��H;L�H;a�H;��H;B�H;խH;A�H;��H;��H;��H;�H;�H;��H;p�H;t�H;*�H;~�H;��H;A�H;��H;�H;�H;��H;��H;A�H;��H;��H;<�H;e�H;��H;��H;��H;e�H;<�H;��H;��H;B�H;��H;��H;�H;�H;��H;D�H;��H;|�H;*�H;s�H;p�H;��H;�H;�H;��H;��H;��H;A�H;ԭH;B�H;��H;b�H;I�H;��H;;�H;�H;��H;\�H;��H;      i�H;ΚH;ϛH;t�H;��H;{�H;��H;q�H;L�H;b�H;��H;�H;6�H;c�H;X�H;�H;��H;��H;��H;��H;��H;��H;��H;�H;��H;.�H;!�H;��H;��H;?�H;��H;��H;?�H;w�H;��H;��H;��H;��H;��H;w�H;<�H;��H;��H;?�H;��H;��H;�H;-�H;��H;�H;��H;��H;��H;��H;��H;��H;��H;�H;U�H;b�H;5�H;�H;��H;c�H;L�H;p�H;��H;�H;��H;t�H;ϛH;ǚH;      ҩH;"�H;ժH;"�H;�H;�H;��H;��H;��H;�H;P�H;��H; �H;_�H;��H;��H;_�H;	�H;q�H;��H;��H;�H;��H;��H; �H;�H;��H;��H;�H;��H;��H;;�H;p�H;��H;��H;��H;��H;��H;��H;��H;o�H;=�H;��H;��H; �H;��H;��H;�H;!�H;��H;��H;�H;��H;��H;q�H;�H;]�H;��H;��H;_�H; �H;��H;O�H;�H;��H;��H;��H;�H;ۭH;"�H;֪H;�H;      �H;d�H;��H;�H;��H;<�H;a�H;ǽH;O�H;��H;��H;��H;S�H; �H;��H;R�H;��H;��H;��H;��H;8�H;��H;��H;�H;��H;��H;n�H;�H;��H;��H;�H;h�H;��H;��H;��H;��H;��H;��H;��H;��H;��H;i�H;�H;��H;��H;�H;m�H;��H;��H;�H;��H;��H;5�H;��H;��H;��H;��H;R�H;��H; �H;S�H;��H;��H;��H;P�H;ĽH;c�H;@�H;��H;�H;��H;[�H;      ��H;3�H;ҺH;˻H;�H;��H;i�H;z�H;��H;�H;}�H;��H;j�H;��H;(�H;a�H;n�H;Q�H;�H;��H;'�H;��H;��H;��H;X�H;�H;��H;A�H;��H;�H;I�H;��H;��H;��H;��H;��H;��H;��H;��H;��H;��H;��H;I�H;�H;��H;A�H;��H;�H;Y�H;��H;��H;��H;%�H;��H;�H;S�H;m�H;a�H;(�H;��H;k�H;��H;{�H;�H;��H;x�H;i�H;��H;�H;˻H;պH;+�H;      ��H;�H;��H;��H;ʾH;<�H;�H;�H;9�H;}�H;��H;$�H;v�H;��H;��H;�H;��H;��H;��H;1�H;��H;��H;��H;��H;��H;D�H;��H;X�H;��H;�H;h�H;��H;��H;��H;��H;��H;��H;��H;��H;��H;��H;��H;h�H;�H;��H;X�H;��H;E�H;��H;��H;��H;��H;��H;1�H;��H;��H;��H;�H;��H;��H;v�H;$�H;��H;��H;:�H;�H;�H;A�H;��H;��H;��H;�H;      ��H;3�H;ҺH;˻H;�H;��H;i�H;z�H;��H;�H;}�H;��H;k�H;��H;(�H;a�H;n�H;Q�H;�H;��H;(�H;��H;��H;��H;Y�H;�H;��H;A�H;��H;�H;I�H;��H;��H;��H;��H;��H;��H;��H;��H;��H;��H;��H;I�H;�H;��H;A�H;��H;�H;X�H;��H;��H;��H;%�H;��H;�H;S�H;m�H;a�H;(�H;��H;j�H;��H;}�H;
�H;��H;w�H;i�H;��H;�H;˻H;ѺH;(�H;      �H;d�H;��H;�H;��H;<�H;c�H;ɽH;O�H;��H;��H;��H;S�H; �H;��H;R�H;��H;��H;��H;��H;9�H;��H;��H;�H;��H;��H;n�H;�H;��H;��H;�H;f�H;��H;��H;��H;��H;��H;��H;��H;��H;��H;l�H;�H;��H;��H;�H;m�H;��H;��H;	�H;��H;��H;5�H;��H;��H;��H;��H;R�H;��H; �H;S�H;��H;��H;��H;O�H;ĽH;c�H;@�H;��H;�H;��H;[�H;      ԩH;"�H;ժH;"�H;�H;�H;��H;��H;��H;�H;P�H;��H; �H;_�H;��H;��H;_�H;	�H;q�H;��H;��H;�H;��H;��H;!�H;�H;��H;��H;�H;��H;��H;;�H;p�H;��H;��H;��H;��H;��H;��H;��H;o�H;=�H;��H;��H; �H;��H;��H;�H; �H;��H;��H;�H;��H;��H;q�H;�H;]�H;��H;��H;_�H; �H;��H;P�H;�H;��H;��H;��H;�H;حH;"�H;֪H;�H;      k�H;ΚH;ЛH;v�H;��H;|�H;��H;p�H;L�H;b�H;��H;�H;5�H;c�H;V�H;�H;��H;��H;��H;��H;��H;��H;��H;�H;��H;.�H;!�H;��H;��H;>�H;��H;��H;=�H;v�H;��H;��H;��H;��H;��H;v�H;<�H;��H;��H;?�H;��H;��H; �H;-�H;��H;~�H;��H;��H;��H;��H;��H;��H;��H;�H;X�H;b�H;5�H;�H;��H;c�H;L�H;m�H;��H;�H;��H;v�H;͛H;˚H;      ��H;��H;\�H;��H;��H;9�H;��H;J�H;a�H;��H;B�H;խH;A�H;��H;��H;��H;�H;�H;��H;q�H;w�H;*�H;~�H;��H;D�H;��H;�H;�H;��H;��H;B�H;��H;��H;<�H;e�H;��H;��H;��H;e�H;<�H;��H;��H;A�H;��H;��H;�H;�H;��H;A�H;��H;|�H;*�H;s�H;p�H;��H;�H;�H;��H;��H;��H;@�H;ԭH;B�H;��H;b�H;H�H;��H;9�H;|�H;��H;]�H;��H;      gH;�gH;liH;QlH;<pH;uH;�zH;��H;ŇH;�H;.�H;��H;��H;��H;A�H;v�H;J�H;��H;��H;��H;��H;[�H;j�H;��H;�H;��H;��H;��H;�H;��H;��H;C�H;��H;��H;�H;J�H;f�H;J�H;�H;��H;��H;E�H;��H;��H;�H;��H;��H;��H;�H;��H;g�H;]�H;��H;��H;��H;��H;J�H;v�H;A�H;��H;��H;��H;+�H;�H;ŇH;��H;�zH;uH;:pH;PlH;miH;�gH;      B@H;AH;mCH;7GH;lLH;�RH;5ZH;ubH;]kH;�tH;D~H;�H;^�H;��H;S�H;��H;�H;��H;B�H;��H;�H;c�H;6�H;��H;e�H;��H;��H;��H;��H;�H;��H;��H;5�H;��H;��H;�H;�H;�H;��H;��H;5�H;��H;��H;�H;��H;��H;��H;��H;b�H;��H;4�H;a�H;�H;��H;A�H;��H;�H;��H;S�H;��H;_�H;�H;D~H;�tH;^kH;ubH;5ZH;�RH;kLH;6GH;mCH;AH;      PH;OH;~H;�H;vH;�%H;�/H;�:H;�FH;�RH;{_H;lH;gxH;o�H;�H;��H;��H;��H;��H;�H;��H;<�H;�H;T�H;��H;�H;��H;��H;a�H;��H;�H;��H;��H; �H;��H;��H;��H;��H;��H; �H;��H;��H;�H;��H;a�H;��H;��H; �H;��H;T�H;�H;<�H;��H;�H;��H;��H;��H;��H;�H;n�H;gxH;lH;{_H;�RH;�FH;�:H;�/H;�%H;qH;�H;{H;NH;      �G;�G;��G;�G;�G;5�G;$�G;�H;H;k'H;
8H;�HH;�XH;]hH;@wH;5�H;6�H;�H;s�H;�H;"�H;j�H;��H;�H;��H;��H;��H;{�H;��H;��H;��H;�H;��H;��H;�H;B�H;V�H;B�H;�H;��H;��H;�H;��H;��H;��H;{�H;��H;��H;��H;�H;��H;l�H;�H;�H;s�H;�H;5�H;6�H;>wH;ZhH;�XH;�HH;8H;k'H;H;�H;&�G;1�G;(�G;�G;��G;��G;      �nG;.qG;xG;قG;�G;U�G;x�G;��G;%�G;M�G;�H;{H;�0H;	EH;QXH;OjH;�zH;�H;ȗH;��H;��H;ͷH;׿H;��H;h�H;_�H;~�H;��H;��H;��H;��H;�H;!�H;��H;r�H;��H;��H;��H;t�H;��H;!�H;�H;��H;��H;��H;��H;}�H;_�H;g�H;��H;ֿH;ͷH;��H;��H;ȗH;�H;�zH;NjH;QXH;	EH;�0H;{H;�H;L�G;%�G;��G;x�G;U�G;��G;قG;xG;"qG;      �F;دF;�F;��F;�F;�!G;�FG;UjG;c�G;)�G;+�G;	�G;A�G;�H;�1H;�HH;N^H;�qH;�H;��H;`�H;�H;%�H;��H;�H;M�H;\�H;��H; �H;��H;��H;��H;.�H;�H;��H;�H;K�H;�H;��H;�H;-�H;��H;��H;��H;��H;��H;\�H;M�H;�H;��H;%�H;�H;Z�H;��H;�H;�qH;M^H;�HH;�1H;�H;A�G;�G;+�G;(�G;b�G;SjG;�FG;�!G;�F;��F;�F;ѯF;      ��D;#�D;�D;�9E;��E;P�E;qPF;�F;��F;<:G;coG;ښG;�G;��G;�H;�H;�:H;�SH;�iH;�}H;ĎH;ɝH;��H;M�H;z�H;!�H;l�H;��H;��H;m�H;"�H;F�H;��H;'�H;��H;_�H;��H;_�H;��H;(�H;��H;J�H;"�H;l�H;��H;��H;k�H;!�H;x�H;L�H;��H;ɝH;��H;�}H;�iH;�SH;�:H;�H;�H;��G;�G;ؚG;aoG;::G;��F;�F;qPF;P�E;��E;�9E;�D;%�D;      �@;cA@;?�@;%RA;�"B;C;Y�C;��D;>�E;�@F;��F;�!G;0hG;��G;a�G;�G;�H;//H;AKH;�cH;�yH;W�H;r�H;�H;F�H;��H;��H;�H;O�H;��H;��H;��H;z�H;��H;�H;��H;��H;��H;	�H;��H;z�H;��H;��H;��H;M�H;�H;��H;��H;D�H;�H;p�H;X�H;�yH;�cH;AKH;2/H;�H;�G;a�G;��G;-hG;�!G;��F;�@F;>�E;��D;Y�C;C;�"B;'RA;>�@;YA@;      �46;��6;1l7;N�8;��:;t�<;W�>;s�@;�tB;��C;�,E;�F;�F;�,G;�xG;W�G;��G;�H;/&H;LEH;H`H;�wH;n�H;s�H;��H;(�H;ٿH;��H;�H;;�H;j�H;~�H;��H;��H;��H;��H;��H;��H;��H;��H;��H;~�H;j�H;9�H;�H;��H;ֿH;)�H;��H;r�H;m�H;�wH;C`H;MEH;.&H;�H;��G;W�G;�xG;�,G;�F;�F;�,E;~�C;�tB;r�@;W�>;v�<;��:;N�8;&l7;|�6;      ��";�M#;.%;x�';H�+;`�/;��3;� 8;�;;??; �A;ԻC;":E;�@F;)�F;�UG;��G;V�G;��G;� H;'BH;�^H;�wH;Z�H;ƝH;�H;ͷH;l�H;=�H;e�H;^�H;'�H;��H;�H;��H;��H;��H;��H;��H;�H;��H;'�H;^�H;a�H;9�H;l�H;˷H;�H;ĝH;X�H;�wH;�^H;$BH;� H;��G;X�G;��G;�UG;*�F;�@F;":E;ԻC;�A;>?;�;;� 8;��3;`�/;\�+;x�';+%;�M#;      ���:H% ;r�;�;)�;Q;Gm;]d';�.;�=5;�:;��>;B;5BD;��E;x�F; 7G;��G;��G;S�G;�H;'BH;F`H;�yH;��H;a�H;��H; �H;��H;�H;��H;o�H;��H;{�H;/�H;�H;��H;�H;/�H;|�H;��H;p�H;��H;�H;��H;!�H;��H;a�H;��H;�yH;F`H;%BH;�H;S�G;��G;��G;7G;x�F;��E;5BD;B;��>;�:;�=5;�.;\d';Fm;Q;.�;�;o�;?% ;      �Y�:�o�:�W�:R�:[&�:���:���:U�	;1Q;�M#;�n-;s�5;�;;�A@;�PC;JGE;vF;"G;��G;
�G;S�G;� H;JEH;�cH;z}H;��H;��H;ޱH;�H;��H;��H;i�H;��H;��H;��H;��H;+�H;��H;��H;��H;��H;j�H;��H;��H;��H;߱H;�H;��H;z}H;�cH;FEH;� H;M�G;�G;��G;"G;vF;IGE;�PC;�A@;�;;r�5;�n-;�M#;1Q;U�	;���:���:g&�:P�:�W�:vo�:      ��	������i���Z���5u9�:k~:L��:�[�:��;��;~%;u0;��8;��>;.�B;��D;�XF;hG;��G;��G;��G;0&H;EKH;�iH;"�H;ȗH;v�H;��H;F�H;��H;��H;��H;o�H;��H;�H;��H;�H;��H;o�H;��H;��H;��H;C�H;��H;v�H;ŗH;#�H;�iH;@KH;+&H;��G;��G;��G;hG;�XF;��D;.�B;��>;��8;u0;}%;��;��;�[�:J��:k~:�:6u9�Z���i������      �A?��9�9)��Z��ܺ~p��H����;9B�@:��:^�:t�	;�Y;Y,;�6;��=;I#B;��D;�XF;"G;��G;V�G;�H;2/H;�SH;�qH;�H;��H;��H;��H;��H;�H;��H;�H;��H;W�H;��H;X�H;��H;�H;��H;!�H;��H;��H;��H;��H;�H;�qH;�SH;,/H;�H;V�G;��G;"G;�XF;�D;H#B;��=;�6;V,;�Y;t�	;\�:��:J�@:�;9H���rp���ܺ�Z�9)��9�      �EֻM�ѻ��ĻmT���񕻶.o�̝.�(ܺ\�B����8\:�&�:���:[Q;);�=5;;=;J#B;��D;vF;!7G;��G;��G;�H;�:H;O^H;�zH;7�H;��H;�H;G�H;	�H;��H;[�H;��H;h�H;��H;h�H;��H;[�H;��H;	�H;G�H;�H;��H;7�H;�zH;Q^H;�:H;�H;��G;��G; 7G;vF;��D;M#B;;=;�=5;);ZQ;���:�&�:\:���8T�B�+̝ܺ.��.o���nT����ĻR�ѻ      ZFB�@�>���4�X�$�v��[�����ݎ�]A?�XӺ����<4�9�q�:�X�:s;��';�=5;��=;.�B;NGE;z�F;�UG;Z�G;�G;�H; IH;OjH;5�H;��H;��H;p�H;��H;�H;|�H;K�H;[�H;�H;[�H;K�H;}�H;�H;��H;p�H;��H;��H;5�H;MjH; IH;�H;�G;W�G;�UG;z�F;NGE;.�B;��=;�=5;��';s;�X�:�q�:,4�9����ZӺ\A?��ݎ����[�v��Y�$���4�B�>�      my��Dݜ��A���I����s���P��%+������Ļ����6|���o��;u9tX�:,�:q;�);��6;��>;�PC;��E;)�F;�xG;e�G;�H;�1H;SXH;>wH;�H;S�H;@�H;��H;X�H;��H;��H;%�H;��H;%�H;��H;��H;V�H;��H;@�H;P�H;�H;>wH;QXH;�1H;�H;b�G;�xG;)�F;��E;�PC;��>;�6;�);q;,�:tX�:�;u9��o�6|�������Ļ����%+���P���s��I���A��Eݜ�      u�����W�Жռ ־�.Ϥ��I����[�
(��Z����9��{���<9xX�:�X�:\Q;\,;��8;�A@;5BD;�@F;�,G;��G;��G;�H;EH;ZhH;o�H;��H;��H;��H;`�H;[�H;�H;��H;��H;��H;�H;[�H;]�H;��H;��H;��H;o�H;[hH;	EH;�H;��G;��G;�,G;�@F;6BD;�A@;��8;],;ZQ;�X�:vX�:�<9�{����9���Z�	(���[��I��.Ϥ� ־�Жռ�W���      6�6�J�3���+�	��e�o�����μ���}���VFB�hs�AT��$�D��{���;u9�q�:���:�Y;u0;�;;B;$:E;�F;4hG;�G;D�G;�0H;�XH;hxH;[�H;��H;>�H;5�H;�H;O�H;g�H;t�H;i�H;O�H;�H;3�H;>�H;��H;[�H;gxH;�XH;�0H;H�G;�G;.hG;�F;":E;B;�;;u0;�Y;���:�q�:�;u9�{��$�D�AT��hs�VFB�}��������μo���e�	����+�K�3�      r₽�؀���u��Xc���K�|1�������վ��]����P����@T����9���o�<4�9�&�:w�	;}%;v�5;��>;ԻC;�F;�!G;ךG;�G;{H;�HH;lH;هH;��H;ͭH;�H;��H;��H;��H;�H;��H;��H;��H;�H;ЭH;��H;هH;lH;�HH;xH;�G;ښG;�!G;�F;һC;��>;v�5;}%;w�	;�&�:,4�9��o���9�AT�������P��]���վ�����|1���K��Xc���u��؀�      <S���r��t�����ԓ����u���N���(��i�Ό˼�A����P�hs��4|�����\:^�:��;�n-;�:;�A;�,E;��F;doG;.�G;�H;8H;|_H;=~H;)�H;>�H;��H;K�H;��H;v�H;��H;v�H;��H;L�H;��H;?�H;)�H;=~H;y_H;8H;�H;0�G;foG;��F;�,E;�A;�:;�n-;��;`�:�\:����6|��is���P��A��Ό˼�i���(���N���u�ԓ�����t���r��      �o��s��置�ս9@��tĥ�{^���Xc�G�3���	�Ό˼�]��VFB��Z򻭜��XӺ���8��:��;�M#;�=5;=?;��C;�@F;=:G;+�G;P�G;m'H;�RH;�tH;�H;��H;c�H;�H;��H;	�H;}�H;
�H;��H;�H;b�H;��H;�H;�tH;�RH;k'H;O�G;,�G;@:G;�@F;��C;=?;�=5;�M#;��;��:`��8ZӺ�����Z�VFB��]��Ό˼��	�G�3��Xc�{^��tĥ�9@����ս���s�      �#�X� �b'������gٽ:S��+l��S�j�G�3��i��վ�}���
(���Ļ^A?�T�B�B�@:�[�:5Q;�.;�;;�tB;?�E;��F;g�G;)�G;H;�FH;UkH;��H;^�H;I�H;��H;I�H;��H;2�H;��H;H�H;��H;F�H;^�H;��H;UkH;�FH;H;&�G;g�G;��F;;�E;�tB;�;;"�.;2Q;�[�:J�@:d�B�]A?���Ļ
(�}����վ��i�G�3�S�j�+l��:S���gٽ����b'�X� �      �S�*�O��E��5�X� �Z�
���罨9��*l���Xc���(��������[�����ݎ�&ܺ <9P��:X�	;[d';� 8;s�@;��D;�F;YjG;��G;�H;�:H;nbH;�H;E�H;j�H;��H;��H;q�H;�H;r�H;��H;��H;h�H;E�H;�H;nbH;�:H;�H;��G;XjG;�F;��D;s�@;� 8;]d';W�	;P��:0<9-ܺ�ݎ������[��������(��Xc�*l���9�����Z�
�X� ��5��E�*�O�      �~��*��,�v��9b�~�H�#,�OZ����:S��z^����N������μ�I���%+����Н.�0���k~:���:?m;��3;P�>;Y�C;rPF;�FG;v�G;#�G;�/H;/ZH;�zH;��H;��H;��H;]�H;b�H;�H;b�H;]�H;��H;��H;��H;�zH;.ZH;�/H;#�G;u�G;�FG;uPF;T�C;P�>;��3;Am;���:k~:0���ӝ.�����%+��I����μ�����N�z^��:S�����OZ�#,�~�H��9b�,�v�*��      ����+����:���M��H�r�*�O�#,�Z�
��gٽtĥ���u�|1�o���.Ϥ���P�[�.o�bp���:���:Q;X�/;o�<;C;L�E;�!G;V�G;7�G;�%H;�RH;uH;7�H;~�H;�H;@�H;��H;>�H;��H;@�H;�H;{�H;9�H;uH;�RH;�%H;7�G;U�G;�!G;M�E;C;p�<;Y�/;Q;���:�:^p���.o�[򻯎P�.Ϥ�o���|1���u�tĥ��gٽZ�
�#,�*�O�I�r��M���:��+���      :���v��O;������UP��I�r�~�H�X� ���8@��ԓ����K�e� ־���s�u���񕻘ܺ�5u9W&�:+�;H�+;��:;�"B;��E;�F;�G;�G;tH;dLH;3pH;|�H;��H;ۭH;t�H;�H;��H;�H;r�H;ܭH;��H;�H;3pH;aLH;qH;�G;��G;�F;��E;�"B;��:;H�+;.�;W&�:�5u9�ܺ��u����s� ־�e���K�ԓ��8@����X� �~�H�I�r�UP������O;���v��      XVھ�*־25ʾu��������M���9b��5�����ս����Xc�	��Жռ�I��Y�$�kT���Z� [��T�:�;��';X�8;.RA;�9E;��F;݂G;!�G;�H;6GH;LlH;��H;p�H;�H;�H;˻H;��H;˻H;�H;�H;o�H;��H;JlH;3GH;�H;"�G;݂G;��F;�9E;)RA;[�8;��';�;R�:�Z���Z�lT��X�$��I��Жռ	���Xc������ս���5��9b��M������u���25ʾ�*־      ���쾶�޾25ʾO;���:��,�v��E�b'����t����u���+��W��A����4���Ļ9)�j���W�:f�;%;!l7;5�@; �D;�F;xG;��G;zH;jCH;ciH;R�H;ɛH;ڪH;��H;˺H;��H;˺H;��H;ڪH;ƛH;R�H;ciH;gCH;wH;��G;xG;�F; �D;0�@;#l7;%;g�;�W�:j��9)���Ļ��4��A���W缇�+���u�t�����b'��E�,�v��:��O;��25ʾ��޾��      Yh���b���쾪*־�v��+���*��*�O�X� �s��r���؀�K�3���Dݜ�@�>�R�ѻ�9�x���ho�:A% ;�M#;}�6;[A@;!�D;ԯF;,qG;~�G;VH;	AH;�gH;�H;ŚH;�H;Q�H;.�H;�H;.�H;S�H;�H;ĚH;��H;�gH;AH;TH;~�G;+qG;ԯF;!�D;XA@;��6;�M#;A% ;fo�:x���ޡ9�S�ѻ@�>�Dݜ���K�3��؀��r��s�X� �*�O�*��+����v���*־���b��      3�$��� ����%��C��*�þ�*��6Dx���=�����Pν	���''K��c�"��r�V����
E^�T�S�,x[:���:'e;j�4;U`?;�mD;��F;dvG;M�G;�H;�OH;�sH;��H;��H;��H;/�H;��H;^�H;��H;.�H;��H;��H;��H;�sH;�OH;�H;M�G;bvG;��F;�mD;R`?;m�4;'e;���:(x[:T�S�	E^����r�V�"���c�''K�	����Pν�����=�6Dx��*��*�þC��%������� �      �� ����T��P��2��
����0��8�s�ڀ:�i9� �ʽ4Z���G��8�.���5S�����/X�4�D�Cd:�B�: ;1�4;؈?;D;]�F;'yG;��G;� H;VPH;QtH;K�H;�H;�H;k�H;��H;o�H;��H;m�H;�H;�H;L�H;QtH;SPH;� H;��G;'yG;_�F;D;Ԉ?;7�4; ;�B�:Cd:4�D��/X���껰5S�.���8��G�4Z�� �ʽi9�ڀ:�8�s��0��
���2��P��T�����      ���T��:�
������Yؾ"���॒���f���0�\[�R8��Ґ����>�����MȤ��6H�^�ܻ rF������}:��:{";l�5;�?;��D;�F;#�G;��G;{#H;�RH;�uH;��H;��H;��H;�H;)�H;��H;)�H;�H;��H;��H;��H;�uH;�RH;x#H;��G;#�G;�F;��D;�?;o�5;{";��:��}:����qF�_�ܻ�6H�MȤ�������>�Ґ��R8��\[���0���f�॒�"����Yؾ����:�
�T��      %��P������AI�*�þ�R��=���xS��Q"��s������}��0��켋�����6�C�ƻ0}*�����-�:�x;r%;m7;�@;�D;�F;��G;��G;;(H;VH;�xH;��H;~�H;ܲH;�H;��H;��H;��H;�H;ܲH;}�H;��H;�xH;VH;:(H;��G;��G;�F;�D;�@;m7;r%;�x;+�:����.}*�D�ƻ��6��������0���}�����s��Q"�xS�=����R��*�þAIᾦ���P��      C��2�很Yؾ*�þĪ�~쏾�k�ڀ:���~�ؽ�����c�`y���Ҽ����D� �d�"�� 5(7��:��
;�(;�_9;˘A;�\E;��F;ݝG;��G;�.H;�ZH;&|H;-�H;��H;��H;L�H;�H;��H;�H;J�H;��H;�H;/�H;&|H;�ZH;�.H;��G;ޝG;��F;�\E;ǘA;�_9;
�(;��
;��: 5(7 ��e�D� �������Ҽ`y��c�����~�ؽ��ڀ:��k�~쏾Ī�*�þ�Yؾ2��      *�þ
���"����R��~쏾8�s��H�����������ѐ����D��c�����@�f�S,�����P����9$��:�;Aj-;��;;��B;�E;�G;��G;��G;�6H;�`H;��H;��H;�H;��H;߾H;��H;�H;��H;߾H;��H;�H;��H;��H;�`H;�6H;��G;��G;�G;�E;��B;��;;Aj-;�; ��:��9�P�����T,�@�f������c���D�ѐ�������������H�8�s�~쏾�R��"���
���      �*���0��॒�=����k��H��#%�\[��Pν
t��d�f�6/%���伈���w�=��?ػ|FL�t�D�R:N�:I�;V2;��=;ښC;�0F;�GG;��G;ZH; @H;�gH;��H;l�H;�H;иH;��H;*�H;��H;*�H;��H;иH;�H;n�H;��H;�gH;@H;ZH;��G;�GG;�0F;ךC;��=;U2;J�;F�:R:h�D�|FL��?ػw�=��������6/%�d�f�
t���Pν\[��#%��H��k�=���॒��0��      6Dx�8�s���f�xS�ڀ:����\[��7ս�榽��}���;��8�W�����r����7G����� ˬ�X��:8�;�}$;�6;8�?;�D;�F;�pG;��G; H;cJH;ooH;y�H;��H;5�H;t�H;��H;��H;b�H;��H;��H;t�H;5�H;��H;y�H;ooH;bJH;H;��G;�pG;��F;�D;8�?;�6;�}$;7�;Z��:�ʬ����7G�������r�W����8���;���}��榽�7ս\[����ڀ:�xS���f�8�s�      ��=�ڀ:���0��Q"��������Pν�榽B����G�4����Ҽ ��JE:�;�ܻ�D^������i:z��:�;T|,;֡:;��A;giE;��F;[�G;��G;�(H;tUH;�wH;��H;b�H;˳H;/�H;�H;��H;N�H;��H;�H;/�H;̳H;e�H;��H;�wH;qUH;�(H;��G;]�G;��F;diE;��A;֡:;U|,;�;~��:�i:�����D^�;�ܻJE:� ����Ҽ4����G�B���榽�Pν�������Q"���0�ڀ:�      ���j9�\[��s�~�ؽ���
t����}� �G������2c��Y�V�F,��*�����`����:R��: ;��3;�0>;��C;F;9G;n�G;�H;)8H;�`H;:�H;*�H;6�H;��H;&�H;��H;�H;O�H;�H;��H;&�H;�H;9�H;*�H;:�H;�`H;'8H;�H;p�G;9G;F;��C;�0>;��3; ;R��:��:�������*��F,�Y�V�2c���������G���}�
t�����~�ؽ�s�\[�j9�      �Pν �ʽR8���������ѐ��d�f���;�4�����EȤ�6�f�)��Kߵ�Ko5���D���-:u��:�>;�+;�_9;�A;��D;N�F;�vG;�G;QH;�GH;�lH;��H;ϞH;2�H;d�H;1�H;��H;?�H;c�H;?�H;��H;1�H;c�H;6�H;ўH;��H;�lH;�GH;PH;�G;�vG;I�F;��D;�A;�_9;�+;�>;}��:��-:��D�Ko5�Jߵ�)��6�f�EȤ����4����;�d�f�ѐ���������R8�� �ʽ      	���4Z��Ґ����}��c���D�6/%��8���Ҽ2c��6�f�����ƻu/X�:���@��9@�:U�;�";��3;c>;oYC;��E;G;&�G;��G;�,H;>WH;OxH;��H;m�H;%�H;K�H;)�H;o�H;}�H;n�H;}�H;p�H;)�H;K�H;'�H;o�H;đH;MxH;>WH;�,H;��G;$�G;G;��E;oYC;c>;��3;�";Z�;>�:@��9:���t/X��ƻ���6�f�2c����Ҽ�8�6/%���D��c���}�Ґ��4Z��      ''K��G���>��0�`y��c����X��� ��Y�V�)���ƻ�od�f�º �(7�4�:���:¡;Q.;�:;:zA;\�D; �F;�nG;w�G;,H;�@H;_fH;��H;f�H;�H;�H;%�H;)�H;��H;��H;w�H;��H;��H;)�H;#�H;�H;�H;g�H;��H;_fH;�@H;.H;t�G;}nG;��F;\�D;<zA;�:;Q.;ġ;���:�4�: �(7f�º�od��ƻ)��Y�V� ��X�����众c�`y��0���>��G�      �c��8���������Ҽ����������r�IE:�E,�Jߵ�s/X�f�º�Ĭ���}:;�:;f�);Lm7;B�?;��C;8F;�)G;E�G;��G;@*H;�SH;�tH;��H;��H;.�H;�H;��H;�H;M�H;��H;��H;��H;M�H;�H;��H;�H;.�H;��H;��H;�tH;�SH;C*H;��G;E�G;�)G;8F;��C;B�?;Mm7;i�);;;�:��}:�Ĭ�d�ºr/X�Jߵ�E,�IE:���r�����������Ҽ�켺����8�      "��.��MȤ����� ���A�f�w�=����=�ܻ�*��Ko5�<��� �(7��}:�n�:H�;�>&;��4;�=;��B;�E;F�F;ʁG;)�G;kH;�AH;�eH;x�H;�H;��H;�H;��H;\�H;��H;��H;��H;��H;��H;��H;��H;\�H;��H;�H;��H;�H;z�H;�eH;�AH;jH;&�G;ƁG;F�F;�E;��B;�=;��4;�>&;H�;�n�:��}: �(7<���Ko5��*��<�ܻ���w�=�@�f� �������MȤ�.��      q�V��5S��6H���6�E� �U,��?ػ9G���D^������D�8��9�4�:3�:I�;%;��3;>�<;�B;�E;2�F;�XG;;�G;� H;�0H;�WH;�vH;,�H;��H;��H;νH;�H;��H;��H;��H;��H;w�H;��H;��H;��H;��H;�H;νH;��H;��H;-�H;�vH;�WH;�0H;| H;8�G;�XG;/�F;�E;�B;?�<;��3;%;I�;9�:�4�:@��9��D�����D^�9G���?ػT,�E� ���6��6H��5S�      ��ﻪ��`�ܻE�ƻe󩻴��wFL��������`����-:>�:���:;�>&;��3;z9<;9�A;�D;{ZF;S5G;2�G;�G;�!H;nJH;nkH;߅H;��H;��H;ظH;&�H;��H;��H;�H;��H;��H;0�H;��H;��H;�H;��H;��H;&�H;׸H;��H;��H;܅H;okH;nJH;�!H;�G;2�G;S5G;{ZF;�D;<�A;|9<;��3;�>&;;���:>�:��-:`���������wFL����d�E�ƻ`�ܻ���      E^��/X��qF�.}*�&���P��x�D�@ˬ��i:��:w��:T�;¡;b�);��4;;�<;7�A;L�D;�9F;G;��G;|�G;wH;V?H;�aH;P}H;��H;��H;ֳH;�H;��H;��H;��H;Y�H;��H;`�H;��H;`�H;��H;Y�H;��H;��H;��H;�H;ӳH;��H;��H;S}H;�aH;R?H;uH;|�G;��G;G;�9F;N�D;6�A;;�<;��4;f�);¡;U�;w��:��:�i:�ˬ�x�D��P����.}*��qF�0X�      D�S�@�D�T������ 2(7�9ҍR:T��:x��:P��:�>;�";Q.;Lm7;�=;B;
�D;�9F;OG;T�G;��G;�H;�6H;�YH;vH;[�H;,�H;;�H;>�H;��H;`�H;��H;V�H;t�H;��H;��H;2�H;��H;��H;t�H;U�H;��H;`�H;��H;;�H;:�H;*�H;_�H;vH;�YH;�6H;�H;��G;U�G;QG;�9F;�D;B;�=;Lm7;Q.;�";�>;P��:~��:R��:֍R:H�9 8(7����T��<�D�      0x[:PCd:��}:+�:��:��:D�:2�;�; ;�+;��3;�:;;�?;��B;�E;tZF; G;O�G;��G;zH;�1H;TH;�pH;�H;��H;#�H;��H;��H;��H;<�H;�H;��H;^�H;4�H;R�H;��H;T�H;4�H;^�H;��H;�H;<�H;��H;��H;��H;"�H;��H;�H;�pH;TH;�1H;wH;��G;O�G;G;uZF;�E;��B;;�?;�:;��3;�+;} ;�;4�;D�: ��:��:-�:��}:0Cd:      ��:�B�:��:�x;��
;�;I�;�}$;Q|,;��3;�_9;_>;9zA;��C;�E;.�F;Q5G;��G;��G;{H;�/H;.QH;@mH;��H;ۗH;ЧH;��H;:�H;��H;U�H;��H;��H;��H;!�H;��H;��H;��H;��H;��H;!�H;��H;��H;��H;R�H;��H;9�H;��H;ҧH;ۗH;��H;?mH;.QH;�/H;}H;��G;��G;Q5G;/�F;�E;��C;9zA;_>;�_9;��3;T|,;�}$;J�;�;��
;�x;��:�B�:      0e;9 ;�";i%;�(;Hj-;^2;�6;ء:;�0>;�A;oYC;\�D;5F;F�F;�XG;0�G;|�G;�H;�1H;.QH;
lH;��H;��H;t�H;k�H;�H;��H;��H;M�H;��H; �H;��H;��H;��H;��H;��H;��H;��H;��H;��H; �H;��H;H�H;��H;��H;�H;m�H;v�H;��H;��H;
lH;-QH;�1H;�H;~�G;/�G;�XG;G�F;5F;\�D;oYC;�A;�0>;١:;�6;^2;Kj-; �(;k%;�";3 ;      p�4;7�4;o�5;m7;�_9;��;;��=;8�?;��A;��C;��D;��E;��F;�)G;ǁG;8�G;�G;vH;�6H;TH;?mH;��H;�H;H�H;��H;��H;e�H;q�H;�H;��H;U�H;*�H;r�H;��H;�H;��H;��H;��H;�H;��H;p�H;)�H;U�H;��H;�H;q�H;b�H;��H;��H;E�H;�H;��H;;mH;TH;�6H;wH;�G;7�G;ǁG;�)G;��F;��E;��D;��C;��A;7�?;��=;��;;�_9;m7;p�5;*�4;      g`?;�?;�?;�@;͘A;��B;ߚC;�D;eiE;F;K�F;G;{nG;E�G;&�G;| H;�!H;U?H;�YH;�pH;��H;��H;F�H;��H;̺H;h�H;��H;F�H;��H;��H;��H;��H;��H;�H;��H;u�H;��H;t�H;��H;�H;��H;��H;��H;��H;��H;E�H;��H;g�H;κH;��H;E�H;��H;��H;�pH;�YH;V?H;�!H;| H;(�G;E�G;{nG;G;K�F;F;giE;�D;ݚC;��B;ԘA;�@;�?;ڈ?;      �mD;	D;v�D;�D;�\E;�E;�0F;��F;��F;9G;�vG;$�G;t�G;��G;mH;�0H;tJH;�aH;$vH; �H;ݗH;x�H; �H;պH;*�H;	�H;��H;Q�H;&�H;7�H;��H;}�H;��H;�H;��H;%�H;h�H;#�H;��H;�H;��H;�H;��H;6�H;%�H;P�H;��H;	�H;,�H;ҺH;��H;x�H;ݗH;#�H;$vH;�aH;qJH;�0H;mH;��G;r�G;%�G;�vG;9G;��F;��F;�0F;�E;�\E;�D;u�D;	D;      ��F;j�F;ܮF;�F;��F;�G;�GG;�pG;W�G;j�G;�G;��G;(H;?*H;�AH;�WH;mkH;M}H;X�H;��H;ͧH;i�H;��H;g�H;�H;u�H;��H;��H;��H;Q�H;O�H;��H;��H;��H;v�H;��H;�H;��H;x�H;��H;��H;��H;O�H;Q�H;��H;��H;��H;u�H;�H;e�H;��H;i�H;ɧH;��H;X�H;P}H;kkH;�WH;�AH;?*H;(H;��G;�G;i�G;X�G;�pG;�GG;�G;��F;�F;ٮF;`�F;      uvG;(yG;#�G;��G;�G;��G;�G;��G;��G;�H;OH;�,H;�@H;�SH;�eH;�vH;߅H;��H;*�H;&�H;��H;�H;d�H;��H;��H;�H;��H;��H; �H;�H;��H;��H;��H;��H;�H;d�H;d�H;b�H;�H;��H;��H;��H;��H;�H;�H;��H;��H; �H;��H;��H;b�H;�H;��H;&�H;*�H;��H;ޅH;�vH;�eH;�SH;�@H;�,H;PH;�H;��G;��G;�G;��G;�G;��G;!�G;(yG;      >�G;��G;��G;��G;��G;��G;[H;$H;�(H;)8H;�GH;AWH;_fH;�tH;z�H;,�H;��H;��H;9�H;��H;9�H;��H;r�H;I�H;L�H;��H;��H;��H;�H;��H;��H;��H;��H;�H;��H;��H;��H;��H;��H;�H;��H;��H;��H;��H; �H;��H;��H;��H;M�H;I�H;q�H;��H;6�H;��H;9�H;��H;��H;,�H;z�H;�tH;]fH;BWH;�GH;*8H;�(H;$H;[H;��G;��G;��G;��G;��G;      �H;� H;x#H;<(H;�.H;�6H;"@H;dJH;qUH;�`H;�lH;QxH;��H;��H;�H;��H;��H;ҳH;>�H;��H;��H;��H;�H;��H; �H;��H;�H;�H;s�H;��H;��H;��H;.�H;��H;��H;�H;1�H;�H;��H;��H;*�H;��H;��H;��H;r�H;�H;�H;��H;"�H;��H;�H;��H;��H;��H;>�H;ԳH;��H;��H;�H;��H;��H;OxH;�lH;�`H;sUH;bJH;"@H;�6H;�.H;<(H;v#H;� H;      �OH;ZPH;�RH;VH;�ZH;�`H;�gH;toH;�wH;?�H;��H;͑H;j�H;��H;��H;��H;ڸH;�H;��H;��H;U�H;J�H;��H;��H;/�H;M�H;�H;��H;��H;��H;��H;)�H;��H;	�H;<�H;a�H;v�H;a�H;<�H;	�H;��H;,�H;��H;��H;��H;��H;�H;M�H;0�H;��H;��H;J�H;T�H;��H;��H;�H;ظH;��H;��H;��H;k�H;͑H;��H;?�H;�wH;uoH;�gH;�`H;�ZH;VH;�RH;WPH;      �sH;atH;�uH;�xH;1|H;��H;ƅH;��H;��H;,�H;ҞH;v�H;�H;2�H;�H;սH;,�H;��H;^�H;A�H;��H;��H;T�H;��H;��H;O�H;��H;��H;��H;��H;�H;��H;�H;Q�H;��H;��H;��H;��H;��H;Q�H;�H;��H;�H;��H;��H;��H;��H;O�H;��H;��H;S�H;��H;��H;B�H;`�H;��H;*�H;ԽH;�H;2�H;�H;t�H;ӞH;.�H;��H;��H;ƅH;��H;-|H;�xH;�uH;atH;      �H;W�H;��H;��H;1�H;��H;n�H;��H;f�H;7�H;7�H;-�H;�H;�H;��H;�H;�H;��H;��H;�H;��H;"�H;*�H;��H;x�H;��H;��H;��H;��H;,�H;��H;�H;M�H;��H;��H;��H;��H;��H;��H;��H;J�H;�H;��H;-�H;��H;��H;��H;��H;{�H;��H;*�H;"�H;��H;�H;��H;��H;�H;�H;��H;�H;�H;,�H;7�H;7�H;h�H;��H;n�H;��H;/�H;��H;��H;S�H;      ��H;�H; �H;��H;��H;	�H;�H;<�H;гH;��H;e�H;R�H;&�H;��H;]�H;��H;��H;��H;X�H;��H;��H;��H;q�H;��H;��H;��H;��H;��H;1�H;��H;	�H;Q�H;��H;��H;��H;��H;	�H;��H;��H;��H;��H;Q�H;	�H;��H;3�H;��H;��H;��H;��H;��H;p�H;��H;��H;��H;X�H;��H;��H;��H;]�H;��H;%�H;P�H;g�H;��H;гH;<�H;�H;�H;�H;��H;�H;�H;      ǰH;�H;��H;�H;��H;��H;ӸH;}�H;3�H;'�H;5�H;-�H;)�H;�H;��H;��H;�H;V�H;v�H;e�H;'�H;��H;��H;�H;�H;��H;}�H;�H;��H;�H;M�H;��H;��H;��H;��H;�H;�H;�H;��H;��H;��H;��H;M�H;	�H;��H;�H;}�H;��H;�H;�H;��H;��H;&�H;d�H;v�H;W�H;�H;��H;��H;�H;)�H;-�H;4�H;'�H;3�H;|�H;ӸH;��H;��H;�H;��H;�H;      (�H;~�H;�H;��H;b�H;ܾH;��H;��H;�H;��H;��H;y�H;��H;S�H;��H;��H;��H;��H;��H;;�H;��H;��H;��H;�H;��H;r�H;�H;��H;��H;=�H;��H;��H;��H;��H;�H;�H;�H;�H;�H;��H;��H;��H;��H;?�H;��H;��H;�H;r�H;��H;�H;��H;��H;��H;9�H;��H;��H;��H;��H;��H;Q�H;��H;y�H;��H;��H;�H;��H;��H;�H;X�H;��H;�H;u�H;      ��H;��H;.�H;��H;)�H;��H;1�H;�H; �H;�H;F�H;��H;��H;��H;��H;��H;��H;Z�H;��H;[�H;��H;��H;��H;x�H;�H;��H;`�H;��H;�H;a�H;��H;��H;��H;�H;�H;0�H;'�H;0�H;�H;�H;��H;��H;��H;a�H;�H;��H;^�H;��H;�H;w�H;��H;��H;��H;[�H;��H;\�H;��H;��H;��H;��H;��H;��H;D�H;�H; �H; �H;1�H;��H;�H;��H;0�H;��H;      \�H;s�H;��H;��H;��H;�H;��H;h�H;U�H;O�H;i�H;u�H;z�H;��H;��H;~�H;6�H;��H;2�H;��H;��H;��H;��H;��H;a�H;�H;`�H;��H;1�H;z�H;��H;��H;�H;�H;�H;)�H;3�H;)�H;�H;�H;�H;��H;��H;{�H;4�H;��H;^�H;�H;a�H;��H;��H;��H;��H;��H;2�H;��H;5�H;~�H;��H;��H;z�H;u�H;i�H;Q�H;V�H;e�H;��H;�H;��H;��H;��H;i�H;      ��H;��H;.�H;��H;)�H;��H;1�H;�H; �H;�H;F�H;��H;��H;��H;��H;��H;��H;Z�H;��H;[�H;��H;��H;��H;x�H;�H;��H;`�H;��H;�H;a�H;��H;��H;��H;�H;�H;0�H;'�H;0�H;�H;�H;��H;��H;��H;a�H;�H;��H;^�H;��H;�H;w�H;��H;��H;��H;[�H;��H;\�H;��H;��H;��H;��H;��H;��H;F�H;�H; �H; �H;1�H;��H;�H;��H;-�H;��H;      '�H;~�H;
�H;��H;b�H;ܾH;��H;��H;�H;��H;��H;y�H;��H;S�H;��H;��H;��H;��H;��H;;�H;��H;��H;��H;�H;��H;r�H;�H;��H;��H;=�H;��H;��H;��H;��H;�H;�H;�H;�H;�H;��H;��H;��H;��H;?�H;��H;��H;�H;r�H;��H;��H;��H;��H;��H;9�H;��H;��H;��H;��H;��H;S�H;��H;y�H;��H;��H;�H;��H;��H;�H;X�H;��H;
�H;t�H;      ɰH;�H;��H;�H;��H;��H;ӸH;|�H;2�H;'�H;5�H;-�H;)�H;�H;��H;��H;�H;V�H;v�H;e�H;*�H;��H;��H;�H;�H;��H;}�H;�H;��H;�H;M�H;��H;��H;��H;��H;�H;�H;�H;��H;��H;��H;��H;M�H;	�H;��H;�H;}�H;��H;�H;�H;��H;��H;&�H;d�H;v�H;W�H;�H;��H;��H;�H;)�H;-�H;5�H;'�H;3�H;{�H;ӸH;��H;��H;�H;��H;�H;      ��H;�H;�H;��H;��H;�H;�H;<�H;гH;��H;g�H;P�H;%�H;��H;]�H;��H;��H;��H;X�H;��H;��H;��H;q�H;��H;��H;��H;��H;��H;1�H;��H;	�H;P�H;��H;��H;��H;��H;	�H;��H;��H;��H;��H;T�H;	�H;��H;3�H;��H;��H;��H;��H;��H;p�H;��H;��H;��H;X�H;��H;��H;��H;_�H;��H;%�H;R�H;e�H;��H;ϳH;:�H;�H;�H;}�H;��H;��H;
�H;      �H;W�H;��H;��H;1�H;��H;p�H;��H;f�H;7�H;7�H;-�H;�H;�H;��H;�H;�H;��H;��H;�H;��H;"�H;,�H;��H;{�H;��H;��H;��H;��H;,�H;��H;�H;L�H;��H;��H;��H;��H;��H;��H;��H;J�H;�H;��H;-�H;��H;��H;��H;��H;x�H;��H;)�H;"�H;��H;�H;��H;��H;�H;�H;��H;�H;�H;,�H;7�H;7�H;h�H;��H;p�H;��H;.�H;��H;��H;R�H;      �sH;atH;�uH;�xH;0|H;��H;ƅH;��H;��H;-�H;ҞH;t�H;�H;5�H;�H;սH;*�H;��H;`�H;B�H;��H;��H;U�H;��H;��H;P�H;��H;��H;��H;��H;�H;��H;�H;Q�H;��H;��H;��H;��H;��H;Q�H;�H;��H;�H;��H;��H;��H;��H;N�H;��H;��H;Q�H;��H;��H;A�H;^�H;��H;*�H;սH;�H;2�H;�H;v�H;ўH;-�H;��H;��H;ƅH;��H;-|H;�xH;�uH;atH;      �OH;ZPH;�RH;VH;�ZH;�`H;�gH;uoH;�wH;?�H;��H;ΑH;k�H;��H;��H;��H;ڸH;�H;��H;��H;X�H;J�H;��H;��H;0�H;N�H;�H;��H;��H;��H;��H;*�H;��H;�H;<�H;a�H;v�H;a�H;<�H;	�H;��H;*�H;��H;��H;��H;��H;�H;L�H;/�H;��H;��H;J�H;T�H;��H;��H;�H;ظH;��H;��H;��H;j�H;͑H;��H;>�H;�wH;uoH;�gH;�`H;�ZH;VH;�RH;XPH;      �H;� H;}#H;;(H;�.H;�6H;%@H;fJH;qUH;�`H;�lH;QxH;��H;��H;�H;��H;��H;ҳH;>�H;��H;��H;��H;�H;��H;"�H;��H;�H;�H;s�H;��H;��H;��H;-�H;��H;��H;�H;1�H;�H;��H;��H;-�H;��H;��H;��H;s�H;�H;�H;��H; �H;��H;�H;��H;��H;��H;>�H;ӳH;��H;��H;�H;��H;��H;QxH;�lH;�`H;sUH;dJH;%@H;�6H;�.H;7(H;{#H;� H;      >�G;��G;��G;��G;��G;��G;[H;'H;�(H;*8H;�GH;BWH;]fH;�tH;z�H;,�H;��H;��H;9�H;��H;;�H;��H;r�H;I�H;M�H;��H;��H;��H;�H;��H;��H;��H;��H;�H;��H;��H;��H;��H;��H;�H;��H;��H;��H;��H; �H;��H;��H;��H;L�H;I�H;q�H;��H;7�H;��H;9�H;��H;��H;-�H;z�H;�tH;_fH;AWH;�GH;)8H;�(H;$H;[H;��G;��G;��G;��G;��G;      ovG;(yG; �G;��G;ݝG;��G; �G;��G;��G;�H;PH;�,H;�@H;�SH;�eH;�vH;߅H;��H;*�H;(�H;��H;�H;d�H;��H;��H;�H;��H;��H; �H;�H;��H;��H;��H;��H;�H;b�H;d�H;b�H;�H;��H;��H;��H;��H;�H;�H;��H;��H;�H;��H;��H;b�H;�H;��H;%�H;*�H;��H;ޅH;�vH;�eH;�SH;�@H;�,H;PH;�H;��G;��G; �G;��G;��G;��G; �G;yG;      ��F;b�F;�F;�F;��F;�G;�GG;�pG;W�G;j�G;�G;��G;(H;?*H;�AH;�WH;mkH;N}H;X�H;��H;ϧH;i�H;��H;g�H;�H;u�H;��H;��H;��H;S�H;O�H;��H;��H;��H;u�H;��H;�H;��H;x�H;��H;��H;��H;O�H;P�H;��H;��H;��H;u�H;�H;e�H;��H;i�H;ɧH;��H;X�H;N}H;kkH;�WH;�AH;?*H;(H;��G;�G;i�G;W�G;�pG;�GG;�G;��F;�F;�F;Z�F;      �mD;	D;v�D;�D;�\E;�E;�0F;��F;��F;9G;�vG;%�G;r�G;��G;mH;�0H;rJH;�aH;$vH;#�H;��H;x�H; �H;պH;,�H;	�H;��H;P�H;&�H;7�H;��H;}�H;��H;�H;��H;#�H;h�H;#�H;��H;�H;��H;��H;��H;6�H;#�H;Q�H;��H;	�H;*�H;ӺH;��H;x�H;ݗH;"�H;$vH;�aH;qJH;�0H;mH;��G;t�G;$�G;�vG;9G;��F;��F;�0F;�E;�\E;�D;u�D;	D;      m`?;�?;�?;�@;ƘA;��B;ۚC;�D;giE;F;L�F;G;}nG;E�G;(�G;| H;�!H;S?H;�YH;�pH;��H;��H;F�H;��H;κH;h�H;��H;E�H;��H;��H;��H;��H;��H;�H;��H;u�H;��H;u�H;��H;�H;��H;��H;��H;��H;��H;F�H;��H;h�H;̺H;��H;E�H;��H;��H;�pH;�YH;V?H;�!H;| H;(�G;E�G;{nG;G;I�F;F;giE;�D;ۚC;��B;՘A;�@;�?;׈?;      m�4;B�4;}�5;
m7;�_9;��;;��=;8�?;��A;��C;��D;��E;��F;�)G;ǁG;8�G;�G;uH;�6H;TH;BmH;��H;�H;H�H;��H;��H;e�H;q�H;�H;��H;U�H;*�H;r�H;��H;�H;��H;��H;��H;�H;��H;q�H;*�H;U�H;��H;�H;q�H;b�H;��H;��H;E�H;�H;��H;<mH;TH;�6H;wH;�G;8�G;ȁG;�)G;��F;��E;��D;��C;��A;7�?;��=;��;;�_9;m7;s�5;1�4;      0e;9 ;�";k%;
�(;Jj-;^2;�6;ء:;�0>;�A;oYC;\�D;5F;F�F;�XG;/�G;|�G;�H;�1H;/QH;
lH;��H;��H;v�H;k�H;�H;��H;��H;M�H;��H; �H;��H;��H;��H;��H;��H;��H;��H;��H;��H; �H;��H;H�H;��H;��H;�H;m�H;t�H;��H;��H;
lH;-QH;�1H;�H;~�G;/�G;�XG;G�F;5F;\�D;qYC;�A;�0>;ۡ:;�6;^2;Hj-;�(;i%;�";3 ;      ���:�B�:��:�x;��
;�;M�;�}$;Q|,;��3;�_9;_>;9zA;��C;�E;/�F;S5G;��G;��G;{H;�/H;.QH;@mH;��H;ۗH;ҧH;��H;9�H;��H;U�H;��H;��H;��H; �H;��H;��H;��H;��H;��H;!�H;��H;��H;��H;R�H;��H;:�H;��H;ЧH;ۗH;��H;?mH;.QH;�/H;}H;��G;��G;P5G;.�F;�E;��C;9zA;^>;�_9;��3;T|,;�}$;M�;�;��
;�x;��:�B�:      (x[:TCd:��}:)�:��:��:F�:4�;�; ;�+;��3;�:;;�?;��B;�E;uZF; G;O�G;��G;}H;�1H;TH;�pH;�H;��H;%�H;��H;��H;��H;<�H;�H;��H;^�H;4�H;T�H;��H;T�H;4�H;^�H;��H;�H;<�H;��H;��H;��H;!�H;��H;�H;�pH;TH;�1H;xH;��G;O�G;G;tZF;�E;��B;;�?;�:;��3;�+;} ;�;5�;F�: ��:��:'�:��}:(Cd:      D�S�@�D�T������ 1(7�9֍R:T��:z��:P��:�>;�";Q.;Lm7;�=;B;
�D;�9F;QG;T�G;��G;�H;�6H;�YH;vH;^�H;-�H;:�H;>�H;��H;`�H;��H;X�H;t�H;��H;��H;2�H;��H;��H;t�H;U�H;��H;`�H;��H;;�H;;�H;)�H;^�H;vH;�YH;�6H;�H;��G;U�G;OG;�9F;�D;B;�=;Lm7;Q.;�";�>;P��:~��:R��:ҍR:@�9 7(7����T��@�D�      
E^��/X��qF�.}*�'���P��|�D��ˬ��i:��:w��:T�;¡;e�);��4;;�<;7�A;L�D;�9F;G;��G;|�G;wH;V?H;�aH;Q}H;��H;��H;ֳH;�H;��H;��H;��H;Y�H;��H;`�H;��H;`�H;��H;Y�H;��H;��H;��H;�H;ӳH;��H;��H;S}H;�aH;R?H;uH;|�G;��G;G;�9F;L�D;6�A;;�<;��4;b�);¡;T�;w��:��:�i:�ˬ�|�D��P��!��.}*��qF�0X�      ��ﻪ��`�ܻE�ƻf󩻴��xFL��������`����-:>�:���:;�>&;��3;~9<;9�A;�D;yZF;T5G;2�G;�G;�!H;nJH;nkH;��H;��H;��H;ظH;&�H; �H;��H;�H;��H;��H;0�H;��H;��H;�H;��H; �H;&�H;׸H;��H;��H;ۅH;okH;nJH;�!H;�G;2�G;Q5G;{ZF;�D;<�A;z9<;��3;�>&;;���:>�:��-:p���������xFL����e�F�ƻ`�ܻ���      r�V��5S��6H���6�E� �U,��?ػ9G���D^������D�@��9�4�:7�:I�;%;��3;>�<;�B;�E;2�F;�XG;9�G;� H;�0H;�WH;�vH;-�H;��H;��H;νH;�H;��H;��H;��H;��H;w�H;��H;��H;��H;��H;�H;νH;��H;��H;,�H;�vH;�WH;�0H;| H;8�G;�XG;1�F;�E;�B;?�<;��3;%;K�;3�:�4�:8��9��D�����D^�9G���?ػT,�E� ���6��6H��5S�      "��.��MȤ����� ���A�f�w�=����=�ܻ�*��Lo5�<��� �(7��}:�n�:H�;�>&;��4;�=;��B;�E;F�F;ʁG;+�G;jH;�AH;�eH;z�H;�H;��H;�H;��H;_�H;��H;��H;��H;��H;��H;��H;��H;\�H;��H;�H;��H;�H;x�H;�eH;�AH;kH;&�G;āG;F�F;�E;��B;�=;��4;�>&;H�;�n�:��}: �(7>���Lo5��*��<�ܻ���w�=�@�f� �������MȤ�.��      �c��8���������Ҽ����������r�JE:�E,�Iߵ�s/X�d�º�Ĭ���}:;�:;g�);Mm7;@�?;��C;8F;�)G;H�G;��G;@*H;�SH;�tH;��H;��H;.�H;�H;��H;�H;M�H;��H;��H;��H;M�H;�H;��H;�H;.�H;��H;��H;�tH;�SH;C*H;��G;C�G;�)G;8F;��C;@�?;Lm7;i�);;9�:��}:�Ĭ�f�ºs/X�Jߵ�E,�IE:���r�����������Ҽ�켻����8�      ''K��G���>��0�`y��c����X��� ��Y�V�)���ƻ�od�f�º �(7�4�:���:¡;Q.;�:;:zA;\�D; �F;�nG;t�G;,H;�@H;_fH;��H;g�H;�H;�H;#�H;)�H;��H;��H;w�H;��H;��H;)�H;#�H;�H;�H;f�H;��H;_fH;�@H;.H;w�G;}nG;��F;\�D;:zA;�:;Q.;¡;���:�4�: �(7f�º�od��ƻ)��X�V� ��X�����众c�`y��0���>��G�      	���4Z��Ґ����}��c���D�6/%��8���Ҽ2c��6�f�����ƻt/X�:���@��9@�:X�;�";��3;`>;oYC;��E;G;$�G;��G;�,H;>WH;OxH;đH;o�H;%�H;L�H;*�H;p�H;�H;n�H;�H;o�H;)�H;I�H;&�H;m�H;ÑH;MxH;>WH;�,H;��G;&�G;G;��E;oYC;e>;��3;�";W�;<�:0��9:���u/X��ƻ���6�f�2c����Ҽ�8�6/%���D��c���}�Ґ��4Z��      �Pν �ʽR8���������ѐ��d�f���;�4�����EȤ�6�f�)��Kߵ�Ko5���D���-:y��:�>;�+;�_9;�A;��D;N�F;�vG;�G;SH;�GH;�lH;��H;ўH;3�H;e�H;1�H;��H;?�H;c�H;?�H;��H;1�H;c�H;3�H;ϞH;��H;�lH;�GH;OH;�G;�vG;I�F;��D;�A;�_9;�+;�>;y��:��-:��D�Ko5�Kߵ�)��6�f�EȤ����4����;�d�f�ѐ���������R8�� �ʽ      ���j9�\[��s�~�ؽ���
t����}���G������2c��Y�V�F,��*�����`����:R��:� ;��3;�0>;��C;F;9G;n�G;�H;'8H;�`H;:�H;*�H;7�H;��H;&�H;��H;�H;O�H;�H;��H;&�H;�H;6�H;*�H;:�H;�`H;)8H;�H;p�G;9G;F;��C;�0>;��3;} ;R��:��:�������*��F,�Y�V�2c���������G���}�
t�����~�ؽ�s�\[�j9�      ��=�ڀ:���0��Q"��������Pν�榽B����G�4����Ҽ ��JE:�;�ܻ�D^������i:~��:�;S|,;֡:;��A;giE;��F;[�G;��G;�(H;tUH;�wH;��H;c�H;ϳH;/�H;�H;��H;N�H;��H;�H;/�H;ɳH;b�H;��H;�wH;qUH;�(H;��G;]�G;��F;diE;��A;֡:;U|,;�;z��:�i:�����D^�;�ܻJE:� ����Ҽ4����G�B���榽�Pν�������Q"���0�ڀ:�      5Dx�8�s���f�xS�ڀ:����\[��7ս�榽��}���;��8�W�����r����7G���� ˬ�Z��:8�;�}$;�6;8�?;�D;��F;�pG;��G;H;dJH;ooH;y�H;��H;7�H;u�H;��H;��H;b�H;��H;��H;u�H;4�H;��H;y�H;ooH;bJH; H;��G;�pG;�F;�D;8�?;�6;�}$;7�;X��:�ʬ����7G�������r�W����8���;���}��榽�7ս\[����ڀ:�xS���f�8�s�      �*���0��॒�=����k��H��#%�\[��Pν
t��d�f�6/%���伈���w�=��?ػ|FL�p�D�R:H�:G�;U2;��=;ۚC;�0F;�GG;��G;ZH; @H;�gH;��H;l�H;�H;ѸH;��H;*�H;��H;*�H;��H;иH;�H;l�H;��H;�gH;@H;ZH;��G;�GG;�0F;ךC;��=;V2;J�;H�:R:l�D�~FL��?ػw�=��������6/%�d�f�
t���Pν\[��#%��H��k�=���॒��0��      *�þ
���"����R��~쏾8�s��H�����������ѐ����D��c�����@�f�T,�����P����9 ��:�;Aj-;��;;��B;�E;�G;��G;��G;�6H;�`H;��H;��H;�H;��H;߾H;��H;�H;��H;߾H;��H;�H;��H;��H;�`H;�6H;��G;��G;�G;�E;��B;��;;Aj-;�; ��:��9�P�����T,�@�f������c���D�ѐ�������������H�8�s�~쏾�R��"���
���      C��2�很Yؾ*�þĪ�~쏾�k�ڀ:���~�ؽ�����c�`y���Ҽ����D� �d�"�� 4(7��:��
;
�(;�_9;͘A;�\E;��F;ݝG;��G;�.H;�ZH;&|H;-�H;��H;��H;L�H;�H;��H;�H;J�H;��H;�H;/�H;&|H;�ZH;�.H;��G;ޝG;��F;�\E;ɘA;�_9;�(;��
;��: 5(7 ��e�D� �������Ҽ`y��c�����~�ؽ��ڀ:��k�~쏾Ī�*�þ�Yؾ2��      %��P������AI�*�þ�R��=���xS��Q"��s������}��0��켋�����6�C�ƻ.}*�����-�:�x;r%;m7;�@;�D;�F;��G;��G;<(H;VH;�xH;��H;~�H;ܲH;�H;��H;��H;��H;�H;ܲH;}�H;��H;�xH;VH;8(H;��G;��G;�F;�D;�@;m7;r%;�x;+�:����/}*�D�ƻ��6��������0���}�����s��Q"�xS�=����R��*�þAIᾦ���P��      ���T��:�
������Yؾ"���॒���f���0�\[�R8��Ґ����>�����MȤ��6H�^�ܻ rF������}:��:{";l�5;�?;��D;�F;#�G;��G;{#H;�RH;�uH;��H;��H;��H;�H;)�H;��H;)�H;�H;��H;��H;��H;�uH;�RH;x#H;��G;#�G;�F;��D;�?;o�5;{";��:��}:����qF�_�ܻ�6H�MȤ�������>�Ґ��R8��\[���0���f�॒�"����Yؾ����:�
�T��      �� ����T��P��2��
����0��8�s�ڀ:�i9� �ʽ4Z���G��8�.���5S�����/X�4�D�Cd:�B�: ;1�4;ڈ?;D;]�F;'yG;��G;� H;VPH;QtH;K�H;�H;�H;k�H;��H;o�H;��H;m�H;�H;�H;L�H;QtH;SPH;� H;��G;&yG;_�F;D;ֈ?;7�4; ;�B�:Cd:4�D��/X���껰5S�.���8��G�4Z�� �ʽi9�ڀ:�8�s��0��
���2��P��T�����      HEb�c]��N���7����u� ���˾��,�j��!,�t���O��Gm�-��9,˼��x�W���1��⥥��:��:�;Y�1;H,>;��C;�wF;	�G;� H;?H;iH;g�H;��H;P�H;3�H;��H;A�H;��H;A�H;��H;3�H;O�H;��H;g�H;iH;	?H;� H;	�G;�wF;��C;E,>;\�1;�;��:�:⥥��1��X����x�:,˼-��Gm�O��t����!,�,�j�����˾u� ������7��N�c]�      c]�f�W��TI�v3� E�������Ǿx����f�:)�'��t;���Fi��k���Ǽ�[t�J�	�$Ȅ��W����:$��:��;qJ2;fZ>;[	D;�F;W�G;-H;�?H;�iH;��H;��H;��H;O�H;��H;l�H;��H;l�H;��H;O�H;��H;��H;��H;�iH;�?H;-H;W�G;�F;[	D;aZ>;vJ2;��; ��:��:�W��#Ȅ�J�	��[t���Ǽ�k��Fi�t;��(��:)��f�x�����Ǿ���� E�v3��TI�g�W�      �N��TI���;�1�'�l��쾂���z󐾶Z��K ��s�C����&^���"����g����Ĩu�� ���3<:7��:;}g3;	�>;�BD;ɖF;��G;�H;]BH;�kH;j�H;��H;?�H;�H;��H;��H;[�H;��H;��H;�H;=�H;��H;j�H;�kH;ZBH;�H;��G;ʖF;�BD;�>;�g3;;7��:�3<:� ��¨u������g��"����&^�C����s潧K ��Z�z󐾂�����l�1�'���;��TI�      ��7�v3�1�'����u� ��{Ծ!���J���|�F�����ӽ���a�L�Kv��뮼PT�ߘ껾PV�<�=�$*i:���:�z ;�$5;��?; �D;�F;
�G;�H;�FH;�nH;��H;��H;��H;��H;J�H;i�H;�H;i�H;J�H;��H;��H;��H;��H;�nH;�FH;�H;
�G;�F;�D;��?;�$5;�z ;���:*i:<�=��PV����PT��뮼Kv�a�L�����ӽ���|�F�J���!����{Ծu� ����1�'�v3�      ��� E�l�u� �X�ݾm���X͓��f��>/�����'���섽Q�6��t�w��]�:�Tʻk.�`ڷ��t�:�;��$;�Y7;n�@;
E;2�F;M�G;�H;OLH;�rH;ƏH;ݤH;5�H;3�H;D�H;\�H;��H;\�H;C�H;3�H;3�H;ߤH;ƏH;�rH;MLH;�H;N�G;0�F;
E;j�@;�Y7;��$;�;�t�:`ڷ�i.�Tʻ]�:�w���t�Q�6��섽�'������>/��f�X͓�m���Y�ݾu� �l� E�      u� ��������{Ծm���x���^�x��SC��^��޽A���{�e�)��E�Ѽ&G������R����� �8)��:�Y;i�);�9;�A;҄E;�G;2�G;z!H;SSH;�wH;��H;��H;R�H;��H;��H;��H;��H;��H;��H;��H;R�H;��H;��H;�wH;OSH;y!H;1�G;�G;τE;�A;�9;i�);�Y;#��: �8����R�����&G��E�Ѽ)��{�e�A����޽�^��SC�^�x�x���m����{Ծ�쾣���      ��˾��Ǿ����!���X͓�^�x���J��K �q��� ������?����뮼+�[�����2|�pW����:��:�';�/;~g<;�C;�F;�NG;��G;@-H;�[H;�}H;חH;تH;͸H;��H;�H;��H;�H;��H;�H;��H;͸H;٪H;ٗH;�}H;}[H;@-H;��G;�NG;~F;�C;|g<;�/;�';��:��:jW�� 3|����+�[��뮼���?���� ��q����K ���J�^�x�X͓�!���������Ǿ      ��x���z�J����f��SC��K �qn���Ž����Z��k�!}ռ-X��_y-�$���V.�����P�:�+�:��;64;O�>;D;�wF;I�G;��G;�9H;kdH;��H;��H;q�H;�H;��H;��H;d�H;��H;d�H;��H;��H;}�H;t�H;��H;��H;hdH;�9H;��G;I�G;�wF;D;O�>;64;��;�+�:�P�:���W.�$���_y-�-X��!}ռ�k��Z�����Žqn���K ��SC��f�J���z�x���      +�j��f��Z�|�F��>/��^�q����ŽH ���Fi��Q+�}t�oT��n�W�����1���Ⱥ�X�9�P�:�Y;��(;"�8;A;�E;�F;�G;�H;GH;�mH;��H;ҡH;O�H;~�H;��H;��H;�H;�H;�H;��H;��H;~�H;Q�H;ҡH;��H;�mH;GH;�H;��G;�F;�E;A;"�8;��(;�Y;�P�: Y�9�Ⱥ�1�����n�W�oT��}t�Q+��Fi�H ���Žq����^��>/�|�F��Z��f�      �!,�;)��K ��������޽ ������Fi��0����鷼��x�����.��>�(�|��p+i:���:X�;��0;e�<;�C;��E;%=G;�G;%H;wTH;�wH;��H;)�H;]�H;��H;P�H;��H;��H;��H;��H;��H;P�H;��H;_�H;)�H;��H;�wH;wTH;%H;�G;"=G;��E;�C;e�<;��0;W�;���:x+i:���>�(��.�������x�鷼����0��Fi���� ���޽�������K �;)�      t���'��s��ӽ�'��A�������Z��Q+�����"��G����0���׻��b�W���Y�9
��:B`;�*';Z7;&$@;@�D;�F;,�G;��G;L8H;bH;�H;j�H;��H;��H;��H;��H;��H;^�H;J�H;^�H;��H;��H;��H;��H;��H;i�H;�H;bH;K8H;��G;(�G;�F;=�D;&$@;Z7;�*';F`;��:�Y�9W����b���׻��0�G���"������Q+��Z����A����'���ӽ�s�(��      O��u;��C�������섽{�e��?��k�}t�鷼G���e7�����Ǆ�F0�@�t�bu�:9,�:�;�1;l�<;{�B;>�E;G;	�G;tH;�JH;ooH;�H;��H;'�H;��H;��H;.�H;��H;�H;��H;�H;��H;0�H;��H;��H;'�H;��H;�H;qoH;�JH;vH;�G;G;<�E;{�B;l�<;�1;�;?,�:`u�: �t�F0��Ǆ���껃e7�G��鷼}t��k��?�{�e��섽���C���u;��      Gm��Fi��&^�b�L�R�6�)����!}ռoT����x���0�����������׷�do`:��:6�;C�*;R�8;)�@;Q�D;~�F;~G;��G;�1H;�[H;�|H;ѕH;�H;��H;��H;��H;��H;��H;��H;��H;��H;��H;��H;��H;��H;��H;�H;ЕH;�|H;�[H;�1H;��G;~G;{�F;Q�D;)�@;R�8;C�*;:�;��:ho`:�׷���������껿�0���x�oT��!}ռ��)��R�6�b�L��&^��Fi�      -���k��Kv��t�D�Ѽ�뮼-X��m�W������׻�Ǆ���X��v5<:���:�Y;�t%;%5;�Z>;aC;��E;L*G;z�G;+H;HH;�lH;�H;�H;֯H;�H;��H;��H;�H;��H;��H;@�H;��H;��H;�H;��H;��H;�H;ԯH;�H;�H;~lH;HH;*H;y�G;I*G;��E;aC;�Z>;%5;�t%;�Y;���:~5<:H�����Ǆ���׻���m�W�-X���뮼D�Ѽ�t�Kv���k�      9,˼��Ǽ�"���뮼w��&G��+�[�`y-�����.����b�J0��׷�r5<:#M�:];��!;�J2;�g<;j0B;CCE;A�F;e�G;�G;�4H;�\H;|H;��H;��H;m�H;��H;R�H;��H;a�H;d�H;�H;��H; �H;e�H;e�H;��H;U�H;��H;j�H;��H;��H;|H;�\H;�4H;�G;`�G;A�F;BCE;k0B;�g<;�J2;��!;];)M�:r5<:�׷�J0㺺�b��.�����ay-�+�[�&G��w���뮼�"����Ǽ      ��x��[t���g�PT�]�:�������&����1��>�(�W����t�`o`:���:];%{ ;��0;v;;=A;0�D;�wF;�cG;l�G;�!H;�MH;�oH;��H;��H;ׯH;��H;x�H;��H;k�H;��H;�H;��H;8�H;��H;�H;��H;k�H;��H;z�H;��H;ӯH;��H;��H;�oH;�MH;�!H;i�G;�cG;�wF;/�D;=A;w;;��0;&{ ;];���:`o`:@�t�W��?�(��1��&���������^�:�PT���g��[t�      X��H�	������Tʻ�R���2|�X.��Ⱥ����Y�9^u�:��:�Y;��!;��0;�:;ȵ@; CD;�2F;�8G;��G;�H;@H;;dH;؀H;��H;Z�H;]�H;`�H;��H;�H;��H;��H;��H;�H;��H;�H;��H;��H;��H;�H;��H;_�H;Z�H;Z�H;��H;ڀH;:dH;{@H;�H;��G;�8G;�2F; CD;̵@;�:;��0;��!;�Y;��:`u�:�Y�9����ȺX.��2|��R��Tʻ�����J�	�      �1��&Ȅ�Ĩu��PV�p.����rW������X�9p+i:
��:7,�:6�;�t%;�J2;s;;ȵ@;�D;"F;?G;��G;�H;�5H;�ZH;IxH;S�H;>�H;+�H;(�H;n�H;��H;-�H;B�H;=�H;P�H;m�H;��H;m�H;Q�H;=�H;B�H;0�H;��H;n�H;%�H;+�H;;�H;V�H;IxH;�ZH;�5H;�H;��G;@G;"F;�D;ȵ@;s;;�J2;�t%;6�;9,�:
��:l+i: Y�9���rW�����j.��PV�Ĩu�*Ȅ�      ڥ���W��� ��8�=��ڷ�`�8 �:�P�:�P�:���:B`;�;@�*;
%5;�g<;=A;CD;"F;�G;��G;}�G;�-H;/SH;mqH;��H;ԝH;��H;)�H;M�H;�H;�H;��H;g�H;��H;��H;��H;��H;��H;��H;��H;g�H;��H;�H;�H;L�H;)�H;��H;՝H;��H;iqH;,SH;�-H;z�G;��G;�G;$F;CD;=A;�g<;
%5;B�*;�;D`;���:�P�:�P�:�:@�8Pڷ�8�=�� ���W��       �:ȡ:�3<:*i:�t�:��:��:�+�:�Y;W�;�*';�1;N�8;�Z>;f0B;)�D;�2F;:G;��G;2�G;�)H;�NH;�lH;a�H;}�H;��H;��H;D�H;��H;�H;L�H;=�H;F�H;n�H;��H;��H;��H;��H;��H;n�H;E�H;?�H;M�H;�H;��H;C�H;��H;��H;}�H;\�H;�lH;�NH;�)H;2�G;��G;<G;�2F;)�D;g0B;�Z>;P�8;�1;�*';T�;�Y;�+�:��:#��:�t�:*i:�3<:��:      ��:<��:?��:���:�;�Y;�';��;��(;��0;�Y7;f�<;%�@;aC;BCE;�wF;�8G;��G;|�G;�)H;�LH;jH;J�H;q�H;��H;�H;ѾH;y�H;:�H;��H;)�H;h�H;��H;��H;��H;��H;��H;��H;��H;��H;��H;k�H;*�H;��H;7�H;x�H;ϾH;�H;��H;m�H;H�H;jH;�LH;�)H;|�G;��G;�8G;�wF;BCE;aC;&�@;f�<;�Y7;��0;��(;��;�';�Y;�;���:?��:��:      �;��;(;�z ;��$;p�);�/;:4;$�8;d�<;'$@;z�B;P�D;��E;C�F;�cG;��G;�H;�-H;�NH;jH;^�H;ʔH;ƤH;�H;ּH;��H;��H;`�H;�H;��H;D�H;`�H;��H;��H;��H;��H;��H;��H;��H;]�H;F�H;��H; �H;\�H;��H;��H;׼H;�H;¤H;ǔH;\�H;jH;�NH;�-H;�H;��G;�cG;D�F;��E;P�D;z�B;&$@;d�<;&�8;:4;�/;s�);��$;�z ;';��;      \�1;sJ2;}g3;�$5;�Y7;�9;|g<;N�>;A;�C;<�D;=�E;{�F;I*G;a�G;g�G;�H;�5H;-SH;�lH;J�H;ʔH;A�H;�H;��H;��H;v�H;I�H;�H;��H;��H;��H;��H;��H;��H;A�H;��H;A�H;��H;��H;��H;��H;��H;��H;�H;I�H;u�H;��H;��H;�H;?�H;ʔH;F�H;�lH;-SH;�5H;�H;g�G;c�G;J*G;{�F;=�E;?�D;�C;A;N�>;|g<;�9;�Y7;�$5;�g3;hJ2;      Z,>;uZ>;�>;��?;n�@;�A;�C;D;�E;��E;�F;G;~G;y�G;�G;�!H;{@H;�ZH;jqH;_�H;m�H;äH;�H;3�H;��H;��H;`�H;+�H;	�H;�H;�H;O�H;��H;��H;|�H;��H;�H;��H;|�H;��H;��H;P�H;~�H;�H;�H;+�H;`�H;��H;��H;/�H;�H;äH;j�H;_�H;jqH;�ZH;{@H;�!H;�G;y�G;~G;G;�F;��E;�E;D;�C;�A;v�@;��?;�>;gZ>;      ��C;b	D;yBD;!�D;
E;҄E;}F;�wF;�F;=G;'�G;	�G;��G;-H;�4H;�MH;?dH;JxH;��H;��H;��H;�H;��H;��H;`�H;�H;��H;��H;��H;��H;��H;��H;��H;r�H;�H;w�H;~�H;v�H;�H;r�H;��H;��H;��H;��H;��H;��H;��H;�H;`�H;��H;��H;�H;��H;��H;��H;MxH;<dH;�MH;�4H;+H;��G;	�G;'�G;=G;�F;�wF;}F;҄E;
E;!�D;xBD;a	D;      �wF;�F;��F;�F;-�F;�G;�NG;C�G;y�G;�G;��G;sH;�1H;HH;�\H;�oH;؀H;Q�H;НH;��H;�H;ӼH;}�H;��H;�H;��H;Q�H;O�H;��H;��H;L�H;��H;h�H;,�H;��H;��H;��H;��H;��H;,�H;e�H;��H;J�H;��H;��H;N�H;Q�H;��H;�H;��H;}�H;ԼH;޳H;��H;НH;S�H;րH;�oH;�\H;HH;�1H;sH;��G;
�G;{�G;B�G;�NG;�G;4�F;�F;��F;�F;      �G;W�G;��G;
�G;P�G;4�G;��G;��G;�H;%H;I8H;�JH;�[H;~lH;|H;��H;��H;;�H;��H;��H;ѾH;��H;u�H;d�H;��H;V�H;6�H;��H;}�H;*�H;k�H;D�H;�H;��H;�H;;�H;I�H;;�H;�H;��H;�H;D�H;j�H;(�H;|�H;��H;6�H;S�H;��H;b�H;t�H;��H;ξH;��H;��H;=�H;��H;��H;|H;~lH;�[H;�JH;K8H;%H;�H;��G;��G;1�G;U�G;�G;��G;U�G;      � H;.H;�H;�H;�H;w!H;C-H;�9H; GH;yTH;bH;toH;�|H;	�H;��H;��H;W�H;'�H;%�H;F�H;v�H;��H;J�H;.�H;��H;O�H;��H;��H;�H;:�H;;�H;�H;��H;�H;N�H;��H;��H;��H;N�H;�H;��H;�H;;�H;7�H;�H;��H;��H;O�H;��H;.�H;I�H;��H;t�H;D�H;'�H;(�H;W�H;��H;��H;�H;�|H;toH;bH;yTH;GH;�9H;C-H;y!H;�H;�H;�H;;H;      ?H;�?H;ZBH;�FH;LLH;OSH;�[H;idH;�mH;�wH;�H;�H;ѕH;�H;��H;ׯH;]�H;$�H;L�H;��H;:�H;\�H;�H;�H;��H;��H;y�H;�H;X�H;(�H;��H;��H;	�H;m�H;��H;��H;��H;��H;��H;m�H;�H;��H;��H;(�H;X�H;�H;|�H;��H;��H;�H;�H;\�H;7�H;��H;L�H;'�H;]�H;ׯH;��H;�H;ѕH;�H;�H;�wH;�mH;kdH;�[H;NSH;SLH;�FH;ZBH;�?H;      iH;�iH;�kH;�nH;�rH; xH;�}H;��H;��H; �H;p�H;͡H;�H;ݯH;m�H;��H;b�H;h�H;�H;#�H;��H; �H;��H;�H;��H;��H;'�H;:�H;(�H;�H;��H;�H;Z�H;��H;��H;��H;��H;��H;��H;��H;W�H;�H;��H;�H;&�H;9�H;&�H;��H;��H;�H;��H; �H;��H;"�H;�H;j�H;`�H;��H;m�H;گH;�H;ˡH;r�H;�H;��H;��H;�}H; xH;�rH;�nH;�kH;�iH;      h�H;�H;u�H;��H;ЏH;��H;ݗH;ƜH;סH;*�H;��H;/�H;��H;�H;��H;�H;��H;�H;�H;Q�H;-�H;��H;��H;��H;��H;L�H;f�H;;�H;��H;��H;�H;f�H;��H;��H;�H;�H; �H; �H;�H;��H;��H;i�H;�H;��H;��H;=�H;i�H;J�H;��H;��H;��H;��H;*�H;Q�H;�H;�H;��H;~�H;��H;�H;��H;/�H;��H;/�H;סH;ƜH;ݗH;��H;͏H;��H;t�H;�H;      ��H;�H;��H;��H;�H;��H;٪H;z�H;R�H;]�H;��H;��H;��H;��H;X�H;��H;�H;-�H;��H;D�H;n�H;F�H;��H;Q�H;��H;��H;A�H;�H;��H;�H;e�H;��H;��H;�H;�H;<�H;X�H;<�H;�H;�H;��H;��H;e�H;�H;��H;�H;B�H;��H;��H;S�H;��H;G�H;n�H;D�H;��H;0�H;	�H;��H;X�H;��H;��H;��H;��H;`�H;U�H;w�H;ڪH;��H;�H;��H;��H;��H;      S�H;��H;F�H;��H;<�H;O�H;͸H;��H;��H;��H;��H;��H;��H;��H;��H;q�H;��H;<�H;g�H;I�H;��H;]�H;��H;��H;��H;g�H;�H;��H;�H;^�H;��H;��H;�H;0�H;U�H;J�H;=�H;J�H;T�H;0�H;�H;��H;��H;_�H;�H;��H;�H;g�H;��H;��H;��H;^�H;��H;J�H;i�H;?�H;��H;q�H;��H;��H;��H;��H;��H;��H;��H;��H;͸H;T�H;5�H;��H;F�H;��H;      <�H;W�H;�H;��H;9�H;��H;��H;��H;��H;P�H;��H;3�H;��H;�H;e�H;��H;��H;:�H;��H;t�H;��H;��H;��H;��H;j�H;'�H;��H;�H;j�H;��H;��H;�H;)�H;=�H;i�H;t�H;T�H;t�H;i�H;=�H;(�H;	�H;��H;��H;m�H;�H;��H;)�H;m�H;��H;��H;��H;��H;t�H;��H;=�H;��H;��H;f�H;�H;��H;5�H;��H;P�H;��H;��H;��H;��H;/�H;��H;�H;P�H;      ��H;�H;��H;P�H;\�H;��H;�H;��H;��H;��H;��H;��H;��H;��H;h�H;�H;��H;L�H;��H;��H;��H;��H;��H;}�H;�H;��H;��H;M�H;��H;��H;�H;�H;R�H;j�H;M�H;j�H;��H;j�H;M�H;j�H;O�H; �H;�H;��H;��H;M�H;��H;��H;�H;|�H;��H;��H;��H;��H;��H;M�H;��H;�H;h�H;��H;��H;��H;��H;��H;��H;��H;�H;��H;R�H;N�H;��H;�H;      8�H;r�H;��H;l�H;k�H;��H;��H;m�H;�H;��H;e�H;'�H;��H;��H;!�H;��H;�H;f�H;��H;��H;��H;�H;>�H;��H;n�H;��H;6�H;��H;��H;��H;�H;?�H;H�H;x�H;j�H;`�H;q�H;`�H;j�H;u�H;F�H;A�H;�H;��H;��H;��H;6�H;��H;p�H;��H;>�H;�H;��H;��H;��H;g�H;�H;��H;"�H;��H;��H;(�H;d�H;��H;�H;j�H;��H;��H;`�H;l�H;��H;i�H;      ��H;��H;g�H;�H;��H;��H;�H;��H;�H;��H;S�H;��H;��H;I�H;��H;?�H;��H;��H;��H;��H;��H;��H;��H;�H;u�H;��H;D�H;��H;��H;�H;!�H;]�H;=�H;X�H;��H;r�H;_�H;r�H;��H;X�H;:�H;_�H;!�H;�H;��H;��H;D�H;��H;u�H;�H;��H;��H;��H;��H;��H;��H;��H;?�H;��H;I�H;��H;��H;S�H;��H;�H;��H;�H;��H;��H;�H;g�H;��H;      8�H;r�H;��H;l�H;k�H;��H;��H;m�H;�H;��H;e�H;(�H;��H;��H;$�H;��H;�H;f�H;��H;��H;��H;�H;>�H;��H;p�H;��H;6�H;��H;��H;��H;�H;?�H;H�H;x�H;j�H;`�H;q�H;`�H;j�H;u�H;F�H;A�H;�H;��H;��H;��H;6�H;��H;n�H;��H;>�H;�H;��H;��H;��H;g�H;�H;��H;!�H;��H;��H;'�H;e�H;��H;�H;j�H;��H;��H;`�H;l�H;��H;h�H;      ��H;�H;��H;P�H;\�H;��H;�H;��H;��H;��H;��H;��H;��H;��H;h�H;�H;��H;L�H;��H;��H;��H;��H;��H;}�H;�H;��H; �H;M�H;��H;��H;�H;�H;R�H;j�H;M�H;j�H;��H;j�H;M�H;j�H;O�H;!�H;�H;��H;��H;M�H;��H;��H;�H;{�H;��H;��H;��H;��H;��H;M�H;��H;�H;h�H;��H;��H;��H;��H;��H;��H;��H;�H;��H;R�H;P�H;��H;�H;      >�H;W�H;�H;��H;9�H;��H;��H;��H;��H;P�H;��H;5�H;��H;�H;f�H;��H;��H;;�H;��H;t�H;��H;��H;��H;��H;m�H;*�H;��H;�H;j�H;��H;��H;�H;)�H;=�H;i�H;t�H;T�H;t�H;i�H;=�H;(�H;�H;��H;��H;m�H;�H;��H;)�H;j�H;��H;��H;��H;��H;t�H;��H;;�H;��H;��H;e�H;�H;��H;3�H;��H;P�H;��H;��H;��H;��H;/�H;��H;�H;P�H;      V�H;��H;G�H;��H;:�H;Q�H;͸H;��H;��H;��H;��H;��H;��H;��H;��H;q�H;��H;<�H;i�H;I�H;��H;^�H;��H;��H;��H;h�H;�H;��H;�H;^�H;��H;��H;�H;/�H;T�H;J�H;=�H;J�H;U�H;/�H;�H;��H;��H;_�H;�H;��H;�H;e�H;��H;��H;��H;]�H;��H;J�H;g�H;<�H;��H;q�H;��H;��H;��H;��H;��H;��H;��H;��H;̸H;T�H;3�H;��H;F�H;��H;      ��H;�H;��H;��H;�H;��H;ܪH;x�H;R�H;`�H;��H;��H;��H;��H;X�H;��H;�H;-�H;��H;F�H;r�H;G�H;��H;S�H;��H;��H;B�H;�H;��H;�H;e�H;��H;��H;�H;�H;<�H;X�H;<�H;�H;�H;��H;��H;e�H;�H;��H;�H;A�H;��H;��H;Q�H;��H;F�H;m�H;D�H;��H;.�H;	�H;��H;X�H;��H;��H;��H;��H;_�H;T�H;w�H;ܪH;��H;ޤH;��H;��H;��H;      h�H;�H;t�H;��H;ЏH;��H;ݗH;ƜH;סH;-�H;��H;/�H;��H;�H;��H;�H;��H;~�H;�H;S�H;.�H;��H;��H;��H;��H;L�H;i�H;=�H;��H;��H;�H;h�H;��H;��H;�H; �H; �H;�H;�H;��H;��H;h�H;�H;��H;��H;;�H;g�H;J�H;��H;��H;��H;��H;*�H;Q�H;�H;�H;��H;�H;��H;�H;��H;/�H;��H;,�H;סH;ƜH;ݗH;��H;͏H;��H;u�H;�H;      iH;�iH;�kH;�nH;�rH;�wH;�}H;��H;��H; �H;q�H;ˡH;�H;ݯH;m�H;��H;b�H;h�H;�H;%�H;��H; �H;��H;�H;��H;��H;'�H;9�H;(�H;�H;��H;�H;X�H;��H;��H;��H;��H;��H;��H;��H;X�H;�H;��H;�H;(�H;:�H;&�H;��H;��H;�H;��H; �H;��H;"�H;�H;j�H;`�H;��H;m�H;ۯH;�H;ˡH;p�H;��H;��H;��H;�}H;�wH;�rH;�nH;�kH;�iH;      ?H;�?H;`BH;�FH;PLH;KSH;�[H;ndH;�mH;�wH;�H;�H;ѕH;�H;��H;ׯH;^�H;%�H;L�H;��H;=�H;\�H;�H;�H;��H;��H;y�H;�H;X�H;)�H;��H;��H;�H;m�H;��H;��H;��H;��H;��H;m�H;�H;��H;��H;&�H;X�H;�H;|�H;��H;��H;�H;�H;\�H;7�H;��H;L�H;%�H;\�H;ٯH;��H;�H;ѕH;�H;�H;�wH;�mH;kdH;�[H;NSH;MLH;�FH;]BH;�?H;      � H;.H;�H;�H;�H;y!H;C-H;�9H;GH;yTH;bH;toH;�|H;	�H;��H;��H;X�H;'�H;'�H;F�H;y�H;��H;J�H;.�H;��H;O�H;��H;��H;�H;:�H;;�H;�H;��H;�H;M�H;��H;��H;��H;N�H;�H;��H;�H;;�H;7�H;�H;��H;��H;O�H;��H;.�H;I�H;��H;t�H;D�H;%�H;'�H;U�H;��H;��H;�H;�|H;toH;bH;yTH;GH;�9H;C-H;u!H;�H;�H;�H;9H;      �G;U�G;��G;�G;L�G;/�G;��G;��G;�H;%H;K8H;�JH;�[H;~lH;|H;��H;��H;;�H;��H;��H;ӾH;��H;u�H;d�H;��H;V�H;7�H;��H;}�H;*�H;j�H;D�H;�H;��H;�H;;�H;I�H;9�H;�H;��H;�H;E�H;k�H;(�H;|�H;��H;6�H;T�H;��H;b�H;t�H;��H;ξH;��H;��H;=�H;��H;��H;|H;~lH;�[H;�JH;K8H;%H;�H;��G;��G;.�G;N�G;�G;��G;J�G;      �wF;�F;ĖF;�F;/�F;�G;�NG;C�G;x�G;�G;��G;rH;�1H;HH;�\H;�oH;؀H;Q�H;НH;��H;�H;ԼH;|�H;��H;�H;��H;Q�H;N�H;��H;��H;J�H;��H;g�H;,�H;��H;��H;��H;��H;��H;,�H;e�H;��H;L�H;��H;��H;O�H;Q�H;��H;�H;��H;}�H;ӼH;�H;��H;НH;S�H;րH;�oH;�\H;HH;�1H;sH;��G;
�G;y�G;@�G;�NG;�G;3�F;�F;ƖF;�F;      ��C;b	D;xBD;!�D;
E;҄E;}F;�wF;�F;!=G;(�G;	�G;��G;+H;�4H;�MH;>dH;JxH;��H;��H;æH;�H;��H;��H;`�H;�H;��H;��H;��H;��H;��H;��H;��H;r�H;�H;v�H;~�H;w�H;�H;q�H;��H;��H;��H;��H;��H;��H;��H;�H;`�H;��H;��H;�H;��H;��H;��H;MxH;<dH;�MH;�4H;+H;��G;	�G;'�G;=G;�F;�wF;}F;҄E;
E;!�D;xBD;b	D;      `,>;qZ>;�>;��?;h�@;�A;�C;D;�E;��E;�F;G;~G;y�G;�G;�!H;|@H;�ZH;jqH;_�H;n�H;äH;�H;3�H;��H;��H;a�H;+�H;	�H;�H;~�H;O�H;��H;��H;y�H;��H;�H;��H;}�H;��H;��H;P�H;�H;�H;�H;+�H;`�H;��H;��H;2�H;�H;äH;j�H;_�H;jqH;�ZH;y@H;�!H;�G;y�G;~G;G;�F;��E;�E;D;�C;�A;x�@;��?;�>;cZ>;      Y�1;�J2;�g3;�$5;�Y7;�9;�g<;N�>;A;�C;=�D;=�E;z�F;J*G;c�G;i�G;�H;�5H;-SH;�lH;K�H;ʔH;A�H;�H;��H;��H;x�H;I�H;�H;��H;��H;��H;��H;��H;��H;A�H;��H;A�H;��H;��H;��H;��H;��H;��H;�H;I�H;t�H;��H;��H;�H;?�H;ʔH;F�H;�lH;-SH;�5H;�H;g�G;c�G;I*G;z�F;=�E;<�D;�C;A;L�>;�g<;
�9;�Y7;�$5;�g3;nJ2;      �;��;(;�z ;��$;q�);�/;:4;$�8;d�<;'$@;z�B;P�D;��E;C�F;�cG;��G;�H;�-H;�NH;jH;\�H;ʔH;ƤH;�H;ּH;��H;��H;`�H;�H;��H;F�H;^�H;��H;��H;��H;��H;��H;��H;��H;^�H;D�H;��H;��H;\�H;��H;��H;׼H;�H;äH;ǔH;^�H;jH;�NH;�-H;�H;��G;�cG;D�F;��E;P�D;{�B;$$@;d�<;&�8;94;�/;p�);��$;�z ;(;��;      ��:4��:E��:���:�;�Y;�';��;��(;��0;�Y7;f�<;(�@;aC;BCE;�wF;�8G;��G;|�G;�)H;�LH;jH;J�H;q�H;��H;�H;ѾH;x�H;:�H;��H;*�H;j�H;��H;��H;��H;��H;��H;��H;��H;��H;��H;j�H;)�H;��H;7�H;y�H;ϾH;�H;��H;m�H;H�H;jH;�LH;�)H;|�G;��G;�8G;�wF;BCE;aC;%�@;f�<;�Y7;��0;��(;��;�';�Y;�;���:E��:��:      �:С:�3<:*i:�t�:��:��:�+�:�Y;V�;�*';�1;N�8;�Z>;g0B;)�D;�2F;:G;��G;2�G;�)H;�NH;�lH;a�H;}�H;��H;��H;C�H;��H; �H;M�H;=�H;H�H;n�H;��H;��H;��H;��H;��H;n�H;E�H;?�H;L�H;�H;��H;D�H;��H;��H;}�H;\�H;�lH;�NH;�)H;2�G;��G;<G;�2F;)�D;f0B;�Z>;N�8;�1;�*';V�;�Y;�+�:��:!��:�t�:*i:�3<:��:      ڥ���W��� ��8�=��ڷ�`�8�:�P�:�P�:���:D`;�;B�*;
%5;�g<;=A;CD;"F;�G;��G;}�G;�-H;/SH;mqH;��H;ԝH;��H;)�H;O�H;�H;�H;��H;i�H;��H;��H;��H;��H;��H;��H;��H;f�H;��H;�H;�H;J�H;)�H;��H;՝H;��H;iqH;,SH;�-H;z�G;��G;�G;$F;CD;=A;�g<;
%5;@�*;�;B`;���:�P�:�P�: �: �8Xڷ�8�=�� ���W��      �1��&Ȅ�¨u��PV�r.����vW������X�9l+i:
��:9,�:6�;�t%;�J2;s;;ɵ@;�D;"F;?G;��G;�H;�5H;�ZH;IxH;S�H;>�H;+�H;(�H;o�H;��H;.�H;C�H;=�H;Q�H;m�H;��H;m�H;P�H;=�H;A�H;.�H;��H;m�H;%�H;+�H;;�H;V�H;IxH;�ZH;�5H;�H;��G;@G;"F;�D;Ƶ@;s;;�J2;�t%;6�;7,�:
��:t+i: Y�9 ��vW�����k.��PV�¨u�*Ȅ�      X��H�	������Tʻ�R���2|�W.��Ⱥ����Y�9`u�:��:�Y;��!;��0;�:;ɵ@; CD;�2F;�8G;��G;�H;@H;:dH;؀H;��H;Z�H;]�H;b�H;��H;�H;��H;��H;��H;�H;��H;�H;��H;��H;��H;�H;��H;]�H;Z�H;Z�H;��H;ڀH;;dH;|@H;�H;��G;�8G;�2F; CD;˵@;�:;��0;��!;�Y;��:^u�:�Y�9����ȺY.��2|��R��Tʻ�����J�	�      ��x��[t���g�PT�^�:�������&����1��>�(�W��@�t�`o`:���:];&{ ;��0;v;;=A;/�D;�wF;�cG;j�G;�!H;�MH;�oH;��H;��H;ٯH;��H;z�H;��H;m�H;��H;�H;��H;8�H;��H;�H;��H;j�H;��H;x�H;��H;ӯH;��H;��H;�oH;�MH;�!H;i�G;�cG;�wF;/�D;=A;w;;��0;%{ ;];���:`o`:��t�W��>�(��1��&���������]�:�PT���g��[t�      9,˼��Ǽ�"���뮼w��&G��,�[�`y-�����.����b�H0��׷�r5<:)M�:];��!;�J2;�g<;j0B;CCE;A�F;e�G;�G;�4H;�\H;|H;��H;��H;m�H;��H;T�H;��H;e�H;e�H; �H;��H;�H;d�H;b�H;��H;U�H;��H;k�H;��H;��H;|H;�\H;�4H;�G;`�G;A�F;CCE;k0B;�g<;�J2;��!;];#M�:r5<:�׷�J0㺺�b��.�����ay-�+�[�&G��w���뮼�"����Ǽ      -���k��Kv��t�D�Ѽ�뮼-X��m�W������׻�Ǆ���X��~5<:���:�Y;�t%;%5;�Z>;aC;��E;M*G;z�G;*H;HH;�lH;�H;�H;֯H;�H;��H;��H;�H;��H;��H;@�H;��H;��H;�H;��H;��H;�H;֯H;�H;�H;~lH;HH;+H;y�G;G*G;��E;aC;�Z>;%5;�t%;�Y;���:v5<:X�����Ǆ���׻���m�W�-X���뮼D�Ѽ�t�Kv���k�      Gm��Fi��&^�b�L�R�6�)����!}ռoT����x���0�����������׷�do`:��:8�;C�*;P�8;(�@;Q�D;�F;	~G;��G;�1H;�[H;�|H;ѕH;�H;��H;��H;��H;��H;��H;��H;��H;��H;��H;��H;��H;��H;��H;�H;ΕH;�|H;�[H;�1H;��G;~G;z�F;Q�D;)�@;R�8;C�*;:�;��:do`:�׷���������껿�0���x�oT��!}ռ��)��R�6�b�L��&^��Fi�      O��u;��C�������섽{�e��?��k�}t�鷼G���e7�����Ǆ�F0� �t�`u�:;,�:�;�1;j�<;{�B;>�E;G;�G;tH;�JH;qoH;�H;��H;'�H;��H;��H;2�H;��H;�H;��H;�H;��H;.�H;��H;��H;'�H;��H;�H;ooH;�JH;vH;	�G;G;<�E;{�B;l�<;�1;�;?,�:^u�:��t�F0��Ǆ���껃e7�G��鷼}t��k��?�{�e��섽���C���u;��      t���'��s��ӽ�'��B�������Z��Q+�����"��G����0���׻��b�W���Y�9��:F`;�*';Z7;&$@;@�D;�F;(�G;��G;L8H;bH;�H;j�H;��H;��H;��H;��H;��H;^�H;J�H;^�H;��H;��H;��H;��H;��H;j�H;�H;bH;K8H;��G;,�G;�F;=�D;&$@;Z7;�*';B`;��:�Y�9W����b���׻��0�G���"������Q+��Z����A����'���ӽ�s�(��      �!,�;)��K ��������޽ ������Fi��0����鷼��x�����.��>�(�|��p+i:���:X�;��0;e�<;�C;��E;"=G;�G;%H;wTH;�wH;��H;)�H;]�H;��H;P�H;��H;��H;��H;��H;��H;P�H;��H;]�H;)�H;��H;�wH;wTH;%H;�G;%=G;��E;�C;e�<;��0;W�;���:x+i:���?�(��.�������x�鷼����0��Fi���� ���޽�������K �;)�      ,�j��f��Z�|�F��>/��^�q����ŽH ���Fi��Q+�}t�oT��n�W�����1���Ⱥ�X�9�P�:�Y;��(;"�8;A;�E;�F;�G;�H;GH;�mH;��H;ҡH;O�H;�H;��H;��H;�H;�H;�H;��H;��H;|�H;O�H;ҡH;��H;�mH;GH;�H;��G;�F;�E;A;"�8;��(;�Y;�P�: Y�9�Ⱥ�1�����n�W�oT��}t�Q+��Fi�H ���Žq����^��>/�|�F��Z��f�      ��x���z�J����f��SC��K �qn���Ž����Z��k�!}ռ-X��_y-�$���U.�����P�:�+�:��;64;O�>;D;�wF;I�G;��G;�9H;kdH;��H;��H;r�H;��H;��H;��H;d�H;��H;f�H;��H;��H;}�H;r�H;��H;��H;hdH;�9H;��G;G�G;�wF;D;O�>;64;��;�+�:�P�:���X.�%���_y-�-X��!}ռ�k��Z�����Žqn���K ��SC��f�J���z�x���      ��˾��Ǿ����!���X͓�^�x���J��K �q��� ������?����뮼+�[�����2|�nW����:��:�';�/;~g<;�C;~F;�NG;��G;@-H;�[H;�}H;ٗH;تH;θH;��H;�H;��H;�H;��H;�H;��H;̸H;تH;חH;�}H;[H;@-H;��G;�NG;�F;�C;|g<;�/;�';��:��:jW�� 3|����+�[��뮼���?���� ��q����K ���J�^�x�X͓�!���������Ǿ      u� ��������{Ծm���x���^�x��SC��^��޽A���{�e�)��E�Ѽ&G������R����� �8#��:�Y;i�);�9;�A;τE;�G;2�G;y!H;SSH;�wH;��H;��H;T�H;��H;��H;��H;��H;��H;��H;��H;Q�H;��H;��H;�wH;OSH;z!H;1�G;�G;҄E;�A;�9;i�);�Y;'��: �8����R�����&G��E�Ѽ)��{�e�A����޽�^��SC�^�x�x���m����{Ծ�쾣���      ��� E�l�u� �X�ݾm���X͓��f��>/�����'���섽Q�6��t�w��]�:�Tʻk.�`ڷ��t�:�;��$;�Y7;n�@;
E;2�F;M�G;�H;PLH;�rH;ƏH;ޤH;5�H;3�H;D�H;\�H;��H;\�H;C�H;3�H;3�H;ޤH;ƏH;�rH;MLH;�H;N�G;0�F;
E;k�@;�Y7;��$;�;�t�:`ڷ�i.�Tʻ]�:�w���t�Q�6��섽�'������>/��f�X͓�m���X�ݾu� �l� E�      ��7�v3�1�'����u� ��{Ծ!���J���|�F�����ӽ���a�L�Kv��뮼PT�ߘ껾PV�<�=�$*i:���:�z ;�$5;��?;�D;�F;
�G;�H;�FH;�nH;��H;��H;��H;��H;J�H;i�H;�H;i�H;J�H;��H;��H;��H;��H;�nH;�FH;�H;
�G;�F; �D;��?;�$5;�z ;���: *i:<�=��PV����PT��뮼Kv�a�L�����ӽ���|�F�J���!����{Ծu� ����1�'�v3�      �N��TI���;�1�'�l��쾂���z󐾶Z��K ��s�C����&^���"����g����Ĩu�� ���3<:5��:;}g3;	�>;�BD;ɖF;��G;�H;]BH;�kH;j�H;��H;?�H;�H;��H;��H;[�H;��H;��H;�H;=�H;��H;j�H;�kH;ZBH;�H;��G;ʖF;�BD;�>;�g3;;7��:�3<:� ��Ĩu������g��"����&^�C����s潧K ��Z�z󐾂�����l�1�'���;��TI�      c]�f�W��TI�v3� E�������Ǿx����f�:)�'��t;���Fi��k���Ǽ�[t�J�	�$Ȅ��W����:$��:��;qJ2;fZ>;[	D;�F;W�G;-H;�?H;�iH;��H;��H;��H;O�H;��H;l�H;��H;l�H;��H;O�H;��H;��H;��H;�iH;�?H;-H;U�G;�F;[	D;cZ>;vJ2;��; ��:��:�W��#Ȅ�J�	��[t���Ǽ�k��Fi�t;��(��:)��f�x�����Ǿ���� E�v3��TI�f�W�      �?��~h��?v��� ��9�X��O/�1y�C�;Ⱆ��+X����ѽ����an;�\�������B(�К���� �e9>�:;�Y.;h�<;�WC;7[F;�G;;0H;�jH;d�H;��H;ǵH;_�H;��H;��H;��H;��H;��H;��H;��H;]�H;ɵH;��H;b�H;~jH;;0H;�G;9[F;�WC;g�<;�Y.;;B�: �e9��Κ���B(�����\��an;������ѽ���+X�Ⱆ�C�;1y��O/�9�X�� ��?v��~h��      ~h��1���c�����y�YvS�rM+��v�9ɾ�����T�!]�\ν����y\8�����x���%�B���:��8�9�-�:��;��.;2�<;oC;�dF;�G;�1H;0kH;֌H;�H;�H;��H;�H;��H;�H;��H;�H;��H;�H;��H;�H;�H;ӌH;,kH;�1H;�G;�dF;oC;-�<;��.;��;�-�:0�98��B����%��x�����z\8�����\ν!]��T�����9ɾ�v�rM+�YvS���y�c���1���      ?v��c���X ��c�h�9E�Y��l���}㼾~���nH�Ո�{�ý�Ȅ��s/��o��#�����J���к@�9~g�:m;l0;7]=;�C;1�F;��G;W6H;lmH;V�H;ߥH;ŶH;6�H;}�H;�H;?�H;�H;?�H;	�H;}�H;3�H;ŶH;ߥH;R�H;imH;W6H;��G;2�F;�C;5]=;o0;m;|g�:(�9�кJ������#���o��s/��Ȅ�{�ýՈ��nH�~��}㼾l���Y��9E�c�h�X ��c���      � ����y�c�h��N��O/����D�߾B���*|��6�r}�䳽kSt�>�!�prμ=F{��_��X������4 :W��:[;�2;�O>;�D;~�F;��G;S=H;�pH;��H;��H;�H;�H;�H;��H;��H;��H;��H;��H;�H;�H;�H;��H;��H;�pH;S=H;��G;}�F;�D;�O>;�2;[;W��:0 :�����X���_�=F{�prμ>�!�kSt�䳽r}��6��*|�B��D�߾����O/��N�c�h���y�      9�X�YvS�9E��O/��S�KW����������NS\��� ���<����Y�{��Ѓ����]�v����b��Y�0�Y:��:�`;z�4;
�?;u�D;�F;0�G;>FH;�uH;�H;ʩH;ĹH;M�H;�H;]�H;S�H;3�H;S�H;\�H;�H;L�H;ǹH;ʩH;�H;�uH;>FH;1�G;�F;t�D;�?;~�4;�`;��:$�Y:�Y�
�b�w�����]�Ѓ��{���Y�<����当� �NS\���������KW���S��O/�9E�YvS�      �O/�rM+�Y�����KW��9ɾB���Mw�� :�k��y�ý�L��^n;�_���sv���E<��˻��-����y�:�^;�%;��7;��@;P5E;�"G;1�G;tPH;D{H;�H;��H;��H;��H;2�H;I�H;�H;��H;�H;I�H;2�H;��H;��H;��H;�H;@{H;sPH;0�G;�"G;O5E;��@;��7;�%;�^;�y�:����-��˻�E<�sv��_���^n;��L��y�ýk��� :��Mw�B��9ɾKW�����Y��rM+�      1y��v�l���D�߾����B��@����nH���E὞u����d�0O�jrμH"��������l�뺐t89�;�:�;�+;�|:;�7B;&�E;GbG;�H;)[H;��H;Z�H;֯H;2�H;��H;�H;B�H;�H;��H;�H;B�H;��H;��H;3�H;֯H;X�H;��H;)[H;�H;IbG;#�E;�7B;�|:;�+;��;�;�:�t89f��������I"��jrμ0O���d��u��E����nH�@���B������D�߾l����v�      C�;9ɾ}㼾B�������Mw��nH�����Z�䳽˕��r\8�p#������^N�B���b��Hx��5:P��:P�;�0;\]=;i�C;�[F; �G;*H;fH;��H;T�H;y�H;��H;R�H;�H;h�H;�H;��H;�H;h�H;�H;R�H;��H;{�H;T�H;��H;fH;*H; �G;�[F;f�C;\]=;�0;R�;N��:�5:�Hx��b�A��^N�����p#��r\8�˕��䳽�Z񽲯��nH��Mw�����B��}㼾9ɾ      Ⱆ�����~���*|�NS\�� :����Z�m$�������K�v���Oļ����������&�����/�:�^;��#;�G6;v�?;#�D;��F;��G;2@H;�pH;�H;��H;L�H;��H;d�H;��H;��H;�H;��H;�H;��H;��H;e�H;��H;L�H;��H;�H;�pH;0@H;��G;��F;"�D;u�?;�G6;��#;�^;�/�:���&������������Oļv���K�����m$���Z���� :�NS\��*|�~������      �+X��T��nH��6��� �k��E�䳽�����mR����ټ�����E<��?ݻd\�~���|!:e�:��;P�,;��:;�7B;ǲE;�LG;sH;�SH;�{H;��H;�H;N�H;w�H;��H;F�H; �H;)�H;��H;+�H; �H;H�H;��H;{�H;O�H;�H;��H;�{H;�SH;sH;�LG;ĲE;�7B;��:;P�,;��;e�:�!:����d\��?ݻ�E<�����ټ����mR�����䳽E�k���� ��6��nH��T�      ��!]�Ո�r}���y�ý�u��˕���K�����o�iv���&R���H^��<�� �=�D��:�B;s";��4;��>;}D;��F;1�G;*H;�dH;��H;L�H;��H;d�H;f�H;��H;�H;Z�H;E�H;�H;E�H;Z�H;�H;��H;i�H;e�H;��H;I�H;��H;�dH;*H;.�G;��F;zD;��>;��4;r";�B;H��: �=�<��H^�����&R�iv���o�����K�˕���u��y�ý��r}�Ո�!]�      �ѽ\ν{�ý䳽<����L����d�r\8�v��ټhv����Y��_�������,[�@�Y:���:xm;�r-;7�:;��A;koE;�"G;��G;�GH;�sH; �H;ŦH;!�H;c�H;P�H;��H;��H;��H;`�H;$�H;`�H;��H;��H;��H;S�H;d�H;�H;ĦH; �H;�sH;�GH;��G;�"G;ioE;��A;7�:;�r-;ym;���:<�Y:([��������_���Y�hv��ټv��r\8���d��L��<���䳽{�ý\ν      ���������Ȅ�kSt��Y�^n;�0O�p#���Oļ�����&R��_������N3�P�Y�|4:Z�:��;@&;
H6;�X?;�D;exF;�G;m!H;�^H;��H;(�H;�H;w�H;=�H;3�H;�H;G�H;�H;��H;G�H;��H;�H;I�H;�H;4�H;>�H;y�H;�H;(�H;��H;�^H;k!H;�G;axF;�D;�X?;	H6;@&;��;Z�:�4:P�Y��N3������_��&R������Oļp#��0O�^n;��Y�kSt��Ȅ�����      an;�y\8��s/�>�!�{��^���irμ��������E<��������N3��Gx���9<�:_;z ;X2;��<;"�B;߲E;i5G;<�G;jFH;�qH;َH;��H;�H;��H;��H;��H;4�H;��H;Q�H;��H;A�H;��H;Q�H;��H;4�H;��H;��H;��H;�H;��H;؎H;�qH;jFH;9�G;e5G;߲E;"�B;��<;X2;| ;_;>�:��9�Gx��N3��������E<��������irμ^���{��>�!��s/�y\8�      \������o�prμу��sv��I"��^N�����?ݻH^��#��X�Y���94�:$��:�;w�.;�|:;$?A;��D;_�F;�G;*H;SaH;M�H;��H;�H;o�H;R�H;p�H;��H;/�H;P�H;��H;��H;�H;��H;��H;Q�H;/�H;��H;p�H;Q�H;m�H;�H;��H;O�H;QaH;*H;�G;_�F;��D;&?A;�|:;z�.;�;$��:4�:��9X�Y�#��H^���?ݻ���^N�I"��sv��у��prμ�o����      �����x���#��=F{���]��E<����C�뻜���d\�>��,[�x4:8�:*��:�[;��,;�8;K!@;1D;�[F;V{G;*H;zPH;NvH;�H;v�H;2�H;c�H;��H;��H;�H;�H;��H;��H;��H;��H;��H;��H;��H;�H;�H;��H;��H;_�H;2�H;t�H; �H;MvH;vPH;&H;T{G;�[F;1D;K!@;�8;��,;�[;*��:<�:x4:,[�>��d\�����C�뻞���E<���]�=F{��#���x��      �B(��%�����_�x����˻����b�&����� �=�<�Y:T�:_;�;��,;:`8;��?;��C;�F;!GG;}�G;'@H;^kH;7�H;:�H;(�H;��H;��H;��H;��H;P�H;��H;�H;��H;��H;��H;��H;��H;�H;��H;Q�H;��H;��H;��H;��H;&�H;?�H;7�H;ZkH;"@H;�G; GG;�F;��C;��?;;`8;��,;�;_;T�:<�Y: �=�����&��b�����˻x����_�����%�      Қ��E���J���X���b���-�p�뺘Hx����|!:D��:���:��;v ;x�.;�8;��?;'�C;�E;l#G;�G;2H;#bH;~�H;��H;��H;�H;�H;��H;N�H;m�H;n�H;"�H;M�H;��H;p�H;��H;p�H;��H;M�H;!�H;o�H;m�H;M�H;��H;�H;޷H;��H;��H;|�H; bH;2H;�G;n#G;�E;)�C;��?;�8;x�.;x ;��;���:D��:t!:����Hx�n����-�
�b��X��J��H���      ��<���к����,�Y�����t89�5:�/�:e�:�B;vm;@&;X2;�|:;J!@;�C;�E;�G;�G;�(H;1[H;�zH;r�H;�H;ֳH;��H;��H;��H;��H;��H;1�H;��H;e�H;��H;3�H;��H;4�H;��H;e�H;��H;2�H;��H;��H;��H;��H;��H;ٳH;�H;q�H;�zH;1[H;�(H;�G;�G;�E;�C;J!@;�|:;Z2;@&;xm;�B;e�:�/�:�5:�t89����Y������к<��       �e9��9H�9$ :$�Y:�y�:�;�:B��:�^;��;o";�r-;H6;��<;"?A;�0D;�F;g#G;
�G;%H;�WH;�vH;��H;w�H;}�H;��H;F�H;��H;��H;p�H;�H;��H;��H;b�H;E�H;��H;1�H;��H;E�H;b�H;��H;��H;�H;n�H;��H;��H;D�H;��H;}�H;t�H;��H;�vH;�WH;%H;
�G;j#G;�F; 1D;"?A;��<;H6;�r-;o";��;�^;H��:�;�:�y�:P�Y:( :@�9X�9      L�:�-�:�g�:C��:��:�^;�;L�;��#;P�,;��4;2�:;�X?;�B;��D;�[F; GG;�G;�(H;�WH;�uH;ÌH;K�H;2�H;[�H;1�H;��H;%�H;�H;��H;��H;�H;��H;(�H;�H;��H;��H;��H;�H;(�H;��H;�H;��H;��H;�H;%�H;��H;1�H;Y�H;.�H;L�H;ŌH;�uH;�WH;�(H;�G; GG;�[F;��D;�B;�X?;2�:;��4;N�,;��#;L�;�;�^;��:I��:�g�:�-�:      ;��;m;
[;�`;�%;�+;�0;�G6;��:;��>;��A;�D;ݲE;_�F;Q{G;}�G;2H;0[H;�vH;H;��H;��H;�H;��H;��H;��H;��H;��H;!�H;x�H;q�H;��H;��H;��H;��H;�H;��H;��H;��H;��H;q�H;v�H;�H;��H;��H;��H;��H;��H;�H;��H;��H;H;�vH;0[H;2H;|�G;Q{G;`�F;߲E;�D;��A;��>;��:;�G6;�0;�+;�%;�`;[;m;��;      �Y.;��.;l0;�2;t�4;��7;�|:;Y]=;u�?;�7B;xD;joE;axF;g5G;�G;&H;&@H;"bH;�zH;��H;K�H;��H;��H;�H;��H;��H;�H;1�H;X�H;��H;��H;��H;��H;��H;'�H;Z�H;��H;Z�H;'�H;��H;��H;��H;��H;��H;V�H;1�H; �H;��H;��H;�H;��H;��H;G�H;��H;�zH;#bH;$@H;$H;�G;g5G;axF;joE;zD;�7B;v�?;[]=;�|:;��7;z�4;�2;l0;��.;      y�<;@�<;>]=;�O>;
�?;��@;�7B;e�C;"�D;ŲE;��F;�"G;�G;9�G;*H;vPH;[kH;��H;p�H;v�H;.�H;�H;�H;q�H;n�H;r�H;��H;��H;[�H;v�H;6�H;I�H;F�H;�H;}�H;��H;��H;��H;~�H;�H;C�H;K�H;6�H;s�H;Y�H;��H;��H;r�H;n�H;m�H;�H;�H;+�H;w�H;q�H;��H;ZkH;wPH;*H;:�G;�G;�"G;��F;ĲE;"�D;f�C;�7B;��@;�?;�O>;>]=;0�<;      �WC;oC;��C;�D;u�D;P5E;!�E;�[F;��F;�LG;-�G;��G;i!H;kFH;SaH;NvH;<�H;��H;�H;��H;]�H;��H;��H;t�H;0�H;B�H;{�H;�H;#�H;��H;�H;��H;��H;q�H;��H;�H;�H;�H;��H;p�H;��H; �H;�H;��H;"�H;�H;{�H;B�H;3�H;r�H;��H;��H;\�H;��H;�H;��H;:�H;NvH;SaH;jFH;i!H;��G;-�G;�LG;��F;�[F;!�E;P5E;x�D;�D;��C;oC;      @[F;�dF;$�F;x�F;�F;�"G;CbG;�G;��G;nH;	*H;�GH;�^H;�qH;J�H;�H;:�H;��H;ӳH;��H;.�H;��H;��H;p�H;;�H;e�H;��H;��H;��H;��H;��H;��H;a�H;��H;�H;O�H;O�H;O�H;�H;��H;^�H;��H;��H;��H;��H;��H;��H;e�H;>�H;p�H;��H;��H;*�H;��H;ӳH;��H;9�H;�H;J�H;�qH;�^H;�GH;
*H;oH;��G;�G;CbG;�"G; �F;x�F;"�F;�dF;      "�G;�G;��G;��G;4�G;1�G;�H;*H;0@H;�SH;�dH;�sH;��H;֎H;��H;v�H;)�H;޷H;��H;H�H;��H;��H; �H;��H;u�H;��H;��H;}�H;��H;��H;��H;4�H;��H;�H;A�H;r�H;��H;r�H;@�H;�H;��H;2�H;��H;��H;��H;{�H;��H;��H;x�H;��H;��H;��H;��H;G�H;��H;�H;(�H;t�H;��H;؎H;��H;�sH;�dH;�SH;1@H;*H;�H;.�G;:�G;��G;��G;�G;      .0H;�1H;]6H;I=H;@FH;qPH;)[H;"fH;�pH;�{H;��H;$�H;(�H;��H;�H;2�H;��H;�H;��H;��H;$�H;��H;/�H;��H;��H;��H;z�H;��H;��H;��H;;�H;��H;��H;J�H;~�H;��H;��H;��H;~�H;J�H;��H;��H;;�H;��H;��H;��H;z�H;��H;��H;��H;.�H;��H;!�H;��H;��H;�H;��H;2�H;�H;��H;%�H;$�H;��H;�{H;�pH;#fH;)[H;sPH;KFH;J=H;[6H;�1H;      �jH;/kH;hmH;�pH;�uH;?{H;��H;��H;�H;��H;K�H;ȦH;�H;�H;n�H;b�H;��H;��H;��H;��H;�H;��H;T�H;]�H;�H;��H;��H;��H;��H;(�H;��H;��H;0�H;m�H;��H;��H;��H;��H;��H;m�H;.�H;��H;��H;'�H;��H;��H;��H;��H;�H;]�H;S�H;��H;�H;��H;��H;��H;��H;c�H;o�H;�H;�H;ǦH;I�H;��H;�H;��H;��H;?{H;�uH;�pH;hmH;#kH;      o�H;ڌH;\�H;��H;��H;�H;]�H;W�H;��H; �H;��H;*�H;}�H;��H;T�H;��H;��H;H�H;��H;r�H;��H;�H;��H;v�H;��H;��H;��H;��H;'�H;��H;��H;6�H;m�H;��H;��H;��H;��H;��H;��H;��H;j�H;7�H;��H;��H;&�H;��H;��H;��H;��H;u�H;��H;�H;��H;r�H;��H;J�H;��H;��H;U�H;��H;}�H;)�H;��H;"�H;��H;Z�H;]�H;�H;��H;��H;X�H;֌H;      ��H;�H;�H;��H;թH;��H;ۯH;��H;P�H;O�H;j�H;m�H;A�H;��H;q�H;��H;��H;k�H;��H;�H;��H;u�H;��H;7�H;�H;��H;��H;=�H;��H;��H;2�H;c�H;��H;��H;��H;��H;��H;��H;��H;��H;��H;d�H;2�H;��H;��H;=�H;��H;��H;�H;7�H;��H;u�H;��H;�H;��H;k�H;��H;��H;q�H;��H;A�H;k�H;j�H;S�H;S�H;��H;ۯH;��H;ҩH;��H;�H;�H;      յH;!�H;̶H;�H;ɹH;��H;2�H;��H;��H;x�H;m�H;Z�H;7�H;��H;��H;�H;W�H;n�H;4�H;��H;�H;t�H;��H;L�H;��H;��H;/�H;��H;��H;6�H;`�H;{�H;��H;��H;��H;��H;��H;��H;��H;��H;��H;~�H;b�H;:�H;��H;��H;2�H;��H;��H;L�H;��H;t�H;�H;��H;4�H;o�H;U�H;�H;��H;��H;7�H;X�H;m�H;z�H;��H;��H;3�H;��H;ǹH;�H;˶H;�H;      `�H;��H;;�H;�H;T�H;��H;~�H;X�H;h�H;��H;��H;��H;�H;:�H;2�H;�H;��H;�H;��H;��H;��H;��H;��H;I�H;��H;\�H;��H;��H;2�H;p�H;��H;��H;��H;��H;��H;��H;��H;��H;��H;��H;��H;��H;��H;t�H;5�H;��H;��H;^�H;��H;J�H;��H;��H;��H;��H;��H; �H;��H;�H;1�H;:�H;	�H;��H;��H;��H;k�H;X�H;~�H;��H;M�H;�H;:�H;��H;      ��H;�H;u�H;�H;	�H;)�H;��H;�H;��H;H�H;�H;��H;J�H;��H;S�H;��H;�H;L�H;e�H;f�H;*�H;��H;|�H;�H;h�H;��H;�H;J�H;k�H;��H;��H;��H;��H;��H;��H;��H;��H;��H;��H;��H;��H;��H;��H;��H;p�H;J�H;�H;��H;i�H;�H;}�H;��H;*�H;g�H;f�H;M�H;�H;��H;S�H;��H;J�H;��H;�H;I�H;��H;�H;��H;/�H; �H;�H;u�H;�H;      ��H;��H;�H;��H;t�H;B�H;I�H;s�H;��H;�H;a�H;��H;�H;X�H;��H;��H;��H;��H;��H;I�H;�H;��H;!�H;~�H;��H;�H;:�H;|�H;��H;��H;��H;��H;��H;��H;��H;��H;��H;��H;��H;��H;��H;��H;��H;��H;��H;~�H;:�H;	�H;��H;~�H;$�H;��H;�H;I�H;��H;��H;��H;��H;��H;X�H;�H;��H;_�H;�H;��H;q�H;H�H;G�H;j�H;��H;�H;��H;      ��H;�H;F�H;��H;_�H;�H;�H;�H;�H;)�H;N�H;i�H;��H;��H;��H;��H;��H;j�H;4�H;��H;��H;��H;U�H;��H;�H;K�H;n�H;��H;��H;��H;��H;��H;��H;��H;��H;��H;��H;��H;��H;��H;��H;��H;��H;��H;��H;��H;n�H;J�H;�H;��H;W�H;��H;��H;��H;6�H;k�H;��H;��H;��H;��H;��H;i�H;L�H;.�H;�H;�H;�H;�H;T�H;��H;F�H;�H;      ��H;��H;(�H;��H;A�H;��H;��H;��H;��H;��H;�H;.�H;K�H;H�H;�H;�H;��H;��H;��H;4�H;��H;�H;~�H;��H;�H;J�H;��H;��H;��H;��H;��H;��H;��H;��H;��H;��H;��H;��H;��H;��H;��H;��H;��H;��H;��H;��H;��H;K�H;�H;��H;~�H;�H;��H;4�H;��H;��H;��H;�H;�H;H�H;K�H;.�H;�H;��H;��H;��H;��H;��H;5�H;��H;(�H;��H;      ��H;�H;F�H;��H;_�H;�H;�H;�H;�H;)�H;N�H;i�H;��H;��H;��H;��H;��H;j�H;6�H;��H;��H;��H;W�H;��H;�H;K�H;p�H;��H;��H;��H;��H;��H;��H;��H;��H;��H;��H;��H;��H;��H;��H;��H;��H;��H;��H;��H;n�H;J�H;�H;��H;U�H;��H;��H;��H;4�H;k�H;��H;��H;��H;��H;��H;i�H;N�H;+�H;�H;�H;�H;�H;T�H;��H;B�H;�H;      ��H;��H;�H;��H;u�H;B�H;I�H;t�H;��H;�H;_�H;��H;�H;X�H;��H;��H;��H;��H;��H;I�H;
�H;��H;#�H;�H;��H;	�H;:�H;~�H;��H;��H;��H;��H;��H;��H;��H;��H;��H;��H;��H;��H;��H;��H;��H;��H;��H;|�H;:�H;�H;��H;{�H;#�H;��H;�H;I�H;��H;��H;��H;��H;��H;X�H;�H;��H;_�H;�H;��H;p�H;I�H;G�H;j�H;��H;�H;��H;      ��H;�H;u�H;�H;	�H;)�H;��H;�H;��H;I�H;�H;��H;J�H;��H;S�H;��H;�H;L�H;f�H;g�H;0�H;��H;}�H;�H;i�H;��H;�H;J�H;m�H;��H;��H;��H;��H;��H;��H;��H;��H;��H;��H;��H;��H;��H;��H;��H;n�H;J�H;�H;��H;h�H;�H;|�H;��H;*�H;f�H;e�H;M�H;�H;��H;T�H;��H;J�H;��H;�H;H�H;��H;�H;��H;.�H; �H;�H;u�H;�H;      c�H;��H;=�H;�H;Q�H;��H;~�H;X�H;i�H;��H;��H;��H;	�H;:�H;1�H;�H;��H;�H;��H;��H;�H;��H;��H;J�H;��H;_�H;��H;��H;3�H;r�H;��H;��H;��H;��H;��H;��H;��H;��H;��H;��H;��H;��H;��H;q�H;3�H;��H;��H;\�H;��H;H�H;��H;��H;��H;��H;��H;�H;��H;�H;2�H;:�H;	�H;��H;��H;��H;h�H;U�H;~�H;��H;L�H;�H;:�H;��H;      ׵H;!�H;ζH;�H;ǹH;��H;5�H;��H;��H;{�H;m�H;Z�H;7�H;��H;��H;�H;X�H;n�H;4�H;��H;�H;t�H;��H;N�H;��H;��H;1�H;��H;��H;9�H;b�H;|�H;��H;��H;��H;��H;��H;��H;��H;��H;��H;|�H;`�H;7�H;��H;��H;1�H;��H;��H;L�H;��H;t�H;�H;��H;4�H;o�H;U�H;�H;��H;��H;7�H;X�H;m�H;z�H;��H;��H;5�H;��H;ĹH;�H;ζH;�H;      ��H;�H;�H;��H;թH;��H;ۯH;��H;R�H;R�H;j�H;k�H;A�H;��H;r�H;��H;��H;j�H;��H;�H;��H;u�H;��H;9�H;�H;��H;��H;=�H;��H;��H;2�H;c�H;��H;��H;��H;��H;��H;��H;��H;��H;��H;d�H;2�H;��H;��H;=�H;��H;��H;�H;7�H;��H;u�H;��H;�H;��H;k�H;��H;��H;q�H;��H;A�H;m�H;h�H;P�H;P�H;��H;ۯH;��H;ѩH;��H;�H;�H;      h�H;ڌH;[�H;��H;��H;�H;^�H;Z�H;��H; �H;��H;*�H;|�H;��H;U�H;��H;��H;H�H;��H;s�H;��H;�H;��H;v�H;��H;��H;��H;��H;'�H;��H;��H;6�H;k�H;��H;��H;��H;��H;��H;��H;��H;k�H;7�H;��H;��H;'�H;��H;��H;��H;��H;u�H;��H;�H;��H;r�H;��H;J�H;��H;��H;T�H;��H;|�H;*�H;��H;�H;��H;X�H;^�H;�H;��H;��H;\�H;،H;      �jH;*kH;mmH;�pH;�uH;:{H;��H;��H;�H;��H;K�H;ȦH;�H;�H;o�H;c�H;��H;��H;��H;��H;�H;��H;T�H;]�H;�H;��H;��H;��H;��H;(�H;��H;��H;/�H;m�H;��H;��H;��H;��H;��H;m�H;/�H;��H;��H;'�H;��H;��H;��H;��H;�H;]�H;S�H;��H;�H;��H;��H;��H;��H;c�H;n�H;�H;�H;ȦH;K�H;��H;�H;��H;��H;<{H;�uH;�pH;lmH;*kH;      .0H;�1H;[6H;J=H;>FH;sPH;)[H;$fH;�pH;�{H;��H;$�H;%�H;��H;�H;2�H;��H;�H;��H;��H;'�H;��H;/�H;��H;��H;��H;z�H;��H;��H;��H;;�H;��H;��H;H�H;|�H;��H;��H;��H;~�H;J�H;��H;��H;;�H;��H;��H;��H;z�H;��H;��H;��H;.�H;��H;!�H;��H;��H;�H;��H;4�H;�H;��H;(�H;$�H;��H;�{H;�pH;"fH;)[H;oPH;HFH;I=H;[6H;�1H;      �G;�G;��G;��G;0�G;-�G;�H;*H;0@H;�SH;�dH;�sH;��H;؎H;��H;v�H;)�H;޷H;��H;J�H;��H;��H;��H;��H;x�H;��H;��H;{�H;��H;��H;��H;4�H;��H;�H;@�H;r�H;��H;q�H;A�H;�H;��H;5�H;��H;��H;��H;}�H;��H;��H;u�H;��H;��H;��H;��H;G�H;��H;�H;(�H;t�H;��H;֎H;��H;�sH;�dH;�SH;0@H;*H;�H;+�G;4�G;��G;��G;��G;      G[F;�dF;+�F;x�F;�F;�"G;EbG;�G;��G;pH;
*H;�GH;�^H;�qH;H�H;�H;:�H;��H;ӳH;��H;0�H;��H;��H;r�H;>�H;e�H;��H;��H;��H;��H;��H;��H;_�H;��H;�H;O�H;O�H;O�H;�H;��H;^�H;��H;��H;��H;��H;��H;��H;e�H;;�H;o�H;��H;��H;*�H;��H;ӳH;��H;9�H;�H;J�H;�qH;�^H;�GH;	*H;nH;��G;�G;FbG;�"G; �F;{�F;.�F;�dF;      �WC;oC;��C;�D;u�D;P5E;!�E;�[F;��F;�LG;.�G;��G;i!H;jFH;SaH;OvH;<�H;��H;�H;��H;_�H;��H;��H;u�H;3�H;B�H;{�H;�H;%�H;��H;�H;��H;��H;p�H;��H;�H;�H;�H;��H;p�H;��H;�H;�H;��H; �H;�H;{�H;B�H;0�H;r�H;��H;��H;\�H;��H;�H;��H;8�H;NvH;SaH;jFH;i!H;��G;-�G;�LG;��F;�[F;!�E;P5E;t�D;�D;��C;oC;      }�<;=�<;D]=;�O>;�?;��@;�7B;e�C;#�D;ǲE;��F;�"G;�G;:�G;*H;wPH;[kH;~�H;q�H;w�H;/�H;�H;�H;q�H;n�H;r�H;��H;��H;\�H;v�H;6�H;I�H;E�H;�H;{�H;��H;��H;��H;~�H;�H;E�H;K�H;6�H;s�H;X�H;��H;��H;r�H;n�H;o�H;�H;�H;+�H;v�H;p�H;��H;ZkH;vPH;*H;9�G;�G;�"G;��F;ĲE;#�D;e�C;�7B;��@;�?;�O>;G]=;/�<;      �Y.; �.;y0;�2;p�4;ā7;�|:;[]=;u�?;�7B;zD;joE;_xF;g5G;�G;&H;&@H; bH;�zH;��H;L�H;��H;��H;�H;��H;��H;�H;1�H;X�H;��H;��H;��H;��H;��H;'�H;Z�H;��H;Z�H;'�H;��H;��H;��H;��H;��H;V�H;1�H; �H;��H;��H;�H;��H;��H;G�H;��H;�zH;#bH;&@H;&H;�G;g5G;_xF;ioE;xD;�7B;v�?;X]=;�|:;Ł7;v�4;�2;p0;��.;      ;��;m;[;�`;�%;�+;�0;�G6;��:;��>;��A;�D;߲E;_�F;S{G;|�G;2H;0[H;�vH;ŌH;��H;��H;�H;��H;��H;��H;��H;��H;!�H;v�H;q�H;��H;��H;��H;��H;�H;��H;��H;��H;��H;q�H;x�H;�H;��H;��H;��H;��H;��H;�H;��H;��H;��H;�vH;0[H;2H;|�G;Q{G;`�F;ݲE;�D;��A;��>;��:;�G6;�0;�+;�%;�`;
[;m;��;      B�:�-�:�g�:I��:��:�^;��;N�;��#;N�,;��4;2�:;�X?;�B;��D;�[F;!GG;�G;�(H;�WH;�uH;ŌH;L�H;3�H;Y�H;1�H;��H;%�H;�H;��H;��H;�H;��H;&�H;�H;��H;��H;��H;�H;(�H;��H;�H;��H;��H;�H;%�H;��H;1�H;[�H;.�H;K�H;ÌH;�uH;�WH;�(H;�G;GG;�[F;��D;�B;�X?;2�:;��4;L�,;��#;N�;��;�^;��:I��:�g�:�-�:      �e9��9X�9$ :0�Y:�y�:�;�:F��:�^;��;o";�r-;H6;��<;"?A; 1D;�F;i#G;
�G;%H;�WH;�vH;��H;z�H;}�H;��H;G�H;��H;��H;p�H;�H;��H;��H;b�H;E�H;��H;1�H;��H;E�H;b�H;��H;��H;�H;n�H;��H;��H;D�H;��H;}�H;s�H;��H;�vH;�WH;%H;
�G;i#G;�F;�0D;"?A;��<;H6;�r-;m";��;�^;H��:�;�:�y�:@�Y: :H�9P�9      ��<���к����0�Y� ���t89�5:�/�:e�:�B;xm;@&;Z2;�|:;J!@;�C;�E;�G;�G;�(H;1[H;�zH;u�H;�H;׳H;��H;��H;��H;��H;��H;1�H;��H;e�H;��H;3�H;��H;3�H;��H;e�H;��H;2�H;��H;��H;��H;��H;��H;ٳH;�H;n�H;�zH;1[H;�(H;�G;�G;�E;�C;J!@;�|:;X2;@&;vm;�B;e�:�/�:�5:�t89����Y������к<��      К��E���J���X���b���-�r�뺠Hx����t!:D��:���:��;v ;x�.;�8;��?;'�C;�E;m#G;�G;2H;#bH;~�H;��H;��H;�H;�H;��H;N�H;m�H;n�H;$�H;M�H;��H;p�H;��H;p�H;��H;M�H;!�H;o�H;m�H;M�H;��H;�H;޷H;��H;��H;|�H; bH;2H;�G;l#G;�E;(�C;��?;�8;x�.;v ;��;���:F��:|!:����Hx�r����-��b��X��J��H���      �B(��%�����_�y����˻����b�&����� �=�<�Y:T�:_;�;��,;=`8;��?;��C;�F;!GG;�G;'@H;^kH;7�H;=�H;)�H;��H;��H;��H;��H;Q�H;��H;�H;��H;��H;��H;��H;��H;�H;��H;Q�H;��H;��H;��H;��H;#�H;=�H;7�H;ZkH;"@H;}�G; GG;�F;��C;��?;:`8;��,;�;_;T�:<�Y: �=�����&��b�����˻x����_�����%�      �����x���#��=F{���]��E<����C�뻜���d\�>��,[�x4:8�:*��:�[;��,;�8;K!@;1D;�[F;T{G;(H;zPH;MvH;�H;w�H;2�H;c�H;��H;��H;�H;�H;��H;��H;��H;��H;��H;��H;��H;�H;�H;��H;��H;_�H;2�H;s�H;�H;NvH;wPH;&H;V{G;�[F;1D;K!@;�8;��,;�[;*��:8�:x4:,[�>��d\�����D�뻞���E<���]�=F{��#���x��      \������o�prμу��sv��I"��^N�����?ݻH^��"��X�Y���94�:$��:�;w�.;�|:;%?A;��D;_�F;�G;*H;QaH;N�H;��H;�H;r�H;R�H;p�H;��H;1�H;Q�H;��H;��H;�H;��H;��H;Q�H;/�H;��H;p�H;Q�H;m�H;�H;��H;O�H;SaH;*H;�G;_�F;��D;%?A;�|:;z�.;	�;$��:4�:��9X�Y�#��H^���?ݻ���^N�I"��sv��у��prμ�o����      an;�y\8��s/�>�!�{��^���irμ��������E<��������N3��Gx���9>�:_;z ;X2;��<;"�B;߲E;i5G;<�G;jFH;�qH;َH;��H;�H;��H;��H;��H;6�H;��H;Q�H;��H;A�H;��H;Q�H;��H;3�H;��H;��H;��H;�H;��H;؎H;�qH;jFH;:�G;e5G;߲E;"�B;��<;X2;z ;_;<�:��9�Gx��N3��������E<��������irμ^���{��>�!��s/�y\8�      ���������Ȅ�kSt��Y�^n;�0O�p#���Oļ�����&R��_������N3�P�Y�|4:^�:��;@&;	H6;�X?;�D;exF;�G;k!H;�^H;��H;(�H;	�H;y�H;>�H;4�H;�H;I�H;�H;��H;G�H;��H;�H;G�H;�H;4�H;=�H;w�H;�H;(�H;��H;�^H;m!H;�G;axF;�D;�X?;	H6;@&;��;X�:|4:P�Y��N3������_��&R������Oļp#��0O�]n;��Y�kSt��Ȅ�����      �ѽ\ν{�ý䳽<����L����d�r\8�v��ټhv����Y��_�������([�@�Y:���:ym;�r-;5�:;��A;koE;�"G;��G;�GH;�sH; �H;ŦH;!�H;d�H;P�H;��H;��H;��H;a�H;$�H;a�H;��H;��H;��H;Q�H;c�H;�H;ĦH; �H;�sH;�GH;��G;�"G;ioE;��A;7�:;�r-;xm;���:<�Y:0[��������_���Y�hv��ټv��s\8���d��L��<���䳽{�ý\ν      ��!]�Ո�r}���y�ý�u��˕���K�����o�iv���&R���H^��<�� �=�F��:�B;s";��4;��>;}D;��F;.�G;*H;�dH;��H;L�H;��H;e�H;f�H;��H;�H;Z�H;E�H;�H;E�H;Z�H;�H;��H;h�H;d�H;��H;I�H;��H;�dH;*H;1�G;��F;zD;��>;��4;r";�B;F��: �=�>��H^�����&R�iv���o�����K�˕���u��y�ý��r}�Ո�!]�      �+X��T��nH��6��� �k��E�䳽�����mR����ټ�����E<��?ݻd\�����|!:e�:��;N�,;��:;�7B;ǲE;�LG;sH;�SH;�{H;H;�H;O�H;z�H;��H;H�H; �H;)�H;��H;+�H; �H;F�H;��H;w�H;N�H;�H;��H;�{H;�SH;sH;�LG;ĲE;�7B;��:;P�,;��;e�:�!:����d\��?ݻ�E<�����ټ����mR�����䳽E�k���� ��6��nH��T�      Ⱆ�����~���*|�NS\�� :����Z�m$�������K�v���Oļ����������&�����/�:�^;��#;�G6;v�?;#�D;��F;��G;2@H;�pH;�H;��H;L�H;��H;g�H;��H;��H;�H;��H;�H;��H;��H;b�H;��H;L�H;��H;�H;�pH;0@H;��G;��F;"�D;u�?;�G6;��#;�^;�/�:���&������������Oļv���K�����m$���Z���� :�NS\��*|�~������      C�;9ɾ}㼾B�������Mw��nH�����Z�䳽˕��r\8�p#������^N�B���b��Hx��5:N��:N�;�0;\]=;h�C;�[F; �G;*H;fH;��H;T�H;{�H;��H;T�H;�H;i�H;�H;��H;�H;h�H;�H;Q�H;��H;y�H;T�H;��H;fH;*H;�G;�[F;f�C;\]=;�0;R�;N��:�5:�Hx��b�B��^N�����p#��r\8�˕��䳽�Z񽲯��nH��Mw�����B��}㼾9ɾ      1y��v�l���D�߾����B��@����nH���E὞u����d�0O�jrμI"��������h�뺐t89�;�:�;�+;�|:;�7B;#�E;IbG;�H;)[H;��H;Z�H;֯H;2�H;��H;��H;B�H;�H;��H;�H;B�H;�H;~�H;2�H;֯H;X�H;��H;)[H;�H;IbG;&�E;�7B;�|:;�+;��;�;�:�t89h��������H"��jrμ0O���d��u��E����nH�@���B������D�߾l����v�      �O/�rM+�Y�����KW��9ɾB���Mw�� :�k��y�ý�L��^n;�_���sv���E<��˻��-����y�:�^;�%;��7;��@;O5E;�"G;2�G;sPH;D{H;�H;��H;��H;��H;2�H;I�H;�H;��H;�H;I�H;2�H;��H;��H;��H;�H;@{H;tPH;0�G;�"G;P5E;��@;��7;�%;�^;�y�:����-��˻�E<�sv��_���^n;��L��y�ýk��� :��Mw�B��9ɾKW�����Y��rM+�      9�X�YvS�9E��O/��S�KW����������NS\��� ���<����Y�{��Ѓ����]�v����b��Y�$�Y:��:�`;z�4;
�?;t�D;�F;0�G;>FH;�uH;�H;ʩH;ƹH;M�H;�H;]�H;S�H;3�H;S�H;[�H;�H;L�H;ǹH;ʩH;�H;�uH;>FH;1�G;�F;u�D;�?;~�4;�`;��:$�Y:�Y�
�b�x�����]�Ѓ��{���Y�<����当� �NS\���������KW���S��O/�9E�YvS�      � ����y�c�h��N��O/����D�߾B���*|��6�r}�䳽kSt�>�!�prμ=F{��_��X������4 :U��:[;�2;�O>;�D;}�F;��G;S=H;�pH;��H;��H;�H;�H;�H;��H;��H;��H;��H;��H;�H;�H;�H;��H;��H;�pH;S=H;��G;~�F;�D;�O>;�2;[;W��:0 :�����X���_�=F{�prμ>�!�kSt�䳽r}��6��*|�B��D�߾����O/��N�c�h���y�      ?v��c���X ��c�h�9E�Y��l���}㼾~���nH�Ո�{�ý�Ȅ��s/��o��#�����J���к(�9|g�:m;l0;7]=;�C;1�F;��G;W6H;lmH;U�H;ߥH;ŶH;6�H;}�H;�H;?�H;�H;?�H;�H;}�H;3�H;ŶH;ߥH;T�H;imH;W6H;��G;2�F;�C;3]=;o0;m;|g�:8�9�кJ������#���o��s/��Ȅ�{�ýՈ��nH�~��}㼾l���Y��9E�c�h�X ��c���      ~h��1���c�����y�YvS�rM+��v�9ɾ�����T�!]�\ν����z\8�����x���%�B���8��8�9�-�:��;��.;2�<;oC;�dF;�G;�1H;0kH;֌H;�H;�H;��H;�H;��H;�H;��H;�H;��H;�H;��H;�H;�H;ӌH;,kH;�1H;�G;�dF;oC;/�<;��.;��;�-�:0�9:��B����%��x�����y\8�����\ν!]��T�����9ɾ�v�rM+�YvS���y�c���1���      gܿ5�ֿ�aǿ?^��1���[o���7����iþ�(���-=��` �A���_�1]�,p���I�C�ѻ]�)�`�R���:V�
;�*;4�:;�B;UIF;C�G;�lH;E�H;��H;{�H;��H;��H;��H;��H;D�H;��H;D�H;��H;��H;��H;��H;{�H;��H;B�H;�lH;C�G;VIF;�B;2�:;�*;V�
;��:��R�]�)�B�ѻ�I�,p��1]��_�A���` ��-=��(���iþ����7�[o�1���?^���aǿ5�ֿ      5�ֿEpѿ�¿������bXi�ѕ3��
�WD��Gl��C�9��.���R��!\� �bx��)�E��ͻ��$� ��	��:d�;��*;L�:;*�B;4UF;��G;enH;ߡH;�H;��H;��H;��H;��H;��H;X�H;��H;X�H;��H;��H;��H;��H;��H;�H;ܡH;enH;��G;6UF;*�B;I�:;��*;d�;	��:0����$��ͻ*�E�bx�� �!\��R���.��C�9�Gl��WD���
�ѕ3�bXi��������¿Fpѿ      �aǿ�¿����������"Y��f'�����8o���.}��k/����&ڟ�#<Q�.#�
ע��(;������ #7�-�:�;�,;��;;�C;UwF;5�G;�rH;l�H;ѸH;P�H;4�H;1�H;��H;��H;��H;�H;��H;��H;��H;0�H;5�H;P�H;θH;i�H;�rH;5�G;UwF;�C;��;;�,;�;-�: %7�������(;�
ע�.#�#<Q�&ڟ�����k/��.}�8o�������f'��"Y�����������¿      ?^������l���[o���@�*�&�޾����<ce�1����ڽ����g@������R���O*�8G��ƛ���G^9b��:/;�d.;�<;ՐC;H�F;��G;�yH;֥H;H�H;^�H;��H;��H;�H;,�H;��H;R�H;��H;,�H;�H;��H;��H;^�H;G�H;ӥH;�yH;��G;H�F;ԐC;�<;�d.;/;f��:�G^9ƛ��7G���O*��R������g@�������ڽ1��<ce�����&�޾*���@�[o�l�������      1����������[o��!J�M�#��\��XD������|PH�����b��!C��� +���ټ&����ܿ��Ȭ��p�:c��:t�;�Y1;)>;�0D;��F;�H;��H;�H;<�H;��H;��H;C�H;��H;��H;��H;��H;��H;��H;��H;B�H;��H;��H;:�H;�H;��H;�H;��F;�0D;&>;�Y1;t�;g��:h�:Ƭ��ۿ����&����ټ� +�!C���b�����|PH�����XD���\��M�#��!J�[o��������      [o�bXi��"Y���@�M�#��
��о�A���i���(����wr���_��5��ɺ�j�`��<��B�d���\�L�X:�P�:a;�4;ާ?;��D;�8G;�0H;֋H;��H;��H;B�H;��H;��H;5�H;��H;H�H;��H;H�H;��H;5�H;��H;��H;B�H;��H;��H;֋H;�0H;�8G;��D;ۧ?;�4;a;�P�:H�X:��\�A�d��<��j�`��ɺ��5��_�wr�������(��i��A���о�
�M�#���@��"Y�bXi�      ��7�ѕ3��f'�*��\���о�����.}��-=�|
���Ľ\��+:�����������7�GĻ��$��M��A��:�{;�D&;6,8;>JA;6�E;�G;�LH;#�H;��H;e�H;�H;B�H;��H;��H;Z�H;��H;R�H;��H;Z�H;��H;��H;C�H;�H;c�H;��H;#�H;�LH;�G;3�E;;JA;5,8;�D&;�{;9��:�M����$�GĻ��7���������+:�\����Ľ|
��-=��.}������о�\��*��f'�ѕ3�      ���
�����&�޾XD���A���.}�*�D�it���ڽ�!��\����Z�ļ�
v�5�������IɺhT�9=��:C(;�-;Ƌ;;��B;�IF;��G;NfH;ٝH;-�H;`�H;�H;��H;��H;��H;��H;)�H;��H;*�H;��H;��H;��H;��H;�H;`�H;*�H;ٝH;MfH;��G;�IF;��B;Ƌ;;�-;E(;;��:hT�9�Iɺ����5���
v�Z�ļ���\��!����ڽit�*�D��.}��A��XD��&�޾�����
�      �iþWD��8o�����������i��-=�jt����R��iys�{ +����v񗼍(;��ѻ�s@�<�!��4j:.Q�:�;�D3;u�>;EFD;��F;�	H;n|H;ͥH;��H;j�H;.�H;0�H;��H;V�H;k�H;��H;�H;��H;n�H;W�H;��H;1�H;1�H;h�H;��H;ϥH;l|H;�	H;��F;BFD;t�>;�D3;�;*Q�:�4j:0�!��s@��ѻ�(;�v����{ +�iys��R�� ��jt��-=��i���������8o��WD��      �(��Gl���.}�<ce�|PH���(�}
���ڽ�R���{�C�6�� �*p��X�`�Ũ��,���HҺ O^9:�;�~(;f�8;JA;6|E;OjG;�=H;{�H;�H;`�H;��H;c�H;��H;��H;�H;��H;,�H;��H;,�H;��H;�H;��H;��H;e�H;��H;]�H;�H;{�H;>H;LjG;5|E;JA;d�8;�~(;�;:O^9�HҺ�,��Ũ�X�`�*p��� �C�6��{��R����ڽ}
���(�|PH�<ce��.}�Gl��      �-=�C�9��k/�1��������Ľ�!��iys�C�6�%#��ɺ��vz����/^��B�$�P}���r:b��:�;�Y1;4I=;ixC;\wF;_�G;AfH;~�H;��H;��H;��H;��H;�H;�H;��H;��H;��H;��H;��H;��H;��H;�H;�H;��H;��H;��H;��H;}�H;CfH;\�G;YwF;fxC;2I=;�Y1;�;b��:��r:X}�A�$�/^������vz��ɺ�%#�C�6�iys��!����Ľ����1���k/�C�9�      �` ��.�������ڽ�b��wr��\��\�{ +�� ��ɺ�=��O*�4ͻ�5R��ƅ���:���:��;�);*u8;��@;�*E;�8G;$H;��H;z�H;2�H;d�H;��H;��H;��H;:�H;��H;,�H;�H;\�H;�H;-�H;��H;;�H;��H;��H;��H;d�H;2�H;y�H;��H;$H;�8G;�*E;��@;*u8;�);��;���:��:�ƅ��5R�4ͻ�O*�=��ɺ�� �{ +�\�\��wr���b����ڽ��.��      A���R��&ڟ�����!C���_�,:�������*p���vz��O*��4ֻ�k�ګ����09��:41;�� ;�D3;z�=;�C;!lF;��G;]H;חH;��H;>�H;}�H;��H;��H;�H;6�H;G�H;��H;��H;��H;��H;��H;G�H;8�H;�H;��H;��H;|�H;?�H;��H;ڗH; ]H;��G;lF;�C;{�=;�D3;�� ;61;��:��09ګ���k��4ֻ�O*��vz�*p����輤��,:��_�!C������&ڟ��R��      �_�!\�"<Q�g@�� +��5�����Z�ļv�X�`����4ͻ�k��Hɺ ]6���::Q�:U�;e.;��:;V�A;d|E;�NG;'H;?�H;�H;��H;��H;j�H;��H;��H;o�H;5�H;�H;L�H;��H;<�H;��H;L�H;�H;5�H;t�H;��H;��H;h�H;��H;��H;
�H;>�H;'H;�NG;d|E;V�A;��:;e.;X�;8Q�:��: Z6��Hɺ�k�3ͻ���X�`�v�Z�ļ�����5�� +�g@�"<Q�!\�      0]� �.#�������ټ�ɺ������
v��(;�ƨ�/^���5R�ޫ�� _6���:?��:*�;S�*;,8;�!@;��D;��F;5�G;fH;H;ͰH;޿H;��H;!�H;�H;_�H;��H;	�H;��H;��H;f�H;��H;f�H;��H;��H;	�H;��H;b�H;�H;�H;��H;޿H;аH;ęH;fH;1�G;��F;��D;�!@;,8;V�*;*�;?��: ��: _6�ޫ���5R�/^��ƨ��(;��
v������ɺ���ټ����.#� �      ,p��bx��	ע��R��&��l�`���7�6���ѻ�,��B�$��ƅ���09��:E��:�;(;�Z6;��>;�C;,IF;�G;)EH;��H;��H;�H;N�H;k�H;T�H;7�H;�H;��H;��H;N�H;)�H;��H;��H;��H;)�H;N�H;��H;��H;�H;9�H;Q�H;k�H;N�H;�H;��H;��H;%EH;�G;)IF;�C;��>;�Z6;(;�;E��:��:��09�ƅ�B�$��,���ѻ6����7�j�`�&���R��	ע�bx��      �I�'�E��(;��O*����<��GĻ�����s@��HҺX}�:��:4Q�:,�; (;@�5;�>;nC;r�E;�cG;z$H;8|H;x�H;^�H;��H;��H;{�H;�H;_�H;��H;��H;��H;��H;��H;�H;2�H;�H;��H;��H;��H;��H;��H;^�H;�H;|�H;��H;��H;^�H;t�H;3|H;z$H;�cG;t�E;oC;>;@�5;(;,�;4Q�:��:��:`}��HҺ�s@�����GĻ�<�����O*��(;�*�E�      F�ѻ�ͻ���8G��޿��P�d���$��Iɺ<�!��N^9��r:}��:21;S�;S�*;�Z6;�>;k�B;��E;9G;�	H;>nH;W�H;��H;�H;��H;��H;�H;��H;@�H;��H;��H;?�H;:�H;��H;D�H;g�H;D�H;��H;<�H;=�H;��H;��H;@�H;��H;�H;��H;��H;�H;��H;U�H;@nH;�	H; 9G;��E;n�B;�>;�Z6;U�*;T�;41;}��:��r:�N^94�!��Iɺ��$�L�d�ڿ��8G������ͻ      Y�)���$�	����Ԭ����\��M��8T�9�4j:釶:Z��:��;�� ;e.;,8;��>;nC;��E;�)G;��G;QdH;��H;ثH;��H;��H;x�H;�H;�H;��H;��H;��H;��H;��H;��H;@�H;u�H;��H;u�H;@�H;��H;��H;��H;��H;��H;��H;�H;�H;{�H;��H;��H;ӫH;��H;OdH;��G;�)G;êE;nC;��>;,8;e.;�� ;��;`��:燶:�4j:8T�9�M����\�Ȭ��ě��	����$�      P�R�P�� 7��G^9d�:0�X:/��:/��:Q�:�;�;�);�D3;~�:;�!@;�C;p�E;9G;��G;�`H;��H;X�H;^�H;��H;��H;u�H;��H;��H;��H;�H;��H;L�H;+�H;��H;o�H;��H;��H;��H;o�H;��H;)�H;M�H;��H;�H;��H;��H;��H;x�H;��H;��H;[�H;X�H;��H;�`H;��G;9G;p�E;�C;�!@;~�:;�D3;�);�;�; Q�:1��:3��:@�X:��:�G^9  7����      ��:'��:3�:R��:S��:�P�:�{;?(;�;�~(;�Y1;%u8;w�=;R�A;��D;(IF;�cG;�	H;OdH;��H;��H;�H;t�H;7�H;�H;��H;��H;��H;h�H;&�H;��H;��H;��H;)�H;��H;��H;��H;��H;��H;)�H;��H;��H;��H;#�H;e�H;��H;��H;��H;�H;3�H;r�H;�H;��H;��H;QdH;�	H;�cG;(IF;��D;S�A;x�=;%u8;�Y1;�~(;�;@(;�{;Q�:U��:X��:9�:��:      ]�
;��;)�;";r�;a;�D&;�-;�D3;d�8;4I=;��@;ߐC;c|E;��F;�G;x$H;>nH;��H;Y�H;�H;��H;{�H;a�H;��H;��H;%�H;��H;��H;J�H;c�H;7�H;��H;a�H;��H;��H;��H;��H;��H;a�H;��H;7�H;c�H;F�H;��H;��H;$�H;��H;��H;\�H;z�H;��H;�H;[�H;��H;@nH;x$H;�G;��F;c|E;ߐC;��@;2I=;c�8;�D3;�-;�D&;a;��;$;*�;|�;      �*;��*;�,;�d.;�Y1;�4;5,8;��;;t�>;JA;cxC;�*E;lF;�NG;2�G;%EH;6|H;W�H;֫H;^�H;t�H;|�H;�H;<�H;:�H;��H;O�H;,�H;��H;�H;��H;��H;(�H;|�H;��H;��H;��H;��H;��H;|�H;%�H;��H;��H;�H;��H;,�H;L�H;��H;<�H;9�H;�H;~�H;p�H;`�H;իH;Y�H;3|H;%EH;2�G;�NG;lF;�*E;fxC;JA;t�>;Ë;;5,8;�4;�Y1;�d.;�,;��*;      H�:;[�:;��;;�<;)>;ڧ?;DJA;��B;BFD;3|E;YwF;�8G;��G;~'H;fH;��H;w�H;��H;��H;��H;2�H;^�H;:�H;%�H;[�H;��H;��H;u�H;��H;��H;Y�H;��H;^�H;��H;��H;��H;�H;��H;��H;��H;\�H;��H;[�H;��H;��H;v�H;��H;��H;\�H;"�H;9�H;^�H;0�H;��H;��H;��H;u�H;��H;fH;~'H;��G;�8G;XwF;2|E;CFD;��B;BJA;ۧ?;1>;�<;��;;L�:;      �B;3�B;�C;אC;�0D;��D;2�E;�IF;��F;HjG;Z�G;$H;�\H;?�H;ęH;��H;e�H;�H;��H;��H;�H;��H;@�H;b�H;��H;��H;;�H;��H;j�H;7�H;��H;�H;q�H;��H;��H;��H;��H;��H;��H;��H;o�H;�H;��H;7�H;i�H;��H;:�H;��H;��H;_�H;?�H;��H;�H;��H;��H;�H;a�H;��H;řH;?�H;�\H;�$H;\�G;IjG;��F;�IF;2�E;��D;�0D;אC;�C;3�B;      ^IF;AUF;HwF;E�F;��F;�8G;��G;��G;�	H;�=H;<fH;��H;ԗH;�H;ɰH;�H;��H;��H;t�H;u�H;}�H;��H;��H;��H;��H;9�H;h�H;L�H;�H;��H;�H;a�H;v�H;��H;��H;��H;��H;��H;��H;��H;u�H;c�H;�H;��H;��H;L�H;g�H;:�H;��H;��H;��H;��H;y�H;t�H;u�H;��H;��H;�H;ʰH;�H;ԗH;��H;=fH;�=H;�	H;��G;��G;�8G;��F;E�F;HwF;6UF;      N�G;��G;2�G;��G;�H;�0H;�LH;KfH;m|H;u�H;}�H;z�H;��H;��H;ݿH;N�H;��H;��H;�H;��H;��H;%�H;L�H;��H;6�H;k�H;=�H;��H;��H;��H;"�H;o�H;��H;��H;��H;��H;��H;��H;��H;��H;��H;o�H;!�H;��H;��H;��H;<�H;i�H;:�H;��H;L�H;%�H;��H;��H;�H;��H;��H;N�H;ݿH;��H;��H;{�H;~�H;w�H;n|H;KfH;�LH;�0H;�H;��G;1�G;��G;      �lH;hnH;�rH;�yH;��H;ՋH;"�H;ܝH;ͥH;�H;��H;3�H;>�H;��H;��H;j�H;y�H;�H;�H;��H;��H;��H;+�H;x�H;}�H;M�H;��H;u�H;��H;*�H;K�H;y�H;��H;��H;��H;��H;��H;��H;��H;��H;��H;x�H;I�H;(�H;��H;u�H;��H;M�H;~�H;v�H;+�H;��H;��H;��H;�H;�H;x�H;j�H;��H;��H;<�H;6�H;��H;�H;ϥH;ݝH;"�H;֋H;��H;�yH;�rH;snH;      U�H;�H;f�H;֥H;�H;��H;��H;+�H;��H;]�H;��H;g�H;|�H;g�H;!�H;T�H;�H;��H;��H;��H;e�H;��H;��H;��H;c�H;�H;��H;��H;�H;P�H;n�H;��H;��H;��H;��H;��H;��H;��H;��H;��H;��H;��H;m�H;O�H;�H;��H;��H;�H;f�H;��H;��H;��H;b�H;��H;��H;��H;�H;T�H;!�H;h�H;}�H;g�H;��H;]�H;��H;-�H;��H;��H;�H;ץH;f�H;֡H;      ��H;�H;׸H;F�H;F�H;��H;f�H;a�H;n�H;��H;��H;��H;��H;��H;�H;9�H;a�H;;�H;��H;�H;%�H;E�H;�H;��H;/�H;��H;��H;*�H;O�H;d�H;��H;��H;��H;��H;��H;��H;��H;��H;��H;��H;��H;��H;��H;c�H;N�H;*�H;��H;��H;0�H;��H;�H;E�H;%�H;�H;��H;>�H;_�H;:�H;�H;��H;��H;��H;��H;��H;q�H;d�H;f�H;��H;F�H;G�H;ԸH;�H;      ~�H;��H;Z�H;g�H;��H;=�H;�H;�H;5�H;g�H;��H;��H;��H;��H;b�H;�H;��H;��H;��H;��H;��H;a�H;��H;\�H;��H;�H;�H;L�H;k�H;��H;��H;��H;}�H;��H;��H;��H;n�H;��H;��H;��H;|�H;��H;��H;��H;m�H;L�H;�H;�H;��H;\�H;��H;a�H;��H;��H;��H;��H;��H;�H;c�H;��H;��H;��H;��H;j�H;5�H;�H;�H;>�H;��H;g�H;Y�H;��H;      ��H;��H;9�H;��H;��H;��H;B�H;��H;1�H;��H;!�H;��H;�H;v�H;��H;��H;��H;��H;��H;S�H;��H;:�H;��H;��H;�H;`�H;k�H;y�H;��H;��H;��H;��H;}�H;x�H;��H;o�H;e�H;n�H;��H;x�H;y�H;��H;��H;��H;��H;{�H;n�H;`�H;�H;��H;��H;:�H;��H;S�H;��H;��H;��H;��H;��H;x�H;�H;��H;"�H;��H;5�H;��H;D�H;��H;��H;��H;9�H;��H;      ��H;��H;7�H;��H;L�H;��H;��H;��H;��H;��H;�H;E�H;;�H;:�H;�H;��H;��H;;�H;��H;/�H;��H;��H;"�H;`�H;h�H;u�H;��H;��H;��H;��H;�H;�H;��H;��H;^�H;]�H;��H;]�H;^�H;��H;}�H;��H;�H;��H;��H;��H;��H;u�H;k�H;a�H;"�H;��H;��H;0�H;��H;<�H;��H;��H;�H;<�H;;�H;C�H;�H;��H;��H;��H;��H;��H;D�H;��H;7�H;��H;      ��H;��H;��H;�H;��H;,�H;��H;��H;X�H;�H;��H;��H;I�H;�H;��H;W�H;��H;:�H;��H;��H;-�H;^�H;x�H;��H;��H;��H;��H;��H;��H;��H;}�H;x�H;{�H;j�H;Y�H;`�H;d�H;`�H;Y�H;j�H;y�H;{�H;}�H;��H;��H;��H;��H;��H;��H;��H;{�H;`�H;,�H;��H;��H;<�H;��H;W�H;��H;
�H;K�H;��H;��H;�H;[�H;��H;��H;0�H;��H;�H;��H;��H;      ��H;��H;��H;3�H;��H;��H;_�H;��H;t�H;�H;��H;:�H;��H;S�H;��H;2�H;��H;��H;@�H;q�H;��H;��H;��H;��H;��H;��H;��H;��H;��H;��H;��H;��H;]�H;Z�H;d�H;Z�H;=�H;Z�H;d�H;Z�H;Z�H;��H;��H;��H;��H;��H;��H;��H;��H;��H;��H;��H;��H;r�H;@�H;��H;��H;2�H;��H;S�H;��H;:�H;��H;�H;u�H;��H;_�H;��H;��H;1�H;��H;��H;      8�H;_�H;��H;��H;��H;@�H;��H;3�H;��H;,�H;��H;*�H;��H;��H;j�H;��H;�H;>�H;v�H;��H;��H;��H;��H;��H;��H;��H;��H;��H;��H;��H;��H;r�H;]�H;d�H;Z�H;V�H;G�H;V�H;Z�H;a�H;\�H;u�H;��H;��H;��H;��H;��H;��H;��H;��H;��H;��H;��H;��H;v�H;@�H;�H;��H;k�H;��H;��H;*�H;��H;.�H;��H;3�H;��H;D�H;��H;��H;��H;X�H;      ��H;�H;�H;Q�H;��H;��H;S�H;��H;&�H;��H;��H;h�H;��H;F�H;��H;��H;7�H;`�H;��H;��H;��H;��H;��H;�H;��H;��H;��H;��H;��H;��H;q�H;k�H;��H;g�H;=�H;G�H;A�H;G�H;=�H;g�H;��H;m�H;q�H;��H;��H;��H;��H;��H;��H;�H;��H;��H;��H;��H;��H;a�H;6�H;��H;��H;F�H;��H;h�H;��H;��H;'�H;��H;S�H;��H;��H;Q�H;�H;��H;      8�H;_�H;��H;��H;��H;@�H;��H;4�H;��H;,�H;��H;*�H;��H;��H;k�H;��H;�H;>�H;v�H;��H;��H;��H;��H;��H;��H;��H;��H;��H;��H;��H;��H;r�H;]�H;d�H;Z�H;V�H;G�H;V�H;Z�H;a�H;\�H;u�H;��H;��H;��H;��H;��H;��H;��H;��H;��H;��H;��H;��H;v�H;@�H;�H;��H;j�H;��H;��H;*�H;��H;-�H;��H;2�H;��H;D�H;��H;��H;��H;W�H;      ��H;��H;��H;3�H;��H;��H;_�H;��H;t�H;�H;��H;:�H;��H;T�H;��H;2�H;��H;��H;@�H;t�H;��H;��H;��H;��H;��H;��H;��H;��H;��H;��H;��H;��H;]�H;Z�H;d�H;Z�H;=�H;Z�H;d�H;Z�H;Z�H;��H;��H;��H;��H;��H;��H;��H;��H;��H;��H;��H;��H;q�H;@�H;��H;��H;2�H;��H;S�H;��H;:�H;��H;�H;t�H;��H;_�H;��H;��H;1�H;��H;��H;      ��H;��H;��H;�H;��H;,�H;��H;��H;Z�H;�H;��H;��H;K�H;
�H;��H;W�H;��H;:�H;��H;��H;0�H;`�H;y�H;��H;��H;��H;��H;��H;��H;��H;}�H;x�H;{�H;j�H;Y�H;`�H;d�H;`�H;Y�H;j�H;y�H;{�H;}�H;��H;��H;��H;��H;��H;��H;��H;y�H;^�H;,�H;��H;��H;<�H;��H;W�H;��H;�H;I�H;��H;��H;�H;Z�H;��H;��H;0�H;��H;�H;��H;��H;      ��H;��H;8�H;��H;J�H;��H;��H;��H;��H;��H;�H;C�H;;�H;<�H;�H;��H;��H;;�H;��H;/�H;��H;��H;#�H;a�H;k�H;v�H;��H;��H;��H;��H;�H;�H;��H;�H;^�H;]�H;��H;]�H;^�H;�H;}�H;��H;�H;��H;��H;��H;��H;t�H;h�H;^�H;!�H;��H;��H;/�H;��H;;�H;��H;��H;�H;:�H;9�H;C�H;�H;��H;��H;��H;��H;��H;C�H;��H;5�H;��H;      ��H;��H;<�H;��H;��H;��H;F�H;��H;3�H;��H;!�H;��H;�H;x�H;��H;��H;��H;��H;��H;T�H;��H;:�H;��H;��H;�H;a�H;n�H;{�H;��H;��H;��H;��H;|�H;x�H;��H;n�H;e�H;n�H;��H;x�H;y�H;��H;��H;��H;��H;y�H;m�H;^�H;�H;��H;��H;:�H;��H;S�H;��H;��H;��H;��H;��H;v�H;�H;��H;"�H;��H;3�H;��H;C�H;��H;��H;��H;;�H;��H;      ~�H;��H;Z�H;g�H;��H;=�H;�H;�H;5�H;h�H;��H;��H;��H;��H;c�H;!�H;��H;��H;��H;��H;��H;a�H;��H;]�H;��H;�H;�H;L�H;m�H;��H;��H;��H;}�H;��H;��H;��H;n�H;��H;��H;��H;{�H;��H;��H;��H;m�H;L�H;�H;�H;��H;[�H;��H;a�H;��H;��H;��H;��H;��H;�H;b�H;��H;��H;��H;��H;h�H;5�H;�H;�H;>�H;��H;g�H;Z�H;��H;      ��H;�H;ָH;G�H;C�H;��H;h�H;b�H;q�H;��H;��H;��H;��H;��H;�H;:�H;a�H;;�H;��H;�H;)�H;E�H;�H;��H;0�H;��H;��H;*�H;O�H;d�H;��H;��H;��H;��H;��H;��H;��H;��H;��H;��H;��H;��H;��H;c�H;O�H;*�H;��H;��H;/�H;��H;�H;E�H;#�H;�H;��H;;�H;_�H;:�H;�H;��H;��H;��H;��H;��H;q�H;b�H;h�H;��H;C�H;F�H;׸H;�H;      M�H;ݡH;l�H;ԥH;�H;��H;��H;.�H;��H;]�H;��H;h�H;}�H;h�H;!�H;T�H;�H;��H;��H;��H;h�H;��H;��H;��H;f�H;�H;��H;��H;�H;P�H;m�H;��H;��H;��H;��H;��H;��H;��H;��H;��H;��H;��H;n�H;N�H;�H;��H;��H;�H;c�H;��H;��H;��H;b�H;��H;��H;��H;�H;U�H;!�H;g�H;|�H;g�H;��H;\�H;��H;-�H;��H;��H;�H;ҥH;j�H;ߡH;      �lH;fnH;�rH;�yH;��H;֋H;"�H;ߝH;ͥH;�H;��H;6�H;<�H;��H;��H;j�H;y�H;�H;�H;��H;��H;��H;+�H;x�H;~�H;M�H;��H;u�H;��H;*�H;I�H;x�H;��H;��H;��H;��H;��H;��H;��H;��H;��H;{�H;K�H;(�H;��H;u�H;��H;M�H;}�H;v�H;+�H;��H;��H;��H;�H;�H;x�H;k�H;��H;��H;>�H;5�H;��H;�H;ϥH;ܝH;"�H;ҋH;��H;�yH;�rH;snH;      H�G;��G;1�G;��G;�H;�0H;�LH;KfH;m|H;x�H;~�H;{�H;��H;��H;ݿH;O�H;��H;��H;�H;��H;��H;%�H;L�H;��H;:�H;k�H;=�H;��H;��H;��H;!�H;o�H;��H;��H;��H;��H;��H;��H;��H;��H;��H;q�H;"�H;��H;��H;��H;<�H;k�H;6�H;��H;J�H;%�H;��H;��H;�H;��H;��H;M�H;ݿH;��H;��H;z�H;~�H;w�H;m|H;JfH;�LH;�0H;�H;��G;/�G;��G;      fIF;:UF;QwF;G�F;��F;�8G;��G;��G;�	H;�=H;<fH;��H;ԗH;�H;ɰH;�H;��H;��H;u�H;t�H;�H;��H;��H;��H;��H;:�H;h�H;L�H;�H;��H;�H;a�H;v�H;��H;��H;��H;��H;��H;��H;��H;t�H;c�H;�H;��H;��H;L�H;g�H;:�H;��H;��H;��H;��H;y�H;t�H;t�H;��H;��H;�H;ɰH;�H;ԗH;��H;<fH;�=H;�	H;��G;��G;�8G;��F;H�F;RwF;1UF;      �B;3�B;�C;אC;�0D;��D;2�E;�IF;��F;KjG;]�G;�$H;�\H;?�H;řH;��H;b�H;�H;��H;��H;�H;��H;?�H;b�H;��H;��H;;�H;��H;m�H;9�H;��H;�H;q�H;��H;��H;��H;��H;��H;��H;��H;o�H;�H;��H;6�H;h�H;��H;:�H;��H;��H;a�H;?�H;��H;�H;��H;��H;�H;a�H;��H;ęH;>�H;�\H;$H;Z�G;FjG;��F;�IF;2�E;��D;�0D;אC;�C;3�B;      K�:;X�:;��;;�<;">;�?;@JA;��B;EFD;5|E;ZwF;�8G;��G;'H;fH;��H;w�H;��H;��H;��H;4�H;^�H;:�H;%�H;\�H;��H;��H;v�H;��H;��H;[�H;��H;]�H;��H;��H;��H;�H;��H;��H;��H;]�H;��H;Y�H;��H;��H;u�H;��H;��H;[�H;$�H;9�H;^�H;/�H;��H;��H;��H;u�H;��H;fH;'H;��G;�8G;XwF;3|E;CFD;��B;@JA;�?;1>;�<;��;;J�:;      �*;��*;�,;�d.;�Y1;�4;9,8;��;;t�>;JA;fxC;�*E;lF;�NG;2�G;&EH;6|H;V�H;իH;^�H;u�H;~�H;�H;<�H;<�H;��H;O�H;,�H;��H;�H;��H;��H;(�H;|�H;��H;��H;��H;��H;��H;|�H;%�H;��H;��H;�H;��H;,�H;L�H;��H;:�H;9�H;�H;|�H;p�H;`�H;֫H;W�H;5|H;%EH;4�G;�NG;lF;�*E;cxC;JA;t�>;��;;9,8;�4;�Y1;�d.;�,;��*;      ]�
;��;)�;$;p�;a;�D&;�-;�D3;c�8;4I=;��@;ߐC;c|E;��F;�G;x$H;?nH;��H;Y�H;�H;��H;|�H;a�H;��H;��H;'�H;��H;��H;J�H;c�H;7�H;��H;a�H;��H;��H;��H;��H;��H;a�H;��H;7�H;c�H;F�H;��H;��H;$�H;��H;��H;\�H;x�H;��H;�H;[�H;��H;?nH;w$H;�G;��F;c|E;ߐC;��@;2I=;d�8;�D3;�-;�D&;a;��;";*�;z�;      ��:��:9�:T��:S��:�P�:�{;C(;�;�~(;�Y1;%u8;x�=;S�A;��D;(IF;�cG;�	H;QdH;��H;��H;�H;t�H;7�H;�H;��H;��H;��H;h�H;&�H;��H;��H;��H;(�H;��H;��H;��H;��H;��H;)�H;��H;��H;��H;#�H;c�H;��H;��H;��H;�H;3�H;r�H;�H;��H;��H;OdH;�	H;�cG;(IF;��D;S�A;w�=;%u8;�Y1;�~(;�;B(;�{; Q�:[��:T��:9�:��:      `�R� �� 7��G^9p�:8�X:3��:1��: Q�:�;�;�);�D3;~�:;�!@;�C;p�E;9G;��G;�`H;��H;X�H;^�H;��H;��H;x�H;��H;��H;��H;�H;��H;L�H;+�H;��H;o�H;��H;��H;��H;o�H;��H;)�H;M�H;��H;�H;��H;��H;��H;u�H;��H;��H;[�H;X�H;��H;�`H;��G;9G;p�E;�C;�!@;~�:;�D3;�);�;�; Q�:1��:3��:<�X:��:�G^9  7����      Y�)���$�	��ě��֬����\��M��8T�9�4j:燶:`��:��;�� ;e.;,8;��>;oC;��E;�)G;��G;RdH;��H;ثH;��H;��H;z�H;�H;�H;��H;��H;��H;��H;��H;��H;@�H;t�H;��H;u�H;@�H;��H;��H;��H;��H;��H;��H;�H;	�H;z�H;��H;��H;ӫH;��H;NdH;��G;�)G;êE;mC;��>;,8;e.;�� ;��;Z��:釶:�4j:0T�9�M����\�ʬ����	����$�      D�ѻ�ͻ���8G��޿��R�d���$��Iɺ<�!��N^9��r:}��:41;T�;U�*;�Z6;�>;m�B;��E;9G;�	H;@nH;W�H;��H;�H;��H;��H;�H;��H;A�H;��H;��H;?�H;<�H;��H;D�H;g�H;D�H;��H;:�H;=�H;��H;��H;>�H;��H;�H;��H;��H;�H;��H;U�H;>nH;�	H;9G;��E;k�B;�>;�Z6;S�*;S�;21;}��:��r:�N^9<�!��Iɺ��$�K�d�ܿ��8G������ͻ      �I�'�E��(;��O*����<��GĻ�����s@��HҺX}�:��:4Q�:,�;(;C�5;�>;oC;r�E;�cG;z$H;9|H;x�H;^�H;��H;��H;|�H;�H;_�H;��H;��H;��H;��H;��H;�H;2�H;�H;��H;��H;��H;��H;��H;\�H;�H;{�H;��H;��H;^�H;t�H;2|H;z$H;�cG;t�E;nC; >;@�5; (;,�;4Q�:��:��:X}��HҺ�s@�����GĻ�<�����O*��(;�)�E�      ,p��bx��	ע��R��&��k�`���7�6���ѻ�,��B�$��ƅ���09��:E��:�;(;�Z6;��>;�C;,IF;�G;(EH;��H;��H;�H;Q�H;k�H;U�H;9�H;�H;��H;��H;N�H;)�H;��H;��H;��H;)�H;N�H;��H;��H;�H;7�H;O�H;k�H;M�H;�H;��H;��H;%EH;�G;)IF;�C;��>;�Z6;(;�;E��:��:��09�ƅ�B�$��,���ѻ6����7�j�`�&���R��	ע�bx��      0]� �.#�������ټ�ɺ������
v��(;�ƨ�0^���5R�ޫ�� _6���:?��:*�;S�*;,8;�!@;��D;��F;6�G;fH;ęH;ΰH;޿H;��H;#�H;�H;b�H;��H;�H;��H;��H;f�H;��H;f�H;��H;��H;	�H;��H;_�H; �H;�H;��H;ݿH;ΰH;H;fH;/�G;��F;��D;�!@;,8;V�*;*�;?��:��: _6�ޫ���5R�0^��ƨ��(;��
v������ɺ���ټ����.#� �      �_�!\�"<Q�g@�� +��5�����Z�ļv�X�`����4ͻ�k��Hɺ \6���::Q�:W�;e.;��:;V�A;d|E;�NG;�'H;>�H;	�H;��H;��H;j�H;��H;��H;q�H;6�H;�H;L�H;��H;<�H;��H;L�H;�H;3�H;q�H;��H;��H;g�H;��H;��H;	�H;?�H;~'H;�NG;d|E;V�A;��:;e.;X�;8Q�:��: ]6��Hɺ�k�4ͻ���W�`�v�Z�ļ�����5�� +�g@�"<Q�!\�      A���R��&ڟ�����!C���_�,:�������*p���vz��O*��4ֻ�k�ګ����09��:61;�� ;�D3;{�=;�C;"lF;��G; ]H;ؗH;��H;?�H;}�H;��H;��H;�H;8�H;G�H;��H;��H;��H;��H;��H;G�H;5�H;�H;��H;��H;{�H;>�H;��H;ۗH;]H;��G;lF;�C;z�=;�D3;�� ;61;��:��09ګ���k��4ֻ�O*��vz�*p����輤��,:��_�!C������&ڟ��R��      �` ��.�������ڽ�b��wr��\��\�{ +�� ��ɺ�=��O*�4ͻ�5R��ƅ���:���:��;�);'u8;��@;�*E;�8G;$H;��H;z�H;2�H;e�H;��H;��H;��H;<�H;��H;-�H; �H;\�H; �H;,�H;��H;8�H;��H;��H;��H;c�H;2�H;y�H;��H;$H;�8G;�*E;��@;*u8;�);��;���:��:�ƅ��5R�4ͻ�O*�=��ɺ�� �{ +�\�\��wr���b����ڽ��.��      �-=�C�9��k/�1��������Ľ�!��jys�C�6�%#��ɺ��vz����/^��A�$�P}���r:b��:�;�Y1;2I=;ixC;]wF;\�G;AfH;~�H;��H;��H;��H;��H;�H;�H;��H;��H;��H;��H;��H;��H;��H;�H;�H;��H;��H;��H;��H;}�H;AfH;_�G;YwF;fxC;4I=;�Y1;�;b��:��r:X}�D�$�/^������vz��ɺ�%#�C�6�iys��!����Ľ����1���k/�C�9�      �(��Gl���.}�<ce�|PH���(�}
���ڽ�R���{�C�6�� �*p��X�`�Ũ��,���HҺ O^9:�;�~(;d�8;JA;7|E;LjG;�=H;{�H;�H;`�H;��H;e�H;��H;��H;�H;��H;,�H;��H;,�H;��H;�H;��H;��H;c�H;��H;]�H;�H;y�H;�=H;OjG;5|E;JA;f�8;�~(;�;:O^9�HҺ�,��Ũ�X�`�*p��� �C�6��{��R����ڽ}
���(�|PH�<ce��.}�Gl��      �iþWD��8o�����������i��-=�jt� ���R��iys�{ +����v񗼍(;��ѻ�s@�4�!��4j:,Q�:�;�D3;u�>;EFD;��F;�	H;n|H;ϥH;��H;h�H;1�H;0�H;��H;W�H;n�H;��H;�H;��H;k�H;V�H;��H;0�H;.�H;h�H;��H;ͥH;l|H;�	H;��F;CFD;t�>;�D3;�;*Q�:�4j:4�!��s@��ѻ�(;�v����{ +�iys��R�� ��jt��-=��i���������8o��WD��      ���
�����&�޾XD���A���.}�*�D�it���ڽ�!��\����Z�ļ�
v�5�������IɺhT�9;��:C(;�-;Ƌ;;��B;�IF;��G;NfH;ٝH;-�H;`�H;�H;��H;��H;��H;��H;)�H;��H;*�H;��H;��H;��H;��H;�H;`�H;*�H;ٝH;MfH;��G;�IF;��B;Ƌ;;�-;E(;7��:hT�9�Iɺ����6���
v�Z�ļ���\��!����ڽit�*�D��.}��A��XD��&�޾�����
�      ��7�ѕ3��f'�*��\���о�����.}��-=�|
���Ľ\��+:�����������7�GĻ��$��M��;��:�{;�D&;6,8;@JA;3�E;�G;�LH;#�H;��H;e�H;�H;B�H;��H;��H;Z�H;��H;R�H;��H;Z�H;��H;��H;B�H;�H;c�H;��H;#�H;�LH;�G;6�E;=JA;5,8;�D&;�{;9��:�M����$�GĻ��7���������+:�\����Ľ|
��-=��.}������о�\��*��f'�ѕ3�      [o�bXi��"Y���@�M�#��
��о�A���i���(����wr���_��5��ɺ�j�`��<��B�d���\�H�X:�P�:a;�4;ާ?;��D;�8G;�0H;֋H;��H;��H;B�H;��H;�H;5�H;��H;H�H;��H;J�H;��H;5�H;��H;��H;B�H;��H;��H;֋H;�0H;�8G;��D;ۧ?;�4;a;�P�:H�X:��\�A�d��<��j�`��ɺ��5��_�wr�������(��i��A���о�
�M�#���@��"Y�bXi�      1����������[o��!J�M�#��\��XD������|PH�����b��!C��� +���ټ&����ܿ��Ȭ��h�:c��:t�;�Y1;)>;�0D;��F;�H;��H;�H;<�H;��H;��H;C�H;��H;��H;��H;��H;��H;��H;��H;B�H;��H;��H;:�H;�H;��H;�H;��F;�0D;'>;�Y1;t�;g��:h�:Ȭ��ۿ����&����ټ� +�!C���b�����|PH�����XD���\��M�#��!J�[o��������      ?^������l���[o���@�*�&�޾����<ce�1����ڽ����g@������R���O*�8G��ƛ���G^9`��:/;�d.;�<;ԐC;H�F;��G;�yH;֥H;J�H;^�H;��H;��H;�H;,�H;��H;R�H;��H;,�H;�H;��H;��H;^�H;G�H;ӥH;�yH;��G;H�F;ՐC;�<;�d.;/;f��:�G^9ƛ��7G���O*��R������g@�������ڽ1��<ce�����&�޾*���@�[o�l�������      �aǿ�¿����������"Y��f'�����8o���.}��k/����&ڟ�#<Q�.#�
ע��(;������ %7�+�:�;�,;��;;�C;UwF;5�G;�rH;l�H;ѸH;P�H;5�H;1�H;��H;��H;��H;�H;��H;��H;��H;0�H;4�H;P�H;θH;i�H;�rH;5�G;UwF;�C;��;;�,;�;-�: %7�������(;�
ע�.#�#<Q�&ڟ�����k/��.}�8o�������f'��"Y�����������¿      5�ֿEpѿ�¿������bXi�ѕ3��
�WD��Gl��C�9��.���R��!\� �bx��)�E��ͻ��$� ��	��:d�;��*;L�:;*�B;4UF;��G;enH;ߡH;�H;��H;��H;��H;��H;��H;X�H;��H;X�H;��H;��H;��H;��H;��H;�H;ܡH;enH;��G;6UF;*�B;I�:;��*;d�;	��:0����$��ͻ*�E�bx�� �!\��R���.��C�9�Gl��WD���
�ѕ3�bXi��������¿Epѿ      ��"$������꿱�ſ�ޞ�(3s��2�@����� j���{HͽƸ����'�@<ͼh�n�R���Q^��,.����:�W;�S%;|o8;��A;uDF;�H;��H;�H;	�H;a�H;V�H;a�H;��H;�H;��H;F�H;��H;�H;��H;`�H;X�H;a�H;�H;�H;��H;�H;uDF;��A;{o8;�S%;�W;���:�,.�Q^�Q���i�n�@<ͼ��'�Ƹ��{Hͽ�� j���@����2�(3s��ޞ���ſ������"$�      "$�������忉�����!cm�W�-�����Rh��Xde�#-�٪ɽ�v��'�$�}�ɼpmj�%����X����(Ɔ:�x;]�%;J�8;�B;�RF;H;E�H;i�H;�H;��H;[�H;R�H;��H;��H;��H;A�H;��H;��H;��H;P�H;[�H;��H;�H;f�H;E�H;H;�RF;�B;G�8;c�%;�x;(Ɔ: ���X�$���pmj�}�ɼ'�$��v��٪ɽ#-�Xde�Rh������W�-�!cm��������忞����      ��������� �ԿNw�����<�\�"����l��[0X�����;����w����������]��黟F����0ʒ:�;U�';׏9;9pB;�zF;�!H;��H;L�H;4�H;��H;b�H;V�H;��H;��H;��H;-�H;��H;��H;��H;U�H;`�H;��H;1�H;I�H;��H;�!H;�zF;9pB;ԏ9;X�';�;0ʒ:��깟F��黣�]����������w��;�����[0X�l�����"�<�\����Nw�� �Կ��𿞏�      ����� �Կp���ޞ�bF�i�C�.E�$�;�I���D���"��g�c�{��֯���J��ѻ��)�P{K�b��:7�
;	N*;��:;�C;#�F;�8H;k�H;��H;��H;��H;[�H;V�H;��H;��H;��H;�H;��H;��H;��H;U�H;[�H;��H;��H;��H;m�H;�8H;$�F;�C;��:;N*;7�
;d��:p{K���)��ѻ��J��֯�{�g�c�"�����D��I��$�;.E�i�C�bF��ޞ�p�� �Կ��      ��ſ���Nw���ޞ�����A�W�6�%�����iɰ��|x�g{+�ӱ����J��  �ʶ��P�1�����*��$
9<�:̅;-�-;��<;��C;�G;�TH;c�H;�H;�H;��H;q�H;O�H;��H;��H;��H;�H;��H;��H;��H;N�H;r�H;��H;�H;�H;c�H;�TH;�G;��C;��<;.�-;̅;@�:�$
9�*����P�1�ʶ���  ��J���ӱ�g{+��|x�iɰ�����6�%�A�W������ޞ�Nw�����      �ޞ�������bF�A�W�X�-����AKɾ�G����O����ƽȸ��΄-���ۼㄼ*4�ǐ��ζ�0^:C��:�;Ɩ1;d>;��D;�\G;\sH;��H;��H;z�H;<�H;��H;E�H;��H;��H;��H;��H;��H;��H;��H;E�H;��H;<�H;w�H;~�H;��H;[sH;�\G;��D;d>;Ɩ1;�;E��:(^:�ζ�ǐ�*4�ㄼ��ۼ΄-�ȸ��ƽ�����O��G��AKɾ���X�-�A�W�bF�������      (3s�!cm�<�\�j�C�7�%�����TҾl�� j��C(����_P����[�{������Y�#��9X���<��k:���:� ;�5;`R@;}uE;�G;J�H;]�H;��H;�H;_�H;��H;@�H;�H;��H;r�H;��H;r�H;��H;�H;A�H;��H;_�H;�H;��H;_�H;I�H;�G;yuE;\R@;�5;� ;���:�k:��<�6X�#����Y����{���[�_P����콬C(� j�l���TҾ���7�%�j�C�<�\�!cm�      �2�W�-�"�.E�����AKɾl����s�:�5���w㻽�v��	z0��;��+���*����6�@5S��M�:|�	;��(;5�9;�/B;�DF;kH;�H;��H;��H;��H;��H;��H;*�H;N�H;\�H;W�H;v�H;W�H;\�H;N�H;,�H;��H;��H;��H;��H;��H;�H;kH;�DF;�/B;5�9;��(;~�	;�M�:@5S�6�����*��+���;�	z0��v��w㻽��:�5���s�l��AKɾ����.E�"�W�-�      @����������$�;iɰ��G�� j�:�5��	�ЪɽZ����J�r���沼��]�����	x�����n:��:�v;��/;�-=;��C;^�F;6IH;��H;;�H;��H;8�H;��H;��H;�H;"�H;)�H;/�H;@�H;0�H;)�H;"�H;�H;��H;��H;7�H;��H;;�H;��H;7IH;[�F;��C;�-=;��/;�v;	��:�n:����	x������]��沼r���J�Z���Ѫɽ�	�:�5� j��G��jɰ�$�;��徹���      ��Rh��l���I���|x���O��C(���Ѫɽ����RDX�G��$<ͼㄼ�X!��s���W��rK����:�y;0�#;"I6;OR@;�PE;��G;��H;��H;H�H;�H;��H;��H;��H;��H;�H;��H;��H;��H;��H;��H;�H;��H;��H;��H;��H;�H;H�H;��H;��H;��G;�PE;NR@;$I6;0�#;�y;���:�rK��W��s���X!�ㄼ$<ͼG��RDX�����Ѫɽ���C(���O��|x��I��l��Rh��       j�Xde�[0X��D�g{+�������w㻽Z���RDX������ۼȾ��}�;�2>ۻ�X���y��?":��:��;��-;��;;�B;�zF;�H;��H;��H;:�H; �H;�H;�H;��H;��H;��H;��H;��H;��H;��H;��H;��H;��H;��H;�H;�H;��H;;�H;��H;��H;�H;�zF;�B;��;;��-;��;��:�?":��y��X�2>ۻ|�;�Ⱦ����ۼ���RDX�Z���w㻽��콃��g{+��D�[0X�Xde�      ��#-������ӱ�ƽ_P���v���J�G����ۼ	��Z�J�����p+��.rѺ�+
9,N�:�;� $;%�5;�?;��D;y\G;fH;
�H;��H;��H;��H;8�H;�H;p�H;��H;x�H;q�H;~�H;V�H;�H;u�H;{�H;��H;r�H;�H;8�H;��H;��H;��H;�H;fH;y\G;��D;�?;%�5;� $;�;4N�:`+
9,rѺp+������Z�J�	����ۼG���J��v��_P��ƽӱ轄����#-�      {Hͽ٪ɽ�;��"����ȸ����[�	z0�r��$<ͼǾ��Z�J����j��M*���V��:�b�:p�;�/;�L<;*C;GmF;��G;"�H;#�H;)�H;)�H;^�H;o�H;�H;D�H;O�H;:�H;5�H;$�H;�H;$�H;5�H;<�H;O�H;F�H;�H;p�H;^�H;)�H;&�H;&�H;�H;��G;CmF;*C;�L<;
�/;p�;�b�:T��:��M*��j����Z�J�Ǿ��$<ͼr��	z0���[�ȸ����"���;��٪ɽ      Ƹ���v����w�g�c��J�΄-�{��;缃沼ㄼ|�;������j��z5��깸?Q:���:�i;N*;��8;��@;�PE;�uG;YiH;��H;��H;.�H;>�H;��H;��H;�H;�H;��H;��H;��H;��H;��H;��H;��H;��H;��H;�H;�H;��H;��H;@�H;-�H;��H;��H;ViH;�uG;�PE;��@;��8;N*;�i;���:�?Q:��y5��j������|�;�ㄼ�沼�;�{�΄-��J�g�c���w��v��      ��'�'�$����{��  ���ۼ����+����]��X!�3>ۻr+��O*� �까�>:#��:2�;P�%;�5;��>;�(D;+�F;�!H;P�H;p�H;�H;��H;��H;	�H;��H;��H;��H;��H;��H;��H;o�H;��H;p�H;��H;��H;��H;��H;��H;��H;�H;��H;��H;�H;p�H;M�H;�!H;+�F;�(D;��>;�5;V�%;/�;'��:��>: ��O*�r+��2>ۻ�X!���]��+�������ۼ�  �{����(�$�      ?<ͼ|�ɼ�����֯�ʶ��ㄼ��Y��*�����s���X�.rѺ���?Q:)��:��
;l�#;��3;�c=; $C;BDF; �G;/�H;�H;.�H;V�H;�H;w�H;D�H;��H;��H;��H;X�H;q�H;-�H;�H;*�H;�H;-�H;q�H;X�H;��H;��H;��H;@�H;w�H;�H;Z�H;.�H; �H;-�H;"�G;?DF; $C;�c=;��3;l�#;��
;+��:�?Q:��.rѺ�X��s������*���Y�ㄼʶ���֯�����}�ɼ      i�n�nmj���]���J�Q�1�*4� ������	x��W���y�P+
9N��:���:2�;h�#;t�2;�<;�pB;G�E;΍G;�eH;�H;T�H;��H;�H;��H;��H;\�H;j�H;Z�H;1�H;�H;��H;��H;��H;��H;��H;��H;��H;�H;4�H;[�H;j�H;[�H;��H;��H;�H;��H;Q�H;�H;�eH;΍G;H�E;�pB;�<;t�2;h�#;2�;���:N��:`+
9��y��W��	x���� ��)4�Q�1���J���]�pmj�      U���&������ѻ���ǐ�<X�6�����rK��?":,N�:�b�:|i;S�%;|�3;�<;a0B;��E;�\G;�HH;e�H;��H;}�H;�H;W�H;`�H;��H;9�H;<�H;�H;��H;��H;��H;v�H;u�H;T�H;u�H;v�H;��H;��H;��H;	�H;<�H;8�H;��H;^�H;Z�H;�H;{�H;��H;e�H;�HH;�\G;E;c0B;�<;~�3;S�%;�i;�b�:,N�:�?":�rK����6�<X�ǐ�����ѻ��*���      Q^��X��F���)��*��ζ���<��6S��n:z��:��:�;l�;N*;�5;�c=;�pB;��E;�JG;s8H;��H;��H;3�H;M�H;��H;�H;��H;�H;�H;��H;��H;��H;z�H;'�H;�H;�H;��H;�H;�H;)�H;y�H;��H;��H;��H;�H;�H;��H;�H;��H;I�H;0�H;��H;��H;t8H;�JG;E;�pB;�c=;�5;N*;n�;�;��:z��:�n:@6S���<��ζ��*���)��F��X�      �,.�̪���김{K��$
9^:��k:�M�:���:�y;��;� $;�/;��8;��>;$C;D�E;�\G;p8H;�H;'�H;B�H;��H;Y�H;��H;w�H;��H;��H;��H;��H;a�H;7�H;�H;��H;��H;��H;��H;��H;��H;��H;�H;8�H;a�H;��H;��H;��H;��H;y�H;��H;T�H;��H;B�H;%�H;�H;p8H;�\G;D�E;$C;��>;��8;�/;� $;��;�y;���:�M�:��k:$^: %
9�{K������      ���:HƆ:0ʒ:P��:*�:I��:���:u�	;�v;.�#;�-;�5;�L<;��@;�(D;>DF;΍G;�HH;��H;%�H;��H;o�H;��H;��H;F�H;��H;��H;��H;��H;H�H;,�H;��H;��H;��H;Y�H;I�H;K�H;K�H;Y�H;��H;��H;��H;,�H;E�H;��H;��H;��H;��H;F�H;�H;��H;o�H;��H;(�H;��H;�HH;̍G;?DF;�(D;��@;�L<; �5;�-;-�#;�v;w�	;���:O��:,�:V��:6ʒ:$Ɔ:      �W;�x;&�;,�
;̅;�; � ;��(;��/; I6;��;;�?;%C;�PE;+�F;�G;�eH;d�H;��H;D�H;n�H;��H;V�H;�H;��H;��H;��H;��H;�H;��H;��H;n�H;E�H;4�H;��H;��H;��H;��H;��H;4�H;B�H;n�H;��H;��H;�H;��H;��H;��H;��H;�H;S�H;��H;m�H;E�H;��H;e�H;�eH;�G;.�F;�PE;'C;�?;��;; I6;��/;��(;"� ;�;��;.�
;(�;�x;      �S%;^�%;T�'; N*;&�-;1;�5;2�9;�-=;KR@;�B;��D;CmF;�uG;�!H;+�H;�H;��H;1�H;��H;��H;W�H;*�H;��H;��H;��H;a�H;�H;��H;��H;O�H;�H;��H;��H;��H;��H;�H;��H;��H;��H;��H;�H;N�H;��H;��H;�H;^�H;��H;��H;��H;)�H;W�H;��H;��H;3�H;��H;�H;+�H;�!H;�uG;CmF;��D;�B;JR@;�-=;2�9;�5;Ŗ1;-�-; N*;T�';R�%;      �o8;W�8;ޏ9;��:;��<;
d>;cR@;�/B;��C;�PE;�zF;y\G;��G;ViH;M�H; �H;T�H;~�H;L�H;V�H;�H;�H;��H;��H;��H;s�H;�H;��H;��H;=�H;��H;��H;��H;[�H;U�H;J�H;%�H;J�H;X�H;[�H;��H;��H;��H;9�H;��H;��H;�H;u�H;��H;��H;��H;�H;|�H;V�H;J�H;��H;S�H;�H;N�H;WiH;��G;y\G;�zF;�PE;��C;�/B;bR@;d>;��<;��:;ޏ9;G�8;      ��A;�B;"pB;�C;��C;��D;yuE;�DF;X�F;��G;�H;fH;�H;��H;q�H;/�H;��H; �H;��H;��H;H�H;��H;��H;��H;T�H;��H;��H;��H;3�H;��H;��H;p�H;?�H;�H;��H;��H;��H;��H;��H;�H;<�H;q�H;��H;��H;0�H;��H;��H;��H;T�H;��H;��H;��H;E�H;��H;��H;#�H;��H;.�H;q�H;��H;�H;fH;�H;��G;Y�F;�DF;yuE;��D;��C;�C;$pB;�B;      DF;�RF;�zF;�F;�G;�\G;�G;bH;0IH;��H;��H;�H; �H;��H;�H;T�H;�H;W�H; �H;u�H;��H;��H;��H;s�H;��H;��H;��H;,�H;��H;��H;M�H;�H;��H;��H;��H;��H;��H;��H;��H;��H;��H;�H;K�H;��H;��H;,�H;��H;��H;��H;o�H;��H;��H;��H;v�H; �H;Y�H;�H;T�H;�H;��H;"�H;
�H;��H;��H;1IH;dH;�G;�\G;�G;�F;�zF;�RF;      H;H;�!H;�8H;�TH;[sH;M�H;�H;��H;��H;��H;��H;$�H;,�H;��H;�H;��H;[�H;��H;��H;��H;��H;^�H;�H;��H;��H;�H;��H;{�H;J�H;�H;��H;��H;{�H;_�H;<�H;P�H;<�H;^�H;z�H;��H;��H;�H;H�H;z�H;��H;�H;��H;��H;�H;^�H;��H;��H;��H;��H;^�H;��H;�H;��H;-�H;&�H;��H;��H;��H;��H;�H;L�H;XsH;�TH;�8H;�!H;H;      ��H;H�H;��H;d�H;c�H;��H;_�H;��H;:�H;G�H;=�H;��H;)�H;A�H;��H;v�H;��H;��H;�H;��H;��H;��H;�H;��H;��H;,�H;��H;��H;:�H;��H;��H;}�H;W�H;$�H;�H;�H;�H;�H;�H;$�H;T�H;}�H;��H;��H;9�H;��H;��H;,�H;��H;��H;�H;��H;��H;��H;�H;��H;��H;w�H;��H;@�H;'�H;��H;=�H;H�H;=�H;��H;_�H;��H;o�H;d�H;��H;S�H;      �H;j�H;H�H;��H;�H;|�H;��H;��H;��H;�H;��H;��H;]�H;��H;�H;C�H;_�H;6�H;�H;��H;��H;�H;��H;��H;,�H;��H;x�H;:�H;��H;��H;p�H;8�H;�H;��H;��H;��H;��H;��H;��H;��H; �H;9�H;o�H;��H;��H;<�H;x�H;��H;/�H;��H;��H;�H;��H;��H;�H;8�H;^�H;D�H;	�H;��H;^�H;��H;��H;�H;��H;��H;��H;|�H;�H;��H;H�H;`�H;      �H;!�H;;�H;��H;�H;z�H;�H;��H;>�H;��H;�H;B�H;q�H;��H;��H;��H;m�H;8�H;��H;��H;E�H;��H;��H;>�H;��H;��H;D�H;��H;��H;e�H;5�H;��H;��H;��H;��H;��H;z�H;��H;��H;��H;��H;��H;6�H;e�H;��H;��H;F�H;��H;��H;;�H;��H;��H;E�H;��H;��H;9�H;l�H;��H;��H;��H;t�H;C�H;�H;��H;?�H;��H;�H;{�H;�H;��H;6�H;�H;      b�H;��H;��H;��H;�H;6�H;e�H;��H;��H;��H;	�H;�H;�H;	�H;��H;��H;_�H;�H;��H;d�H;.�H;��H;L�H;��H;��H;K�H;��H;��H;l�H;6�H;��H;��H;��H;y�H;W�H;a�H;a�H;a�H;W�H;z�H;��H;��H;��H;5�H;m�H;��H;��H;M�H;��H;��H;I�H;��H;,�H;d�H;��H;�H;_�H;��H;��H;�H;�H;�H;�H;��H;��H;��H;e�H;8�H;�H;��H;��H;��H;      `�H;i�H;d�H;`�H;t�H;��H;��H;��H;��H;��H;��H;z�H;F�H;�H;��H;��H;9�H;��H;��H;>�H;��H;q�H;�H;��H;k�H;�H;��H;}�H;5�H;��H;��H;��H;z�H;H�H;3�H;0�H;4�H;0�H;3�H;H�H;v�H;��H;��H;��H;6�H;~�H;��H;�H;p�H;��H;�H;q�H;��H;>�H;��H;��H;9�H;��H;��H;�H;G�H;z�H;��H;��H;��H;��H;��H;��H;r�H;_�H;d�H;d�H;      `�H;^�H;\�H;^�H;W�H;A�H;@�H;3�H;	�H;��H;��H;��H;R�H;��H;��H;\�H;�H;��H;}�H;�H;��H;B�H;��H;��H;6�H;��H;��H;X�H;�H;��H;��H;|�H;5�H;*�H;*�H;�H;��H;�H;*�H;*�H;3�H;}�H;��H;��H;�H;Z�H;��H;��H;9�H;��H;��H;D�H;��H;�H;}�H;��H;�H;_�H;��H;��H;T�H;��H;��H;��H;	�H;3�H;A�H;D�H;R�H;^�H;\�H;Y�H;      ��H;��H;��H;��H;��H;�H;��H;V�H;%�H;�H;��H;��H;=�H;��H;��H;x�H; �H;��H;)�H;��H;��H;2�H;��H;\�H;�H;��H;t�H;!�H;��H;��H;y�H;H�H;&�H;�H;�H;��H;��H;��H;�H;�H;%�H;L�H;y�H;��H;��H;#�H;t�H;��H;�H;\�H;��H;3�H;��H;��H;)�H;��H;��H;{�H;��H;��H;?�H;��H;��H;�H;&�H;W�H;��H;��H;��H;��H;��H;��H;      �H;�H;��H;��H;��H;��H;��H;g�H;0�H;��H;��H;��H;=�H;��H;��H;5�H;��H;s�H;�H;��H;]�H;��H;��H;V�H;��H;��H;[�H;�H;��H;��H;W�H;5�H;)�H;�H;��H;��H;��H;��H;��H;�H;&�H;8�H;W�H;��H;��H;�H;[�H;��H;��H;U�H;��H;��H;Z�H;��H;�H;u�H;��H;6�H;��H;��H;?�H;��H;��H;��H;0�H;e�H;��H;��H;��H;��H;��H;�H;      ��H;��H;��H;��H;��H;��H;x�H;a�H;:�H;��H;��H;��H;)�H;��H;t�H;�H;��H;p�H;�H;��H;N�H;��H;��H;K�H;��H;��H;8�H;�H;��H;��H;b�H;4�H;�H;��H;��H;��H;��H;��H;��H;��H;�H;7�H;b�H;��H;��H;�H;9�H;��H;��H;K�H;��H;��H;L�H;��H;�H;r�H;��H;�H;t�H;��H;+�H;��H;��H;��H;;�H;`�H;y�H;��H;��H;��H;��H;��H;      B�H;H�H;;�H;�H;�H;��H;��H;}�H;G�H;��H;��H;b�H;�H;��H;��H;1�H;��H;J�H;��H;��H;I�H;��H;z�H;%�H;��H;��H;J�H;�H;��H;|�H;b�H;:�H;��H;��H;��H;��H;��H;��H;��H;��H;��H;;�H;b�H;}�H;��H;�H;J�H;��H;��H;"�H;z�H;��H;H�H;��H;��H;L�H;��H;1�H;��H;��H;�H;b�H;��H;��H;H�H;|�H;��H;��H;�H;�H;:�H;A�H;      ��H;��H;��H;��H;��H;��H;y�H;a�H;:�H;��H;��H;��H;+�H;��H;v�H;�H;��H;p�H;�H;��H;O�H;��H;��H;M�H;��H;��H;;�H;�H;��H;��H;b�H;4�H;�H;��H;��H;��H;��H;��H;��H;��H;�H;7�H;b�H;��H;��H;�H;8�H;��H;��H;H�H;��H;��H;L�H;��H;�H;r�H;��H;�H;t�H;��H;)�H;��H;��H;��H;:�H;`�H;x�H;��H;��H;��H;��H;��H;      �H;�H;��H;��H;��H;��H;��H;g�H;0�H;��H;��H;��H;?�H;��H;��H;6�H;��H;s�H;�H;��H;`�H;��H;��H;V�H;��H;��H;\�H;�H;��H;��H;W�H;5�H;)�H;�H;��H;��H;��H;��H;��H;�H;&�H;:�H;W�H;��H;��H;�H;Z�H;��H;��H;T�H;��H;��H;Y�H;��H;�H;u�H;��H;5�H;��H;��H;=�H;��H;��H;��H;0�H;e�H;��H;��H;��H;��H;��H;�H;      ��H;��H;��H;��H;��H;��H;��H;V�H;%�H;�H;��H;��H;?�H;��H;��H;{�H; �H;��H;)�H;��H;��H;3�H;��H;]�H;�H;��H;t�H;#�H;��H;��H;y�H;I�H;&�H;�H;�H;��H;��H;��H;�H;�H;%�H;L�H;y�H;��H;��H;!�H;t�H;��H;�H;[�H;��H;2�H;��H;��H;)�H;��H;��H;x�H;��H;��H;=�H;��H;��H;�H;&�H;V�H;��H;��H;��H;��H;��H;��H;      d�H;`�H;]�H;`�H;V�H;@�H;@�H;2�H;	�H;��H;��H;��H;T�H;��H;��H;_�H;�H;��H;}�H;�H;��H;D�H;��H;��H;9�H;��H;��H;Z�H;�H;��H;��H;|�H;4�H;)�H;*�H;�H;��H;�H;*�H;)�H;3�H;~�H;��H;��H;�H;X�H;��H;��H;6�H;��H;��H;B�H;��H;�H;}�H;��H;�H;\�H;��H;��H;Q�H;��H;��H;��H;	�H;0�H;>�H;B�H;N�H;^�H;Z�H;^�H;      `�H;i�H;g�H;_�H;r�H;��H;��H;��H;��H;��H;��H;{�H;G�H;�H;��H;��H;;�H;��H;��H;?�H;��H;q�H;�H;��H;p�H;�H;��H;~�H;5�H;��H;��H;��H;y�H;H�H;3�H;0�H;4�H;0�H;3�H;H�H;v�H;��H;��H;��H;6�H;}�H;��H;	�H;k�H;��H;�H;q�H;��H;>�H;��H;��H;8�H;��H;��H;�H;F�H;x�H;��H;��H;��H;��H;��H;��H;p�H;]�H;g�H;f�H;      b�H;��H;��H;��H;�H;8�H;e�H;��H;��H;��H;�H;�H;�H;�H;��H;��H;_�H;�H;��H;d�H;0�H;��H;L�H;��H;��H;N�H;��H;��H;l�H;6�H;��H;��H;��H;z�H;W�H;a�H;a�H;a�H;W�H;y�H;��H;��H;��H;5�H;m�H;��H;��H;J�H;��H;��H;I�H;��H;,�H;d�H;��H;�H;^�H;��H;��H;	�H;�H;�H;�H;��H;��H;��H;e�H;8�H;�H;��H;��H;��H;      �H;#�H;8�H;��H;�H;x�H;�H;��H;?�H;��H;�H;C�H;t�H;��H;��H;��H;m�H;8�H;��H;��H;J�H;��H;��H;>�H;��H;��H;F�H;��H;��H;f�H;6�H;��H;��H;��H;��H;��H;z�H;��H;��H;��H;��H;��H;5�H;c�H;��H;��H;C�H;��H;��H;=�H;��H;��H;C�H;��H;��H;9�H;l�H;��H;��H;��H;q�H;B�H;�H;��H;?�H;��H;�H;z�H;�H;��H;9�H;!�H;      �H;f�H;L�H;��H;�H;z�H;��H; �H;��H;�H;��H;��H;^�H;��H;	�H;D�H;_�H;6�H;�H;��H;��H;�H;��H;��H;/�H;��H;w�H;<�H;��H;��H;o�H;6�H;�H;��H;��H;��H;��H;��H;��H;��H;�H;9�H;p�H;��H;��H;:�H;z�H;��H;,�H;��H;��H;�H;��H;��H;�H;8�H;^�H;D�H;�H;��H;]�H;��H;��H;�H;��H;��H;��H;z�H;�H;��H;L�H;f�H;      ��H;F�H;��H;d�H;b�H;��H;_�H;��H;;�H;H�H;>�H;��H;'�H;A�H;��H;w�H;��H;��H;�H;��H;��H;��H;�H;��H;��H;,�H;��H;��H;<�H;��H;��H;}�H;U�H;#�H;�H;�H;�H;�H;�H;$�H;U�H;~�H;��H;��H;9�H;��H;��H;,�H;��H;��H;�H;��H;��H;��H;�H;��H;��H;w�H;��H;@�H;)�H;��H;;�H;G�H;;�H;��H;_�H;��H;l�H;d�H;��H;S�H;      �H;H;�!H;�8H;�TH;XsH;J�H;�H;��H;��H;��H;��H;'�H;-�H;��H;�H;��H;]�H;��H;��H;��H;��H;^�H;�H;��H;��H;�H;��H;{�H;J�H;�H;��H;��H;z�H;^�H;<�H;P�H;;�H;_�H;z�H;��H;��H;�H;H�H;z�H;��H;�H;��H;��H;�H;^�H;��H;��H;��H;��H;]�H;��H;�H;��H;,�H;$�H;��H;��H;��H;��H;�H;J�H;UsH;�TH;�8H;�!H;H;      �DF;�RF;�zF;!�F;�G;�\G;�G;dH;0IH;��H;��H;�H;"�H;��H;�H;V�H;�H;W�H; �H;v�H;��H;��H;��H;r�H;��H;��H;��H;,�H;��H;��H;K�H;�H;��H;��H;��H;��H;��H;��H;��H;��H;��H;�H;M�H;��H;��H;,�H;��H;��H;��H;p�H;��H;��H;��H;u�H; �H;Y�H;�H;T�H;�H;��H; �H;�H;��H;��H;/IH;aH;�G;�\G;�G; �F;�zF;�RF;      ��A;�B;"pB;�C;��C;��D;yuE;�DF;Y�F;��G;�H;fH;�H;��H;q�H;/�H;��H; �H;��H;��H;I�H;��H;��H;��H;T�H;��H;��H;��H;3�H;��H;��H;p�H;=�H;�H;��H;��H;��H;��H;��H;�H;=�H;r�H;��H;��H;0�H;��H;��H;��H;T�H;��H;��H;��H;E�H;��H;��H;#�H;��H;/�H;q�H;��H;�H;fH;�H;��G;X�F;�DF;yuE;��D;��C;�C;$pB;�B;      �o8;U�8;�9;��:;��<;d>;_R@;�/B;��C;�PE;�zF;z\G;��G;WiH;N�H;�H;U�H;~�H;J�H;V�H;��H;�H;��H;��H;��H;s�H;�H;��H;��H;=�H;��H;��H;��H;Y�H;T�H;J�H;%�H;J�H;V�H;[�H;��H;��H;��H;:�H;��H;��H;�H;u�H;��H;��H;��H;�H;|�H;V�H;L�H;�H;Q�H; �H;M�H;ViH;��G;y\G;�zF;�PE;��C;�/B;_R@;d>;��<;��:;�9;G�8;      �S%;l�%;b�';N*;"�-;Ȗ1;�5;2�9;�-=;KR@;�B;��D;BmF;�uG;�!H;-�H;�H;��H;3�H;��H;��H;W�H;*�H;��H;��H;��H;a�H;�H;��H;��H;N�H;�H;��H;��H;��H;��H;�H;��H;��H;��H;��H;�H;O�H;��H;��H;�H;`�H;��H;��H;��H;)�H;W�H;��H;��H;1�H;��H;�H;+�H;�!H;�uG;BmF;��D;�B;HR@;�-=;1�9;�5;Ȗ1;)�-;N*;Y�';\�%;      �W;�x;&�;.�
;ȅ;�;"� ;��(;��/; I6;��;;�?;'C;�PE;-�F;�G;�eH;d�H;��H;D�H;o�H;��H;V�H;�H;��H;��H;��H;��H;�H;��H;��H;n�H;D�H;4�H;��H;��H;��H;��H;��H;4�H;D�H;n�H;��H;��H;�H;��H;��H;��H;��H;�H;S�H;��H;m�H;E�H;��H;e�H;�eH;�G;-�F;�PE;%C;�?;��;; I6;��/;��(; � ;�;ޅ;,�
;(�;�x;      ���:@Ɔ:8ʒ:T��:*�:7��:���:z�	;�v;,�#;�-; �5;�L<;��@;�(D;?DF;΍G;�HH;��H;'�H;��H;o�H;��H;��H;F�H;��H;��H;��H;��H;H�H;,�H;��H;��H;��H;Y�H;I�H;K�H;I�H;Y�H;��H;��H;��H;,�H;E�H;��H;��H;��H;��H;F�H;�H;��H;o�H;��H;'�H;��H;�HH;̍G;>DF;�(D;��@;�L<;�5;�-;*�#;�v;x�	;���:K��:2�:T��::ʒ:&Ɔ:      �,.������김{K��$
9^:��k:�M�:���:�y;��;� $;�/;��8;��>;$C;E�E;�\G;p8H;�H;*�H;B�H;��H;X�H;��H;y�H;��H;��H;��H;��H;a�H;8�H;�H;��H;��H;��H;��H;��H;��H;��H;�H;8�H;a�H;��H;��H;��H;��H;y�H;��H;T�H;��H;B�H;$�H;�H;p8H;�\G;B�E;$C;��>;��8;�/;� $;��;�y;���:�M�:��k: ^: %
9�{K������      Q^��X��F���)��*��ζ���<��6S��n:z��:��:�;n�;N*;	�5;�c=;�pB;E;�JG;s8H;��H;��H;4�H;M�H;��H;�H;��H;�H;�H;��H;��H;��H;|�H;)�H;�H;�H;��H;�H;�H;'�H;y�H;��H;��H;��H;�H;�H;��H;�H;��H;I�H;.�H;��H;��H;t8H;�JG;��E;�pB;�c=;	�5;N*;l�;�;��:z��:�n:�6S���<��ζ��*���)��F��X�      T���&������ѻ���ǐ�<X�6�����rK��?":,N�:�b�:i;S�%;~�3;�<;a0B;E;�\G;�HH;e�H;��H;�H;�H;Y�H;`�H;��H;<�H;=�H;	�H;��H;��H;��H;v�H;u�H;T�H;u�H;v�H;��H;��H;��H;�H;;�H;6�H;��H;]�H;Z�H;�H;x�H;��H;e�H;�HH;�\G;��E;b0B;�<;|�3;S�%;~i;�b�:*N�:�?":�rK����6�=X�
ǐ�����ѻ��*���      i�n�nmj���]���J�R�1�*4�!������	x��W���y�`+
9N��:���:2�;h�#;v�2;�<;�pB;G�E;ύG;�eH;�H;U�H;��H;�H;��H;��H;^�H;m�H;[�H;4�H;�H;��H;��H;��H;��H;��H;��H;��H;�H;2�H;Z�H;i�H;X�H;��H;��H;�H;��H;P�H;�H;�eH;̍G;H�E;�pB;�<;t�2;h�#;2�;���:N��:P+
9��y��W��	x����!��*4�Q�1���J���]�pmj�      ?<ͼ|�ɼ�����֯�ʶ��ㄼ��Y��*�����s���X�.rѺ���?Q:+��:��
;n�#;��3;�c=; $C;BDF;"�G;/�H;�H;.�H;X�H;�H;w�H;F�H;��H;��H;��H;Z�H;q�H;-�H;�H;*�H;�H;-�H;q�H;W�H;��H;��H;��H;@�H;w�H;�H;X�H;.�H; �H;+�H; �G;?DF; $C;�c=;��3;k�#;��
;)��:�?Q:��.rѺ�X��s�� ����*���Y�ㄼʶ���֯�����}�ɼ      ��'�'�$����{��  ���ۼ����+����]��X!�2>ۻr+��O*� �까�>:'��:2�;S�%;�5;��>;�(D;+�F;�!H;Q�H;p�H;�H;��H;��H;�H;��H;��H;��H;��H;��H;��H;o�H;��H;o�H;��H;��H;��H;��H;��H;��H;�H;��H;��H;�H;p�H;K�H;�!H;+�F;�(D;��>;�5;S�%;1�;#��:��>: ��O*�r+��3>ۻ�X!���]��+�������ۼ�  �{����(�$�      Ƹ���v����w�g�c��J�΄-�{��;缃沼ㄼ|�;������j��z5��깸?Q:���:�i;N*;��8;��@;�PE;�uG;YiH;��H;��H;.�H;@�H;��H;��H;�H;�H;��H;��H;��H;��H;��H;��H;��H;��H;��H;�H;�H;��H;��H;>�H;-�H;��H;��H;ViH;�uG;�PE;��@;��8;N*;�i;���:�?Q:��z5��j������|�;�ㄼ�沼�;�{�΄-��J�g�c���w��v��      {Hͽ٪ɽ�;��"����ȸ����[�	z0�r��$<ͼǾ��Z�J����j��M*���V��:�b�:p�;
�/;�L<;*C;GmF;��G;�H;&�H;)�H;)�H;a�H;p�H;�H;D�H;O�H;<�H;5�H;$�H;�H;$�H;5�H;:�H;N�H;D�H;�H;o�H;[�H;)�H;&�H;&�H;"�H;��G;CmF;*C;�L<;
�/;p�;�b�:T��:��M*��j����Z�J�Ǿ��$<ͼr��	z0���[�Ǹ����"���;��٪ɽ      ��#-������ӱ�ƽ_P���v���J�G����ۼ	��Z�J�����p+��,rѺ�+
92N�:�;� $;#�5;�?;��D;z\G;fH;�H;��H;��H;��H;8�H;�H;p�H;��H;|�H;u�H;�H;V�H;�H;q�H;x�H;��H;q�H;�H;8�H;��H;��H;��H;�H;fH;w\G;��D;�?;%�5;� $;�;2N�:`+
92rѺp+������Z�J�	����ۼG���J��v��_P��ƽӱ轄����#-�       j�Xde�[0X��D�g{+�������w㻽Z���RDX������ۼȾ��}�;�2>ۻ�X���y��?":��:��;�-;��;;�B;�zF;�H;��H;��H;;�H;�H;�H;�H;��H;��H;��H;��H;��H;��H;��H;��H;��H;��H;��H;�H;�H;��H;:�H;��H;��H;�H;�zF;�B;��;;�-;��;��:�?":��y��X�2>ۻ|�;�Ⱦ����ۼ���RDX�Z���w㻽��콃��g{+��D�[0X�Xde�      ��Rh��l���I���|x���O��C(���Ѫɽ����RDX�G��$<ͼㄼ�X!��s���W��rK����:�y;.�#;$I6;OR@;�PE;��G;��H;��H;H�H;�H;��H;��H;��H;��H;�H;��H;��H;��H;��H;��H;�H;��H;��H;��H;��H;�H;H�H;��H;��H;��G;�PE;NR@;"I6;0�#;�y;���:�rK��W��s���X!�ㄼ$<ͼG��RDX�����Ѫɽ���C(���O��|x��I��l��Rh��      @����������$�;iɰ��G�� j�:�5��	�ѪɽZ����J�r���沼��]�����	x�����n:��:�v;��/;�-=;��C;[�F;7IH;��H;;�H;��H;7�H;��H;��H;�H;"�H;)�H;0�H;@�H;/�H;)�H;"�H; �H;��H;��H;7�H;��H;;�H;��H;6IH;^�F;��C;�-=;��/;�v;	��:�n:����	x������]��沼r���J�Z���Ъɽ�	�:�5� j��G��jɰ�$�;��徹���      �2�W�-�"�.E�����AKɾl����s�:�5���w㻽�v��	z0��;��+���*����6�@5S��M�:{�	;��(;5�9;�/B;�DF;kH;�H;��H;��H;��H;��H;��H;-�H;O�H;]�H;W�H;v�H;Y�H;\�H;O�H;)�H;��H;��H;��H;��H;��H;�H;iH;�DF;�/B;5�9;��(;~�	;�M�:@5S�6�����*��+���;�	z0��v��w㻽��:�5���s�l��AKɾ����.E�"�W�-�      (3s�!cm�<�\�j�C�7�%�����TҾl�� j��C(����_P����[�{������Y�"��8X���<��k:���:� ;�5;`R@;yuE;�G;J�H;_�H;��H;�H;_�H;��H;B�H;��H;��H;r�H;��H;r�H;��H;�H;>�H;��H;_�H;�H;��H;]�H;I�H;�G;}uE;]R@;�5;� ;���:�k:��<�6X�$����Y����{���[�_P����콬C(� j�l���TҾ���7�%�j�C�<�\�!cm�      �ޞ�������bF�A�W�X�-����AKɾ�G����O����ƽȸ��΄-���ۼㄼ*4�ǐ��ζ�(^:=��:�;Ŗ1;d>;��D;�\G;\sH;��H;��H;z�H;<�H;��H;G�H;��H;��H;��H;��H;��H;��H;��H;D�H;��H;<�H;w�H;~�H;��H;[sH;�\G;��D;d>;Ɩ1;�;E��:(^:�ζ�ǐ�*4�ㄼ��ۼ΄-�ȸ��ƽ�����O��G��AKɾ���X�-�A�W�bF�������      ��ſ���Nw���ޞ�����A�W�6�%�����iɰ��|x�g{+�ӱ����J��  �ʶ��P�1�����*��$
9:�:̅;,�-;��<;��C;�G;�TH;c�H;�H;�H;��H;q�H;O�H;��H;��H;��H;�H;��H;��H;��H;N�H;q�H;��H;�H;�H;c�H;�TH;�G;��C;��<;0�-;̅;@�:p$
9�*����P�1�ʶ���  ��J���ӱ�g{+��|x�iɰ�����6�%�A�W������ޞ�Nw�����      ����� �Կp���ޞ�bF�i�C�.E�$�;�I���D���"��g�c�{��֯���J��ѻ��)�P{K�^��:7�
;
N*;��:;�C;$�F;�8H;m�H;��H;��H;��H;[�H;V�H;��H;��H;��H;�H;��H;��H;��H;U�H;Y�H;��H;��H;��H;k�H;�8H;$�F;�C;��:;N*;7�
;d��:p{K���)��ѻ��J��֯�{�g�c�"�����D��I��$�;.E�i�C�bF��ޞ�p�� �Կ��      ��������� �ԿNw�����<�\�"����l��[0X�����;����w����������]��黟F����0ʒ:�;U�';׏9;9pB;�zF;�!H;��H;L�H;4�H;��H;`�H;W�H;��H;��H;��H;-�H;��H;��H;��H;U�H;`�H;��H;/�H;I�H;��H;�!H;�zF;9pB;ԏ9;X�';�;0ʒ:��깟F��黣�]����������w��;�����[0X�l�����"�<�\����Nw�� �Կ��𿞏�      "$�������忉�����!cm�W�-�����Rh��Xde�#-�٪ɽ�v��'�$�}�ɼpmj�$����X����(Ɔ:�x;]�%;J�8;�B;�RF;H;E�H;i�H;�H;��H;[�H;R�H;��H;��H;��H;A�H;��H;��H;��H;P�H;[�H;��H;�H;f�H;E�H;H;�RF;�B;I�8;c�%;�x;(Ɔ: ���X�$���pmj�}�ɼ'�$��v��٪ɽ#-�Xde�Rh������W�-�!cm��������忞����      �>���8���*�O������˿p��G�b�E\�6m־^��S�:��J�)��D�B�9��}������/������t�>:�t�:kp ;�J6;%EA;�IF;�NH; �H;"I;�I;.I;�I;�I;I;� I;��H;G�H;��H;� I;I;�I;�I;.I;�I;"I; �H;�NH;�IF;%EA;�J6;np ;�t�:x�>:����/�����}���9��D�B�)���J�S�:�^��6m־E\�G�b�p���˿����O���*���8�      ��8��4��g&�7��>����<ƿ򲗿�>]�î�Q�Ѿ�p���*7����%W��KR?��|�k8�������8����G:� �:!;/�6;8lA;�YF;�TH;��H;6"I;�I;
I;�I;dI;I;� I;��H;0�H;��H;� I;I;cI;�I;I;�I;3"I;��H;�TH;�YF;8lA;,�6;
!;� �:�G::��������k8���|�KR?�%W�����*7��p��Q�Ѿî��>]�򲗿�<ƿ>���7���g&��4�      ��*��g&��#�v�V[�sL�������M�s5��>ľ����,��D�钐��5�.�ݼ
���q
���x��sk�d�b:�l�:$#;�7;��A;�F;�dH;�I;t"I;I;�I;^I;I;�I;> I;��H;��H;��H;< I;�I;I;]I;�I;I;s"I;�I;�dH;�F;��A;�7;(#;�l�:d�b:�sk���x��q
�
��.�ݼ�5�钐��DὬ�,����>ľs5���M����sL��V[�v��#��g&�      O�7��v����˿B1��:�y�Ŏ6��z �����4�l�+��ͽ#�����&���˼5�k�
�����X�̘ �ȵ�:l�;1&;�9;��B;-�F;�}H;
I;�"I;KI;�I;�I;�I;fI;��H;A�H;��H;A�H;��H;dI;�I;�I;�I;II;}"I;
I;�}H;-�F;��B;�9;3&;l�;̵�:Ԙ ���X�
���5�k���˼��&�#����ͽ+�4�l������z �Ŏ6�:�y�B1���˿���v�7��      ����>���V[忸˿�T���}�R�®��E۾ԗ����M���	������j��3�d����O�#�׻|�/�������:� 
;,*;{;;kC;�'G;�H;I;$"I;I;�I;�
I;�I;�I;d�H;��H;�H;��H;c�H;�I;�I;�
I;�I;I;""I;I;�H;�'G;kC;v;;0*;� 
;���:��|�/�"�׻��O�d���3���j������	���M�ԗ���E۾®�}�R���T���˿V[�>���      �˿�<ƿsL��B1����>]���)�%��ֳ���{���,�r��'��P`I��J���,���3/��+��� ��1695�:
�;p.;A.=;�aD;
�G;��H; I;\!I;wI;kI;�	I;�I;	I;��H;/�H;��H;/�H;��H;	I;�I;�	I;kI;uI;Y!I;I;��H;	�G;�aD;<.=;p.;
�;5�:�169� ��+���3/��,���J��P`I�'��r�齦�,���{�ֳ�%����)��>]��B1��sL���<ƿ      p��򲗿���:�y�}�R���)�ov��>ľ^���I�Yl����������&�ЮҼ��}�$B�����������!:I+�:[z;�3;{j?;�\E;�G;��H;�I;�I;�I;�I;�I;�I;8 I;��H;��H;��H;��H;��H;: I;�I;�I;�I;�I;�I;�I;��H;�G;�\E;xj?;�3;[z;K+�:��!:��������%B���}�ЮҼ��&��������Yl��I�^���>ľov���)�}�R�:�y����򲗿      G�b��>]���M�Ŏ6�®�%���>ľ$q��{�Z�+�R9ݽ!W����L����F����G��׻�;�xm�Ɋ:�i;=P$;��7;��A;1JF;PCH;
�H;� I;�I;�I;6I;II;�I;3�H;�H;��H;-�H;��H;�H;6�H;�I;LI;6I;�I;�I;� I;
�H;PCH;.JF;��A;��7;=P$;�i;
Ɋ:pm��;��׻��G�F�������L�!W��R9ݽ+�{�Z�$q���>ľ%��®�Ŏ6���M��>]�      E\�î�s5��z ��E۾ֳ�^��{�Z�M?#����A����j�$��Aϼ����������xlۺ8;�9�4�:x�;��,;��;;V�C;�G;j�H;�I;�!I;�I;_I;EI;�I;[I;9�H;#�H;��H;@�H;��H;#�H;:�H;\I;�I;EI;]I;�I;�!I;�I;l�H;�G;T�C;��;;��,;y�;�4�:8;�9vlۺ����������Aϼ$����j��A�����M?#�{�Z�^��ֳ��E۾�z �s5�î�      6m־Q�Ѿ�>ľ����ԗ����{��I�+�����V���{�=�/�"���,��4=�+�һ3�@�h� ���k:M�:-b;��3;Qj?;�2E;�G;��H;SI;� I;�I;�I;=	I;I;��H;�H;�H;��H;v�H;��H;�H;�H;��H;I;?	I;�I;�I;� I;QI;��H;�G;�2E;Qj?;��3;-b;M�:��k:d� �4�@�+�һ4=��,��"��=�/��{��V�����+��I���{�ԗ�������>ľQ�Ѿ      ^���p����4�l���M���,�Yl�R9ݽ�A���{���5��J��;���T[�?������O���Q�9�:��;G*;B�9;|kB;�F;�NH;��H;: I;�I;�I;9I;,I;]I;~�H;��H;��H;��H;��H;��H;��H;��H;~�H;bI;,I;9I;�I;�I;: I;��H;�NH;�F;{kB;B�9;F*;��;�:�Q�9�O������?��T[�;���J����5��{��A��R9ݽYl���,���M�4�l����p��      S�:��*7���,�+���	�r�齃���!W����j�=�/��J���I����k�`��-��2��`���4Ɋ:�o�:4;~r3;@�>;K�D;��G;i�H;'I;L!I;�I;�I;�
I;I;} I;��H;��H;��H;��H;��H;��H;��H;��H;��H;� I;I;�
I;�I;�I;K!I;(I;i�H;��G;I�D;@�>;~r3;4;�o�::Ɋ:x���2���-��`���k��I���J��=�/���j�!W������r�齃�	�+���,��*7�      �J�����D��ͽ���'�������L�$��"��;����k����SI����/��/��>:���:�B;��,;��:;M�B;�xF;�<H;�H;&I;�I;I;bI;�I;�I;��H;��H;U�H;��H;��H;��H;��H;��H;W�H;��H;��H;�I;�I;`I;I;�I;'I;�H;�<H;�xF;O�B;��:;��,;�B;���:�>:�/���/�SI�������k�;��"��$����L����'������ͽ�D����      )��%W��钐�"�����j�P`I���&����@ϼ�,���T[�`�SI��0;��mk�H:f5�:�;*&;��6;�!@;W2E;��G;��H;I;!I;nI;/I;I;WI;� I;��H;$�H;��H;��H;��H;f�H;��H;��H;��H;%�H;��H;� I;ZI;I;/I;nI;!I;I;��H;�G;W2E;�!@;��6;*&;�;`5�:H:�mk�0;�SI��`��T[��,��@ϼ�����&�P`I���j�#���钐�%W��      D�B�KR?��5���&��3��J��ѮҼF�����4=�?��-����/��mk�x��9�׳:��;R!;z3;�=;��C;@�F;4dH;�H;�I;/I;�I;CI;�I;�I;d�H;�H;��H;��H;b�H;��H;X�H;��H;c�H;��H;��H;"�H;d�H;�I;�I;DI;�I;1I;�I;�H;/dH;@�F;��C;�=;z3;W!;��;�׳:x��9�mk���/��-��?�5=����F��ѮҼ�J���3���&��5�LR?�      9���|�-�ݼ��˼d���,��ߟ}���G����,�һ����4���/�@:�׳:$�;�b;ѣ0;�<;ȮB;�IF;�H;G�H;�I;� I;9I;XI;{
I;�I;B I;P�H;t�H;-�H;F�H;B�H;��H;\�H;��H;C�H;I�H;-�H;w�H;P�H;B I;�I;|
I;WI;<I;� I;�I;C�H;�H;�IF;ȮB;�<;ӣ0;�b;&�;�׳:H:�/�2������,�һ�����G�ߟ}��,��d����˼-�ݼ�|�      }���j8����5�k���O��3/�#B��׻����3�@��O��x����>:`5�:��;�b;��/;L;;]�A;��E;�G;�H;�
I;� I;!I;I;�I;�I;�I;��H;_�H;��H;��H;�H;7�H;��H;T�H;��H;7�H;"�H;��H;��H;_�H;��H;�I;�I;�I;I;!I;� I;�
I;�H;�G;��E;^�A;N;;��/;�b;��;`5�:�>:p����O��4�@������׻#B��3/���O�5�k���k8��      ������q
�	���$�׻�+�������;�zlۺt� ��Q�9.Ɋ:���:�;U!;̣0;M;;ޓA;�pE;��G;�H;�H;�I;YI;zI;DI;�I;�I;%�H;e�H;��H;%�H;B�H;�H;"�H;��H;_�H;��H;"�H;�H;B�H;)�H;��H;d�H;"�H;�I;�I;EI;zI;VI;�I;�H;�H;��G;�pE;�A;L;;ϣ0;U!;�;���:0Ɋ:�Q�9|� �zlۺ�;������+��"�׻
����q
���      /�������x���X���/�� ������m�(;�9t�k:�:�o�:�B;+&;z3;�<;]�A;�pE;�tG;}H;K�H;KI;�I;eI;I;�
I;I;u I;s�H;F�H;��H;��H;��H;��H;�H;��H;��H;��H;�H;��H;��H;��H;��H;D�H;p�H;v I;I;�
I;I;bI;�I;KI;H�H;}H;�tG;�pE;\�A;�<;|3;+&;�B;�o�:�:x�k:8;�9�m칪���ݺ ��/���X���x����      ��������sk�ؘ ��� 169��!:�Ȋ:�4�:I�:��;.;~�,;�6;�=;��B;��E;��G;}H;��H;�I;7 I;�I;|I;�I;MI;�I;l�H;�H;`�H;	�H;6�H;��H;��H;�H;��H;��H;��H;�H;��H;��H;7�H;	�H;]�H;�H;l�H;�I;MI;�I;xI;�I;7 I;�I;��H;}H;��G;��E;®B;�=;�6;��,;0;��;C�:�4�: Ɋ:��!:P169���ؘ ��sk�,���      ��>:X�G:l�b:���:���:5�:G+�:�i;t�;+b;A*;wr3;��:;�!@;��C;�IF;�G;�H;K�H;�I;? I;eI;]I;�I;7I;�I;D�H;��H;��H;��H;o�H;��H;��H;��H;9�H;��H;��H;��H;9�H;��H;��H;��H;o�H;��H;��H;��H;C�H;�I;7I;�I;]I;eI;< I;�I;K�H;��H;�G;�IF;��C;�!@;��:;wr3;@*;+b;u�;�i;G+�:5�:���:���:t�b:�G:      �t�:�:�l�:c�;� 
;�;az;=P$;��,;��3;B�9;?�>;L�B;V2E;@�F;�H;�H;�H;KI;8 I;dI;�I;\I;�I;I;��H;G�H;r�H;��H;��H;�H;��H;��H;��H;[�H;�H;��H;�H;[�H;��H;��H;��H;�H;��H;��H;r�H;E�H;��H;I;�I;ZI;�I;bI;9 I;KI;	�H;�H;�H;A�F;V2E;L�B;?�>;B�9;��3;��,;@P$;az;�;� 
;c�;�l�:�:      op ;!;$#;(&;$*;p.;�3;�7;��;;Nj?;xkB;I�D;�xF;��G;1dH;C�H;�
I;�I;�I;�I;]I;^I;I;{I;W�H;��H;��H;M�H;�H;:�H;��H;��H;��H;�H;z�H;@�H;-�H;@�H;z�H;�H;��H;��H;��H;7�H;�H;M�H;��H;��H;Y�H;xI;I;^I;YI;�I;�I;�I;�
I;C�H;3dH;��G;�xF;K�D;{kB;Mj?;��;;�7;�3;p.;+*;*&;&#;�!;      �J6;;�6;�7;�9;z;;:.=;~j?;��A;T�C;�2E;�F;��G;�<H;��H;�H;�I;� I;ZI;dI;{I;�I;�I;{I;o�H;��H;��H;��H;S�H;`�H;��H;��H;��H;��H;N�H;��H;��H;p�H;��H;��H;P�H;��H;��H;��H;��H;]�H;S�H;��H;��H;��H;m�H;yI;�I;�I;{I;eI;\I;� I;�I;�H;��H;�<H;��G;�F;�2E;T�C;��A;}j?;<.=;�;;�9;�7;,�6;      -EA;BlA;��A;��B;kC;�aD;�\E;*JF;�G;��G;�NH;i�H;�H;I;�I;� I;&I;zI;I;�I;:I;!I;]�H;��H;�H;��H;[�H;p�H;��H;��H;��H;��H; �H;��H; �H;��H;��H;��H;"�H;��H;��H;��H;��H;��H;��H;p�H;X�H;��H;�H;��H;\�H;!I;9I;�I;I;~I;#I;� I;�I;I;�H;i�H;�NH;��G;�G;*JF;�\E;�aD;kC;��B;��A;BlA;      �IF;�YF;�F;'�F;�'G;��G;��G;ICH;g�H;��H;��H;'I;!I;!I;-I;6I;I;BI;�
I;JI;I;��H;��H;��H;��H;��H;��H;��H;��H;��H;��H;��H;[�H;��H;v�H;Y�H;H�H;Y�H;x�H;��H;W�H;��H;��H;��H;��H;��H;��H;��H;��H;��H;��H;��H;zI;JI;�
I;BI;I;8I;-I;!I;!I;'I;��H;��H;g�H;ICH;��G; �G;�'G;'�F;��F;�YF;      OH;�TH;�dH;�}H;�H;��H;��H;�H;�I;LI;7 I;K!I;�I;nI;�I;XI;I;�I;I;�I;D�H;H�H;��H;��H;V�H;��H;�H;��H;��H;��H;��H;�H;��H;0�H; �H;��H;��H;��H;��H;/�H;��H;�H;��H;��H;��H;��H; �H;��H;W�H;��H;��H;H�H;@�H;�I;I;�I; I;WI;�I;nI;�I;L!I;9 I;LI;�I;�H;��H;��H;
�H;�}H;�dH;�TH;      �H;��H;�I;�	I;I;I;�I; !I;�!I;� I;�I;�I;I;/I;CI;z
I;�I;�I;r I;m�H;��H;r�H;M�H;T�H;k�H;��H;��H;��H;��H;��H;�H;r�H;�H;��H;r�H;C�H;:�H;C�H;r�H;��H;
�H;r�H;�H;��H;��H;��H;��H;��H;m�H;T�H;K�H;r�H;��H;m�H;s I;�I;�I;{
I;CI;/I;I;�I;�I;� I;�!I;!I;�I;I;I;�	I;�I;��H;      ."I;8"I;p"I;�"I;"I;W!I;�I;�I;�I;�I;�I;�I;_I;I;�I;�I;�I;!�H;r�H;�H;��H;��H;�H;c�H;��H;��H;��H;��H;��H;�H;e�H;��H;��H;5�H;��H;��H;��H;��H;��H;5�H;��H;��H;g�H;�H;��H;��H;��H;��H;��H;c�H;�H;��H;��H;�H;p�H;#�H;�I;�I;�I;I;_I;�I;�I;�I;�I;�I;�I;U!I;&"I;�"I;p"I;/"I;      �I;�I;$I;HI;I;yI;�I;�I;bI;�I;=I;�
I;�I;_I;�I;C I;��H;`�H;C�H;`�H;��H;��H;3�H;��H;��H;��H;��H;��H;
�H;V�H;��H;|�H;�H;��H;��H;��H;s�H;��H;��H;��H;�H;�H;��H;U�H;�H;��H;��H;��H;��H;��H;2�H;��H;��H;a�H;C�H;a�H;��H;E I;�I;_I;�I;�
I;@I;�I;dI;�I;�I;yI;I;II; I;�I;      1I;I;�I;�I;�I;gI;�I;<I;KI;@	I;2I; I;�I;� I;g�H;V�H;f�H;��H;��H;�H;r�H;�H;��H;��H;��H;��H;��H; �H;d�H;��H;`�H;��H;��H;v�H;D�H;&�H;�H;'�H;D�H;w�H;��H;�H;_�H;��H;e�H; �H;��H;��H;��H;��H;��H;�H;o�H;�H;��H;��H;c�H;V�H;g�H;� I;�I; I;3I;D	I;LI;?I;�I;hI;�I;�I;�I;I;      �I;�I;`I;�I;�
I;�	I;�I;PI;�I;I;bI;� I;��H;��H;#�H;{�H;��H;'�H;��H;=�H;��H;��H;��H;��H;��H;��H;�H;r�H;��H;|�H;��H;��H;[�H;4�H;��H;��H;��H;��H;��H;4�H;X�H;��H;��H;~�H;��H;r�H;�H;��H;��H;��H;��H;��H;��H;=�H;��H;)�H;��H;}�H;&�H;��H;��H;� I;cI;I;�I;OI;�I;�	I;�
I;�I;`I;�I;      �I;tI;I;�I;�I;�I;�I;�I;bI;��H;��H;�H;��H;(�H;��H;0�H;��H;>�H;��H;��H;��H;��H;��H;��H;��H;X�H;��H;�H;��H;�H;��H;\�H;�H;��H;��H;��H;��H;��H;��H;��H;�H;^�H;��H;�H;��H;�H;��H;W�H;��H;��H;��H;��H;��H;��H;��H;?�H;��H;3�H;��H;)�H;��H;�H;��H;��H;bI;�I;�I;�I;�I;�I;I;mI;      (I;I;�I;jI;�I; I;8 I;=�H;=�H;�H;��H;��H;X�H;��H;��H;N�H;'�H;�H;��H;��H;��H;��H;�H;N�H;|�H;��H;)�H;��H;0�H;��H;t�H;4�H;��H;��H;��H;��H;s�H;��H;��H;��H;��H;6�H;t�H;��H;3�H;��H;)�H;��H;~�H;N�H;�H;��H;��H;��H;��H;�H;&�H;P�H;��H;��H;Z�H;��H;��H;�H;?�H;>�H;8 I;I;�I;jI;�I;I;      � I;� I;F I;��H;{�H;��H;��H;�H;)�H;�H;��H;��H;��H;��H;f�H;J�H;>�H;�H;�H;�H;=�H;Y�H;t�H;��H;�H;r�H;��H;q�H;��H;��H;C�H; �H;��H;��H;n�H;b�H;d�H;b�H;n�H;��H;��H;�H;C�H;��H;��H;q�H;��H;t�H;�H;��H;v�H;[�H;:�H;�H;�H;�H;=�H;L�H;i�H;��H;��H;��H;��H;�H;*�H;�H;��H;��H;q�H;��H;E I;� I;      ��H;��H;��H;C�H;��H;(�H;��H;��H;��H;��H;��H;��H;��H;��H;��H;��H;��H;�H;��H;��H;��H;�H;=�H;��H;��H;S�H;��H;A�H;��H;��H;'�H;��H;��H;��H;b�H;H�H;H�H;H�H;b�H;��H;��H;��H;'�H;��H;��H;A�H;��H;R�H;��H;��H;=�H;�H;��H;��H;��H;��H;��H;��H;��H;��H;��H;��H;��H;��H;��H;��H;��H;-�H;��H;@�H;��H;��H;      A�H;6�H;	�H;��H;+�H;y�H;��H;4�H;D�H;s�H;��H;��H;��H;p�H;]�H;d�H;[�H;W�H;��H;��H;��H;��H;'�H;o�H;��H;B�H;��H;=�H;��H;t�H;�H;��H;��H;v�H;d�H;I�H;F�H;I�H;d�H;v�H;��H;��H;�H;v�H;��H;=�H;��H;D�H;��H;l�H;'�H;��H;��H;��H;��H;X�H;Y�H;d�H;]�H;p�H;��H;��H;��H;v�H;F�H;3�H;��H;}�H; �H;��H;�H;.�H;      ��H;��H;��H;@�H;��H;(�H;��H;��H;��H;��H;��H;��H;��H;��H;��H;��H;��H;�H;��H;��H;��H;�H;=�H;��H;��H;S�H;��H;A�H;��H;��H;'�H;��H;��H;��H;b�H;H�H;H�H;H�H;b�H;��H;��H;��H;'�H;��H;��H;A�H;��H;R�H;��H;��H;=�H;�H;��H;��H;��H;��H;��H;��H;��H;��H;��H;��H;��H;��H;��H;��H;��H;-�H;��H;C�H;��H;��H;      � I;� I;E I;��H;{�H;��H;��H;�H;*�H;�H;��H;��H;��H;��H;i�H;L�H;>�H;�H;�H;�H;>�H;[�H;v�H;��H;�H;r�H;��H;q�H;��H;��H;C�H; �H;��H;��H;n�H;b�H;d�H;b�H;n�H;��H;��H;�H;C�H;��H;��H;q�H;��H;r�H;�H;��H;t�H;Y�H;:�H;�H;�H;�H;=�H;J�H;h�H;��H;��H;��H;��H;�H;)�H;�H;��H;��H;q�H;��H;C I;� I;      )I;I;�I;jI;�I; I;8 I;=�H;=�H;�H;��H;��H;Z�H;��H;��H;P�H;'�H;�H;��H;��H;��H;��H;�H;P�H;~�H;��H;)�H;��H;2�H;��H;t�H;4�H;��H;��H;��H;��H;s�H;��H;��H;��H;��H;6�H;t�H;��H;3�H;��H;)�H;��H;|�H;M�H;�H;��H;��H;��H;��H;�H;%�H;N�H;��H;��H;X�H;��H;��H;�H;?�H;=�H;8 I;I;�I;jI;�I;I;      �I;tI;I;�I;�I;�I;�I;�I;bI;��H;��H;�H;��H;)�H;��H;3�H;��H;>�H;��H;��H;��H;��H;��H;��H;��H;X�H;��H;�H;��H;�H;��H;\�H;�H;��H;��H;��H;��H;��H;��H;��H;�H;_�H;��H;�H;��H;�H;��H;W�H;��H;��H;��H;��H;��H;��H;��H;>�H;��H;0�H;��H;(�H;��H;�H;��H;��H;bI;�I;�I;�I;�I;�I;I;rI;      �I;�I;bI;�I;�
I;�	I;�I;OI;�I;I;cI;� I;��H;��H;&�H;}�H;��H;(�H;��H;>�H;��H;��H;��H;��H;��H;��H;�H;r�H;��H;|�H;��H;��H;Z�H;4�H;��H;��H;��H;��H;��H;4�H;X�H;��H;��H;~�H;��H;r�H;�H;��H;��H;��H;��H;��H;��H;=�H;��H;(�H;��H;{�H;#�H;��H;��H;� I;bI;I;�I;NI;�I;�	I;�
I;�I;bI;�I;      1I;I;�I;�I;�I;gI;�I;=I;LI;C	I;3I; I;�I;� I;g�H;W�H;d�H;��H;��H;�H;t�H;�H;��H;��H;��H;��H;��H; �H;d�H;��H;_�H;��H;��H;w�H;D�H;'�H;�H;&�H;D�H;v�H;��H;�H;`�H;��H;e�H; �H;��H;��H;��H;��H;��H;�H;o�H;�H;��H;��H;c�H;V�H;g�H;� I;�I; I;/I;B	I;KI;<I;�I;hI;�I;�I;�I;I;      �I;�I;#I;II;I;vI;�I;�I;fI;�I;@I;�
I;�I;aI;�I;E I;��H;`�H;C�H;d�H;��H;��H;3�H;��H;��H;��H;��H;��H;�H;V�H;��H;~�H;�H;��H;��H;��H;s�H;��H;��H;��H;�H;~�H;��H;U�H;
�H;��H;��H;��H;��H;��H;2�H;��H;��H;`�H;C�H;a�H;��H;E I;�I;^I;�I;�
I;=I;�I;dI;�I;�I;wI;I;HI;#I;�I;      '"I;3"I;t"I;�"I;$"I;R!I;�I;�I;�I;�I;�I;�I;_I;I;�I;�I;�I;"�H;p�H;�H;��H;��H;�H;c�H;��H;��H;��H;��H;��H;�H;g�H;��H;��H;5�H;��H;��H;��H;��H;��H;5�H;��H;��H;e�H;
�H;��H;��H;��H;��H;��H;c�H;�H;��H;��H;�H;r�H;"�H;�I;�I;�I;I;_I;�I;�I;�I;�I;�I;�I;T!I;!"I;"I;w"I;5"I;      �H;��H;�I;�	I;I;I;�I;!I;�!I;� I;�I;�I;I;0I;DI;{
I;�I;�I;s I;m�H;��H;r�H;M�H;T�H;m�H;��H;��H;��H;��H;��H;�H;r�H;�H;��H;q�H;C�H;:�H;C�H;r�H;��H;�H;t�H;�H;��H;��H;��H;��H;��H;k�H;T�H;K�H;r�H;��H;m�H;r I;�I;�I;{
I;CI;.I;I;�I;�I;� I;�!I;!I;�I;�I;I;�	I;�I;��H;      OH;�TH;�dH;�}H;�H;��H;��H;�H;�I;MI;9 I;L!I;�I;mI;�I;XI;I;�I;I;�I;G�H;H�H;��H;��H;W�H;��H;�H;��H;��H;��H;��H;�H;��H;/�H;��H;��H;��H;��H; �H;/�H;��H;�H;��H;��H;��H;��H; �H;��H;V�H;��H;��H;H�H;@�H;�I;I;�I; I;WI;�I;nI;�I;K!I;7 I;MI;�I;�H;��H;�H;�H;�}H;�dH;�TH;      �IF;�YF;��F;*�F;�'G;�G;��G;ICH;f�H;��H;��H;%I;!I;!I;,I;8I;I;AI;�
I;JI;�I;��H;��H;��H;��H;��H;��H;��H;��H;��H;��H;��H;Z�H;��H;u�H;Y�H;H�H;Y�H;x�H;��H;W�H;��H;��H;��H;��H;��H;��H;��H;��H;��H;��H;��H;zI;JI;�
I;DI;I;6I;-I;!I;!I;'I;��H;��H;f�H;HCH;��G;��G;�'G;(�F; �F;�YF;      -EA;BlA;��A;��B;kC;�aD;�\E;(JF;�G;��G;�NH;i�H;�H;I;�I;� I;%I;{I;I;�I;;I;!I;]�H;��H;�H;��H;Z�H;p�H;��H;��H;��H;��H;��H;��H; �H;��H;��H;��H; �H;��H;��H;��H;��H;��H;��H;p�H;Z�H;��H;�H;��H;\�H;!I;9I;�I;I;|I;"I;� I;�I;I;�H;i�H;�NH;��G;�G;(JF;�\E;�aD;kC;��B;��A;ClA;      �J6;:�6;��7;�9;s;;@.=;{j?;��A;U�C;�2E;�F;��G;�<H;��H;�H;�I;� I;ZI;eI;{I;�I;�I;{I;q�H;��H;��H;��H;S�H;b�H;��H;��H;��H;��H;N�H;��H;��H;p�H;��H;��H;N�H;��H;��H;��H;��H;]�H;S�H;��H;��H;��H;o�H;yI;�I;�I;{I;dI;\I;� I;�I;�H;��H;�<H;��G;�F;�2E;U�C;��A;{j?;@.=;�;;�9;��7;-�6;      kp ;!;4#;*&;!*;"p.;�3;�7;��;;Nj?;{kB;K�D;�xF;��G;3dH;D�H;�
I;�I;�I;�I;`I;^I;I;{I;Y�H;��H;��H;M�H;�H;:�H;��H;��H;��H;�H;z�H;@�H;-�H;@�H;z�H;�H;��H;��H;��H;7�H;�H;M�H;��H;��H;W�H;xI;I;^I;YI;�I;�I;�I;�
I;C�H;3dH;��G;�xF;I�D;ykB;Kj?;��;;�7;�3;!p.;&*;+&;,#;!;      �t�:�:�l�:c�;� 
;�;az;>P$;��,;��3;D�9;?�>;L�B;V2E;@�F;�H;�H;�H;KI;8 I;fI;�I;\I;�I;I;��H;G�H;r�H;��H;��H;�H;��H;��H;��H;[�H;�H;��H;�H;[�H;��H;��H;��H;�H;��H;��H;r�H;D�H;��H;I;�I;ZI;�I;bI;9 I;KI;	�H;�H;�H;A�F;V2E;L�B;@�>;A�9;��3;��,;=P$;az;�;� 
;c�;�l�:�:      l�>:@�G:|�b:���:���:5�:K+�:�i;t�;+b;A*;wr3;��:;�!@;��C;�IF;�G;�H;K�H;�I;? I;eI;]I;�I;7I;�I;D�H;��H;��H;��H;o�H;��H;��H;��H;9�H;��H;��H;��H;9�H;��H;��H;��H;o�H;��H;��H;��H;C�H;�I;7I;�I;\I;eI;< I;�I;K�H;�H;�G;�IF;��C;�!@;��:;wr3;C*;(b;w�;�i;K+�:5�:���:���:��b:�G:      ��������sk��� ����@169��!:�Ȋ:�4�:E�:��;0;~�,;�6;�=;®B;��E;��G;}H;��H;�I;7 I;�I;~I;�I;MI;�I;l�H;�H;`�H;	�H;6�H;��H;��H;�H;��H;��H;��H;�H;��H;��H;7�H;	�H;]�H;�H;l�H;�I;MI;�I;xI;�I;7 I;�I;��H;}H;��G;��E;��B;�=;�6;~�,;-;��;E�:�4�: Ɋ:��!:P169����� ��sk�,���      /�������x���X���/�� ������m�(;�9x�k:�:�o�:�B;+&;z3;�<;^�A;�pE;�tG;}H;L�H;KI;�I;gI;I;�
I;I;v I;s�H;G�H;��H;��H;��H;��H;�H;��H;��H;��H;�H;��H;��H;��H;��H;C�H;o�H;u I;I;�
I;I;aI;�I;KI;H�H;}H;�tG;�pE;Z�A;�<;z3;+&;�B;�o�:�:t�k:8;�9�m칪���ݺ ���/���X���x����      ������q
�
���&�׻�+�������;�zlۺ|� ��Q�90Ɋ:���:�;U!;ϣ0;M;;��A;�pE;��G;�H;�H;�I;ZI;zI;EI;�I;�I;&�H;e�H;��H;(�H;C�H;�H;"�H;��H;_�H;��H;!�H;�H;A�H;(�H;��H;d�H;"�H;�I;�I;EI;zI;UI;�I;�H;�H;��G;�pE;ߓA;L;;̣0;U!;�;���:.Ɋ:�Q�9t� �zlۺ�;������+��#�׻	����q
���      }���j8����5�k���O��3/�$B��׻����4�@��O��p����>:`5�:��;�b;��/;L;;^�A;��E;�G;�H;�
I;� I;!I;I; I;�I;�I;��H;_�H;��H;��H;"�H;7�H;��H;T�H;��H;7�H; �H;��H;��H;_�H;��H;�I;�I;�I;I;!I;� I;�
I;�H;�G;��E;]�A;N;;��/;�b;��;`5�:�>:x����O��4�@������׻$B��3/���O�5�k���k8��      9���|�-�ݼ��˼d���,��ߟ}���G����,�һ����2���/�@:�׳:&�;�b;ң0;�<;ȮB;�IF;�H;F�H;�I;� I;;I;ZI;|
I;�I;B I;P�H;v�H;/�H;I�H;C�H;��H;\�H;��H;B�H;F�H;,�H;w�H;P�H;B I;�I;{
I;UI;;I;� I;�I;C�H;�H;�IF;ȮB;�<;ң0;�b;$�;�׳:@:�/�4������,�һ�����G�ߟ}��,��d����˼-�ݼ�|�      D�B�KR?��5���&��3��J��ѮҼF�����5=�?��-����/��mk�x��9�׳:��;T!;z3;�=;��C;@�F;4dH;�H;�I;1I;�I;DI;�I;�I;d�H;�H;��H;��H;c�H;��H;X�H;��H;b�H;��H;��H;"�H;d�H;�I;�I;CI;�I;0I;�I;�H;-dH;@�F;��C;�=;z3;U!;��;�׳:x��9�mk���/��-��?�4=����F��ѮҼ�J���3���&��5�LR?�      )��%W��钐�#�����j�P`I���&����@ϼ�,���T[�`�SI��0;��mk�H:f5�:�;*&;��6;�!@;W2E;��G;��H;I;!I;oI;/I;!I;ZI;� I;��H;'�H;��H;��H;��H;f�H;��H;��H;��H;"�H;��H;� I;WI;I;/I;nI;!I;I;��H;�G;W2E;�!@;��6;*&;�;d5�:H:�mk�0;�SI��`��T[��,��@ϼ�����&�P`I���j�#���钐�%W��      �J�����D��ͽ���'�������L�$��"��;����k����SI����/��/��>:���:�B;��,;��:;O�B;�xF;�<H;�H;&I;�I;I;bI;�I;�I;��H;��H;W�H;��H;��H;��H;��H;��H;U�H;��H;��H;�I;�I;_I;I;�I;)I;�H;�<H;�xF;M�B;��:;��,;�B;���:�>:�/���/�SI�������k�;��"��$����L����'������ͽ�D����      S�:��*7���,�+���	�r�齃���!W����j�=�/��J���I����k�`��-��2��p���6Ɋ:�o�:3;{r3;@�>;L�D;��G;i�H;*I;L!I;�I;�I;�
I;I;~ I;��H;��H;��H;��H;��H;��H;��H;��H;��H;~ I;I;�
I;�I;�I;K!I;'I;i�H;��G;H�D;@�>;~r3;3;�o�::Ɋ:p���4���-��`���k��I���J��=�/���j�!W������r�齃�	�+���,��*7�      ^���p����4�l���M���,�Yl�R9ݽ�A���{���5��J��;���T[�?������O���Q�9�:��;D*;B�9;|kB;�F;�NH;��H;: I;�I;�I;9I;,I;]I;�H;��H;��H;��H;��H;��H;��H;��H;|�H;_I;,I;9I;�I;�I;: I;��H;�NH;�F;ykB;B�9;D*;��;�:�Q�9�O������?��T[�;���J����5��{��A��R9ݽYl���,���M�4�l����p��      6m־Q�Ѿ�>ľ����ԗ����{��I�+�����V���{�=�/�"���,��4=�+�һ3�@�h� ���k:M�:,b;��3;Rj?;�2E;�G;��H;SI;� I;�I;�I;?	I;I;��H;�H;�H;��H;v�H;��H;�H;�H;��H;I;=	I;�I;�I;� I;QI;��H;�G;�2E;Pj?;��3;-b;K�:��k:d� �4�@�,�һ4=��,��"��=�/��{��V�����+��I���{�ԗ�������>ľQ�Ѿ      E\�î�s5��z ��E۾ֳ�^��{�Z�M?#����A����j�$��Aϼ����������xlۺ8;�9�4�:w�;��,;��;;V�C;�G;l�H;�I;�!I;�I;]I;EI;�I;^I;:�H;#�H;��H;@�H;��H;#�H;9�H;ZI;�I;EI;]I;�I;�!I;�I;j�H;�G;T�C;��;;��,;y�;�4�:8;�9vlۺ����������Aϼ$����j��A�����M?#�{�Z�^��ֳ��E۾�z �s5�î�      G�b��>]���M�Ŏ6�®�%���>ľ$q��{�Z�+�R9ݽ!W����L����F����G��׻�;�pm�Ɋ:�i;=P$;��7;��A;.JF;PCH;�H;� I;�I;�I;6I;KI;�I;7�H;�H;��H;-�H;��H;�H;4�H;�I;II;6I;�I;�I;� I;	�H;OCH;1JF;��A;��7;=P$;�i;
Ɋ:xm��;��׻��G�F�������L�!W��R9ݽ+�{�Z�$q���>ľ%��®�Ŏ6���M��>]�      p��򲗿���:�y�}�R���)�ov��>ľ^���I�Yl����������&�ЮҼ��}�$B�����������!:G+�:[z;�3;}j?;�\E;�G;��H;�I;�I;�I;�I;�I;�I;; I;��H;��H;��H;��H;��H;8 I;�I;�I;�I;�I;�I;�I;��H;�G;�\E;zj?;�3;[z;K+�:��!:��������$B���}�ЮҼ��&��������Yl��I�^���>ľov���)�}�R�:�y����򲗿      �˿�<ƿsL��B1����>]���)�%��ֳ���{���,�r��'��P`I��J���,���3/��+��� �p1695�:
�;p.;@.=;�aD;
�G;��H;I;^!I;yI;kI;�	I;�I;	I;��H;/�H;��H;1�H;��H;	I;�I;�	I;kI;uI;X!I; I;��H;
�G;�aD;=.=;p.;
�;5�:p169� ��+���3/��,���J��P`I�'��r�齦�,���{�ֳ�%����)��>]��B1��sL���<ƿ      ����>���V[忸˿�T���}�R�®��E۾ԗ����M���	������j��3�d����O�"�׻|�/������:� 
;-*;z;;kC;�'G;�H;I;%"I;I;�I;�
I;�I;�I;d�H;��H;�H;��H;c�H;�I;�I;�
I;�I;I;""I;I;�H;�'G;kC;y;;/*;� 
;���:��|�/�"�׻��O�d���3���j������	���M�ԗ���E۾®�}�R���T���˿V[�>���      O�7��v����˿B1��:�y�Ŏ6��z �����4�l�+��ͽ#�����&���˼5�k�
�����X�̘ �Ƶ�:l�;1&;�9;��B;-�F;�}H;
I;�"I;LI;�I;�I;�I;dI;��H;A�H;��H;A�H;��H;fI;�I;�I;�I;II;"I;
I;�}H;-�F;��B;�9;3&;l�;̵�:Ԙ ���X�
���5�k���˼��&�#����ͽ+�4�l������z �Ŏ6�:�y�B1���˿���v�7��      ��*��g&��#�v�V[�sL�������M�s5��>ľ����,��D�钐��5�.�ݼ
���q
���x��sk�`�b:�l�:$#;�7;��A;�F;�dH;�I;v"I;I;�I;^I;I;�I;> I;��H;��H;��H;> I;�I;I;]I;�I;I;r"I;�I;�dH;�F;��A;�7;(#;�l�:d�b:�sk���x��q
�
��.�ݼ�5�钐��DὬ�,����>ľs5���M����sL��V[�v��#��g&�      ��8��4��g&�7��>����<ƿ򲗿�>]�î�Q�Ѿ�p���*7����%W��KR?��|�k8�������8��� �G:� �:!;0�6;8lA;�YF;�TH;��H;6"I;�I;I;�I;dI;I;� I;��H;0�H;��H;� I;I;cI;�I;
I;�I;3"I;��H;�TH;�YF;8lA;-�6;
!;� �:�G::��������k8���|�KR?�%W�����*7��p��Q�Ѿî��>]�򲗿�<ƿ>���7���g&��4�      �Aq���i���U�H:�@�����>���w���|A�e5�� ���^Z�����A���]�����d��>",��5���Ѻ���9@��:y�;|Y4;��@;�VF;��H;�GI;�bI;JOI;[:I;*I;]I;�I;I;�I;�I;�I;I;�I;\I;*I;[:I;HOI;�bI;�GI;��H;�VF;��@;zY4;{�;@��:���9�Ѻ�5��>",��d������]��A������^Z�� ��e5�|A�w���>�������@�H:���U���i�      ��i���b�\�O�.5�2i�������������q<���� f��b
V�HE	�!���IY�g9�>�����(��R��f�Ⱥ��:���:<�;b�4;��@;�hF;חH;MII;�bI;�NI;�9I;�)I;'I;�I;�I;�I;�I;�I;�I;�I;%I;�)I;�9I;�NI;�bI;MII;חH;�hF;��@;^�4;@�;���:�:j�Ⱥ�R����(�>���g9��IY�!��HE	�b
V� f������q<������������2i�.5�\�O���b�      ��U�\�O�J-?�/�'���N�῵欿c�{�ga/���뾞���I����d���ZN�Y5������/H�G ��̈��0�":��:��;��5;�`A;�F;s�H;SMI;5bI;�MI;�8I; )I;�I;$I;}I;EI;EI;EI;|I;$I;I;!)I;�8I;�MI;0bI;UMI;s�H;�F;�`A;��5;��;��:0�":Ј��G ��/H�����Y5���ZN�d������I�������ga/�c�{��欿N����/�'�J-?�\�O�      H:�.5�/�'��������lȿ���n$_���Y�Ҿݕ���6�����*���`=�8�漨)��;G�
6������Q:5�:-0";2�7;�&B;+�F;��H;(SI;�`I;�KI;]7I;�'I;zI;XI;�I;�I;�
I;�I;�I;ZI;zI;�'I;]7I;�KI;�`I;)SI;��H;+�F;�&B;.�7;20";5�:��Q:��
6��:G��)��8���`=��*������6�ݕ��Y�Ҿ��n$_����lȿ�������/�'�.5�      @�2i�������J�ѿl������q<��:��a����q����Wн罅��'�Pb̼�zl��.���X�$��L�:��;"�&;��9;jC;�MG;�H;xYI;�^I;�HI;#5I;&I;!I;HI;�I;�
I;�	I;�
I;�I;HI;I;&I;#5I;�HI;�^I;vYI;�H;�MG;hC;�9;%�&;��;R�:(���X��.���zl�Pb̼�'�罅��Wн����q��a���:��q<���l���K�ѿ������2i�      �������N��lȿl���������O���}]׾{����I�����A��=�d�l�x֮��QH��jλ�$��#�ر�:�N;�+;<;?4D;��G;�I;�^I;�[I;#EI;b2I;�#I;I;�I;�I;�	I;�I;�	I;�I;�I;I;�#I;b2I; EI;�[I;�^I;�I;��G;>4D;<;�+;�N;ڱ�:�#��$��jλ RH�x֮�l�=�d��A������I�{���}]׾����O�����l���lȿN�Ύ��      >��������欿�������O��x����� ���l���"��ܽ���`=����p���k"�R���ۺ��9�?�:�L;й0;�>;�ME;�#H;&I;bI;EWI;�@I;3/I;!I;{I;BI;LI;�I;�I;�I;LI;CI;{I;�!I;3/I;�@I;CWI;bI;&I;�#H;�ME;�>;Ϲ0;�L;�?�:��9�ۺR���k"�p������`=����ܽ��"��l�� ����뾂x���O�������欿����      w�������c�{�n$_��q<������~��	w��
�6�����!���h����ݷ��w d�a.��^^e� H[���Z:υ�:�, ;��5;�A;WF;�H;!AI;�bI;�QI;,<I;+I;�I;LI;xI;�	I;(I;mI;(I;�	I;xI;JI;�I;+I;,<I;�QI;�bI;!AI;�H;WF;�A;��5;�, ;Ӆ�:��Z: H[�\^e�b.��w d�ݷ������h�!������
�6�	w��~��������q<�n$_�c�{�����      |A��q<�ga/����:�}]׾� ��	w��>�DE	�����ڽ����3�\�꼔���",��W��#�� �P���:�M
;�f);��:;a@C;8@G;��H;�TI;
`I;jKI;!7I;�'I;�I;�I;zI;I;�I;�I;�I;I;}I;�I;�I;�'I;7I;gKI;`I;�TI;��H;6@G;^@C;��:;�f);�M
;��:��P�"���W�� ",�����\�꼗�3�ڽ������DE	�>�	w��� ��}]׾�:���ga/��q<�      e5�������Y�Ҿ�a��{����l�
�6�DE	���Ƚk���aG����`֮��W�}��2�k�����d,:��:8�;ד1;��>;zE;k�G;`I;f_I;�ZI;zDI;�1I;q#I;�I;8I;A
I;JI;I;]I;I;KI;C
I;7I;�I;o#I;�1I;wDI;�ZI;e_I;aI;i�G;wE;��>;ד1;8�;��:�d,:���4�k�}���W�`֮�����aG�k����ȽDE	�
�6��l�{����a��Y�Ҿ������      � �� f�����ݕ����q��I���"���������k���ZN�Y�¼E�y��$��Q��M� � |W�C�:b0;e�&;#x8;� B;˛F;�H;�@I;5bI;�RI;\=I;Q,I;I;&I;�I;I;wI;YI;�I;YI;wI;I;�I;(I;I;S,I;Z=I;�RI;5bI;�@I;�H;ǛF;� B;#x8;d�&;`0;C�: lW�O� ��Q���$�E�y�¼Y��ZN�k������������"��I���q�ݕ����� f��      �^Z�b
V��I��6�������ܽ!��ڽ���aG�X��ȼ|)��p�(�K��G5������Z:��:TS;K'1;�=;�D;n�G;2�H;YI;Z^I;�II;76I;�&I;�I;�I;�
I;�I;�I;� I;��H;� I;�I;�I;�
I;�I;�I;�&I;76I;�II;Z^I;YI;1�H;l�G;�D;�=;K'1;TS;��:��Z:���G5�L��p�(�|)���ȼX��aG�ڽ��!���ܽ������6��I�b
V�      ���GE	��������Wн�A�����h���3����¼|)��%x/���һ9�X�#����9���:�>;yf);�`9;�&B;��F;�}H;7I;�aI;�UI;�@I;/I;<!I;�I;fI;"I;�I;� I;��H;<�H;��H;� I;�I;"I;iI;�I;=!I;/I;�@I;�UI;�aI;7I;�}H;�F;�&B;�`9;wf);�>;���:��9�"��9�X���һ%x/�|)��¼�����3��h��󑽢A���Wн��콺��HE	�      �A��!��c���*��潅�=�d��`=����[��_֮�D�y�p�(���һe]e�z����f9$��:o�;�1";`�4;�m?;E;��G;��H;�WI;�^I;JKI;�7I;5(I;�I;gI;�
I;bI;\I;��H;�H;}�H;�H;��H;\I;bI;�
I;iI;�I;4(I;�7I;LKI;�^I;�WI;��H;��G;E;�m?;a�4;�1";q�;"��:�f9t���b]e���һp�(�D�y�_֮�[�꼖���`=�<�d�潅��*��c��!��      �]��IY��ZN��`=���'�l����ݷ�������W��$�N��;�X�|����9���:���:��;�0;�<;��C;eG;@�H;	@I;naI;UI;~@I;S/I;�!I;�I;QI;�I;�I;"�H;��H;L�H;��H;L�H;��H;#�H;�I;�I;QI;�I;�!I;S/I;�@I;UI;maI;@I;:�H;eG;��C;"�<;�0;��;���:���:�9z���:�X�L���$��W�����ݷ�����k���'��`=��ZN��IY�      ���g9�W5��7��Pb̼y֮�o��x d� ",�~���Q��G5�#�� �f9���:	�:M�;	�-;��:;LB;|VF;XKH; I;]I;d\I;�HI;H6I;a'I;\I;�I;[
I;�I;< I;�H;��H;��H;+�H;��H;��H;�H;; I;�I;[
I;�I;ZI;c'I;G6I;�HI;f\I;]I;I;ZKH;zVF;LB;��:;
�-;K�;	�:���:�f9 #��G5��Q��~�� ",�x d�o��x֮�Pb̼7��W5��h9�      �d��=��������)���zl��QH��k"�b.���W��1�k�M� ������9"��:���:I�;�-;�9;�aA;��E;h�G;��H;ESI;W`I;+PI;�<I;�,I;�I;tI;QI;�I;�I;��H;��H;�H;��H;��H;��H;�H;��H;��H;�I;�I;PI;sI;�I;�,I;�<I;,PI;U`I;ASI;��H;h�G;��E;�aA;
�9;�-;J�;���:"��:��9���N� �2�k��W��b.���k"��QH��zl��)������>���      @",���(�/H�:G��.���jλR��b^e�#����� pW�|�Z:���:m�;��;�-;�9;�A;dE;d�G;��H;�GI;7aI;�UI;�BI;�1I;-$I;I;.I;�I;6I;��H;��H;�H;L�H;U�H;(�H;V�H;L�H;�H;��H;��H;6I;�I;,I;I;-$I;�1I;�BI;�UI;6aI;�GI;��H;g�G;dE;�A;�9;�-;��;o�;���:|�Z: xW����%��c^e�R���jλ�.��:G�/H���(�      �5���R��D ��
6���X��$��ۺH[� �P��d,:A�:��:�>;�1";�0;��:;�aA;dE;7�G;��H;>I;p`I;�YI;3GI;%6I;�'I;0I;�I;=I;�I; I;E�H;a�H;7�H;��H;��H;��H;��H;��H;7�H;a�H;H�H; I;�I;;I;�I;-I;�'I;%6I;/GI;�YI;p`I;>I;��H;7�G;dE;�aA;��:;�0;�1";�>;��:C�:�d,:��P�H[��ۺ�$��X�
6��D ���R��      �ѺJ�Ⱥʈ�� ��0��P$�ؕ�9��Z:���:��:`0;NS;sf);Z�4;�<;LB;��E;c�G;��H;�:I;�_I;�[I;dJI;G9I;�*I;I;8I;CI;�I;QI;+�H;��H;R�H;o�H;:�H;t�H;)�H;u�H;;�H;p�H;R�H;��H;-�H;PI;�I;CI;6I;I;�*I;D9I;aJI;�[I;�_I;�:I;��H;d�G;��E;LB;�<;Z�4;sf);PS;`0;	��:���:��Z:���9$���"��ʈ��\�Ⱥ      ���98�:4�":��Q:8�:ڱ�:�?�:Ņ�:�M
;5�;a�&;E'1;�`9;�m?;��C;xVF;i�G;��H;	>I;�_I;T\I;�KI;W;I;-I;!I;4I;�I;)I;�I;�H;x�H;��H;z�H;��H;��H;�H;��H;�H;��H;��H;x�H;��H;x�H;�H;�I;*I;�I;4I;!I;-I;V;I;�KI;Q\I;�_I;	>I;��H;g�G;zVF;��C;�m?;�`9;G'1;a�&;5�;�M
;ǅ�:�?�:౩::�:��Q:4�":��:      F��:���:�:�:��;�N;�L;�, ;�f);ԓ1;%x8;�=;�&B;E;cG;VKH;��H;�GI;p`I;�[I;�KI;�;I;/.I;r"I;yI;VI;\	I;�I;��H;/�H;�H;��H;��H;_�H;��H;��H;��H;��H;��H;_�H;��H;��H;�H;*�H;��H;�I;Z	I;XI;zI;n"I;,.I;�;I;�KI;�[I;p`I;�GI;��H;UKH;fG;E;�&B;�=;#x8;ԓ1;�f);�, ;�L;�N;��;�:�:���:      ~�;<�;��;&0";�&;�+;Ϲ0;��5;��:;��>;� B;�D;�F;��G;=�H;I;BSI;9aI;�YI;eJI;W;I;2.I;�"I;BI;I;?
I;oI;��H;��H;��H;��H;��H;=�H;�H;4�H;��H;��H;��H;5�H;�H;<�H;��H;��H;��H;��H;��H;lI;A
I;I;=I;�"I;2.I;S;I;gJI;�YI;:aI;BSI;I;=�H;��G;�F;�D;� B;��>;��:;��5;͹0;�+; �&;&0";��;.�;      �Y4;n�4;�5;-�7;�9;<;�>;�A;^@C;vE;ǛF;l�G;�}H;��H;@I;]I;W`I;�UI;1GI;C9I;-I;q"I;@I;cI;�
I;�I;. I;*�H;��H;)�H;��H;7�H;��H;��H;�H;��H;��H;��H;	�H;��H;��H;7�H;��H;'�H;��H;*�H;- I;�I;�
I;aI;?I;r"I;-I;C9I;1GI;�UI;U`I;]I;@I;��H;�}H;l�G;ǛF;uE;^@C;�A;�>;<;��9;0�7;�5;`�4;      ��@;��@;�`A;�&B;jC;>4D;�ME;WF;3@G;b�G;�H;1�H;7I;�WI;naI;f\I;2PI;�BI;)6I;�*I;!I;|I;I;�
I;/I;^ I;s�H;&�H;c�H;#�H;C�H;��H;��H;��H;"�H;��H;��H;��H;$�H;��H;��H;��H;C�H; �H;`�H;&�H;p�H;` I;1I;�
I;I;|I;!I;�*I;)6I;�BI;/PI;d\I;naI;�WI;7I;1�H;�H;b�G;3@G;WF;�ME;?4D;jC;�&B;�`A;��@;      �VF;�hF;�F;(�F;�MG;�G;�#H;��H;��H;\I;�@I;YI;�aI;�^I;UI;�HI;�<I;�1I;�'I; I;0I;VI;<
I;�I;W I;��H;X�H;��H;.�H;<�H;��H;��H;��H;��H;F�H;��H;��H;��H;G�H;��H;~�H;��H;��H;:�H;-�H;��H;U�H;��H;X I;�I;<
I;VI;,I; I;�'I;�1I;�<I;�HI;UI;�^I;�aI;YI;�@I;ZI;��H;�H;�#H;��G;�MG;(�F;�F;�hF;      ��H;חH;n�H;��H;�H;�I;&I;AI;�TI;b_I;2bI;[^I;�UI;IKI;~@I;G6I;�,I;*$I;0I;8I;�I;\	I;nI;. I;l�H;Z�H;��H;S�H;k�H;��H;m�H;O�H;}�H;��H;y�H;#�H;�H;%�H;w�H;��H;x�H;O�H;m�H;��H;j�H;S�H;��H;Z�H;o�H;. I;lI;\	I;�I;8I;0I;,$I;�,I;G6I;�@I;IKI;�UI;Z^I;2bI;a_I;�TI;AI;&I;�I;�H;��H;n�H;ؗH;      �GI;OII;VMI;%SI;vYI;�^I;bI;�bI;
`I;�ZI;�RI;�II;�@I;�7I;S/I;`'I;�I;I;�I;CI;)I;�I;��H;*�H;!�H;��H;Q�H;G�H;��H;k�H;D�H;L�H;��H;�H;��H;��H;x�H;��H;��H;�H;��H;L�H;D�H;j�H;��H;H�H;P�H;��H;#�H;*�H;��H;�I;&I;CI;�I;I;�I;`'I;S/I;�7I;�@I;�II;�RI;�ZI;`I;�bI;bI;�^I;�YI;#SI;WMI;YII;      cI;�bI;/bI;�`I;�^I;�[I;DWI;�QI;gKI;vDI;X=I;:6I;/I;3(I;�!I;ZI;vI;*I;=I;�I;�I;��H;��H;��H;\�H;0�H;g�H;��H;^�H;@�H;8�H;z�H;��H;k�H;�H;��H;��H;��H;�H;k�H;��H;}�H;8�H;?�H;^�H;��H;j�H;0�H;_�H;��H;��H;��H;�I;�I;=I;,I;tI;\I;�!I;4(I;/I;:6I;X=I;vDI;gKI;�QI;EWI;�[I;�^I;�`I;/bI;�bI;      ROI;�NI;�MI;�KI;�HI;#EI;�@I;,<I;&7I;�1I;W,I;�&I;@!I;�I;�I;�I;TI;�I;�I;QI;�H;*�H;��H;(�H;�H;7�H;��H;h�H;?�H;@�H;i�H;��H;6�H;��H;��H;b�H;]�H;c�H;��H;��H;4�H;��H;i�H;?�H;=�H;j�H;��H;9�H;�H;(�H;��H;*�H;�H;SI;�I;�I;QI;�I;�I;�I;B!I;�&I;W,I;�1I;&7I;0<I;�@I;$EI;�HI;�KI;�MI;�NI;      ]:I;:I;�8I;h7I;/5I;]2I;9/I;�+I;�'I;t#I;I;�I;�I;mI;TI;`
I;�I;4I; I;.�H;|�H;�H;��H;��H;<�H;��H;h�H;D�H;5�H;k�H;��H;/�H;��H;Q�H;�H;��H;��H;��H;�H;Q�H;��H;0�H;��H;i�H;6�H;D�H;g�H;��H;?�H;��H;��H;�H;z�H;1�H; I;6I;�I;`
I;UI;kI;�I;�I;I;v#I;�'I;�+I;9/I;_2I;-5I;h7I;�8I;:I;      !*I;�)I;#)I;�'I;&I;�#I;!I;�I;�I;�I;(I;�I;iI;I;�I;�I;�I;��H;I�H;��H;��H;��H;��H;:�H;��H;��H;M�H;J�H;w�H;��H;-�H;��H;/�H;��H;��H;��H;x�H;��H;��H;��H;,�H;��H;/�H;��H;y�H;J�H;M�H;��H;��H;:�H;��H;��H;��H;��H;J�H;��H;�I;�I;�I;I;iI;�I;*I;�I;�I;�I;!I;�#I;&I;�'I;#)I;�)I;      \I;2I;�I;�I;)I;{I;xI;MI;�I;5I;�I;�
I;"I;eI;�I;? I;��H;��H;c�H;U�H;~�H;��H;:�H;��H;��H;�H;z�H;��H;��H;9�H;��H;2�H;��H;��H;M�H;C�H;P�H;C�H;M�H;��H;��H;3�H;��H;:�H;��H;��H;w�H;�H;��H;��H;9�H;��H;}�H;V�H;c�H;��H;��H;A I;�I;fI;"I;�
I;�I;8I;�I;NI;xI;}I;"I;�I;�I;+I;      �I;�I;I;^I;NI;�I;BI;~I;~I;A
I;"I;�I;�I;aI;&�H;�H;��H;�H;:�H;t�H;��H;]�H;�H;��H;��H;��H;��H;�H;h�H;��H;N�H;��H;��H;\�H;#�H;�H;��H;�H;#�H;\�H;��H;��H;N�H;��H;k�H;�H;��H;��H;��H;��H;�H;_�H;��H;t�H;:�H;�H;��H;	�H;(�H;bI;�I;�I;"I;D
I;~I;I;BI;�I;BI;^I;I;�I;       I;�I;�I;�I;�I;�I;OI;�	I;"I;KI;}I;�I;� I;��H;��H;��H;�H;H�H;��H;>�H;��H;��H;1�H;	�H;�H;C�H;s�H;��H;�H;��H;�H;��H;M�H;$�H;�H;��H;��H;��H;�H;$�H;J�H;��H;�H;��H;�H;��H;r�H;C�H;�H;�H;0�H;��H;��H;?�H;��H;H�H;�H;��H;��H;��H;� I;�I;~I;MI;#I;�	I;OI;�I;�I;�I;�I;�I;      �I;�I;JI;�I;�
I;�	I;�I;0I;�I;I;`I;� I;��H;�H;O�H;��H;��H;Q�H;��H;x�H;�H;��H;��H;��H;��H;��H;"�H;�H;��H;`�H;��H;��H;C�H;�H;��H;��H;��H;��H;��H;�H;B�H;��H;��H;b�H;��H;�H; �H;��H;��H;��H;��H;��H;�H;y�H;��H;R�H;��H;��H;P�H;�H;��H;� I;]I;I;�I;0I;�I;�	I;�
I;�I;II;�I;      �I;�I;OI;�
I;�	I;�I;�I;qI;�I;ZI;�I;��H;@�H;��H;��H;2�H;��H; �H;��H;,�H;��H;��H;��H;��H;��H;��H;�H;y�H;��H;_�H;��H;~�H;Q�H;��H;��H;��H;��H;��H;��H;��H;N�H;�H;��H;b�H;��H;y�H;�H;��H;��H;��H;��H;��H;��H;,�H;��H;!�H;��H;2�H;��H;��H;@�H;��H;�I;]I;�I;pI;�I;�I;�	I;�
I;OI;�I;      �I;�I;JI;�I;�
I;�	I;�I;0I;�I;I;`I;� I;��H;�H;P�H;��H;��H;Q�H;��H;y�H; �H;��H;��H;��H;��H;��H;"�H;�H;��H;`�H;��H;��H;C�H;�H;��H;��H;��H;��H;��H;�H;B�H;��H;��H;b�H;��H;�H;�H;��H;��H;��H;��H;��H;�H;x�H;��H;R�H;��H;��H;O�H;�H;��H;� I;_I;I;�I;0I;�I;�	I;�
I;�I;FI;�I;       I;�I;�I;�I;�I;�I;OI;�	I;#I;MI;~I;�I;� I;��H;��H;��H;�H;H�H;��H;?�H;��H;��H;1�H;	�H;�H;C�H;u�H;��H;�H;��H;�H;��H;M�H;$�H;�H;��H;��H;��H;�H;$�H;J�H;��H;�H;��H;�H;��H;r�H;C�H;�H;�H;0�H;��H;��H;>�H;��H;H�H;�H;��H;��H;��H;� I;�I;|I;MI;"I;�	I;OI;�I;�I;�I;�I;�I;      �I;�I;I;^I;NI;�I;BI;~I;}I;D
I;"I;�I;�I;bI;(�H;	�H;��H;�H;:�H;t�H;��H;_�H;�H;��H;��H;��H;��H;�H;h�H;��H;N�H;��H;��H;\�H;#�H;�H;��H;�H;#�H;\�H;��H;��H;N�H;��H;k�H;�H;��H;��H;��H;��H;�H;]�H;��H;t�H;:�H;�H;��H;�H;&�H;aI;�I;�I; I;A
I;�I;~I;BI;�I;BI;^I;I;�I;      _I;3I;�I;�I;(I;zI;vI;LI;�I;7I;�I;�
I;"I;fI;�I;A I;��H;��H;c�H;U�H;�H;��H;<�H;��H;��H;��H;z�H;��H;��H;9�H;��H;2�H;��H;��H;M�H;C�H;P�H;C�H;M�H;��H;��H;5�H;��H;:�H;��H;��H;v�H;~�H;��H;��H;9�H;��H;{�H;V�H;c�H;��H;��H;? I;�I;eI; I;�
I;�I;7I;�I;LI;xI;}I;!I;�I;�I;0I;      !*I;�)I;')I;�'I;&I;�#I;�!I;�I;�I;�I;*I;�I;iI;I;�I;�I;�I;��H;J�H;��H;��H;��H;��H;:�H;��H;��H;M�H;J�H;y�H;��H;/�H;��H;/�H;��H;��H;��H;x�H;��H;��H;��H;,�H;��H;-�H;��H;y�H;J�H;K�H;��H;��H;:�H;��H;��H;��H;��H;I�H;��H;�I;�I;�I;I;iI;�I;(I;�I;�I;�I;�!I;�#I;&I;�'I;&)I;�)I;      ]:I;:I;�8I;h7I;.5I;]2I;9/I;�+I;�'I;u#I;I;�I;�I;mI;UI;b
I;�I;4I; I;/�H;~�H;�H;��H;��H;?�H;��H;g�H;D�H;5�H;k�H;��H;0�H;��H;Q�H;�H;��H;��H;��H;�H;Q�H;��H;0�H;��H;i�H;6�H;D�H;g�H;��H;<�H;��H;��H;�H;x�H;/�H; I;4I;�I;`
I;UI;mI;�I;�I;I;u#I;�'I;�+I;9/I;_2I;-5I;h7I;�8I;:I;      HOI;�NI;�MI;�KI;�HI; EI;�@I;-<I;(7I;�1I;W,I;�&I;B!I;�I;�I;�I;SI;�I;�I;TI;�H;*�H;��H;(�H;�H;:�H;��H;j�H;@�H;@�H;i�H;��H;6�H;��H;��H;b�H;]�H;c�H;��H;��H;4�H;��H;i�H;?�H;?�H;h�H;��H;7�H;�H;(�H;��H;*�H;�H;QI;�I;�I;QI;�I;�I;�I;?!I;�&I;W,I;�1I;(7I;.<I;�@I;!EI;�HI;�KI;�MI;�NI;      	cI;�bI;5bI;�`I;�^I;�[I;GWI;�QI;gKI;vDI;[=I;<6I;/I;4(I;�!I;\I;wI;*I;=I;�I;�I;��H;��H;��H;_�H;0�H;g�H;��H;`�H;@�H;8�H;z�H;��H;k�H;�H;��H;��H;��H;�H;k�H;��H;|�H;8�H;?�H;]�H;��H;g�H;0�H;\�H;��H;��H;��H;�I;�I;=I;,I;sI;\I;�!I;4(I;/I;:6I;X=I;uDI;gKI;�QI;EWI;�[I;�^I;�`I;5bI;�bI;      �GI;MII;WMI;#SI;uYI;�^I;bI;�bI;`I;�ZI;�RI;�II;�@I;�7I;S/I;`'I;�I;I;�I;CI;,I;�I;��H;*�H;#�H;��H;P�H;H�H;��H;k�H;D�H;L�H;��H;�H;��H;��H;x�H;��H;��H;�H;��H;M�H;D�H;h�H;��H;G�H;P�H;��H;!�H;,�H;��H;�I;%I;CI;�I;I;�I;a'I;S/I;�7I;�@I;�II;�RI;�ZI;
`I;�bI;bI;�^I;�YI;%SI;WMI;]II;      ��H;֗H;r�H;��H;�H;�I;&I;AI;�TI;b_I;2bI;Z^I;�UI;IKI;�@I;H6I;�,I;,$I;0I;9I;�I;\	I;nI;0 I;o�H;Z�H;��H;S�H;k�H;��H;m�H;O�H;{�H;��H;w�H;#�H;�H;#�H;y�H;��H;{�H;Q�H;m�H;��H;j�H;S�H;��H;[�H;l�H;. I;lI;\	I;�I;8I;0I;,$I;�,I;F6I;~@I;JKI;�UI;[^I;4bI;b_I;�TI;AI;&I;�I;�H;��H;o�H;ϗH;      �VF;�hF;�F;+�F;�MG;��G;�#H;�H;��H;\I;�@I;YI;�aI;�^I;UI;�HI;�<I;�1I;�'I; I;2I;VI;<
I;�I;X I;��H;W�H;��H;0�H;<�H;��H;��H;�H;��H;F�H;��H;��H;��H;G�H;��H;~�H;��H;��H;9�H;-�H;��H;U�H;��H;W I;�I;=
I;VI;,I; I;�'I;�1I;�<I;�HI;UI;�^I;�aI;YI;�@I;YI;��H;��H;�#H;�G;�MG;)�F;�F;�hF;      ��@;��@;�`A;�&B;hC;>4D;�ME;WF;4@G;d�G;�H;1�H;7I;�WI;naI;f\I;0PI;�BI;)6I;�*I;!I;|I;I;�
I;1I;` I;r�H;&�H;c�H;"�H;C�H;��H;��H;��H;"�H;��H;��H;��H;"�H;��H;��H;��H;C�H;�H;`�H;&�H;p�H;^ I;/I;�
I;I;|I;!I;�*I;)6I;�BI;/PI;f\I;naI;�WI;7I;1�H;�H;a�G;3@G;WF;�ME;>4D;fC;�&B;�`A;��@;      �Y4;n�4;�5;-�7;�9;<;�>;�A;`@C;wE;țF;n�G;�}H;��H;@I;]I;W`I;�UI;1GI;C9I;-I;r"I;@I;cI;�
I;�I;. I;*�H;��H;)�H;��H;7�H;��H;��H;�H;��H;��H;��H;	�H;��H;��H;9�H;��H;'�H;��H;*�H;- I;�I;�
I;bI;?I;q"I;-I;C9I;1GI;�UI;V`I;]I;@I;��H;�}H;l�G;śF;uE;`@C;�A;�>;<;��9;+�7;�5;a�4;      z�;H�;��;(0";�&;�+;ҹ0;��5;��:;��>;� B;�D;�F;��G;=�H;I;DSI;7aI;�YI;eJI;Y;I;2.I;�"I;@I;I;@
I;oI;��H;��H;��H;��H;��H;=�H;�H;5�H;��H;��H;��H;4�H;�H;<�H;��H;��H;��H;��H;��H;lI;A
I;I;@I;�"I;2.I;S;I;gJI;�YI;:aI;BSI;I;>�H;��G;�F;�D;� B;��>;��:;��5;ҹ0;�+;�&;(0";��;6�;      F��:���:�:�:��;�N;�L;�, ;�f);ԓ1;%x8;�=;�&B;E;cG;VKH;��H;�GI;p`I;�[I;�KI;�;I;/.I;r"I;zI;WI;[	I;�I;��H;/�H;�H;��H;��H;_�H;��H;��H;��H;��H;��H;_�H;��H;��H;�H;*�H;��H;�I;X	I;XI;yI;p"I;,.I;�;I;�KI;�[I;p`I;�GI;��H;VKH;eG;E;�&B;�=;#x8;ԓ1;�f);�, ;�L;�N;��;�:�:���:      ���9 �:H�":��Q:8�:̱�:�?�:ͅ�:�M
;4�;c�&;G'1;�`9;�m?;��C;zVF;h�G;��H;	>I;�_I;T\I;�KI;W;I;-I;!I;4I;�I;*I;�I;�H;x�H;��H;z�H;��H;��H;�H;��H;�H;��H;��H;z�H;��H;x�H;�H;�I;)I;�I;4I;!I;-I;V;I;�KI;Q\I;�_I;	>I;��H;g�G;xVF;��C;�m?;�`9;E'1;c�&;2�;�M
;˅�:�?�:ޱ�:D�:��Q:L�":��:      �ѺD�ȺĈ��"��$��@$����9��Z:���:��:`0;NS;sf);Z�4;�<;LB;��E;c�G;��H;�:I;�_I;�[I;dJI;I9I;�*I;I;8I;CI;�I;SI;-�H;��H;S�H;p�H;;�H;u�H;)�H;u�H;:�H;o�H;P�H;��H;+�H;MI;�I;CI;5I;I;�*I;C9I;aJI;�[I;�_I;�:I;��H;d�G;��E;LB;�<;\�4;sf);NS;^0;	��:���:��Z:���9 $���"��ʈ��\�Ⱥ      �5���R��D ��
6���X��$��ۺH[���P��d,:C�:��:�>;�1";�0;��:;�aA;dE;7�G;��H;
>I;p`I;�YI;3GI;%6I;�'I;0I;�I;>I;�I; I;F�H;b�H;7�H;��H;��H;��H;��H;��H;7�H;_�H;F�H; I;�I;:I;�I;-I;�'I;%6I;/GI;�YI;p`I;>I;��H;7�G;dE;�aA;��:;�0;�1";�>;��:A�:�d,:@�P�H[��ۺ�$��X�
6��D ���R��      @",���(�/H�;G��.���jλR��e^e�%����� pW�x�Z:���:m�;��;�-;	�9;�A;dE;e�G;��H;�GI;:aI;�UI;�BI;�1I;.$I;I;0I;�I;6I;��H;��H;�H;L�H;U�H;(�H;U�H;L�H;�H;��H;��H;6I;�I;,I;I;*$I;�1I;�BI;�UI;4aI;�GI;��H;e�G;dE;�A;�9;�-;��;m�;���:|�Z: pW����%��h^e�R���jλ�.��:G�/H���(�      �d��=��������)���zl� RH��k"�b.���W��2�k�M� ������9"��:���:J�;�-;�9;�aA;��E;i�G;��H;FSI;Y`I;,PI;�<I;�,I;�I;wI;QI;�I;�I;��H;��H;�H;��H;��H;��H;�H;��H;��H;�I;�I;PI;qI;�I;�,I;�<I;+PI;S`I;?SI;��H;g�G;��E;�aA;
�9;�-;I�;���:"��:��9���M� �2�k��W��b.���k"��QH��zl��)������>���      ���g9�W5��7��Pb̼x֮�o��x d� ",�~���Q��G5� #���f9���:	�:N�;	�-;��:;LB;|VF;ZKH;I;]I;f\I;�HI;J6I;c'I;^I;�I;[
I;�I;< I;�H;��H;��H;+�H;��H;��H;�H;; I;�I;[
I;�I;WI;a'I;G6I;�HI;d\I;]I;I;XKH;zVF;LB;��:;
�-;K�;	�:���: �f9#��G5��Q��~�� ",�x d�o��x֮�Pb̼7��W5��h9�      �]��IY��ZN��`=���'�l����ݷ�������W��$�L��:�X�z����9���:���:��;�0;�<;��C;eG;@�H;	@I;maI;UI;�@I;S/I;�!I;�I;QI;�I;�I;#�H;��H;L�H;��H;L�H;��H;#�H;�I;�I;QI;�I;�!I;S/I;~@I;UI;naI;@I;:�H;eG;��C;!�<;�0;��;���:���:�9|���;�X�N���$��W�����ݷ�����k���'��`=��ZN��IY�      �A��!��c���*��潅�<�d��`=����[��_֮�D�y�p�(���һd]e�t����f9$��:p�;�1";`�4;�m?;E;��G;��H;�WI;�^I;LKI;�7I;7(I;�I;iI;�
I;cI;^I;��H;�H;}�H;�H;��H;[I;aI;�
I;gI;�I;4(I;�7I;IKI;�^I;�WI;��H;��G;E;�m?;_�4;�1";q�;"��:�f9z���d]e���һp�(�D�y�_֮�[�꼖���`=�<�d�罅��*��c��!��      ���GE	��������Wн�A�����h���3����¼|)��%x/���һ9�X� #����9���:�>;wf);�`9;�&B;��F;�}H;7I;�aI;�UI;�@I;/I;=!I;�I;gI;"I;�I;� I;��H;<�H;��H;� I;�I; I;fI;�I;<!I;/I;�@I;�UI;�aI;7I;�}H;�F;�&B;�`9;wf);�>;���:��9#��9�X���һ%x/�|)��¼�����3��h��󑽢A���Wн��콺��HE	�      �^Z�b
V��I��6�������ܽ!��ڽ���aG�X��ȼ|)��q�(�L��G5������Z:��:TS;H'1;�=;�D;o�G;1�H;YI;Z^I;�II;:6I;�&I;�I;�I;�
I;�I;�I;� I;��H;� I;�I;�I;�
I;�I;�I;�&I;66I;�II;X^I;YI;2�H;j�G;�D;�=;K'1;TS;��:��Z:���G5�L��p�(�|)���ȼX��aG�ڽ��!���ܽ������6��I�b
V�      � �� f�����ݕ����q��I���"���������k���ZN�Y�¼E�y��$��Q��M� � pW�C�:b0;c�&;#x8;� B;˛F;�H;�@I;7bI;�RI;\=I;S,I;I;&I;�I;I;wI;YI;�I;YI;wI;I;�I;'I;I;Q,I;Z=I;�RI;4bI;�@I;�H;ǛF;� B;#x8;d�&;`0;C�: lW�N� ��Q���$�E�y�¼Y��ZN�k������������"��I���q�ݕ����� f��      e5�������Y�Ҿ�a��{����l�
�6�DE	���Ƚk���aG����`֮��W�}��2�k�����d,:��:6�;ד1;��>;zE;i�G;aI;f_I;�ZI;zDI;�1I;o#I;�I;8I;C
I;JI;I;]I;I;JI;A
I;7I;�I;q#I;�1I;wDI;�ZI;e_I;`I;k�G;wE;��>;ד1;8�;��:�d,:���2�k�~���W�`֮�����aG�k����ȽDE	�
�6��l�{����a��Y�Ҿ������      |A��q<�ga/����:�}]׾� ��	w��>�DE	�����ڽ����3�\�꼔���",��W��#�� �P���:�M
;�f);��:;a@C;6@G;��H;�TI;`I;jKI;7I;�'I;�I;�I;}I;I;�I;�I;�I;I;zI;�I;�I;�'I;7I;gKI;
`I;�TI;��H;8@G;^@C;��:;�f);�M
;��: �P�"���W��",�����\�꼗�3�ڽ������DE	�>�	w��� ��}]׾�:���ga/��q<�      w�������c�{�n$_��q<������~��	w��
�6�����!���h����ݷ��w d�`.��\^e� H[���Z:ͅ�:�, ;��5;�A;WF;�H;!AI;�bI;�QI;,<I;+I;�I;LI;zI;�	I;(I;mI;)I;�	I;zI;JI;�I;+I;,<I;�QI;�bI;AI;�H;WF;�A;��5;�, ;Ӆ�:��Z:H[�[^e�b.��w d�ݷ������h�!������
�6�	w��~��������q<�n$_�c�{�����      >��������欿�������O��x����� ���l���"��ܽ���`=����p���k"�R���ۺ��9�?�:�L;й0;�>;�ME;�#H;&I;bI;GWI;�@I;3/I;!I;|I;EI;LI;�I;�I;�I;LI;BI;yI;!I;3/I;�@I;DWI;bI;&I;�#H;�ME;�>;Ϲ0;�L;�?�:��9�ۺR���k"�p������`=����ܽ��"��l�� ����뾂x���O�������欿����      �������N��lȿl���������O���}]׾{����I�����A��=�d�l�x֮��QH��jλ�$��#�ұ�:�N;�+;<;>4D;��G;�I;�^I;�[I;#EI;b2I;�#I;�I;�I;�I;�	I;�I;�	I;�I;�I;~I;�#I;b2I; EI;�[I;�^I;�I;��G;?4D;<;�+;�N;ڱ�:�#��$��jλ RH�x֮�l�=�d��A������I�{���}]׾����O�����l���lȿN�Ύ��      @�2i�������J�ѿl������q<��:��a����q����Wн罅��'�Pb̼�zl��.���X�(��L�:��;"�&;��9;hC;�MG;�H;vYI;�^I;�HI;#5I;&I;!I;HI;�I;�
I;�	I;�
I;�I;HI;I;&I;#5I;�HI;�^I;xYI;�H;�MG;jC;�9;%�&;��;N�:(���X��.���zl�Pb̼�'�罅��Wн����q��a���:��q<���l���J�ѿ������2i�      H:�.5�/�'��������lȿ���n$_���Y�Ҿݕ���6�����*���`=�8�漨)��:G�
6������Q:5�:/0";2�7;�&B;+�F;��H;)SI;�`I;�KI;]7I;�'I;|I;ZI;�I;�I;�
I;�I;�I;XI;yI;�'I;]7I;�KI;�`I;(SI;��H;,�F;�&B;.�7;00";5�:��Q:��
6��:G��)��8���`=��*������6�ݕ��Y�Ҿ��n$_����lȿ�������/�'�.5�      ��U�\�O�J-?�/�'���N�῵欿c�{�ga/���뾞���I����d���ZN�Y5������/H�G ��Ј��,�":��:��;��5;�`A;�F;s�H;UMI;3bI;�MI;�8I;!)I;�I;$I;}I;EI;EI;EI;}I;$I;I; )I;�8I;�MI;2bI;SMI;s�H;�F;�`A;��5;��;��:0�":Ј��G ��/H�����Y5���ZN�d������I�������ga/�c�{��欿N����/�'�J-?�\�O�      ��i���b�\�O�.5�2i�������������q<���� f��b
V�HE	�!���IY�g9�>�����(��R��f�Ⱥ�:���::�;b�4;��@;�hF;חH;MII;�bI;�NI;�9I;�)I;'I;�I;�I;�I;�I;�I;�I;�I;%I;�)I;�9I;�NI;�bI;MII;֗H;�hF;��@;`�4;@�;���:��:j�Ⱥ�R����(�>���g9��IY�!��HE	�b
V� f������q<������������2i�.5�\�O���b�      ᶕ�T���Ҭ��/�_���7�|�!}߿����,b��V�.l¾Jx�d.���Ž��t�'��^����?��M��ׯ�P�x9���:��;ȼ2;u@@;�fF;_�H;��I;��I;S|I;\I;�CI;F2I;�%I;�I;�I;oI;�I;�I;�%I;D2I;�CI;\I;Q|I;��I;��I;_�H;�fF;u@@;Ƽ2;��;���:p�x9ٯ��M����?�_��'����t���Žd.�Jx�.l¾�V��,b����!}߿|���7�/�_�Ҭ��T���      T���E���%}��+Y��3�����$ڿ&��Ž\����(���s��3�5����p�`�M���<<���������9���:(�;u%3;�p@;zF;��H;<�I;3�I;�{I;�[I;�CI;�1I;�%I;cI;�I;AI;�I;eI;�%I;�1I;�CI;�[I;�{I;0�I;<�I;��H;zF;�p@;r%3;.�;���:���9������<<�N��`��p�5����3��s�(�����Ž\�&���$ڿ����3��+Y�%}�E���      Ҭ��%}�?tf��lG�آ%��p�0�ʿ\����>M����V�����d�ɤ�̷�-�d��
�~I����1�G������8��9���:r;�U4;��@;0�F;^�H;�I;��I;�yI;�YI;�BI;1I;�$I;�I;I;�I;I;�I;�$I;1I;BI;�YI;�yI;��I;�I;^�H;0�F;��@;�U4;u;���:8��9���G�����1�~I���
�-�d�̷�ɤ���d�V�������>M�\���0�ʿ�p�آ%��lG�?tf�%}�      /�_��+Y��lG� f.�|���꿳���N䂿��5���󾎰��O�N�W��Q���Q�
���u����h!�jg����0
:�
�:A�;�16;��A;�G;/I;v�I;ŘI;�vI;�WI;�@I;�/I;�#I;�I;II;�I;II;�I;�#I;�/I;�@I;�WI;�vI;I;x�I;/I;�G;��A;�16;D�;�
�:4
:��jg���h!�v���
����Q�R��W��O�N���������5�N䂿�������|� f.��lG��+Y�      ��7��3�آ%�|��<����ſ
���Ľ\�=����Ͼ����a�3��轻z��{�9�Y�ἓ���z�\7}�Xct���^:�+�:�#;ٍ8;��B;bsG;�%I;�I;/�I;ArI;STI;$>I;�-I;Q"I;�I;%I;�I;%I;�I;Q"I;�-I;%>I;STI;>rI;/�I;�I;�%I;`sG;��B;Ս8;��#;�+�:��^:\ct�Z7}��z����Y��{�9��z����a�3�������Ͼ=��Ľ\�
�����ſ�<��|�آ%��3�      |�����p������ſ%���Ps���1�3r���d���d�}I�ΈŽ��}�]*�EC���^��B�<�D��D�� �:��;�);Q7;;oD;��G;�HI;�I;�I;�lI;1PI;;I;U+I;Z I;�I;�I;kI;�I;�I;[ I;U+I;;I;0PI;�lI;�I;�I;�HI;��G;mD;L7;;�);��; �:�D�<�D��B��^�EC��]*���}�ΈŽ}I��d��d��3r����1��Ps�%����ſ��꿄p����      !}߿�$ڿ0�ʿ����
����Ps�SX:����'l¾�ǆ���7����85���Q�����t���75�N��^�� %�8Wʼ:��;�.;��=;�EE;ZH;�hI;d�I;��I;bfI;ZKI;e7I;�(I;I;/I;�I;�I;�I;/I;I;�(I;g7I;\KI;`fI;��I;d�I;�hI;ZH;�EE;��=;�.;��;Yʼ:�$�8^��L���75��t������Q�85�������7��ǆ�'l¾���SX:��Ps�
�������0�ʿ�$ڿ      ���&��[���N䂿Ľ\���1�����J˾Ꝓ�E�N�y��I������U�'�_�Ҽ��|��z��n���w����&:Q�:�;�W4;	�@;kgF;��H;N�I;_�I;u�I;W_I;FI;G3I;_%I;�I;�I; I;�I; I;�I;�I;^%I;G3I;FI;W_I;r�I;_�I;N�I;��H;jgF;�@;�W4;�;!Q�:��&:�w���n���z���|�_�ҼU�'����I���y��E�N�Ꝓ��J˾�����1�Ľ\�N䂿[���&��      �,b�Ž\��>M���5�=��3r��'l¾Ꝓ�$&W��3�9Sؽ�z��XG����vI����?�t�̻P�-�������:��;��&;g|9;C;�dG;�I;�I;��I;�vI;�WI;i@I;�.I;�!I;�I;�I;I;�I;I;�I;�I;�!I;�.I;i@I;�WI;�vI;��I;}�I;�I;�dG;
C;g|9;��&;��;���:���O�-�u�̻��?�vI�����XG��z��9Sؽ�3�$&W�Ꝓ�'l¾3r��=����5��>M�Ž\�      �V������������Ͼ�d���ǆ�E�N��3��c�[����\�0��$C���o���	��눻�ﳺ���9���:�h;��/;~�=;�E;>3H;�WI;��I;:�I; lI;�OI;c:I;(*I;_I;�I;0I;�I;�I;�I;1I;�I;]I;)*I;c:I;�OI;�kI;:�I;��I;�WI;<3H;�E;~�=;��/;�h;���:���9�ﳺ�눻��	��o�$C��0����\�[���cཱ3�E�N��ǆ��d����Ͼ���������      .l¾(��V������������d���7�y��9Sؽ[���d�A*�^kּ&\����'���nR�`|����:�Z;�#;z=7;o�A;W�F;��H;��I;*�I;�I;-aI;�GI;14I;c%I;�I;�I;�I;�
I;�	I;�
I;�I;�I;�I;f%I;14I;�GI;*aI;�I;+�I;��I;��H;S�F;n�A;z=7;�#;�Z;��:H|��qR�����'�&\��^kּA*��d�[��9Sؽy����7��d���������V���(��      Jx��s���d�O�N�a�3�}I����I����z����\�A*��ݼB���#<<��ڻїV�Dct��&:	��:�C;�</;�D=;�D;��G;79I;�I;�I;TtI;kVI;�?I;�-I;� I;�I;�I;�
I;5I;RI;5I;�
I;�I;�I;� I;�-I;�?I;mVI;UtI;�I;�I;59I;��G;�D;�D=;�</;�C;	��:(�&:Dct�їV��ڻ#<<�B����ݼA*���\��z��I������}I�a�3�O�N���d��s�      d.��3�ɤ�W����ΈŽ85�����XG�0��^kּB����xC�z>�,6}�������x9ُ�:J	;v�&;�;8;��A;�F;�H;yyI;ӝI;5�I;rfI;LI;�7I;�'I;�I;I;�I;QI;�I;�I;�I;QI;�I;	I;�I;�'I;�7I;LI;rfI;5�I;֝I;wyI;�H;��F;��A;�;8;u�&;J	;ߏ�:��x9����+6}�z>��xC�B���^kּ0��XG����85��ΈŽ��W��ɤ��3�      ��Ž5���̷�Q���z����}��Q�U�'����$C��%\��"<<�z>�hn�����@����:���:P�;�'3;��>;�E;�H;�<I;�I;�I;�vI;YI;�AI;�/I;�!I;I;-I;�	I;�I;aI;�I;aI;�I;�	I;/I;%I;�!I;�/I;�AI;YI;�vI;�I;�I;�<I;�H;�E;��>;�'3;Q�;���:���: ����hn��z>�"<<�&\��$C�����U�'��Q���}��z��Q��̷�5���      ��t��p�,�d��Q�{�9�]*����_�ҼvI���o���'��ڻ,6}�����5�(�:�m�:��;,�.;[<;�oC;�7G;��H;�I;�I;�I;_fI;�LI;:8I;"(I;I;�I;�I;�I;�I;	I;� I;	I;�I;�I;�I;�I; I; (I;88I;�LI;_fI;�I;�I;�I;��H;�7G;�oC;]<;,�.;��;�m�:,�:�5����.6}��ڻ��'��o�vI��_�Ҽ���]*�{�9��Q�,�d��p�      '��`��
�
���Y��EC���t����|���?���	���їV�����@�0�:C�:i;\�+;4�9;��A;�fF;��H;�_I;̛I;ّI;DsI;�VI;�@I;/I;-!I;�I;JI;I;�I;� I;��H;F�H;��H;� I;�I;I;MI;�I;.!I;/I;�@I;�VI;GsI;ّI;ɛI;�_I;��H;�fF;��A;4�9;]�+;i;C�:4�: �����їV�����	���?���|��t��DC��Y��
����
�a�      ^��L��~I��v�������^��75��z�t�̻�눻mR�@ct���x9���:�m�:i;��*;�8;+�@;#�E;z(H;�8I;�I;Y�I;�~I;�`I;�HI;�5I;�&I;�I;wI;:
I;�I;� I;0�H;��H;#�H;��H;2�H;� I;�I;<
I;wI;�I;�&I;�5I;�HI;�`I;�~I;T�I;��I;�8I;y(H;(�E;,�@;�8;��*;i;�m�:���:��x9Dct�mR��눻t�̻�z��75��^����v���~I��M��      ��?��<<���1��h!��z��B�N���n��P�-��ﳺP|���&:ӏ�:���:��;X�+;�8;z�@;0^E;��G;�I;-�I;��I;u�I;�iI;|PI;J<I;�+I;�I;�I;�I;kI;�I;�H;��H;��H;�H;��H;��H;�H;�I;mI;�I;�I;�I;�+I;I<I;}PI;�iI;r�I;��I;-�I;�I;��G;0^E;}�@;�8;Y�+;��;���:ӏ�:�&:P|���ﳺP�-��n��N���B黪z��h!���1��<<�      �M����D���jg��a7}�8�D�[���w��������9��:	��:L	;S�;,�.;2�9;)�@;0^E;��G;�I;�I;I�I;��I;�pI;�VI;�AI;�0I;�"I;�I;-I;1I;�I;��H;��H;��H;��H;�H;��H;��H;��H;��H;�I;1I;*I;�I;�"I;�0I;�AI;�VI;�pI;��I;I�I;�I;�I;��G;2^E;)�@;2�9;/�.;S�;L	;	��:��:���9����w��[��4�D�]7}�jg��D�����      ֯����������hct��D�`$�8��&:���:���:�Z;�C;r�&;�'3;W<;��A;"�E;��G;�I;�|I;�I;�I;�uI;�[I;MFI;�4I;p&I;�I;�I;$
I;3I;x�H;�H;v�H;��H;��H;_�H;��H;��H;v�H;�H;y�H;4I;"
I;�I;�I;m&I;�4I;OFI;�[I;�uI;�I;�I;�|I;�I;��G;"�E;��A;X<;�'3;s�&;�C;�Z;���:���:��&:`$�8�D�@ct������ ���      ��x9H��9P��9
:��^:�:Wʼ:Q�:��;�h;�#;�</;�;8;��>;�oC;�fF;z(H;�I;�I;�I;�I;?xI;�^I;{II;�7I;M)I;MI;�I;�I;�I;� I;��H;��H;x�H;��H;��H;��H;��H;��H;y�H;��H;��H;� I;�I;�I;�I;MI;N)I;�7I;wII;�^I;?xI;�I;�I;�I;�I;y(H;�fF;�oC;��>;�;8;�</;�#;�h;��;Q�:Sʼ:�:��^:
:P��9���9      ���:���:��:�
�:�+�:��;�;�;��&;��/;|=7;�D=;��A;�E;7G;��H;�8I;-�I;G�I;�I;>xI;�_I;%KI;�9I;:+I;AI;zI;}I;�I;I;C�H;��H;\�H;}�H;"�H;O�H;)�H;O�H;"�H;~�H;Z�H;��H;C�H;{I;�I;}I;xI;BI;;+I;�9I;"KI;�_I;;xI;�I;G�I;.�I;�8I;��H;�7G;�E;��A;�D=;|=7;��/;��&;�;�;��;�+�:�
�:��:���:      ��;(�;r;:�;�#;�);�.;�W4;h|9;}�=;m�A;�D;�F;�H;��H;�_I;�I;��I;��I;�uI;�^I;&KI;g:I;b,I;| I;�I;�I;�I;dI;��H;F�H;u�H;L�H;��H;��H;��H;��H;��H;��H;��H;J�H;u�H;F�H;��H;bI;�I;�I;�I;} I;`,I;f:I;(KI;�^I;�uI;��I;��I;�I;�_I;��H;�H;��F;�D;o�A;|�=;g|9;�W4;�.;�);�#;9�;s;�;      ܼ2;�%3;�U4;�16;֍8;L7;;��=;�@;C;�E;T�F;��G;�H;�<I;�I;ɛI;W�I;v�I;�pI;�[I;xII;�9I;`,I;� I;^I;cI;�I;I;��H;��H;��H;j�H;�H;�H;-�H;��H;C�H;��H;.�H;�H;|�H;l�H;��H;��H;��H;I;�I;cI;`I;� I;^,I;�9I;vII;�[I;�pI;y�I;V�I;ɛI;�I;�<I;�H;��G;S�F;}E;C;�@;��=;N7;;ݍ8;�16;�U4;v%3;      @@;�p@;��@;��A;��B;mD;�EE;dgF;�dG;63H;��H;69I;uyI;�I;�I;ۑI;�~I;�iI;�VI;RFI;�7I;=+I;� I;dI;�I;�I;I;��H;�H; �H;a�H;a�H;��H;��H;��H;^�H;=�H;^�H;��H;��H;��H;c�H;a�H;��H;�H;��H;I;�I;�I;aI;� I;=+I;�7I;TFI;�VI;�iI;�~I;ّI;�I;�I;syI;59I;��H;63H;�dG;dgF;�EE;oD;��B;��A;��@;�p@;      �fF;,zF; �F;�G;_sG;{�G;
ZH;��H;�I;�WI;��I;�I;ϝI;�I;�I;BsI;�`I;yPI;�AI;�4I;I)I;>I;�I;`I;�I;�I;-�H;B�H;
�H;��H;t�H;��H;W�H;n�H;��H;N�H;T�H;N�H;��H;n�H;T�H;��H;r�H;��H;�H;B�H;,�H;�I;�I;`I;�I;>I;D)I;�4I;�AI;|PI;�`I;BsI;�I;�I;НI;�I;��I;�WI;�I;��H;
ZH;{�G;csG;�G;!�F;"zF;      i�H;��H;Z�H;2I;�%I;�HI;�hI;H�I;z�I;��I;'�I;�I;2�I;�vI;]fI;�VI;�HI;H<I;�0I;n&I;NI;zI;�I;�I;{I;0�H;H�H;*�H;��H;v�H;��H;5�H;&�H;K�H;��H;S�H;S�H;S�H;��H;K�H;#�H;5�H;��H;u�H;��H;*�H;D�H;/�H;}I;�I;�I;zI;JI;n&I;�0I;I<I;�HI;�VI;_fI;�vI;2�I;�I;'�I;��I;}�I;J�I;�hI;�HI;�%I;1I;Y�H;��H;      ��I;@�I; �I;s�I;�I;�I;d�I;`�I;��I;9�I;��I;XtI;qfI;YI;�LI;�@I;�5I;�+I;�"I;�I;�I;}I;�I;I;��H;D�H;)�H;��H;��H;��H;'�H; �H;�H;B�H;��H;��H;h�H;��H;��H;B�H;�H; �H;)�H;��H;��H;��H;)�H;D�H;��H;I;�I;}I;�I;�I;�"I;�+I;�5I;�@I;�LI;YI;nfI;VtI;��I;9�I;��I;c�I;d�I;�I;��I;r�I;!�I;J�I;      ��I;0�I;�I;ȘI;+�I;�I;��I;r�I;�vI;�kI;*aI;nVI;�KI;�AI;88I;/I;�&I;�I;�I;�I;�I;�I;bI;��H;�H;�H;��H;��H;��H;�H;��H;��H;��H;e�H;�H;��H;��H;��H;�H;g�H;��H;��H;��H;�H;��H;��H;��H;�H;�H;��H;`I;�I;�I;�I;�I;�I;�&I;/I;:8I;�AI; LI;nVI;(aI;�kI;�vI;t�I;��I;�I;2�I;ȘI;�I;(�I;      [|I;�{I;�yI;�vI;MrI;�lI;dfI;Y_I;�WI;�OI;�GI;�?I;�7I;�/I;"(I;.!I;�I;�I;*I;%
I;�I;{I;��H;��H;��H;��H;r�H;��H;�H;��H;��H;��H;>�H;��H;K�H;�H;�H;�H;K�H;��H;;�H;��H;��H;��H;�H;��H;r�H;��H;��H;��H;��H;{I;�I;%
I;*I;�I;�I;.!I;#(I;�/I;�7I;�?I;�GI;�OI;�WI;\_I;dfI;�lI;IrI;�vI;�yI;�{I;      \I;�[I;ZI;�WI;]TI;,PI;`KI;FI;p@I;f:I;74I;�-I;�'I;�!I;"I;�I;~I;�I;3I;7I;� I;B�H;D�H;��H;\�H;r�H;��H;'�H;��H;��H;��H;�H;��H;�H;��H;��H;��H;��H;��H;�H;��H;�H;��H;��H;��H;'�H;��H;r�H;^�H;��H;A�H;B�H;� I;8I;3I;�I;}I;�I;#I;�!I;�'I;�-I;74I;g:I;p@I;FI;^KI;-PI;ZTI;�WI;ZI;�[I;      �CI;�CI;�BI;�@I;%>I;	;I;e7I;K3I;�.I;(*I;f%I;� I;�I;&I;�I;QI;C
I;jI;�I;�H;��H;��H;u�H;m�H;^�H;��H;3�H; �H;��H;��H;
�H;��H;��H;��H;T�H;!�H;�H;!�H;T�H;��H;��H;��H;�H;��H;��H; �H;3�H;��H;a�H;m�H;t�H;��H;��H;�H;�I;mI;C
I;QI;�I;&I;�I;� I;f%I;(*I;�.I;K3I;d7I;
;I;$>I;�@I;�BI;�CI;      F2I;2I;1I;�/I;�-I;P+I;~(I;_%I;"I;\I;�I;�I;
I;2I;�I;I;�I;�I;��H;�H;��H;Z�H;L�H;��H;��H;V�H;#�H;�H;��H;A�H;��H;��H;q�H;,�H;��H;��H;��H;��H;��H;,�H;n�H;��H;��H;B�H;��H;�H;!�H;V�H;��H;��H;J�H;Z�H;��H;�H;��H;�I;�I;"I;�I;2I;	I;�I;�I;]I;"I;a%I;~(I;S+I;�-I;�/I;1I;�1I;      �%I;�%I;�$I;�#I;V"I;P I;I;�I;�I;�I;�I;�I;�I;�	I;�I;�I;� I;�H;��H;z�H;��H;~�H;��H;�H;��H;m�H;G�H;=�H;d�H;��H;�H;��H;'�H;��H;��H;}�H;b�H;}�H;��H;��H;%�H;��H;�H;��H;g�H;?�H;F�H;k�H;��H;�H;��H;~�H;}�H;{�H;��H;�H;� I;�I;�I;�	I;�I;�I;�I;�I;�I;�I;I;T I;K"I;�#I;�$I;�%I;      �I;sI;�I;�I;�I;�I;/I;I;�I;0I;�I;�
I;VI;�I;�I;� I;7�H;��H;��H;��H;��H;"�H;��H;.�H;��H;��H;��H;��H;�H;L�H;��H;V�H;��H;��H;S�H;G�H;P�H;G�H;S�H;��H;��H;Y�H;��H;N�H;�H;��H;��H;��H;��H;.�H;��H;"�H;��H;��H;��H;��H;6�H;� I;�I;�I;WI;�
I;�I;3I;�I;I;0I;�I;�I;�I;�I;jI;      �I;�I;I;KI;0I;�I;I;&I;I;�I;�
I;AI;�I;jI;I;��H;��H;��H;��H;��H;��H;N�H;��H;��H;Z�H;K�H;Q�H;��H;��H;�H;��H;$�H;��H;��H;G�H;/�H;*�H;/�H;G�H;~�H;��H;'�H;��H;�H;��H;��H;P�H;J�H;\�H;��H;��H;O�H;��H;��H;��H;��H;��H;��H;I;hI;�I;AI;�
I;�I;I;&I;I;�I;'I;II;I;�I;      hI;HI;�I;�I;�I;dI;�I;�I;�I;�I;�	I;\I;�I;�I;� I;K�H;)�H;�H;�H;c�H;��H;*�H;��H;C�H;9�H;O�H;N�H;k�H;��H;�H;��H;�H;��H;h�H;P�H;+�H;�H;+�H;P�H;h�H;��H;�H;��H;
�H;��H;k�H;L�H;Q�H;9�H;A�H;��H;*�H;��H;c�H;�H;�H;'�H;K�H;� I;�I;�I;\I;�	I;�I;�I;�I;�I;hI;�I;�I;�I;@I;      �I;�I;I;II;0I;�I;I;&I;I;�I;�
I;AI;�I;jI;I;��H;��H;��H;��H;��H;��H;O�H;��H;��H;\�H;K�H;S�H;��H;��H;�H;��H;$�H;��H;��H;G�H;/�H;*�H;/�H;G�H;~�H;��H;'�H;��H;�H;��H;��H;N�H;J�H;Z�H;��H;��H;N�H;��H;��H;��H;��H;��H;��H;I;hI;�I;AI;�
I;�I;I;&I;I;�I;%I;KI;I;�I;      �I;sI;�I;�I;�I;�I;0I;I;�I;1I;�I;�
I;WI;�I;�I;� I;7�H;��H;��H;��H;��H;"�H;��H;/�H;��H;��H;��H;��H;�H;L�H;��H;V�H;��H;��H;S�H;G�H;P�H;G�H;S�H;��H;��H;[�H;��H;N�H;�H;��H;��H;��H;��H;+�H;��H;"�H;��H;��H;��H;��H;6�H;� I;�I;�I;VI;�
I;�I;1I;�I;I;/I;�I;�I;�I;�I;jI;      �%I;�%I;�$I;�#I;U"I;P I;I;�I;�I;�I;�I;�I;�I;�	I;�I;�I;� I;�H;��H;z�H;��H;~�H;��H;�H;��H;m�H;F�H;?�H;d�H;��H;�H;��H;'�H;��H;��H;}�H;b�H;}�H;��H;��H;%�H;��H;�H;��H;g�H;=�H;F�H;m�H;��H;�H;��H;~�H;}�H;{�H;��H;�H;� I;�I;�I;�	I;�I;�I;�I;�I;�I;�I;I;T I;K"I;�#I;�$I;�%I;      H2I;2I;1I;�/I;�-I;O+I;}(I;^%I;"I;\I;�I;�I;	I;2I;�I;"I;�I;�I;��H;�H;��H;Z�H;L�H;��H;��H;W�H;#�H;�H;��H;A�H;��H;��H;p�H;+�H;��H;��H;��H;��H;��H;+�H;n�H;��H;��H;B�H;��H;�H;!�H;T�H;��H;��H;J�H;Z�H;��H;�H;��H;�I;�I;I;�I;2I;	I;�I;�I;]I;"I;^%I;~(I;R+I;�-I;�/I;1I;2I;      �CI;�CI;�BI;�@I;%>I;;I;g7I;I3I;�.I;(*I;f%I;� I;�I;&I;�I;QI;D
I;mI;�I;��H;��H;��H;u�H;m�H;a�H;��H;3�H; �H;��H;��H;�H;��H;��H;��H;T�H;!�H;�H;!�H;T�H;��H;��H;��H;
�H;��H;��H; �H;3�H;��H;^�H;m�H;t�H;��H;��H;�H;�I;kI;A
I;QI;�I;&I;�I;� I;f%I;)*I;�.I;I3I;g7I;
;I;">I;�@I;�BI;�CI;      \I;�[I;ZI;�WI;]TI;,PI;^KI;FI;p@I;f:I;74I;�-I;�'I;�!I;#I;�I;}I;�I;3I;8I;� I;B�H;D�H;��H;^�H;t�H;��H;'�H;��H;��H;��H;�H;��H;�H;��H;��H;��H;��H;��H;�H;��H;�H;��H;��H;��H;'�H;��H;q�H;\�H;��H;A�H;B�H;� I;7I;3I;�I;}I;�I;"I;�!I;�'I;�-I;54I;g:I;o@I;FI;`KI;-PI;ZTI;�WI;ZI;�[I;      Q|I;�{I;�yI;�vI;HrI;�lI;dfI;Y_I;�WI;�OI;�GI;�?I;�7I;�/I;#(I;.!I;�I;�I;*I;'
I;�I;{I;��H;��H;��H;��H;t�H;��H;�H;��H;��H;��H;<�H;��H;K�H;�H;�H;�H;K�H;��H;<�H;��H;��H;��H;�H;��H;q�H;��H;��H;��H;��H;{I;�I;'
I;*I;�I;�I;/!I;"(I;�/I;�7I;�?I;�GI;�OI;�WI;Z_I;dfI;�lI;IrI;�vI;�yI;�{I;      ��I;,�I;��I;ŘI;1�I;�I;��I;t�I;�vI;�kI;*aI;pVI; LI;�AI;:8I;/I;�&I;�I;�I;�I;�I;�I;bI;��H;�H;�H;��H;��H;��H;�H;��H;��H;��H;g�H;�H;��H;��H;��H;�H;e�H;��H;��H;��H;�H;��H;��H;��H;�H;�H;��H;`I;�I;�I;�I;�I;�I;�&I;/I;88I;�AI;�KI;nVI;*aI;�kI;�vI;u�I;��I;�I;,�I;ØI;��I;,�I;      ��I;=�I;!�I;r�I;�I;�I;d�I;b�I;��I;9�I;��I;VtI;nfI;YI;�LI;�@I;�5I;�+I;�"I;�I;�I;}I;�I;I;��H;D�H;)�H;��H;��H;��H;)�H; �H;�H;@�H;��H;��H;h�H;��H;��H;B�H;�H;�H;'�H;��H;��H;��H;)�H;D�H;��H;I;�I;}I;�I;�I;�"I;�+I;�5I;�@I;�LI;YI;qfI;XtI;�I;9�I;��I;c�I;d�I;�I;��I;s�I;!�I;K�I;      c�H;��H;\�H;,I;�%I;�HI;�hI;H�I;}�I;��I;(�I;�I;2�I;�vI;_fI;�VI;�HI;H<I;�0I;p&I;QI;zI;�I;�I;}I;0�H;G�H;*�H;��H;v�H;��H;5�H;%�H;K�H;��H;S�H;S�H;Q�H;��H;J�H;%�H;7�H;��H;u�H;��H;*�H;D�H;0�H;{I;�I;�I;zI;JI;p&I;�0I;I<I;�HI;�VI;]fI;�vI;2�I;�I;(�I;��I;z�I;H�I;�hI;�HI;�%I;.I;\�H;��H;      �fF;)zF;+�F;�G;`sG;}�G;
ZH;��H;�I;�WI;��I;�I;НI;�I;�I;CsI;�`I;zPI;�AI;�4I;L)I;>I;�I;`I;�I;�I;-�H;B�H;�H;��H;r�H;��H;V�H;n�H;��H;N�H;T�H;N�H;��H;n�H;T�H;��H;t�H;��H;�H;B�H;,�H;�I;�I;`I;�I;>I;D)I;�4I;�AI;zPI;�`I;BsI;�I;�I;НI;�I;��I;�WI;�I;��H;ZH;}�G;csG;�G;+�F;zF;      @@;�p@;��@;��A;��B;mD;�EE;dgF;�dG;73H;��H;59I;syI;�I;�I;ۑI;�~I;�iI;�VI;TFI;�7I;=+I;� I;dI;�I;�I;�I;��H;�H; �H;a�H;a�H;��H;��H;��H;^�H;=�H;^�H;��H;��H;��H;d�H;a�H;��H;�H;��H;}I;�I;�I;cI;� I;=+I;�7I;TFI;�VI;�iI;�~I;ۑI;�I;�I;uyI;69I;��H;53H;�dG;dgF;�EE;mD;��B;��A;��@;�p@;      ߼2;�%3;�U4;�16;ύ8;Q7;;��=;�@;C;�E;S�F;��G;�H;�<I;�I;ɛI;W�I;v�I;�pI;�[I;zII;�9I;`,I;� I;`I;cI;�I;I;��H;��H;��H;j�H;}�H;�H;+�H;��H;C�H;��H;.�H;�H;}�H;l�H;��H;��H;��H;I;�I;cI;^I;� I;^,I;�9I;tII;�[I;�pI;y�I;V�I;țI;�I;�<I;�H;��G;S�F;~E;C;�@;��=;Q7;;ލ8;�16;�U4;u%3;      ��;3�;�;:�;�#;�);�.;�W4;h|9;}�=;n�A;�D;ߟF;�H;��H;�_I;�I;��I;��I;�uI;�^I;(KI;g:I;b,I;} I;�I;�I;�I;dI;��H;F�H;u�H;L�H;��H;��H;��H;��H;��H;��H;��H;J�H;u�H;F�H;��H;bI;�I;�I;�I;| I;`,I;f:I;&KI;�^I;�uI;��I;��I;�I;�_I;��H;�H;��F;�D;n�A;z�=;g|9;�W4;�.;�);�#;;�;y;$�;      ���:���:��:�
�:�+�:��;�;�;��&;��/;}=7;�D=;��A;�E;�7G;��H;�8I;-�I;G�I;�I;?xI;�_I;%KI;�9I;;+I;AI;zI;}I;�I;I;C�H;��H;\�H;~�H;"�H;O�H;)�H;O�H;"�H;}�H;Z�H;��H;C�H;{I;�I;}I;vI;BI;:+I;�9I;"KI;�_I;;xI;�I;G�I;.�I;�8I;��H;�7G;�E;��A;�D=;z=7;��/;��&;�;�;��;�+�:�
�:��:���:      @�x9��9p��9
:��^:� �:Yʼ:Q�:��;�h;�#;�</;�;8;��>;�oC;�fF;z(H;�I;�I;�I;�I;?xI;�^I;{II;�7I;N)I;MI;�I;�I;�I;� I;��H;��H;x�H;��H;��H;��H;��H;��H;x�H;��H;��H;� I;�I;�I;�I;LI;N)I;�7I;wII;�^I;?xI;�I;�I;�I;�I;y(H;�fF;�oC;��>;�;8;�</;�#;�h;��;Q�:[ʼ:�:��^:
:p��9���9      ٯ���������Xct��D�`$�8��&:���:���:�Z;�C;s�&;�'3;X<;��A;"�E;��G;�I;�|I;�I;�I;�uI;�[I;OFI;�4I;p&I;�I;�I;%
I;4I;x�H;�H;v�H;��H;��H;_�H;��H;��H;v�H;�H;y�H;3I;!
I;�I;�I;m&I;�4I;MFI;�[I;�uI;�I;�I;�|I;�I;��G;"�E;��A;W<;�'3;r�&;�C;�Z;���:���:��&:`$�8�D�Dct������ ���      �M����B���jg��c7}�9�D�[���w��������9��:	��:L	;S�;,�.;2�9;+�@;0^E;��G;�I;�I;I�I;��I;�pI;�VI;�AI;�0I;�"I;�I;-I;1I;�I;��H;��H;��H;��H;�H;��H;��H;��H;��H;�I;1I;*I;�I;�"I;�0I;�AI;�VI;�pI;��I;I�I;�I;�I;��G;2^E;(�@;2�9;-�.;S�;L	;	��:��:���9����w��[��4�D�]7}�jg��B�����      ��?��<<���1��h!��z��B�N���n��P�-��ﳺH|���&:ӏ�:���:��;Y�+;�8;{�@;0^E;��G;�I;-�I;��I;v�I;�iI;|PI;J<I;�+I;�I;�I;�I;kI;�I;�H;��H;��H;�H;��H;��H;�H;�I;mI;�I;�I;�I;�+I;H<I;}PI;�iI;q�I;��I;-�I;�I;��G;0^E;{�@;�8;X�+;��;���:׏�:�&:P|���ﳺP�-��n��N���B黫z��h!���1��<<�      ^��L��~I��v�������^��75��z�t�̻�눻kR�Dct���x9���:�m�:i;��*;�8;,�@;%�E;z(H;�8I;�I;Y�I;�~I;�`I;�HI;�5I;�&I;�I;wI;<
I;�I;� I;2�H;��H;#�H;��H;0�H;� I;�I;<
I;wI;�I;�&I;�5I;�HI;�`I;�~I;T�I;��I;�8I;y(H;&�E;+�@;�8;��*;i;�m�:���:��x9@ct�mR��눻t�̻�z��75��^����v���~I��M��      '��`��
�
���Y��EC���t����|���?���	���їV����� �0�:C�:i;\�+;4�9;��A;�fF;��H;�_I;ΛI;ّI;GsI;�VI;�@I;!/I;.!I;�I;KI;I;�I;� I;��H;F�H;��H;� I;�I;I;KI;�I;-!I;/I;�@I;�VI;FsI;ّI;țI;�_I;��H;�fF;��A;4�9;]�+;i;C�:.�:@�����їV�����	���?���|��t��EC��Y��
����
�a�      ��t��p�,�d��Q�{�9�]*����_�ҼvI���o���'��ڻ.6}�����5�,�:�m�:��;,�.;[<;�oC;�7G;��H;�I;�I;�I;`fI;�LI;<8I;"(I; I;�I;�I;�I;�I;	I;� I;	I;�I;�I;�I;�I;I; (I;78I;�LI;]fI;�I;�I;�I;��H;�7G;�oC;]<;,�.;��;�m�:(�:�5����,6}��ڻ��'��o�vI��_�Ҽ���]*�{�9��Q�,�d��p�      ��Ž5���̷�Q���z����}��Q�U�'����$C��%\��"<<�z>�hn����� ����:���:Q�;�'3;��>;�E;�H;�<I;�I;�I;�vI;YI;�AI;�/I;�!I;!I;/I;�	I;�I;aI;�I;aI;�I;�	I;,I;!I;�!I;�/I;�AI;YI;�vI;�I;�I;�<I;�H;�E;��>;�'3;P�;���:���:@����hn��z>�"<<�%\��$C�����U�'��Q���}��z��Q��̷�5���      d.��3�ɤ�W����ΈŽ85�����XG�0��^kּB����xC�z>�+6}�������x9ݏ�:J	;u�&;�;8;��A;�F;��H;wyI;֝I;5�I;rfI;LI;�7I;�'I;�I;	I;�I;QI;�I;�I;�I;QI;�I;I;�I;�'I;�7I; LI;rfI;2�I;֝I;yyI;�H;��F;��A;�;8;u�&;J	;ߏ�:��x9����,6}�z>��xC�B���^kּ0��XG����85��ΈŽ��W��ɤ��3�      Jx��s���d�O�N�a�3�}I����I����z����\�A*��ݼB���#<<��ڻїV�@ct� �&:	��:�C;�</;�D=;�D;��G;59I;�I;�I;UtI;nVI;�?I;�-I;� I;�I;�I;�
I;7I;RI;7I;�
I;�I;�I;� I;�-I;�?I;jVI;TtI;�I;�I;79I;��G;�D;�D=;�</;�C;	��: �&:Lct�ӗV��ڻ#<<�B����ݼA*���\��z��I������}I�a�3�O�N���d��s�      .l¾(��V������������d���7�y��9Sؽ[���d�A*�^kּ&\����'���nR�P|����:�Z;�#;z=7;q�A;W�F;��H;��I;-�I;�I;-aI;�GI;14I;c%I;�I;�I;�I;�
I;�	I;�
I;�I;�I;�I;e%I;14I;�GI;*aI;�I;*�I;��I;��H;Q�F;m�A;z=7;�#;�Z;��:H|��oR�����'�&\��^kּA*��d�[��9Sؽy����7��d���������V���(��      �V������������Ͼ�d���ǆ�E�N��3��c�[����\�0��$C���o���	��눻�ﳺ���9���:�h;��/;~�=;�E;<3H;�WI;��I;:�I;lI;�OI;c:I;(*I;_I;�I;1I;�I;�I;�I;0I;�I;]I;(*I;c:I;�OI;�kI;:�I;��I;�WI;>3H;�E;}�=;��/;�h;���:���9�ﳺ�눻��	��o�$C��0����\�[���cཱ3�E�N��ǆ��d����Ͼ���������      �,b�Ž\��>M���5�=��3r��'l¾Ꝓ�$&W��3�9Sؽ�z��XG����vI����?�t�̻P�-�������:��;��&;g|9;C;�dG;�I;�I;��I;�vI;�WI;i@I;�.I;"I;�I;�I;I;�I;I;�I;�I;�!I;�.I;i@I;�WI;�vI;��I;|�I;�I;�dG;
C;e|9;��&;��;���:���O�-�u�̻��?�vI�����XG��z��9Sؽ�3�$&W�Ꝓ�'l¾3r��=����5��>M�Ž\�      ���&��[���N䂿Ľ\���1�����J˾Ꝓ�E�N�y��I������U�'�_�Ҽ��|��z��n���w����&:Q�:�;�W4;�@;jgF;��H;O�I;_�I;w�I;W_I;FI;G3I;^%I;�I; I; I;�I;!I;�I;�I;^%I;E3I;FI;W_I;r�I;_�I;N�I;��H;kgF;�@;�W4;�;Q�:��&:�w���n���z���|�_�ҼU�'����I���y��E�N�Ꝓ��J˾�����1�Ľ\�N䂿[���&��      !}߿�$ڿ0�ʿ����
����Ps�SX:����'l¾�ǆ���7����85���Q�����t���75�L��^���$�8Sʼ:��;�.;��=;�EE;ZH;�hI;d�I;��I;bfI;\KI;e7I;�(I;I;/I;�I;�I;�I;/I;I;�(I;e7I;ZKI;`fI;��I;d�I;�hI;ZH;�EE;��=;�.;��;Wʼ:�$�8^��L���75��t������Q�85�������7��ǆ�'l¾���SX:��Ps�
�������0�ʿ�$ڿ      |�����p������ſ%���Ps���1�3r���d���d�}I�ΈŽ��}�]*�EC���^��B�<�D��D�� �:��;�);Q7;;mD;��G;�HI;�I;�I;�lI;0PI;;I;V+I;[ I;�I;�I;kI;�I;�I;Z I;S+I;;I;1PI;�lI;�I;�I;�HI;��G;oD;L7;;�);��; �:�D�<�D��B��^�EC��]*���}�ΈŽ}I��d��d��3r����1��Ps�%����ſ��꿄p����      ��7��3�آ%�|��<����ſ
���Ľ\�=����Ͼ����a�3��轻z��{�9�Y�ἓ���z�Z7}�\ct���^:�+�:�#;ٍ8;��B;bsG;�%I;�I;2�I;ArI;STI;$>I;�-I;Q"I;�I;%I;�I;%I;�I;Q"I;�-I;$>I;STI;>rI;.�I;�I;�%I;`sG;��B;֍8;��#;�+�:��^:\ct�\7}��z����Y��{�9��z����a�3�������Ͼ=��Ľ\�
�����ſ�<��|�آ%��3�      /�_��+Y��lG� f.�|���꿳���N䂿��5���󾎰��O�N�W��Q���Q�
���u����h!�jg����,
:�
�:A�;�16;��A;�G;/I;x�I;ŘI;�vI;�WI;�@I;�/I;�#I;�I;II;�I;II;�I;�#I;�/I;�@I;�WI;�vI;I;v�I;.I;�G;��A;�16;D�;�
�:4
:��jg���h!�v���
����Q�Q��W��O�N���������5�N䂿�������|� f.��lG��+Y�      Ҭ��%}�?tf��lG�آ%��p�0�ʿ\����>M����V�����d�ɤ�̷�-�d��
�~I����1�G������0��9���:r;�U4;��@;0�F;^�H;�I;��I;�yI;�YI;�BI;1I;�$I;�I;I;�I;I;�I;�$I;1I;BI;�YI;�yI;��I;�I;^�H;0�F;��@;�U4;u;���:8��9���G�����1�~I���
�-�d�̷�ɤ���d�V�������>M�\���0�ʿ�p�آ%��lG�?tf�%}�      T���E���%}��+Y��3�����$ڿ&��Ž\����(���s��3�5����p�`�M���<<���������9���:(�;u%3;�p@;zF;��H;<�I;3�I;�{I;�[I;�CI;�1I;�%I;cI;�I;AI;�I;eI;�%I;�1I;�CI;�[I;�{I;0�I;<�I;��H;zF;�p@;s%3;.�;���:���9������<<�N��`��p�5����3��s�(�����Ž\�&���$ڿ����3��+Y�%}�E���      ����,������U���K�Q�Ǚ$�6�����>�}�I(�A�׾�T���L+���սj����L���iO���ͻ?�� .m8�o�:��;~�1;�?;/vF;� I;��I;��I;��I;�vI;�WI;BI;22I;(I;"I;. I;"I;(I;22I;BI;�WI;�vI;��I;��I;��I;� I;/vF;�?;z�1;��;�o�:�.m8@����ͻ�iO�L����j����ս�L+��T��A�׾I(�>�}���6���Ǚ$�K�Q�U��������,��      �,��b��$P���{���K��x �����r�����w��$���Ҿg��� (���ѽѷ��$����ҔK�%ɻܟ� ��8��:��;��1;8@;ʊF;NI;�I;V�I;�I;�uI;mWI;�AI;�1I;�'I;�!I; I;�!I;�'I;�1I;�AI;nWI;�uI;��I;S�I;!�I;NI;ʊF;7@;��1;��;��: ��8ݟ�%ɻҔK����$�ѷ����ѽ (�g�����Ҿ�$���w�r��������x ���K��{�$P��b��      ����$P�������d���;�$���㿴���#f�e�� ž��z���=�ƽ#0v�R5�*����o@�f���,i�0du9�K�:j];83;j�@;?�F;yI;��I;��I;��I;tI;VI;�@I;#1I;('I;L!I;oI;L!I;&'I;#1I;�@I;VI;tI;��I;��I;��I;wI;?�F;j�@;83;m];�K�:0du9-i�f����o@�*���R5�#0v�=�ƽ����z� že��#f�������$����;���d����$P��      U����{���d��F�Ǚ$�;����ɿ/蒿��K�R���j�� Zb�G�2���q�a����8�����.�~d����غ���9-Z�:�X;�25;k�A;�!G;|7I;��I;��I;��I;�pI;�SI;�>I;�/I;�%I;b I;qI;b I;�%I;�/I;�>I;�SI;�pI;��I;��I;��I;{7I;�!G;j�A;�25;�X;-Z�:���9��غ~d����.�8������q�a�2���G� Zb��j��R����K�/蒿��ɿ;��Ǚ$��F���d��{�      K�Q���K���;�Ǚ$��;
��޿�����w�s,���澞���(�D������I��"�G����N��v�����������9:ڨ�:o!;¶7;�B;��G;*ZI;n�I;��I;��I;�lI;�PI;V<I;�-I;S$I; I;	I; I;Q$I;�-I;V<I;�PI;�lI;�I;��I;n�I;*ZI;��G;�B;��7;o!;ڨ�:��9:�������u���N�����"�G��I������(�D��������s,���w�����޿�;
�Ǚ$���;���K�      Ǚ$��x �$��;���޿q���˅���F�~�
��~����z��$���ս���>2+���ϼPp�n����]��*����:Y�;'9';ތ:;B�C;QH;�}I;`�I;��I;�I;�gI;�LI;\9I;y+I;f"I;5I;jI;5I;f"I;y+I;\9I;�LI;�gI;�I;��I;b�I;�}I;PH;@�C;ڌ:;'9';Y�;���:�*��]�m���Pp���ϼ>2+������ս�$���z��~��~�
��F�˅��q����޿;��$���x �      6��������㿌�ɿ���˅����P�e��=�׾�`��U�H����@��Q�a���ơ���D��ɻ� ��έ�SX�:�;�I-;p|=;jCE;�H;I�I;�I;��I;�I;�aI;eHI;�5I;�(I; I;I;�I;I; I;�(I;�5I;eHI;�aI;�I;��I;!�I;I�I;�H;iCE;l|=;�I-;�;WX�: ϭ�� ��ɻ�D�ơ����P�a��@����U�H��`��=�׾e����P�˅�������ɿ�㿵���      ��r�������/蒿��w��F�e��̰�!����Yb�*����ѽ�%��D4�ԟ�X��y���G��>潺8��9�r�:1 ;+:3;cQ@;�vF;^�H;I�I;��I;ΤI;�zI;	[I;UCI;�1I;�%I;�I;�I;dI;�I;�I;�%I;�1I;VCI;	[I;�zI;̤I;��I;H�I;^�H;�vF;_Q@;+:3;1 ;�r�:0��9>潺�G��z��X��ԟ�D4��%����ѽ*���Yb�!���̰�e���F���w�/蒿����r���      >�}���w�#f���K�s,�~�
�=�׾!�����k���'�fz꽝I���;V�:M�����iO�JG�.oE�������:�� ;�$;��8;��B;D�G;|KI;U�I;Z�I;��I;GqI;�SI;�=I;�-I;H"I;�I;XI;�I;XI;�I;H"I;�-I;�=I;�SI;GqI;��I;Z�I;S�I;|KI;A�G;��B;��8;�$;�� ;���:���-oE�JGໜiO����:M��;V��I��fz���'���k�!���=�׾~�
�s,���K�#f���w�      I(��$�e��R������~���`���Yb���'��U�H$��B�m�#����ϼ�/��.�������غ�:�9���:3G; H.;\|=;�E; ]H;f�I;��I;��I;=�I;BgI;BLI;'8I;I)I;�I;�I;�I;jI;�I;�I;�I;G)I;)8I;CLI;BgI;:�I;��I;��I;f�I;�\H;�E;[|=; H.;3G;���:�:�9�غ����.���/����ϼ#��B�m�H$���U���'��Yb��`���~�����R��e���$�      A�׾��Ҿž�j��������z�U�H�*��fz�H$���/v�2+�ؐ�����5��ɻ�4�0&��:���:~o!;TP6;PlA;%�F;��H;ַI;��I;!�I;�}I;�\I;�DI;G2I;�$I; I;�I;�I;�I;�I;�I;I;�$I;J2I;�DI;�\I;�}I;!�I;��I;طI;��H;!�F;NlA;TP6;|o!;���::&���4��ɻ��5���ؐ�2+��/v�H$��gz�*��U�H���z������j��ž��Ҿ      �T��g�����z� Zb�(�D��$�����ѽ�I��B�m�2+�������<�K���W�p�����Ȕ�9�T�:0;��-;��<;�zD;�H;�mI;*�I;��I;ҕI;�oI;�RI;�<I;B,I; I;NI;sI;�I;	I;�I;wI;PI; I;E,I;�<I;�RI;�oI;ԕI;��I;,�I;�mI;�H;�zD;��<;��-;0;�T�:���9Ɩ��W�p���<�K�������2+�B�m��I����ѽ���$�(�D� Zb���z�g���      �L+� (���G�������ս�@���%���;V�#��א�����pMS�>�����C�@	o8�q�:;��$;E_7;r�A;��F;=�H;��I;��I;ʭI;#�I;�bI;�HI;P5I;f&I;qI;I;/I;I;H
I;I;/I;�I;oI;g&I;P5I;�HI;�bI;#�I;ɭI;��I;��I;;�H;��F;t�A;E_7;��$;;�q�: 	o8�C���>��pMS�����א�#���;V��%���@����ս����G��� (�      ��ս��ѽ=�ƽ2����I�����P�a�D4�9M���ϼ��<�K�>��-G��f���o�$��:^C�:�Y;&�1;�l>;#E;.0H;aqI;F�I;.�I;�I;GsI;�UI;0?I;�-I;� I;�I;�I;I;TI;vI;TI;I;�I;�I;� I;�-I;2?I;�UI;GsI;�I;0�I;F�I;^qI;,0H;$E;�l>;(�1;�Y;fC�:��:��o�f�,G��>��<�K�����ϼ9M�D4�P�a�����I��2���<�ƽ��ѽ      j��ѷ��#0v�q�a�"�G�>2+���ԟ�����/����5�����f��֬��g:��:K�;[I-;`g;;COC;NSG;�I;�I;c�I;C�I;J�I;NcI;�II;6I;�&I;
I;xI;#I;�I;�I;�I;�I;�I;&I;xI;I;�&I;6I;�II;PcI;J�I;F�I;d�I;	�I;�I;OSG;COC;cg;;[I-;N�;��:�g:�֬�f�������5��/�����ԟ���>2+�"�G�q�a�#0v�ѷ��      ��$�R5���������ϼš��X���iO�.���ɻX�p��C���o��g:u`�:�G;�*;�9;	�A;�uF;a�H;
�I;��I;�I;��I;�pI;yTI;�>I;^-I;�I;�I;:I;�I;�I;�I;I;�I;�I;�I;9I;�I;�I;_-I;�>I;yTI;�pI;��I;�I;��I;�I;c�H;�uF;	�A;�9;�*;�G;u`�:�g:��o��C�X�p��ɻ/���iO�X��š����ϼ������Q5�%�      L�����*���8����N��Pp��D�x��JG໽����4������	o8 ��:��:�G;H�(;޶7;��@;�E;�QH;]mI;��I;=�I;ߢI;j}I;�^I;�FI;4I;&%I;�I;�I;3
I;PI; I;) I;��H;* I;!I;QI;2
I;�I;�I;&%I;4I;�FI;�^I;l}I;�I;:�I;��I;]mI;�QH;�E;��@;�7;H�(;�G;��: ��:�	o8���4�����IG�x���D�Pp��N��8���*������      �iO�ҔK��o@���.�v��r����ɻ�G��*oE��غ&�����9�q�:^C�:K�;�*;޶7;�P@; ]E;5H;JI;ŽI;��I;O�I;��I;�hI;�NI;�:I;*I;�I;�I;I;YI;OI;q�H;��H;�H;��H;q�H;QI;XI;"I;�I;�I;|*I;�:I;�NI;�hI;��I;M�I;��I;ŽI;JI;7H;]E;�P@;ܶ7;�*;M�;^C�:�q�:���9&���غ,oE��G���ɻp���u����.��o@�ԔK�      ��ͻ$ɻa���~d������]�� �D潺���p:�9:�T�:;�Y;[I-;�9;��@; ]E;��G;w5I;��I;��I;�I;��I;�pI;�UI;�@I;x/I;�!I;�I;�I;�I;�I;`�H;��H;W�H;��H;W�H;��H;c�H;�I;�I;�I;�I;�!I;x/I;�@I;�UI;�pI;��I;�I;��I;��I;z5I;��G;]E;��@;�9;^I-;�Y;;�T�::p:�9���B潺� ��]����~d��a���$ɻ      =��˟�-i���غ������*�@ϭ���9���:���:���:0;��$;!�1;^g;;�A;�E;4H;v5I;�I;��I;��I;ڗI;�vI;�[I;�EI;�3I;w%I;�I;�I;�	I;�I;��H;��H;f�H;*�H;��H;+�H;f�H;��H;��H;�I;�	I;�I;�I;x%I;�3I;�EI;�[I;�vI;חI;��I;��I;��I;w5I;5H;�E;�A;^g;;!�1;��$;0;���:���:���:��9@ϭ��*�������غ,i�ԟ�      �/m8���8pdu9X��9\�9:���:WX�:�r�:�� ;1G;zo!;��-;B_7;�l>;BOC;�uF;�QH;JI;��I;��I;��I;��I;�zI;�_I;�II;�7I;�(I;�I;I;`I;(I;i I;��H;��H;B�H;%�H;��H;%�H;B�H;��H;��H;k I;(I;^I;I;�I;�(I;�7I;�II;�_I;�zI;��I;�I;��I;��I;JI;�QH;�uF;BOC;�l>;B_7;��-;zo!;0G;�� ;�r�:SX�:���:d�9:h��9`du9`��8      �o�:!��:�K�:Z�:Ҩ�:`�;�;3 ;�$;H.;VP6;��<;o�A; E;LSG;_�H;[mI;ŽI;��I;��I;��I;'|I;�aI;�KI;�9I;#+I;�I;�I;�I;jI;1I;5�H;�H;��H;0�H;P�H;�H;P�H;0�H;��H;�H;5�H;1I;gI;�I;�I;�I;&+I;�9I;�KI;�aI;)|I;��I;��I;��I;ƽI;ZmI;]�H;OSG;!E;o�A;��<;TP6;H.;�$;6 ;�;a�;���:Z�:�K�:��:      ��;��;k];{X;o!;'9';�I-;':3;��8;[|=;NlA;�zD;��F;00H;�I;�I;��I;��I; �I;ۗI;�zI;�aI;�LI;a;I;�,I;u I;gI;9I;}I;I;��H;?�H;��H;��H;I�H;��H;d�H;��H;J�H;��H;��H;?�H;��H;I;{I;:I;dI;w I;�,I;^;I;�LI;�aI;�zI;ޗI;�I;��I;��I;�I;�I;.0H;��F;�zD;NlA;Y|=;��8;(:3;�I-;)9';o!;{X;m];��;      ��1;��1;83;�25;��7;ڌ:;t|=;\Q@;��B;�E;#�F;�H;8�H;^qI;�I;��I;:�I;P�I;��I;�vI;�_I;�KI;^;I;-I;.!I;]I;I;ZI;�I;:�H;��H;��H;f�H;��H;��H;�H;��H;�H;��H;��H;e�H;��H;��H;9�H;�I;ZI;I;^I;/!I;-I;^;I;�KI;�_I;�vI;��I;R�I;8�I;��I;�I;_qI;6�H;�H;!�F;�E;��B;_Q@;s|=;ی:;ƶ7;�25;83;��1;      �?;?@;U�@;m�A;�B;@�C;fCE;�vF;@�G;�\H;��H;�mI;��I;F�I;c�I;�I;�I;��I;�pI;�[I;�II;�9I;�,I;4!I;�I;�I;�I;9I;��H;��H;��H;j�H;��H;0�H;/�H;��H;p�H;��H;/�H;0�H;��H;m�H;��H;��H;��H;:I;�I;�I;�I;1!I;�,I;�9I;�II;�[I;�pI;��I;�I;�I;c�I;D�I;��I;�mI;��H;�\H;@�G;�vF;eCE;B�C;�B;m�A;S�@;>@;      :vF;ڊF;.�F;�!G;��G;GH;�H;W�H;zKI;c�I;ӷI;*�I;��I;,�I;@�I;��I;j}I;�hI;�UI;�EI;�7I;"+I;r I;ZI;�I;	I;�I;��H;0�H;�H;i�H;}�H;��H;��H;��H;Y�H;*�H;Y�H;��H;��H;��H;�H;i�H;
�H;/�H;��H;�I;	I;�I;ZI;r I;"+I;�7I;�EI;�UI;�hI;i}I;��I;B�I;.�I;��I;*�I;ӷI;a�I;yKI;X�H;�H;GH;��G;�!G;.�F;ϊF;      � I;NI;rI;7I;*ZI;�}I;K�I;B�I;U�I;��I;��I;��I;ŭI;�I;I�I;�pI;�^I;�NI;�@I;�3I;�(I;�I;fI;I;�I;�I;�H;e�H;�H;w�H;g�H;��H;Z�H;\�H;��H;G�H;�H;G�H;��H;Z�H;X�H;��H;g�H;v�H;�H;e�H;�H;�I;�I;I;dI;�I;�(I;�3I;�@I;�NI;�^I;�pI;I�I;�I;ŭI;��I;��I;��I;U�I;D�I;K�I;�}I;.ZI;~7I;tI;PI;      ��I;$�I;��I;��I;k�I;_�I;�I;��I;Z�I;��I;$�I;ՕI;"�I;GsI;OcI;wTI;�FI;�:I;v/I;x%I;�I;�I;:I;[I;6I;��H;d�H;;�H;��H;g�H;��H;"�H;�H;F�H;��H;B�H;1�H;C�H;��H;F�H;�H;"�H;��H;d�H;��H;<�H;d�H;��H;7I;]I;:I;�I;�I;x%I;u/I;�:I;�FI;wTI;NcI;EsI;�I;ՕI;"�I;��I;]�I;��I;�I;_�I;u�I;��I;��I;0�I;      �I;R�I;��I;��I;��I;��I;��I;ˤI;��I;8�I;�}I;�oI;�bI;�UI;�II;�>I; 4I;{*I;�!I;�I;I;�I;{I;�I;��H;2�H;�H;��H;m�H;��H;�H;��H;��H;<�H;��H;u�H;l�H;v�H;��H;<�H;��H;��H;�H;��H;n�H;��H;�H;0�H;��H;�I;yI;�I;I;�I;�!I;|*I;4I;�>I;�II;�UI;�bI;�oI;�}I;8�I;��I;ˤI;��I;��I;��I;��I;��I;H�I;      şI;�I;��I;��I;�I;�I;��I;�zI;MqI;GgI;�\I;�RI;�HI;6?I;6I;_-I;(%I;�I;�I;�I;`I;gI;I;9�H;��H;�H;s�H;d�H;��H;�H;��H;��H;��H;`�H;��H;��H;��H;��H;��H;`�H;��H;��H;��H;�H;��H;e�H;s�H;�H;��H;:�H;I;gI;`I;�I;�I;�I;'%I;_-I;	6I;6?I;�HI;�RI; ]I;GgI;MqI;�zI;��I;�I;��I;��I;��I;�I;      �vI;vI;tI;qI;�lI;�gI;�aI;
[I;�SI;ELI;�DI;�<I;S5I;�-I;�&I;�I;�I;�I;�I;�	I;.I;1I;��H;��H;��H;i�H;c�H;��H;�H;��H;��H;��H;*�H;��H;L�H;�H;��H;�H;L�H;��H;'�H;��H;��H;��H;�H;��H;d�H;i�H;��H;��H;��H;1I;*I;�	I;�I;�I;�I;�I;�&I;�-I;S5I;�<I;�DI;HLI;�SI;[I;�aI;�gI;�lI;qI;tI;vI;      �WI;vWI;VI;�SI;�PI;�LI;aHI;WCI;�=I;'8I;J2I;J,I;g&I;� I;I;�I;�I;I;�I;�I;p I;8�H;@�H;��H;i�H;}�H;��H; �H;��H;��H;��H;&�H;��H;�H;��H;��H;��H;��H;��H;�H;��H;'�H;��H;��H;��H;"�H;��H;|�H;l�H;��H;=�H;8�H;n I;�I;�I;"I;�I;�I;I;� I;f&I;I,I;J2I;'8I;�=I;WCI;`HI;�LI;�PI;�SI;VI;rWI;      BI;�AI;�@I;�>I;[<I;X9I;�5I;�1I;�-I;D)I;�$I;
 I;oI;�I;zI;:I;7
I;RI;�I;��H;��H;�H;��H;i�H;��H;��H;[�H;�H;��H;��H;,�H;��H;��H;��H;K�H;!�H;)�H;!�H;K�H;��H;��H;��H;,�H;��H;��H;�H;X�H;��H;��H;i�H;��H;�H;��H;��H;�I;TI;6
I;<I;zI;�I;nI; I;�$I;F)I;�-I;�1I;�5I;Z9I;T<I;�>I;�@I;�AI;      <2I;�1I;1I;�/I;�-I;q+I;�(I;�%I;K"I;�I;I;UI;�I;�I;'I;�I;WI;NI;e�H;��H;��H;��H;��H;��H;,�H;��H;W�H;C�H;9�H;]�H;��H;�H;��H;2�H;�H;��H;��H;��H;�H;2�H;��H;�H;��H;^�H;<�H;C�H;W�H;��H;/�H;��H;��H;��H;��H;��H;e�H;OI;UI;�I;'I;�I;�I;UI;I;�I;M"I;�%I;�(I;u+I;�-I;�/I;1I;�1I;      (I;�'I;*'I;�%I;e$I;]"I; I;�I;�I;�I;�I;~I;3I;	I; I;�I;'I;m�H;��H;k�H;J�H;2�H;I�H;��H;(�H;��H;��H;��H;��H;��H;L�H;��H;K�H;�H;��H;��H;��H;��H;��H;	�H;H�H;��H;L�H;��H;��H;��H;��H;��H;(�H;��H;H�H;2�H;H�H;k�H;��H;m�H;%I;�I;I;	I;3I;~I;�I;�I;�I;�I; I;`"I;[$I;�%I;*'I;�'I;      "I;�!I;P!I;b I;I;-I;!I;�I;bI;�I;�I;�I;"I;]I;�I;�I;1 I;��H;\�H;/�H;-�H;P�H;��H;�H;��H;W�H;F�H;@�H;v�H;��H;�H;��H; �H;��H;��H;o�H;i�H;o�H;��H;��H;�H;��H;�H;��H;w�H;@�H;F�H;V�H;��H;�H;��H;P�H;,�H;1�H;\�H;��H;. I;�I;�I;[I;"I;�I;�I;�I;bI;�I;!I;1I;I;a I;P!I;�!I;      ' I; I;xI;rI;I;cI;�I;dI;�I;dI;�I;I;J
I;|I;�I;I;��H;�H;��H;��H;��H;�H;c�H;��H;l�H;(�H;�H;4�H;n�H;��H;��H;��H;+�H;��H;��H;j�H;P�H;j�H;��H;��H;'�H;��H;��H;��H;p�H;4�H;	�H;)�H;l�H;��H;c�H;�H;��H;��H;��H;�H;��H;I;�I;|I;J
I;I;�I;gI;�I;dI;�I;hI;I;rI;xI; I;      "I;�!I;P!I;a I;I;-I;!I;�I;cI;�I;�I;�I;"I;]I;�I;�I;1 I;��H;\�H;/�H;/�H;P�H;��H;�H;��H;W�H;G�H;@�H;v�H;��H;�H;��H; �H;��H;��H;o�H;i�H;o�H;��H;��H;�H;��H;�H;��H;w�H;@�H;C�H;V�H;��H;�H;��H;P�H;,�H;1�H;\�H;��H;. I;�I;�I;[I;"I;�I;�I;�I;bI;�I;!I;1I;I;b I;M!I;�!I;      (I;�'I;)'I;�%I;e$I;]"I; I;�I;�I;�I;�I;~I;3I;	I;I;�I;'I;m�H;��H;k�H;L�H;2�H;I�H;��H;(�H;��H;��H;��H;��H;��H;L�H;��H;K�H;	�H;��H;��H;��H;��H;��H;�H;H�H;��H;L�H;��H;��H;��H;��H;��H;(�H;��H;H�H;2�H;H�H;k�H;��H;m�H;%I;�I; I;	I;3I;~I;�I;�I;�I;�I; I;`"I;[$I;�%I;)'I;�'I;      =2I;�1I;1I;�/I;�-I;q+I;�(I;�%I;K"I;�I;I;UI;�I;�I;'I;�I;WI;NI;e�H;��H;�H;��H;��H;��H;/�H;��H;W�H;C�H;;�H;]�H;��H;�H;��H;2�H;�H;��H;��H;��H;�H;2�H;��H;�H;��H;^�H;<�H;C�H;W�H;��H;,�H;��H;��H;��H;��H;��H;e�H;OI;UI;�I;'I;�I;�I;UI;I;�I;M"I;�%I;�(I;u+I;�-I;�/I;1I;�1I;      BI;�AI;�@I;�>I;Z<I;W9I;�5I;�1I;�-I;D)I;�$I; I;nI;�I;zI;<I;9
I;RI;�I;��H;��H;�H;��H;i�H;��H;��H;[�H;�H;��H;��H;,�H;��H;��H;��H;K�H;!�H;)�H;!�H;K�H;��H;��H;��H;,�H;��H;��H;�H;W�H;��H;��H;h�H;��H;�H;��H;��H;�I;RI;5
I;:I;zI;�I;nI;
 I;�$I;F)I;�-I;�1I;�5I;Z9I;T<I;�>I;�@I;�AI;      �WI;vWI;VI;�SI;�PI;�LI;bHI;WCI;�=I;'8I;J2I;I,I;f&I;� I;I;�I;�I; I;�I;�I;s I;8�H;@�H;��H;l�H;}�H;��H;"�H;��H;��H;��H;&�H;��H;�H;��H;��H;��H;��H;��H;�H;��H;'�H;��H;��H;��H; �H;��H;|�H;i�H;��H;?�H;8�H;n I;�I;�I; I;�I;�I;I;� I;g&I;J,I;J2I;)8I;�=I;WCI;bHI;�LI;�PI;�SI;VI;tWI;      �vI;vI;tI;qI;�lI;�gI;�aI;
[I;�SI;FLI;�DI;�<I;S5I;�-I;�&I;�I;�I;�I;�I;�	I;/I;1I;��H;��H;��H;j�H;d�H;��H;�H;��H;��H;��H;)�H;��H;L�H;�H;��H;�H;L�H;��H;'�H;��H;��H;��H;�H;��H;c�H;h�H;��H;��H;��H;1I;*I;�	I;�I;�I;�I;�I;�&I;�-I;S5I;�<I;�DI;FLI;�SI;
[I;�aI;�gI;�lI;qI;tI;vI;      ��I;�I;��I;��I;��I;�I;��I;�zI;NqI;EgI; ]I;�RI;�HI;7?I;	6I;_-I;(%I;�I;�I;�I;dI;gI;I;9�H;��H;�H;t�H;e�H;��H;�H;��H;��H;��H;^�H;��H;��H;��H;��H;��H;`�H;��H;��H;��H;�H;��H;d�H;q�H;�H;��H;:�H;	I;gI;^I;�I;�I;�I;'%I;a-I;6I;6?I;�HI;�RI;�\I;EgI;NqI;�zI;��I;�I;��I;��I;��I;�I;      	�I;N�I;��I;��I;��I;��I;��I;ˤI;��I;8�I;�}I;�oI;�bI;�UI;�II;�>I; 4I;|*I;�!I;�I;I;�I;|I;�I;��H;2�H;�H;��H;n�H;��H;�H;��H;��H;<�H;��H;v�H;l�H;u�H;��H;<�H;��H;��H;�H;��H;m�H;��H;�H;0�H;��H;�I;yI;�I;I;�I;�!I;|*I;4I;�>I;�II;�UI;�bI;�oI;�}I;7�I;��I;ΤI;��I;��I;��I;��I;��I;O�I;      ��I;"�I;��I;��I;h�I;_�I;�I;��I;[�I;��I;$�I;ՕI;�I;GsI;OcI;wTI;�FI;�:I;u/I;x%I;�I;�I;<I;]I;7I;��H;d�H;<�H;��H;g�H;��H;"�H;�H;D�H;��H;B�H;1�H;C�H;��H;F�H;�H;#�H;��H;d�H;��H;;�H;d�H;��H;6I;[I;9I;�I;�I;x%I;v/I;�:I;�FI;yTI;OcI;EsI;"�I;֕I;"�I;��I;Z�I;��I;�I;\�I;v�I;��I;��I;0�I;      � I;MI;uI;z7I;&ZI;�}I;I�I;B�I;U�I;��I;��I;��I;ŭI;�I;I�I;�pI;�^I;�NI;�@I;�3I;�(I;�I;fI;I;�I;�I;�H;e�H;�H;w�H;g�H;��H;Z�H;Z�H;��H;G�H;�H;F�H;��H;Z�H;X�H;��H;g�H;v�H;�H;e�H;�H;�I;�I;I;dI;�I;�(I;�3I;�@I;�NI;�^I;�pI;I�I;�I;ŭI;��I;��I;��I;S�I;B�I;I�I;�}I;*ZI;z7I;tI;DI;      ?vF;ԊF;9�F;�!G;��G;HH;�H;W�H;yKI;c�I;ӷI;)�I;��I;.�I;@�I;��I;j}I;�hI;�UI;�EI;�7I;"+I;r I;ZI;�I;	I;�I;��H;0�H;�H;i�H;}�H;��H;��H;��H;Y�H;*�H;Y�H;��H;��H;��H;�H;i�H;�H;/�H;��H;�I;	I;�I;ZI;r I;"+I;�7I;�EI;�UI;�hI;i}I;��I;@�I;.�I;��I;*�I;ӷI;`�I;wKI;W�H;�H;GH;��G;�!G;9�F;̊F;      �?;?@;U�@;m�A;�B;@�C;eCE;�vF;@�G;�\H;��H;�mI;��I;D�I;c�I;�I;�I;��I;�pI;�[I;�II;�9I;�,I;4!I;�I;�I;�I;:I;��H;��H;��H;l�H;��H;0�H;.�H;��H;p�H;��H;/�H;/�H;��H;m�H;��H;��H;��H;9I;�I;�I;�I;2!I;�,I;�9I;�II;�[I;�pI;��I;�I;�I;c�I;D�I;��I;�mI;��H;�\H;?�G;�vF;fCE;@�C;�B;m�A;S�@;?@;      ��1;��1;83;�25;��7;��:;p|=;]Q@;��B;�E;!�F;�H;9�H;_qI;�I;��I;:�I;P�I;��I;�vI;�_I;�KI;a;I;-I;/!I;^I;I;ZI;�I;<�H;��H;��H;f�H;��H;��H;�H;��H;�H;��H;��H;e�H;��H;��H;7�H;�I;ZI;I;]I;.!I;-I;];I;�KI;�_I;�vI;��I;R�I;8�I;��I;�I;_qI;8�H;�H;!�F;�E;��B;]Q@;p|=;��:;ɶ7;�25;83;��1;      ��;��;|];{X;o!;*9';�I-;':3;��8;[|=;NlA;�zD;��F;.0H;�I;�I;��I;��I;�I;ۗI;�zI;�aI;�LI;a;I;�,I;v I;fI;:I;}I;I;��H;?�H;��H;��H;J�H;��H;d�H;��H;I�H;��H;��H;?�H;��H;I;{I;9I;cI;v I;�,I;^;I;�LI;�aI;�zI;ޗI;�I;��I;��I;�I;�I;00H;��F;�zD;PlA;Y|=;��8;':3;�I-;+9';o!;|X;q];��;      �o�:��:�K�:Z�:Ҩ�:`�;�;3 ;�$;H.;VP6;��<;o�A;!E;NSG;_�H;ZmI;ŽI;��I;��I;��I;)|I;�aI;�KI;�9I;&+I;�I;�I;�I;kI;1I;5�H;�H;��H;0�H;P�H;�H;P�H;0�H;��H;�H;5�H;1I;gI;�I;�I;�I;%+I;�9I;�KI;�aI;'|I;��I;��I;��I;ƽI;ZmI;_�H;NSG;!E;o�A;��<;TP6;H.;�$;5 ;�;`�;���:Z�:�K�:��:      �-m8���8�du9h��9\�9:���:YX�:�r�:�� ;0G;|o!;��-;B_7;�l>;BOC;�uF;�QH;JI;��I;��I;��I;��I;�zI;�_I;�II;�7I;�(I;�I;I;`I;(I;i I;��H;��H;B�H;%�H;��H;%�H;B�H;��H;��H;k I;(I;]I;I;�I;�(I;�7I;�II;�_I;�zI;��I;�I;��I;��I;JI;�QH;�uF;BOC;�l>;B_7;��-;|o!;.G;�� ;�r�:YX�:���:x�9:h��9�du9`��8      ?��ʟ�)i���غ������*�@ϭ� ��9���:���:���:0;��$;!�1;\g;;�A;�E;4H;w5I;�I;��I;��I;ۗI;�vI;�[I;�EI;�3I;x%I;�I;�I;�	I;�I;��H;��H;f�H;+�H;��H;+�H;f�H;��H;��H;�I;�	I;�I;�I;w%I;�3I;�EI;�[I;�vI;חI;��I;��I;��I;v5I;5H;�E;�A;^g;;!�1;��$;0;���:���:���:��9@ϭ��*�������غ,i�՟�      ��ͻ$ɻa���~d������]�� �D潺���p:�9:�T�:;�Y;]I-;�9;��@;]E;��G;y5I;��I;��I; �I;��I;�pI;�UI;�@I;x/I;�!I;�I;�I;�I;�I;c�H;��H;W�H;��H;W�H;��H;`�H;�I;�I;�I;�I;�!I;x/I;�@I;�UI;�pI;��I;�I;��I;��I;y5I;��G;]E;��@;�9;]I-;�Y;;�T�::p:�9���D潺� ��]����~d��a���$ɻ      �iO�ҔK��o@���.�v��s����ɻ�G��,oE��غ&�����9�q�:\C�:M�;�*;޶7;�P@;]E;5H;JI;ŽI;��I;R�I;��I;�hI;�NI;�:I;*I;�I;�I;I;YI;QI;q�H;��H;�H;��H;q�H;OI;XI; I;�I;�I;|*I;�:I;�NI;�hI;��I;I�I;��I;ŽI;JI;7H; ]E;�P@;ݶ7;�*;K�;^C�:�q�:���9&���غ,oE��G���ɻp���u����.��o@�ԔK�      L�����*���8����N��Pp��D�x��JG໾����4����	o8 ��:��:�G;I�(;�7;��@;�E;�QH;]mI;��I;>�I;�I;j}I;�^I;�FI; 4I;'%I;�I;�I;3
I;QI;!I;) I;��H;) I; I;QI;2
I;�I;�I;$%I;4I;�FI;�^I;l}I;ߢI;8�I;��I;]mI;�QH;�E;��@;�7;H�(;�G;��:$��:�	o8�����4�����IG�x���D�Pp��N��8���*������      ��$�R5���������ϼš��X���iO�.���ɻX�p��C���o��g:u`�:�G;�*;�9;	�A;�uF;c�H;	�I;��I;�I;��I;�pI;yTI;�>I;_-I;�I;�I;:I;�I;�I;�I;I;�I;�I;�I;9I;�I;�I;^-I;�>I;yTI;�pI;��I;�I;��I;�I;a�H;�uF;	�A;�9;�*;�G;u`�:�g:��o��C�X�p��ɻ.���iO�X��š����ϼ������R5�%�      j��ѷ��#0v�q�a�"�G�>2+���ԟ�����/����5�����f��֬��g:��:K�;[I-;bg;;COC;OSG;�I;�I;d�I;E�I;L�I;PcI;�II;6I;�&I;I;zI;&I;�I;�I;�I;�I;�I;%I;xI;I;�&I;6I;�II;NcI;I�I;E�I;c�I;�I;�I;NSG;BOC;bg;;[I-;N�;��:�g:�֬�f�������5��/�����ԟ���>2+�"�G�q�a�#0v�ѷ��      ��ս��ѽ=�ƽ2����I�����P�a�D4�9M���ϼ��<�K�>��-G��f���o�$��:dC�:�Y;&�1;�l>;$E;00H;bqI;F�I;/�I;�I;GsI;�UI;0?I;�-I;� I;�I;�I;I;TI;vI;TI;I;�I;�I;� I;�-I;0?I;�UI;GsI;�I;/�I;F�I;^qI;*0H;#E;�l>;&�1;�Y;dC�: ��:��o�f�,G��>��<�K�����ϼ9M�D4�P�a�����I��2���=�ƽ��ѽ      �L+� (���G�������ս�@���%���;V�#��א�����pMS�>�����C⺀	o8�q�:;��$;D_7;t�A;��F;?�H;��I;��I;ʭI;#�I;�bI;�HI;P5I;f&I;oI;�I;/I;I;H
I;I;/I;I;oI;f&I;P5I;�HI;�bI;#�I;ȭI;��I;��I;6�H;��F;r�A;D_7;��$;;�q�:@	o8�C���>��pMS�����א�#���;V��%���@����ս����G��� (�      �T��g�����z� Zb�(�D��$�����ѽ�I��B�m�2+�������<�K���W�p�����Д�9�T�:0;��-;��<;�zD;�H;�mI;,�I;��I;ԕI;�oI;�RI;�<I;B,I; I;RI;wI;�I;	I;�I;sI;NI; I;C,I;�<I;�RI;�oI;ҕI;��I;*�I;�mI;�H;�zD;��<;��-;0;�T�:���9��Z�p���<�K�������2+�B�m��I����ѽ���$�(�D� Zb���z�g���      A�׾��Ҿž�j��������z�U�H�*��gz�H$���/v�2+�ؐ�����5��ɻ�4�(&��:���:|o!;TP6;QlA;%�F;��H;طI;��I;!�I;�}I;�\I;�DI;G2I;�$I;I;�I;�I;�I;�I;�I; I;�$I;H2I;�DI;�\I;�}I;!�I;��I;ַI;��H; �F;NlA;TP6;|o!;���::&���4��ɻ��5���ؐ�2+��/v�H$��fz�*��U�H���z������j��ž��Ҿ      I(��$�e��R������~���`���Yb���'��U�H$��B�m�#����ϼ�/��.�������غ�:�9���:1G; H.;\|=;�E;�\H;g�I;��I;��I;=�I;BgI;CLI;'8I;I)I;�I;�I;�I;jI;�I;�I;�I;G)I;'8I;BLI;BgI;:�I;��I;��I;f�I; ]H;�E;[|=; H.;1G;���:�:�9�غ����.���/����ϼ#��B�m�H$���U���'��Yb��`���~�����R��e���$�      >�}���w�#f���K�s,�~�
�=�׾!�����k���'�fz꽝I���;V�:M�����iO�JG�-oE�������:�� ;�$;��8;��B;A�G;}KI;V�I;Z�I;��I;FqI;�SI;�=I;�-I;H"I;�I;XI;�I;XI;�I;H"I;�-I;�=I;�SI;FqI;��I;Z�I;S�I;|KI;D�G;��B;��8;�$;�� ;���:���,oE�KGໜiO����:M��;V��I��fz���'���k�!���=�׾~�
�s,���K�#f���w�      ��r�������/蒿��w��F�e��̰�!����Yb�*����ѽ�%��D4�ԟ�X��y���G��>潺8��9�r�:1 ;+:3;bQ@;�vF;_�H;I�I;��I;ϤI;�zI;	[I;UCI;�1I;�%I;�I;�I;dI;�I;�I;�%I;�1I;SCI;	[I;�zI;̤I;��I;H�I;\�H;�vF;_Q@;+:3;1 ;�r�: ��9>潺�G��z��X��ԟ�D4��%����ѽ*���Yb�!���̰�e���F���w�/蒿����r���      6��������㿌�ɿ���˅����P�e��=�׾�`��U�H����@��Q�a���ơ���D��ɻ� ��έ�QX�:�;�I-;p|=;iCE;�H;I�I;!�I;��I;�I;�aI;eHI;�5I;�(I; I;I;�I;I; I;�(I;�5I;dHI;�aI;�I;��I;�I;H�I;�H;jCE;m|=;�I-;�;WX�: ϭ�� ��ɻ�D�ơ����P�a��@����U�H��`��=�׾e����P�˅�������ɿ�㿵���      Ǚ$��x �$��;���޿q���˅���F�~�
��~����z��$���ս���>2+���ϼPp�n����]��*����:Y�;&9';ތ:;@�C;QH;�}I;b�I;��I;�I;�gI;�LI;\9I;y+I;f"I;5I;jI;6I;f"I;y+I;[9I;�LI;�gI;�I;��I;`�I;�}I;PH;B�C;ڌ:;'9';Y�;���:�*��]�m���Pp���ϼ>2+������ս�$���z��~��~�
��F�˅��q����޿;��$���x �      K�Q���K���;�Ǚ$��;
��޿�����w�s,���澞���(�D������I��"�G����N��v���������x�9:ڨ�:o!;¶7;�B;��G;(ZI;n�I;��I;��I;�lI;�PI;V<I;�-I;S$I; I;	I; I;Q$I;�-I;T<I;�PI;�lI;�I;��I;n�I;+ZI;��G;�B;��7;o!;ڨ�:��9:�������u���N�����"�G��I������(�D��������s,���w�����޿�;
�Ǚ$���;���K�      U����{���d��F�Ǚ$�;����ɿ/蒿��K�R���j�� Zb�G�2���q�a����8�����.�~d����غ���9-Z�:�X;�25;j�A;�!G;{7I;��I;��I;��I;�pI;�SI;�>I;�/I;�%I;b I;qI;b I;�%I;�/I;�>I;�SI;�pI;��I;��I;��I;|7I;�!G;k�A;�25;�X;-Z�:���9��غ~d����.�8������q�a�2���G� Zb��j��R����K�/蒿��ɿ;��Ǚ$��F���d��{�      ����$P�������d���;�$���㿴���#f�e�� ž��z���=�ƽ#0v�R5�*����o@�f���-i� du9�K�:j];83;j�@;?�F;xI;��I;��I;��I;tI;VI;�@I;#1I;('I;L!I;oI;L!I;('I;#1I;�@I;VI;tI;��I;��I;��I;xI;?�F;j�@;83;m];�K�:0du9-i�f����o@�*���R5�#0v�=�ƽ����z� že��#f�������$����;���d����$P��      �,��b��$P���{���K��x �����r�����w��$���Ҿg��� (���ѽѷ��$����ҔK�%ɻܟ� ��8��:��;��1;7@;ʊF;NI;!�I;U�I;�I;�uI;mWI;�AI;�1I;�'I;�!I; I;�!I;�'I;�1I;�AI;nWI;�uI;��I;U�I;�I;MI;ʊF;8@;��1;��;��: ��8ݟ�%ɻҔK����$�ѷ����ѽ (�g�����Ҿ�$���w�r��������x ���K��{�$P��b��      E(��r'���o��O�d��X1�x�Ŀ����3�x���x����4�l��Y+���'���ü(yY��kٻ�o&���p����:�;�0;Ͷ?;�F;� I;@�I;�I;e�I;��I;�dI;�KI;:I;�.I;�'I;	&I;�'I;�.I;:I;�KI;�dI;��I;d�I;	�I;@�I;� I;�F;Ͷ?;�0;�;���:��p��o&��kٻ(yY���ü�'�Y+��l�ཾ�4��x��x���3����Ŀx��X1�d�O��o��r'��      r'���X��g^�������]]���,�Q9�7g��U�����/����o��h1��hܽ��~-$�Xl���|U�D�Ի0!� �,���:2;�51;�?;��F;q'I;��I;\�I;w�I;�I;dI;�KI;�9I;f.I;�'I;�%I;�'I;g.I;�9I;KI;dI;�I;t�I;Y�I;��I;q'I;��F;�?;�51;8;��: �,�1!�D�Ի�|U�Yl��~-$����hܽh1��o���ྛ�/�U���7g��Q9���,��]]�����g^���X��      �o��g^���ē��4z�6K�i��T��(ﱿV�v��X#���Ѿń��&�p�нb̀�]��n���:�I�jǻx4�&9]�:��;O�2;Ӆ@;(�F;';I;4�I;@�I;ײI;��I;�bI;?JI;�8I;�-I;�&I;%I;�&I;�-I;�8I;=JI;�bI;��I;ԲI;?�I;4�I;';I;(�F;Ӆ@;K�2;��;]�: &9z4�kǻ:�I�n���]��b̀�p�н�&�ń���Ѿ�X#�V�v�(ﱿT��i��6K��4z��ē�g^��      O������4z���V��X1��<�uؿ����RZ��	�*���KUo����^y��,l�W��R��2�7�𻱻n���ǳ9x��:)�;��4;�tA;�2G;�XI;��I;��I;E�I;8�I;`I;<HI;c7I;>,I;�%I;�#I;�%I;>,I;d7I;;HI;`I;8�I;D�I;��I;��I;�XI;�2G;�tA;��4;,�;x��:�ǳ9p��𻱻2�7��R��W�,l�^y�����KUo�*����	��RZ����uؿ�<��X1���V��4z�����      d��]]�6K��X1�[f��oQ��U���]58��A���נ���O���_什�Q����8ߓ��� �rV���尺��":W��:V ;&17;N�B;��G;*|I;&�I;��I;�I;}|I;|\I;�EI;\5I;x*I;o$I;k"I;o$I;w*I;^5I;�EI;|\I;}|I;�I;��I;&�I;+|I;��G;N�B;"17;X ;W��:��":�尺rV���� �8ߓ�����Q�_什����O��נ��A��]58�U���oQ���[f��X1�6K��]]�      �X1���,�i���<��6g��f_���U�΂�׌Ⱦ
ń�+�-�i��P ��$�2�?ټR�{��!�sn��O���u:2Q ;&;f#:;��C;H&H;T�I;g�I;�I;�I;�vI;XI;0BI;�2I;T(I;�"I;� I;�"I;T(I;�2I;0BI;XI;�vI;�I;�I;g�I;S�I;F&H;��C;_#:;&;2Q ;��u:�O�qn��!�S�{�?ټ$�2�P ��i��+�-�
ń�׌Ⱦ΂��U�f_��6g��<�i����,�      x�Q9�T��uؿoQ��f_��8�_��X#�r���f��;�S�{�����l�@�w���M�x�Ի��+�8T��:�e;],;50=;�BE;��H;��I;!�I;��I;��I;�oI;	SI;T>I;�/I;�%I;3 I;�I;3 I;�%I;�/I;U>I;
SI;�oI;�I;��I;!�I;��I;��H;�BE;10=;],;�e; �:@8T���+�v�Ի�M�w��@�l�����{�;�S��f��r���X#�8�_�f_��oQ��uؿT��Q9�      Ŀ7g��(ﱿ���U����U��X#�v��f���JUo��#��hܽ����n<����5���}� ��᝻��Ժw�9��:�V;�2;!@;��F;"I;<�I;��I;o�I;��I;ChI;PMI;�9I;0,I;�"I;�I;I;�I;�"I;0,I;�9I;SMI;ChI;��I;l�I;��I;;�I;"I;��F;!@;�2;�V;��: w�9��Ժ�᝻}� �4�������n<�����hܽ�#�JUo�f���v���X#��U�U������(ﱿ7g��      ���U���V�v��RZ�]58�΂�r��f���hoy�^1�`O��[什�`�L�����`yY���O�T��1���u:���:�#;\98;K�B;��G;:mI;R�I;A�I;q�I;��I;`I;DGI;55I;g(I;�I;�I;NI;�I;�I;h(I;55I;EGI;`I;��I;n�I;C�I;O�I;:mI;��G;H�B;\98;�#;���:��u:�1�N�T���`yY����L���`�[什`O��^1�hoy�f���r��΂�]58��RZ�V�v�U���      �3���/��X#��	��A��׌Ⱦ�f��JUo�^1�̰��|n��Ҽx��'��>ټ�@���k��������P�39=$�:sR;Pe-;0=;
E;�xH;ͯI;S�I;��I;F�I;TvI;�WI;�@I;50I;e$I;�I;�I;zI;�I;�I;g$I;50I;�@I;�WI;UvI;C�I;��I;S�I;ͯI;�xH;
E;0=;Pe-;sR;9$�:P�39��𺬼���k��@���>ټ�'�Ҽx�|n��̰��^1�JUo��f��׌Ⱦ�A���	��X#���/�      x���྅�Ѿ)����נ�
ń�;�S��#�`O��|n��Ì���2����s�>�߾ԻH�B��#�Pm:hH�:� ;޼5;�FA;��F;�I;��I;��I;�I;��I;�jI;�NI;O:I;!+I;< I;I;�I;�I;�I;I;> I;+I;R:I; OI;�jI;��I;�I;��I;��I;�I;��F;�FA;�5;� ;fH�:Pm:�#�I�B�޾Իs�>�������2�Ì�|n��`O���#�;�S�
ń��נ�*�����Ѿ��      �x���o��ń�KUo���O�+�-�{��hܽ[什Ҽx���2�mb��NR��G|U�:2�����鰺�w�9C�:YD;��,;i<;�rD;�%H;�I;��I;#�I;I�I;M�I;_I;JFI;�3I;�%I;I;�I;�I;yI;�I;�I;I;�%I;�3I;KFI;_I;L�I;I�I;$�I;��I;�I;�%H;�rD;i<; �,;XD;C�:�w�9�鰺��:2��G|U�NR��nb����2�Ҽx�[什�hܽ{�+�-���O�KUo�ń��o��      ��4�h1��&������i�ཅ�������`��'���NR��6�]�o���U��tX���6o�,��:��;r#;^�6;�tA;��F;�	I;��I;�I;��I;\�I; qI;�SI;�=I;	-I;� I;�I;I;�I;~I;�I;I;�I;� I;-I;�=I;�SI;!qI;]�I;��I; �I;��I;�	I;��F;�tA;^�6;t#;��;4��:�6o�nX���U��p��6�]�NR����'��`��������i��������&�h1�      k�ླྀhܽp�н]y��_什P ��l��n<�K���>ټ��F|U�o������E1�������u:�l�:M�;�71;�)>;�	E;SJH;��I;��I;��I;+�I;�I;�bI;�HI;j5I;�&I;�I;�I;I;cI;`
I;cI;I;�I;�I;�&I;l5I;�HI;�bI; �I;+�I;��I;��I;��I;RJH;�	E;�)>;�71;M�;�l�:��u:����B1�����p��F|U��𛼺>ټK���n<�l�P ��_什^y��p�н�hܽ      X+����b̀�,l��Q�#�2�@��������@��s�>�:2���U��G1����%R:1��:(;�\,;�;;1<C;�eG;�9I;��I;z�I;�I;��I;�qI;�TI;�>I;z-I;n I;�I;�I;I;SI;RI;SI;I;�I;�I;s I;}-I;�>I;�TI;�qI;��I;�I;z�I;��I;�9I;�eG;0<C;�;;�\,;*;/��:%R:x��G1��U��:2��s�>��@��������@�#�2��Q�,l�b̀���      �'�~-$�\��W� ���?ټw��5���_yY��k�޾Ի��pX������%R:��:�R;�);"�8;ΡA;рF;z�H;p�I;��I;��I;�I;L�I;aI;7HI;�4I;�%I;�I;I;�I;�I;SI;�I;TI;�I;�I;I;�I;�%I;�4I;3HI;aI;J�I;�I;��I;��I;l�I;z�H;΀F;ΡA;"�8;�);�R;��:%R:����tX����޾Ի�k�_yY�5���w��?ټ���W�\��~-$�      ��üWl��n����R��8ߓ�R�{��M�|� � �컪���E�B��鰺�6o���u:1��:�R;u�';Y17;�@;C�E;�lH;v�I;��I;��I;N�I;��I;mI;�QI;l<I;�+I;�I;I;�I;&I;�I;kI;�I;kI;�I;'I;�I;I;�I;�+I;k<I;�QI;	mI;��I;O�I;��I;��I;v�I;�lH;F�E;�@;[17;u�';�R;5��:��u:�6o��鰺F�B����� ��|� ��M�R�{�7ߓ��R��n���Xl��      *yY��|U�:�I�1�7��� ��!�v�Ի�᝻N�T����#��w�9,��:�l�:(;�);W17;o @;]E;%H;�kI;O�I;��I;;�I;r�I;�wI;�ZI;�CI;�1I;�#I;kI;�I;q	I;�I;xI;��H;A�H;��H;xI;�I;q	I;�I;kI;�#I;�1I;�CI;�ZI;�wI;r�I;8�I;��I;Q�I;�kI;	%H;�]E;r @;V17;�);*;�l�:,��:�w�9�#����O�T��᝻x�Ի�!��� �1�7�:�I��|U�      �kٻD�Իfǻ𻱻tV��ln���+���Ժ�1�p�39\m:E�:��;O�;�\,; �8; �@;]E;�
H;�VI;��I;3�I;5�I;��I;I�I;�bI;�JI;h7I;(I;�I;rI;I;{I;xI;��H;&�H;��H;&�H;��H;zI;{I;I;rI;�I;(I;j7I;�JI;�bI;I�I;��I;1�I;3�I;��I;�VI;�
H;�]E;��@;"�8;�\,;O�;��;E�:\m:P�39�1���Ժ��+�gn�qV��𻱻fǻD�Ի      �o&�!�z4�v���尺��O�@8T��v�9��u:9$�:fH�:TD;p#;�71;~;;ǡA;A�E;%H;�VI;U�I;��I;Y�I;ĭI;A�I;SiI;oPI;d<I;;,I;cI;I;I;�I;�I;q�H;�H;��H;H�H;��H;�H;r�H;�I;�I;	I;I;^I;;,I;a<I;oPI;UiI;<�I;��I;Z�I;��I;W�I;�VI;%H;A�E;ȡA;~;;�71;p#;UD;fH�:3$�:��u:�v�9`8T��O��尺x��z4�'!�      @�p� ~,�`&9�ǳ9܍":��u: �:��:���:qR;� ;��,;\�6;�)>;/<C;̀F;�lH;�kI;��I;��I;��I;^�I;��I;�mI;�TI;n@I;�/I;f"I;�I;�I;I;�I;��H;��H;��H;��H;�H;��H;��H;��H;��H;�I;I;�I;�I;g"I;�/I;n@I;�TI;�mI;��I;^�I;��I;��I;��I;�kI;�lH;̀F;/<C;�)>;\�6;��,;� ;pR;���:��:�:��u:��":�ǳ9P&9 �,�      ���:#�:}�:j��:O��::Q ;�e;�V;�#;Oe-;�5;i<;�tA;�	E;�eG;v�H;u�I;N�I;1�I;Z�I;\�I;:�I;LpI;�WI;4CI;�2I;�$I;�I;�I;�	I;�I;:�H;��H;C�H;��H;p�H;�H;p�H;��H;C�H;��H;;�H;�I;�	I;�I;�I;�$I;�2I;6CI;�WI;HpI;<�I;Z�I;\�I;3�I;Q�I;r�I;u�H;�eG;�	E;�tA;i<;�5;Me-;�#;�V;�e;:Q ;y��:j��:}�:�:      �;4;��;#�;N ;&;],;�2;`98;0=;�FA;�rD;��F;SJH;�9I;l�I;��I;��I;5�I;ǭI;��I;MpI;�XI;�DI;-4I;�&I;gI;+I;�
I;�I;��H;��H;-�H;�H;z�H;��H;O�H;��H;{�H;�H;+�H;��H;��H;�I;�
I;+I;dI;�&I;14I;�DI;�XI;MpI;��I;ɭI;5�I;��I;��I;k�I;�9I;SJH;��F;�rD;�FA;0=;_98;�2;],;&;T ;#�;��;&;      #�0;�51;V�2;��4;#17;b#:;:0=; !@;K�B;
E;��F;�%H;�	I;��I;��I;��I;��I;=�I;��I;<�I;�mI;�WI;�DI;�4I;�'I;vI;EI;�I;xI;r I;r�H;#�H;��H;��H;��H;��H;��H;��H;��H;��H;��H;&�H;s�H;r I;xI;�I;DI;vI;�'I;�4I;�DI;�WI;�mI;>�I;��I;?�I;��I;��I;��I;��I;�	I;�%H;��F;
E;K�B;!@;80=;b#:;*17;��4;S�2;�51;      ٶ?;�?;��@;�tA;K�B;��C;�BE;��F;��G;�xH;�I;�I;��I;��I;y�I;��I;R�I;q�I;M�I;WiI;�TI;7CI;34I;�'I;�I;�I;WI;"I;� I;��H;X�H;��H;��H;�H;�H;h�H;4�H;i�H;�H;�H;��H;��H;Z�H;��H;� I;$I;WI;�I;�I;�'I;14I;9CI;�TI;ZiI;M�I;t�I;Q�I;��I;y�I;��I;��I;�I;�I;�xH;��G;��F;�BE;��C;K�B;�tA;��@;�?;      &�F;��F;�F;�2G;��G;?&H;��H;I;8mI;ǯI;��I;��I;�I;��I;�I;�I;��I;�wI;�bI;kPI;h@I;�2I;�&I;uI;�I;�I;cI;BI;�H;��H;��H;��H;��H;i�H;��H;�H;��H;�H;��H;i�H;��H;��H;��H;��H;�H;CI;cI;�I;�I;sI;�&I;�2I;d@I;lPI;�bI;�wI;��I;�I;�I;��I;�I;��I;��I;ƯI;8mI;I;��H;?&H;��G;�2G;�F;��F;      � I;q'I;!;I;�XI;(|I;V�I;��I;5�I;P�I;P�I;��I;$�I;��I;)�I;��I;I�I;mI;�ZI;�JI;b<I;�/I;�$I;eI;EI;SI;fI;JI;.�H;��H;��H;��H;��H;�H;�H;W�H;��H;��H;��H;V�H;�H;�H;��H;��H;��H;��H;/�H;II;dI;XI;EI;dI;�$I;�/I;b<I;�JI;�ZI;mI;G�I;��I;)�I;��I;$�I;��I;N�I;R�I;7�I;��I;S�I;-|I;�XI;!;I;p'I;      4�I;��I;7�I;��I;#�I;d�I;�I;��I;D�I;��I;�I;K�I;Z�I;�I;�qI;aI;�QI;�CI;g7I;;,I;f"I;�I;,I;�I; I;DI;.�H;��H;��H;��H;��H;��H;��H;��H;�H;��H;��H;��H;�H;��H;��H;��H;��H;��H;��H;��H;.�H;DI;"I;�I;,I;�I;c"I;<,I;g7I;�CI;�QI;aI;�qI;�I;Y�I;K�I;�I;��I;D�I;��I;�I;d�I;-�I;��I;5�I;��I;      �I;V�I;8�I;��I;��I;	�I;��I;k�I;o�I;B�I;��I;M�I;qI;�bI;�TI;3HI;o<I;�1I;(I;aI;�I;�I;�
I;{I;� I;�H;��H;��H;��H;��H;��H;��H;��H;��H;*�H;��H;��H;��H;*�H;��H;��H;��H;��H;��H;��H;��H;��H;�H;� I;}I;�
I;�I;�I;aI;(I;�1I;n<I;4HI;�TI;�bI;qI;M�I;��I;@�I;o�I;k�I;��I;	�I;��I;��I;8�I;K�I;      k�I;{�I;ڲI;D�I;��I;!�I;��I;��I;��I;XvI;�jI;%_I;�SI;�HI;�>I;�4I;�+I;�#I;�I;I;�I;�	I;�I;r I;��H;��H;��H;��H;��H;��H;n�H;U�H;x�H;��H;Q�H;�H;��H;�H;Q�H;��H;v�H;V�H;o�H;��H;��H;��H;��H;��H;��H;r I;�I;�	I;�I;	I;�I;�#I;�+I;�4I;�>I;�HI;�SI;&_I;�jI;XvI;��I;��I;��I;!�I;��I;E�I;ֲI;x�I;      ��I;�I;��I;?�I;�|I;�vI;�oI;ChI;#`I;�WI;OI;RFI;�=I;o5I;~-I;�%I;�I;hI;tI;I;I;�I;��H;s�H;T�H;��H;��H;��H;��H;q�H;N�H;Q�H;��H;
�H;��H;r�H;4�H;r�H;��H;
�H;��H;S�H;N�H;o�H;��H;��H;��H;��H;W�H;u�H;��H;�I;I;I;uI;iI;�I;�%I;~-I;m5I;�=I;RFI;OI;�WI;"`I;EhI;�oI;�vI;�|I;?�I;��I;�I;      �dI;#dI;�bI;
`I;z\I;XI;SI;SMI;EGI;�@I;R:I;�3I;-I;�&I;u I;�I;I;�I;#I;�I;�I;>�H; �H;&�H;��H;��H;��H;��H;��H;U�H;N�H;��H;��H;h�H;�H;��H;��H;��H;�H;h�H;��H;��H;P�H;V�H;��H;��H;��H;��H;��H;&�H;��H;>�H;�I;�I;#I;�I;I;�I;u I;�&I;-I;�3I;R:I;�@I;EGI;SMI;SI;XI;y\I;
`I;�bI;dI;      �KI;�KI;@JI;BHI;�EI;,BI;M>I;�9I;85I;10I;!+I;�%I;� I;�I;�I;I;�I;j	I;~I;�I;��H;��H;+�H;��H;��H;��H;�H;��H;��H;{�H;��H;��H;R�H;��H;��H;]�H;k�H;]�H;��H;��H;O�H;��H;��H;}�H;��H;��H;�H;��H;��H;��H;*�H;��H;��H;�I;~I;l	I;�I;I;�I;�I;� I;�%I;!+I;30I;65I;�9I;M>I;.BI;�EI;BHI;@JI;�KI;      :I;�9I;�8I;j7I;a5I;�2I;�/I;3,I;i(I;d$I;A I;I;�I;�I;�I;�I;-I;�I;~I;w�H;��H;C�H;�H;��H;�H;h�H; �H;��H;��H;��H;�H;g�H;��H;{�H;9�H;�H;��H;�H;9�H;{�H;��H;j�H;�H;��H;��H;��H; �H;f�H;�H;��H;�H;C�H;��H;x�H;~I;�I;-I;�I;�I;�I;�I;I;? I;d$I;k(I;5,I;�/I;�2I;W5I;j7I;�8I;�9I;      �.I;t.I;�-I;E,I;�*I;M(I;�%I;�"I;�I;�I;I;�I;I;�I;I;�I;�I;sI;��H;�H;��H;��H;z�H;��H;�H;��H;S�H;�H;(�H;Q�H;��H;�H;��H;:�H;��H;��H;��H;��H;��H;<�H;��H;�H;��H;S�H;+�H;�H;S�H;��H;�H;��H;x�H;��H;��H;�H;��H;tI;�I;�I;I;�I;I;�I;I;�I;�I;�"I;�%I;P(I;�*I;E,I;�-I;k.I;      �'I;�'I; 'I;�%I;|$I;{"I;5 I;�I;�I;�I;�I;�I;�I;kI;WI;WI;rI;��H;+�H;��H;��H;p�H;��H;��H;e�H;�H;��H;��H;��H;�H;r�H;��H;[�H;�H;��H;��H;��H;��H;��H;�H;Y�H;��H;r�H;�H;��H;��H;��H;�H;f�H;��H;��H;p�H;��H;��H;+�H;��H;qI;XI;WI;jI;�I;�I;�I;�I;�I;�I;5 I;"I;r$I;�%I; 'I;�'I;      &I;�%I;%I;�#I;r"I;� I;�I;I;PI;tI;�I;~I;I;f
I;SI;�I;�I;7�H;��H;M�H;�H;�H;M�H;��H;1�H;��H;��H;��H;��H;��H;9�H;��H;m�H;��H;��H;��H;��H;��H;��H;��H;j�H;��H;9�H;��H;��H;��H;��H;��H;1�H;��H;M�H;�H;�H;M�H;��H;9�H;�I;�I;SI;f
I;I;~I;�I;wI;PI;I;�I;� I;g"I;�#I;%I;�%I;      �'I;�'I; 'I;�%I;|$I;z"I;5 I;�I;�I;�I;�I;�I;�I;kI;WI;XI;rI;��H;+�H;��H;��H;p�H;��H;��H;f�H;�H;��H;��H;��H;�H;r�H;��H;[�H;�H;��H;��H;��H;��H;��H;�H;Y�H;��H;r�H;�H;��H;��H;��H;�H;e�H;��H;��H;p�H;��H;��H;+�H;��H;qI;WI;WI;jI;�I;�I;�I;�I;�I;�I;5 I;"I;p$I;�%I;�&I;�'I;      �.I;u.I;�-I;C,I;�*I;M(I;�%I;�"I;�I;�I;I;�I;I;�I;I;�I;�I;sI;��H;�H;��H;��H;z�H;��H;�H;��H;U�H;�H;*�H;Q�H;��H;�H;��H;<�H;��H;��H;��H;��H;��H;:�H;��H;�H;��H;S�H;+�H;�H;R�H;��H;�H;��H;z�H;��H;��H;�H;��H;tI;�I;�I;I;�I;I;�I;I;�I;�I;�"I;�%I;P(I;�*I;E,I;�-I;k.I;      :I;�9I;�8I;j7I;a5I;�2I;�/I;3,I;i(I;d$I;A I;I;�I;�I;�I;�I;.I;�I;~I;w�H;��H;C�H;�H;��H;�H;h�H;�H;��H;��H;��H;�H;g�H;��H;{�H;9�H;�H;��H;�H;9�H;{�H;��H;j�H;�H;��H;��H;��H;��H;h�H;�H;��H;�H;C�H;��H;w�H;~I;�I;,I;�I;�I;�I;�I;I;A I;d$I;k(I;5,I;�/I;�2I;U5I;j7I;�8I;�9I;      �KI;�KI;AJI;CHI;�EI;+BI;M>I;�9I;85I;10I;!+I;�%I;� I;�I;�I;I;�I;j	I;~I;�I;��H;��H;+�H;��H;��H;��H;�H;��H;��H;{�H;��H;��H;P�H;��H;��H;\�H;k�H;]�H;��H;��H;O�H;��H;��H;}�H;��H;��H;�H;��H;��H;��H;*�H;��H;��H;�I;~I;j	I;�I;I;�I;�I;� I;�%I;!+I;30I;85I;�9I;M>I;,BI;�EI;CHI;?JI;�KI;      �dI;#dI;�bI;
`I;z\I;XI;SI;SMI;EGI;�@I;R:I;�3I;-I;�&I;u I;�I;I;�I;#I;�I;�I;>�H; �H;&�H;��H;��H;��H;��H;��H;U�H;P�H;��H;��H;h�H;�H;��H;��H;��H;�H;h�H;��H;��H;N�H;V�H;��H;��H;��H;��H;��H;&�H;��H;>�H;�I;�I;#I;�I;I;�I;u I;�&I;-I;�3I;R:I;�@I;GGI;SMI;SI;XI;w\I;
`I;�bI;dI;      ��I;�I;��I;?�I;�|I;�vI;�oI;ChI;"`I;�WI;OI;RFI;�=I;o5I;~-I;�%I;�I;iI;uI;I;I;�I;��H;u�H;W�H;��H;��H;��H;��H;q�H;N�H;Q�H;��H;
�H;��H;r�H;4�H;r�H;��H;
�H;��H;S�H;N�H;o�H;��H;��H;��H;��H;T�H;u�H;��H;�I;I;I;tI;hI;�I;�%I;~-I;p5I;�=I;RFI;OI;�WI;"`I;EhI;�oI;�vI;�|I;?�I;��I;�I;      b�I;{�I;ٲI;D�I;��I;�I;��I;��I;��I;VvI;�jI;%_I;�SI;�HI;�>I;�4I;�+I;�#I;�I;I;�I;�	I;�I;r I;��H;��H;��H;��H;��H;��H;o�H;U�H;w�H;��H;Q�H;�H;��H;�H;Q�H;��H;w�H;V�H;n�H;��H;��H;��H;��H;��H;��H;r I;�I;�	I;�I;I;�I;�#I;�+I;�4I;�>I;�HI;�SI;&_I;�jI;VvI;��I;��I;��I; �I;��I;D�I;ٲI;|�I;      �I;R�I;?�I;��I;��I;�I;��I;k�I;n�I;B�I;��I;M�I;qI;�bI;�TI;4HI;o<I;�1I;(I;cI;�I;�I;�
I;{I;� I;�H;��H;��H;��H;��H;��H;��H;��H;��H;(�H;��H;��H;��H;*�H;��H;��H;��H;��H;��H;��H;��H;��H;�H;� I;}I;�
I;�I;�I;aI;(I;�1I;n<I;4HI;�TI;�bI;qI;M�I;��I;B�I;o�I;l�I;��I;�I;��I;��I;=�I;R�I;      4�I;��I;7�I;��I;"�I;d�I;�I;��I;D�I;��I;�I;K�I;Y�I; �I;�qI;aI;�QI;�CI;g7I;<,I;i"I;�I;.I;�I;"I;DI;.�H;��H;��H;��H;��H;��H;��H;��H;�H;��H;��H;��H;�H;��H;��H;��H;��H;��H;��H;��H;.�H;DI; I;�I;+I;�I;c"I;<,I;g7I;�CI;�QI;aI;�qI;�I;Z�I;L�I;�I;��I;D�I;��I;�I;a�I;/�I;��I;5�I;��I;      � I;p'I;#;I;�XI;&|I;R�I;��I;5�I;R�I;P�I;��I;$�I;��I;)�I;��I;I�I;mI;�ZI;�JI;d<I;�/I;�$I;gI;GI;XI;fI;JI;/�H;��H;��H;��H;��H;�H;�H;V�H;��H;��H;��H;W�H;�H;�H;��H;��H;��H;��H;.�H;II;fI;SI;DI;cI;�$I;�/I;b<I;�JI;�ZI;mI;G�I;��I;*�I;��I;$�I;��I;P�I;P�I;5�I;��I;P�I;(|I;�XI;!;I;f'I;      *�F;��F;%�F;�2G;��G;A&H;��H;I;7mI;ǯI;��I;��I;�I;��I;�I;�I;��I;�wI;�bI;lPI;i@I;�2I;�&I;sI;�I;�I;dI;CI;�H;��H;��H;��H;��H;i�H;��H;�H;��H;�H;��H;i�H;��H;��H;��H;��H;�H;BI;bI;�I;�I;sI;�&I;�2I;d@I;kPI;�bI;�wI;��I;�I;�I;��I;�I;��I;��I;ƯI;7mI;I;��H;?&H;��G;�2G;$�F;��F;      ٶ?;�?;��@;�tA;K�B;��C;�BE;��F;��G;�xH;�I;�I;��I;��I;y�I;��I;R�I;r�I;M�I;XiI;�TI;9CI;34I;�'I;�I;�I;XI;$I;� I;��H;Z�H;��H;��H;�H;�H;h�H;4�H;i�H;�H;�H;��H;��H;X�H;��H;� I;"I;VI;�I;�I;�'I;14I;7CI;�TI;XiI;M�I;t�I;O�I;��I;y�I;��I;��I;�I;�I;�xH;��G;��F;�BE;��C;H�B;�tA;��@;�?;      '�0;�51;Z�2;��4;17;g#:;50=;!@;L�B;
E;��F;�%H;�	I;��I;��I;��I;��I;=�I;��I;>�I;�mI;�WI;�DI;�4I;�'I;wI;EI;�I;{I;s I;s�H;$�H;��H;��H;��H;��H;��H;��H;��H;��H;��H;$�H;r�H;o I;wI;�I;DI;vI;�'I;�4I;�DI;�WI;�mI;>�I;��I;>�I;��I;��I;��I;��I;�	I;�%H;��F;
E;L�B;!@;40=;f#:;-17;��4;X�2;�51;      �;>;��;#�;L ;&;],;�2;`98;0=;�FA;�rD;��F;SJH;�9I;l�I;��I;��I;5�I;ǭI;��I;MpI;�XI;�DI;14I;�&I;gI;+I;�
I;�I;��H;��H;-�H;�H;{�H;��H;O�H;��H;z�H;�H;+�H;��H;��H;�I;�
I;+I;dI;�&I;-4I;�DI;�XI;MpI;��I;ȭI;5�I;��I;��I;l�I;�9I;UJH;��F;�rD;�FA;0=;_98;�2;],;&;R ;%�;��;,;      ���:�:}�:j��:O��::Q ;�e;�V;�#;Me-;�5;i<;�tA;�	E;�eG;v�H;s�I;O�I;3�I;Z�I;]�I;<�I;LpI;�WI;6CI;�2I;�$I;�I;�I;�	I;�I;;�H;��H;C�H;��H;p�H;�H;p�H;��H;C�H;��H;:�H;�I;�	I;�I;�I;�$I;�2I;4CI;�WI;HpI;:�I;Z�I;\�I;1�I;Q�I;s�I;v�H;�eG;�	E;�tA;i<;�5;Oe-;�#;�V;�e;:Q ;{��:j��:y�:�:      ��p� �,��&9�ǳ9܍":��u:"�:��:���:pR;� ;��,;\�6;�)>;/<C;̀F;�lH;�kI;��I;��I;��I;^�I;��I;�mI;�TI;n@I;�/I;g"I;�I;�I;I;�I;��H;��H;��H;��H;�H;��H;��H;��H;��H;�I;I;�I;�I;f"I;�/I;n@I;�TI;�mI;��I;^�I;��I;��I;��I;�kI;�lH;̀F;/<C;�)>;\�6;��,;� ;pR;���:��:&�:��u:��":�ǳ9�&9 �,�      �o&�!�u4�x���尺��O�@8T��v�9��u:7$�:fH�:UD;p#;�71;~;;ȡA;A�E;%H;�VI;U�I;��I;Z�I;ĭI;A�I;UiI;pPI;b<I;;,I;cI;	I;	I;�I;�I;r�H;�H;��H;H�H;��H;�H;q�H;�I;�I;I;I;]I;;,I;`<I;nPI;SiI;<�I;��I;Y�I;��I;W�I;�VI;%H;A�E;ǡA;~;;�71;p#;RD;bH�:3$�:��u:�v�9@8T��O��尺x��w4�)!�      �kٻD�Իfǻ𻱻tV��ln���+���Ժ�1�P�39\m:E�:��;O�;�\,;"�8; �@;�]E;�
H;�VI;��I;3�I;7�I;��I;I�I;�bI;�JI;j7I;(I;�I;rI;I;}I;zI;��H;&�H;��H;&�H;��H;xI;zI;I;rI;�I;(I;h7I;�JI;�bI;I�I;��I;0�I;3�I;��I;�VI;�
H;�]E;��@; �8;�\,;O�;��;E�:\m:p�39�1���Ժ��+�gn�qV��𻱻fǻD�Ի      *yY��|U�:�I�1�7��� ��!�x�Ի�᝻N�T����#��w�9,��:�l�:(;�);Y17;p @;�]E;%H;�kI;Q�I;��I;=�I;r�I;�wI;�ZI;�CI;�1I;�#I;kI;�I;q	I;�I;xI;��H;A�H;��H;xI;�I;p	I;�I;kI;�#I;�1I;�CI;�ZI;�wI;r�I;7�I;��I;O�I;�kI;	%H;]E;r @;V17;�);(;�l�:,��:�w�9�#����N�T��᝻x�Ի�!��� �1�7�:�I��|U�      ��üWl��n����R��8ߓ�R�{��M�|� � �컫���E�B��鰺�6o���u:5��:�R;x�';Y17;�@;E�E;�lH;v�I;��I;��I;O�I;��I;mI;�QI;n<I;�+I;�I;I;�I;'I;�I;kI;�I;kI;�I;'I;�I;I;�I;�+I;i<I;�QI;	mI;��I;N�I;��I;��I;v�I;�lH;E�E;�@;[17;v�';�R;1��:��u:�6o��鰺E�B����� ��|� ��M�R�{�7ߓ��R��n���Xl��      �'�~-$�\��W� ���?ټw��5���_yY��k�޾Ի��tX������%R:��:�R;�);"�8;ΡA;πF;z�H;o�I;��I;��I;�I;M�I;aI;7HI;�4I;�%I;�I;I;�I;�I;SI;�I;SI;�I;�I;I;�I;�%I;�4I;3HI;aI;I�I;�I;��I;��I;l�I;z�H;΀F;ΡA;"�8;�);�R;��:%R:����pX����޾Ի�k�^yY�5���w��?ټ���W�\��~-$�      X+����b̀�,l��Q�#�2�@��������@��s�>�:2���U��G1�x��%R:1��:(;�\,;�;;0<C;�eG;�9I;��I;z�I;�I;��I;�qI;�TI;�>I;}-I;p I;�I;�I;I;SI;RI;SI;I;�I;�I;p I;z-I;�>I;�TI;�qI;��I;�I;z�I;��I;�9I;�eG;/<C;�;;�\,;,;/��:%R:���G1��U��:2��s�>��@��������@�#�2��Q�,l�b̀���      k�ླྀhܽp�н^y��_什P ��l��n<�K���>ټ��G|U�p������D1�������u:�l�:M�;�71;�)>;�	E;VJH;��I;��I;��I;+�I; �I;�bI;�HI;l5I;�&I;�I;�I;I;cI;`
I;cI;I;�I;�I;�&I;j5I;�HI;�bI;�I;*�I;��I;��I;��I;OJH;�	E;�)>;�71;M�;�l�:��u:����G1�����o��F|U��𛼺>ټK���n<�l�P ��_什^y��p�н�hܽ      ��4�h1��&������i�ཅ�������`��'���NR��6�]�p���U��pX��@6o�0��:��;r#;\�6;�tA;��F;�	I;��I;�I;��I;]�I;#qI;�SI;�=I;	-I;� I;�I;I;�I;~I;�I;I;�I;� I;	-I;�=I;�SI;qI;\�I;��I;�I;��I;�	I;��F;�tA;^�6;t#;��;0��:�6o�tX���U��o��6�]�NR����'��`��������i��������&�h1�      �x���o��ń�KUo���O�+�-�{��hܽ[什Ҽx���2�nb��NR��G|U�:2�����鰺�w�9C�:XD;��,;i<;�rD;�%H;�I;��I;&�I;I�I;M�I;_I;KFI;�3I;�%I;I;�I;�I;yI;�I;�I;I;�%I;�3I;JFI;_I;L�I;I�I;"�I;��I;�I;�%H;�rD;i<;��,;XD;C�:�w�9�鰺��:2��G|U�NR��nb����2�Ҽx�[什�hܽ{�+�-���O�KUo�ń��o��      x���྅�Ѿ)����נ�
ń�;�S��#�`O��|n��Ì���2����s�>�޾ԻH�B��#�Pm:hH�:� ;�5;�FA;��F;�I;��I;��I;�I;��I;�jI; OI;O:I;!+I;> I;I;�I;�I;�I;I;< I;+I;O:I;�NI;�jI;��I;�I;��I;��I;�I;��F;�FA;޼5;� ;fH�:Pm:�#�I�B��Իs�>�������2�Ì�|n��`O���#�;�S�
ń��נ�)�����Ѿ��      �3���/��X#��	��A��׌Ⱦ�f��JUo�^1�̰��|n��Ҽx��'��>ټ�@���k��������P�39=$�:qR;Pe-;0=;
E;�xH;ͯI;T�I;��I;F�I;TvI;�WI;�@I;50I;g$I;�I;�I;zI;�I;�I;e$I;40I;�@I;�WI;TvI;C�I;��I;Q�I;ͯI;�xH;
E;0=;Pe-;sR;9$�:P�39��𺬼���k��@���>ټ�'�Ҽx�|n��˰��^1�JUo��f��،Ⱦ�A���	��X#���/�      ���U���V�v��RZ�]58�΂�r��f���hoy�^1�`O��[什�`�L�����`yY� ��O�T��1���u:���:�#;]98;K�B;��G;;mI;R�I;C�I;q�I;��I;`I;DGI;65I;h(I;�I;�I;NI;�I;�I;g(I;45I;BGI;`I;��I;n�I;A�I;O�I;:mI;��G;F�B;[98;�#;���:��u:�1�N�T���`yY����L���`�[什`O��^1�hoy�f���r��΂�]58��RZ�V�v�U���      Ŀ7g��(ﱿ���U����U��X#�v��f���JUo��#��hܽ����n<����5���|� ��᝻��Ժw�9��:�V;�2;!@;��F;"I;<�I;��I;o�I;��I;ChI;QMI;�9I;1,I;�"I;�I;I;�I;�"I;1,I;�9I;PMI;ChI;��I;l�I;��I;;�I; I;��F;!@;�2;�V;��: w�9��Ժ�᝻}� �5�������n<�����hܽ�#�JUo�f���v���X#��U�U������(ﱿ7g��      x�Q9�T��uؿoQ��f_��8�_��X#�r���f��;�S�{�����l�@�w���M�x�Ի��+�08T��:�e;],;70=;�BE;��H;��I;!�I;��I;��I;�oI;	SI;U>I;�/I;�%I;3 I;�I;3 I;�%I;�/I;R>I;	SI;�oI;�I;��I;!�I;��I;��H;�BE;10=;],;�e; �:@8T���+�v�Ի�M�w��@�l�����{�;�S��f��r���X#�8�_�f_��oQ��uؿT��Q9�      �X1���,�i���<��6g��f_���U�΂�׌Ⱦ
ń�+�-�i��P ��$�2�?ټR�{��!�qn��O���u:2Q ;&;c#:;��C;H&H;T�I;g�I;�I;�I;�vI;XI;2BI;�2I;T(I;�"I;� I;�"I;T(I;�2I;/BI;XI;�vI;�I;�I;g�I;S�I;F&H;��C;`#:;&;2Q ;��u:�O�sn��!�S�{�?ټ$�2�P ��i��+�-�
ń�׌Ⱦ΂��U�f_��6g��<�i����,�      d��]]�6K��X1�[f��oQ��U���]58��A���נ���O���_什�Q����8ߓ��� �rV���尺��":W��:V ;&17;N�B;��G;*|I;&�I;��I;�I;}|I;|\I;�EI;^5I;x*I;o$I;k"I;o$I;w*I;\5I;�EI;|\I;}|I;�I;��I;&�I;+|I;��G;N�B;#17;X ;W��:��":�尺rV���� �8ߓ�����Q�_什����O��נ��A��]58�U���oQ���[f��X1�6K��]]�      O������4z���V��X1��<�uؿ����RZ��	�*���KUo����^y��,l�W��R��2�7�𻱻n��ǳ9x��:)�;��4;�tA;�2G;�XI;��I;��I;G�I;8�I;`I;<HI;d7I;>,I;�%I;�#I;�%I;>,I;c7I;;HI;`I;8�I;D�I;��I;��I;�XI;�2G;�tA;��4;,�;x��:�ǳ9p��𻱻2�7��R��W�,l�^y�����KUo�*����	��RZ����uؿ�<��X1���V��4z�����      �o��g^���ē��4z�6K�i��T��(ﱿV�v��X#���Ѿń��&�p�нb̀�]��n���:�I�jǻz4��%9]�:��;O�2;Ӆ@;(�F;';I;4�I;@�I;ײI;��I;�bI;?JI;�8I;�-I;�&I;%I;�&I;�-I;�8I;=JI;�bI;��I;ԲI;?�I;4�I;';I;(�F;Ӆ@;K�2;��;]�: &9z4�jǻ:�I�n���]��b̀�p�н�&�ń���Ѿ�X#�V�v�(ﱿT��i��6K��4z��ē�g^��      r'���X��g^�������]]���,�Q9�7g��U�����/����o��h1��hܽ��~-$�Xl���|U�D�Ի0!� �,���:2;�51;�?;��F;q'I;��I;\�I;w�I;�I;dI;�KI;�9I;f.I;�'I;�%I;�'I;g.I;�9I;KI;dI;�I;t�I;Y�I;��I;p'I;��F;�?;�51;8;��: �,�1!�D�Ի�|U�Yl��~-$����hܽh1��o���ྛ�/�U���7g��Q9���,��]]�����g^���X��   